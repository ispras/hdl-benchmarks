module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 ;
output n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , 
 n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , 
 n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , 
 n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , 
 n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , 
 n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , 
 n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , 
 n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , 
 n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , 
 n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , 
 n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , 
 n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , 
 n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , 
 n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , 
 n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , 
 n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , 
 n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , 
 n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , 
 n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , 
 n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , 
 n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , 
 n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , 
 n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , 
 n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , 
 n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , 
 n379 , n380 , n381 , n382 , n383 ;
wire n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , 
 n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , 
 n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , 
 n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , 
 n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , 
 n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
 n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , 
 n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , 
 n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , 
 n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , 
 n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , 
 n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , 
 n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , 
 n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , 
 n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , 
 n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , 
 n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , 
 n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , 
 n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , 
 n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , 
 n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , 
 n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
 n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
 n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
 n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
 n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , 
 n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , 
 n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , 
 n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , 
 n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , 
 n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , 
 n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , 
 n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , 
 n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , 
 n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , 
 n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
 n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , 
 n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , 
 n1149 , n1150 , n1151 , n168462 , n168463 , n168464 , n168465 , n168466 , n168467 , n168468 , 
 n168469 , n168470 , n168471 , n168472 , n168473 , n168474 , n168475 , n168476 , n168477 , n168478 , 
 n168479 , n168480 , n168481 , n168482 , n168483 , n168484 , n168485 , n168486 , n168487 , n168488 , 
 n168489 , n168490 , n168491 , n168492 , n168493 , n168494 , n168495 , n168496 , n168497 , n168498 , 
 n168499 , n168500 , n168501 , n168502 , n168503 , n168504 , n168505 , n168506 , n168507 , n168508 , 
 n168509 , n168510 , n168511 , n168512 , n168513 , n168514 , n168515 , n168516 , n168517 , n168518 , 
 n168519 , n168520 , n168521 , n168522 , n168523 , n168524 , n168525 , n168526 , n168527 , n168528 , 
 n168529 , n168530 , n168531 , n168532 , n168533 , n168534 , n168535 , n168536 , n168537 , n168538 , 
 n168539 , n168540 , n168541 , n168542 , n168543 , n168544 , n168545 , n168546 , n168547 , n168548 , 
 n168549 , n168550 , n168551 , n168552 , n168553 , n168554 , n168555 , n168556 , n168557 , n168558 , 
 n168559 , n168560 , n168561 , n168562 , n168563 , n168564 , n168565 , n168566 , n168567 , n168568 , 
 n168569 , n168570 , n168571 , n168572 , n168573 , n168574 , n168575 , n168576 , n168577 , n168578 , 
 n168579 , n168580 , n168581 , n168582 , n168583 , n168584 , n168585 , n168586 , n168587 , n168588 , 
 n168589 , n168590 , n168591 , n168592 , n168593 , n168594 , n168595 , n168596 , n168597 , n168598 , 
 n168599 , n168600 , n168601 , n168602 , n168603 , n168604 , n168605 , n168606 , n168607 , n168608 , 
 n168609 , n168610 , n168611 , n168612 , n168613 , n168614 , n168615 , n168616 , n168617 , n168618 , 
 n168619 , n168620 , n168621 , n168622 , n168623 , n168624 , n168625 , n168626 , n168627 , n168628 , 
 n168629 , n168630 , n168631 , n168632 , n168633 , n168634 , n168635 , n168636 , n168637 , n168638 , 
 n168639 , n168640 , n168641 , n168642 , n168643 , n168644 , n168645 , n168646 , n168647 , n168648 , 
 n168649 , n168650 , n168651 , n168652 , n168653 , n168654 , n168655 , n168656 , n168657 , n168658 , 
 n168659 , n168660 , n168661 , n168662 , n168663 , n168664 , n168665 , n168666 , n168667 , n168668 , 
 n168669 , n168670 , n168671 , n168672 , n168673 , n168674 , n168675 , n168676 , n168677 , n168678 , 
 n168679 , n168680 , n168681 , n168682 , n168683 , n168684 , n168685 , n1217 , n168687 , n1219 , 
 n168689 , n168690 , n1222 , n168692 , n1224 , n168694 , n1226 , n168696 , n168697 , n1229 , 
 n168699 , n168700 , n1232 , n1233 , n1234 , n168704 , n1236 , n1237 , n1238 , n168708 , 
 n1240 , n168710 , n168711 , n1243 , n168713 , n168714 , n1246 , n1247 , n168717 , n1249 , 
 n168719 , n168720 , n168721 , n168722 , n1254 , n168724 , n168725 , n1257 , n168727 , n168728 , 
 n1260 , n168730 , n1262 , n1263 , n168733 , n168734 , n1266 , n168736 , n168737 , n1269 , 
 n1270 , n168740 , n168741 , n1273 , n168743 , n1275 , n168745 , n1277 , n168747 , n168748 , 
 n1280 , n168750 , n168751 , n1283 , n1284 , n168754 , n1286 , n168756 , n168757 , n1289 , 
 n168759 , n168760 , n168761 , n168762 , n1294 , n168764 , n168765 , n1297 , n168767 , n168768 , 
 n1300 , n168770 , n1302 , n1303 , n1304 , n1305 , n1306 , n168776 , n168777 , n1309 , 
 n168779 , n168780 , n1312 , n1313 , n1314 , n1315 , n168785 , n168786 , n1318 , n168788 , 
 n1320 , n1321 , n168791 , n1323 , n168793 , n168794 , n1326 , n168796 , n168797 , n1329 , 
 n1330 , n168800 , n168801 , n1333 , n168803 , n168804 , n1336 , n168806 , n168807 , n1339 , 
 n168809 , n1341 , n168811 , n168812 , n1344 , n168814 , n1346 , n1347 , n1348 , n1349 , 
 n1350 , n168820 , n1352 , n168822 , n168823 , n168824 , n168825 , n1357 , n168827 , n168828 , 
 n1360 , n168830 , n1362 , n168832 , n168833 , n1365 , n1366 , n168836 , n1368 , n168838 , 
 n168839 , n168840 , n1372 , n168842 , n168843 , n1375 , n168845 , n168846 , n168847 , n168848 , 
 n1380 , n168850 , n168851 , n1383 , n1384 , n168854 , n168855 , n1387 , n168857 , n1389 , 
 n168859 , n1391 , n168861 , n168862 , n1394 , n1395 , n168865 , n1397 , n168867 , n168868 , 
 n1400 , n168870 , n168871 , n168872 , n168873 , n1405 , n168875 , n168876 , n1408 , n168878 , 
 n168879 , n1411 , n168881 , n168882 , n1414 , n1415 , n168885 , n1417 , n168887 , n168888 , 
 n1420 , n1421 , n168891 , n168892 , n168893 , n168894 , n1426 , n168896 , n1428 , n1429 , 
 n1430 , n168900 , n168901 , n1433 , n168903 , n1435 , n168905 , n168906 , n1438 , n168908 , 
 n1440 , n168910 , n168911 , n168912 , n168913 , n1445 , n168915 , n168916 , n168917 , n1449 , 
 n168919 , n168920 , n1452 , n168922 , n1454 , n1455 , n1456 , n1457 , n1458 , n168928 , 
 n1460 , n168930 , n168931 , n1463 , n168933 , n168934 , n1466 , n168936 , n168937 , n1469 , 
 n1470 , n1471 , n168941 , n1473 , n1474 , n168944 , n168945 , n1477 , n168947 , n168948 , 
 n1480 , n168950 , n168951 , n168952 , n1484 , n168954 , n168955 , n1487 , n1488 , n1489 , 
 n1490 , n168960 , n1492 , n168962 , n1494 , n168964 , n1496 , n1497 , n168967 , n168968 , 
 n1500 , n168970 , n168971 , n1503 , n168973 , n1505 , n168975 , n1507 , n168977 , n168978 , 
 n1510 , n168980 , n168981 , n1513 , n1514 , n168984 , n1516 , n168986 , n168987 , n1519 , 
 n168989 , n168990 , n168991 , n168992 , n1524 , n168994 , n168995 , n1527 , n168997 , n168998 , 
 n1530 , n169000 , n1532 , n1533 , n1534 , n1535 , n1536 , n169006 , n169007 , n1539 , 
 n169009 , n169010 , n1542 , n169012 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
 n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n169025 , n169026 , n1558 , n169028 , 
 n1560 , n1561 , n1562 , n169032 , n1564 , n169034 , n169035 , n1567 , n169037 , n169038 , 
 n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n169048 , 
 n1580 , n1581 , n169051 , n169052 , n1584 , n169054 , n169055 , n1587 , n169057 , n169058 , 
 n169059 , n1591 , n169061 , n169062 , n1594 , n169064 , n1596 , n1597 , n169067 , n169068 , 
 n169069 , n1601 , n169071 , n169072 , n1604 , n169074 , n169075 , n1607 , n169077 , n1609 , 
 n169079 , n1611 , n169081 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
 n1620 , n1621 , n169091 , n1623 , n169093 , n169094 , n169095 , n1627 , n169097 , n1629 , 
 n1630 , n1631 , n169101 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
 n169109 , n169110 , n1642 , n169112 , n169113 , n169114 , n169115 , n1647 , n169117 , n169118 , 
 n1650 , n169120 , n169121 , n169122 , n1654 , n169124 , n169125 , n1657 , n1658 , n169128 , 
 n1660 , n1661 , n169131 , n169132 , n1664 , n169134 , n169135 , n1667 , n1668 , n1669 , 
 n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
 n169149 , n1681 , n169151 , n169152 , n1684 , n169154 , n169155 , n1687 , n1688 , n169158 , 
 n169159 , n1691 , n169161 , n169162 , n169163 , n169164 , n1696 , n169166 , n169167 , n1699 , 
 n169169 , n169170 , n1702 , n169172 , n169173 , n1705 , n169175 , n1707 , n1708 , n1709 , 
 n169179 , n1711 , n169181 , n169182 , n1714 , n1715 , n169185 , n169186 , n1718 , n169188 , 
 n169189 , n1721 , n169191 , n1723 , n169193 , n169194 , n169195 , n169196 , n1728 , n169198 , 
 n169199 , n169200 , n1732 , n169202 , n169203 , n169204 , n169205 , n1737 , n169207 , n169208 , 
 n1740 , n1741 , n1742 , n169212 , n1744 , n1745 , n169215 , n169216 , n1748 , n169218 , 
 n169219 , n1751 , n169221 , n169222 , n1754 , n169224 , n169225 , n1757 , n169227 , n169228 , 
 n1760 , n169230 , n169231 , n1763 , n169233 , n169234 , n1766 , n1767 , n1768 , n1769 , 
 n169239 , n1771 , n169241 , n169242 , n1774 , n1775 , n169245 , n1777 , n169247 , n169248 , 
 n1780 , n169250 , n169251 , n169252 , n169253 , n1785 , n169255 , n169256 , n1788 , n169258 , 
 n169259 , n1791 , n169261 , n169262 , n1794 , n169264 , n169265 , n1797 , n169267 , n169268 , 
 n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n169276 , n1808 , n1809 , 
 n169279 , n169280 , n1812 , n169282 , n169283 , n1815 , n169285 , n169286 , n1818 , n1819 , 
 n169289 , n1821 , n169291 , n169292 , n1824 , n169294 , n1826 , n169296 , n169297 , n1829 , 
 n1830 , n169300 , n169301 , n1833 , n169303 , n169304 , n1836 , n1837 , n169307 , n169308 , 
 n1840 , n169310 , n1842 , n169312 , n1844 , n169314 , n169315 , n1847 , n1848 , n169318 , 
 n1850 , n169320 , n169321 , n169322 , n169323 , n1855 , n169325 , n169326 , n1858 , n169328 , 
 n169329 , n1861 , n169331 , n169332 , n1864 , n169334 , n169335 , n1867 , n169337 , n169338 , 
 n1870 , n1871 , n169341 , n1873 , n169343 , n1875 , n169345 , n169346 , n1878 , n1879 , 
 n169349 , n169350 , n1882 , n169352 , n169353 , n1885 , n169355 , n1887 , n1888 , n169358 , 
 n169359 , n1891 , n169361 , n169362 , n1894 , n169364 , n169365 , n169366 , n169367 , n1899 , 
 n169369 , n169370 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n169377 , n1909 , 
 n1910 , n169380 , n169381 , n1913 , n169383 , n169384 , n1916 , n169386 , n169387 , n1919 , 
 n169389 , n169390 , n1922 , n169392 , n169393 , n1925 , n1926 , n1927 , n1928 , n1929 , 
 n1930 , n169400 , n1932 , n169402 , n169403 , n169404 , n1936 , n169406 , n1938 , n1939 , 
 n169409 , n1941 , n169411 , n169412 , n1944 , n1945 , n169415 , n1947 , n169417 , n169418 , 
 n1950 , n169420 , n169421 , n1953 , n169423 , n169424 , n169425 , n169426 , n1958 , n169428 , 
 n169429 , n1961 , n169431 , n169432 , n1964 , n169434 , n169435 , n1967 , n1968 , n1969 , 
 n169439 , n169440 , n1972 , n169442 , n169443 , n1975 , n169445 , n169446 , n1978 , n169448 , 
 n169449 , n1981 , n169451 , n169452 , n1984 , n1985 , n1986 , n1987 , n1988 , n169458 , 
 n169459 , n1991 , n169461 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
 n2000 , n2001 , n2002 , n169472 , n169473 , n169474 , n2006 , n169476 , n169477 , n2009 , 
 n169479 , n2011 , n2012 , n2013 , n2014 , n169484 , n169485 , n169486 , n2018 , n169488 , 
 n169489 , n2021 , n169491 , n2023 , n2024 , n2025 , n2026 , n169496 , n2028 , n169498 , 
 n2030 , n2031 , n169501 , n169502 , n169503 , n2035 , n169505 , n169506 , n2038 , n169508 , 
 n169509 , n2041 , n169511 , n2043 , n2044 , n2045 , n169515 , n2047 , n2048 , n2049 , 
 n169519 , n169520 , n2052 , n169522 , n2054 , n2055 , n169525 , n169526 , n2058 , n169528 , 
 n2060 , n2061 , n169531 , n2063 , n169533 , n169534 , n2066 , n169536 , n169537 , n2069 , 
 n169539 , n169540 , n2072 , n169542 , n169543 , n2075 , n169545 , n169546 , n2078 , n2079 , 
 n169549 , n169550 , n2082 , n169552 , n169553 , n169554 , n2086 , n169556 , n169557 , n2089 , 
 n169559 , n2091 , n169561 , n2093 , n2094 , n169564 , n169565 , n2097 , n169567 , n169568 , 
 n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n169578 , 
 n2110 , n2111 , n169581 , n169582 , n169583 , n2115 , n169585 , n169586 , n2118 , n169588 , 
 n169589 , n2121 , n169591 , n169592 , n2124 , n169594 , n169595 , n169596 , n2128 , n169598 , 
 n2130 , n169600 , n169601 , n2133 , n169603 , n169604 , n169605 , n169606 , n2138 , n169608 , 
 n169609 , n2141 , n169611 , n2143 , n2144 , n169614 , n169615 , n2147 , n169617 , n169618 , 
 n2150 , n169620 , n169621 , n2153 , n169623 , n169624 , n2156 , n169626 , n169627 , n2159 , 
 n169629 , n169630 , n2162 , n169632 , n169633 , n2165 , n169635 , n169636 , n2168 , n2169 , 
 n169639 , n2171 , n169641 , n169642 , n169643 , n169644 , n2176 , n169646 , n169647 , n2179 , 
 n169649 , n169650 , n2182 , n169652 , n169653 , n2185 , n2186 , n169656 , n2188 , n169658 , 
 n169659 , n2191 , n169661 , n2193 , n169663 , n169664 , n2196 , n2197 , n2198 , n2199 , 
 n2200 , n2201 , n2202 , n169672 , n2204 , n169674 , n2206 , n2207 , n2208 , n2209 , 
 n169679 , n2211 , n169681 , n2213 , n2214 , n169684 , n2216 , n169686 , n169687 , n2219 , 
 n169689 , n169690 , n2222 , n169692 , n2224 , n2225 , n169695 , n2227 , n169697 , n2229 , 
 n2230 , n169700 , n169701 , n2233 , n2234 , n169704 , n169705 , n2237 , n2238 , n169708 , 
 n169709 , n2241 , n2242 , n169712 , n169713 , n2245 , n2246 , n2247 , n169717 , n169718 , 
 n2250 , n2251 , n2252 , n2253 , n2254 , n169724 , n169725 , n169726 , n2258 , n169728 , 
 n169729 , n2261 , n169731 , n2263 , n169733 , n169734 , n2266 , n169736 , n2268 , n2269 , 
 n169739 , n169740 , n169741 , n2273 , n169743 , n169744 , n2276 , n169746 , n169747 , n2279 , 
 n169749 , n169750 , n2282 , n169752 , n2284 , n169754 , n2286 , n2287 , n169757 , n2289 , 
 n169759 , n169760 , n169761 , n169762 , n2294 , n169764 , n169765 , n2297 , n169767 , n169768 , 
 n2300 , n169770 , n169771 , n2303 , n169773 , n169774 , n169775 , n169776 , n2308 , n169778 , 
 n169779 , n2311 , n169781 , n169782 , n2314 , n2315 , n2316 , n2317 , n169787 , n2319 , 
 n169789 , n2321 , n169791 , n2323 , n169793 , n169794 , n2326 , n2327 , n169797 , n2329 , 
 n169799 , n169800 , n2332 , n169802 , n169803 , n169804 , n169805 , n2337 , n169807 , n169808 , 
 n2340 , n169810 , n169811 , n2343 , n169813 , n169814 , n169815 , n2347 , n169817 , n2349 , 
 n2350 , n169820 , n169821 , n2353 , n169823 , n169824 , n2356 , n169826 , n169827 , n2359 , 
 n169829 , n2361 , n169831 , n2363 , n169833 , n169834 , n2366 , n169836 , n169837 , n2369 , 
 n2370 , n169840 , n2372 , n169842 , n169843 , n2375 , n169845 , n169846 , n169847 , n169848 , 
 n2380 , n169850 , n169851 , n2383 , n169853 , n169854 , n2386 , n169856 , n169857 , n2389 , 
 n169859 , n169860 , n2392 , n169862 , n169863 , n2395 , n2396 , n2397 , n169867 , n169868 , 
 n2400 , n169870 , n169871 , n2403 , n2404 , n169874 , n169875 , n2407 , n2408 , n2409 , 
 n169879 , n2411 , n169881 , n169882 , n2414 , n169884 , n2416 , n2417 , n2418 , n169888 , 
 n2420 , n2421 , n169891 , n169892 , n169893 , n2425 , n169895 , n169896 , n2428 , n169898 , 
 n169899 , n2431 , n169901 , n169902 , n169903 , n2435 , n169905 , n2437 , n2438 , n169908 , 
 n2440 , n169910 , n2442 , n169912 , n169913 , n2445 , n169915 , n169916 , n2448 , n169918 , 
 n2450 , n169920 , n2452 , n169922 , n169923 , n2455 , n2456 , n169926 , n2458 , n169928 , 
 n169929 , n2461 , n169931 , n169932 , n169933 , n169934 , n2466 , n169936 , n169937 , n2469 , 
 n169939 , n169940 , n2472 , n169942 , n169943 , n2475 , n169945 , n169946 , n169947 , n2479 , 
 n169949 , n2481 , n169951 , n169952 , n2484 , n2485 , n169955 , n2487 , n169957 , n169958 , 
 n2490 , n169960 , n2492 , n169962 , n169963 , n2495 , n169965 , n169966 , n169967 , n2499 , 
 n169969 , n2501 , n2502 , n169972 , n169973 , n2505 , n169975 , n169976 , n2508 , n169978 , 
 n169979 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n169986 , n2518 , n169988 , 
 n169989 , n2521 , n169991 , n169992 , n2524 , n169994 , n2526 , n2527 , n169997 , n2529 , 
 n169999 , n170000 , n2532 , n170002 , n2534 , n170004 , n2536 , n2537 , n170007 , n170008 , 
 n2540 , n170010 , n170011 , n2543 , n170013 , n170014 , n170015 , n2547 , n170017 , n2549 , 
 n170019 , n170020 , n2552 , n2553 , n2554 , n170024 , n170025 , n2557 , n170027 , n170028 , 
 n2560 , n170030 , n170031 , n2563 , n170033 , n2565 , n2566 , n170036 , n2568 , n2569 , 
 n170039 , n170040 , n2572 , n170042 , n170043 , n2575 , n170045 , n170046 , n2578 , n170048 , 
 n170049 , n2581 , n170051 , n2583 , n2584 , n170054 , n170055 , n170056 , n2588 , n170058 , 
 n170059 , n2591 , n170061 , n2593 , n2594 , n170064 , n170065 , n2597 , n170067 , n170068 , 
 n2600 , n170070 , n170071 , n2603 , n170073 , n2605 , n170075 , n170076 , n2608 , n170078 , 
 n170079 , n170080 , n170081 , n2613 , n170083 , n170084 , n2616 , n170086 , n2618 , n2619 , 
 n170089 , n170090 , n2622 , n170092 , n170093 , n2625 , n170095 , n170096 , n2628 , n170098 , 
 n2630 , n170100 , n170101 , n2633 , n170103 , n170104 , n170105 , n170106 , n2638 , n170108 , 
 n170109 , n2641 , n170111 , n170112 , n2644 , n170114 , n170115 , n2647 , n170117 , n170118 , 
 n2650 , n2651 , n170121 , n170122 , n2654 , n2655 , n2656 , n170126 , n170127 , n2659 , 
 n2660 , n2661 , n170131 , n170132 , n2664 , n170134 , n170135 , n2667 , n170137 , n170138 , 
 n2670 , n170140 , n2672 , n2673 , n170143 , n170144 , n2676 , n170146 , n170147 , n2679 , 
 n170149 , n170150 , n170151 , n2683 , n170153 , n170154 , n2686 , n170156 , n2688 , n2689 , 
 n170159 , n170160 , n2692 , n170162 , n170163 , n2695 , n170165 , n2697 , n170167 , n170168 , 
 n2700 , n170170 , n170171 , n2703 , n170173 , n2705 , n2706 , n170176 , n170177 , n2709 , 
 n170179 , n170180 , n2712 , n170182 , n2714 , n2715 , n2716 , n2717 , n2718 , n170188 , 
 n170189 , n2721 , n170191 , n2723 , n2724 , n170194 , n170195 , n2727 , n170197 , n2729 , 
 n170199 , n2731 , n170201 , n2733 , n2734 , n2735 , n2736 , n2737 , n170207 , n2739 , 
 n2740 , n170210 , n170211 , n2743 , n170213 , n170214 , n2746 , n170216 , n170217 , n2749 , 
 n170219 , n170220 , n2752 , n170222 , n170223 , n2755 , n2756 , n2757 , n170227 , n2759 , 
 n2760 , n170230 , n170231 , n2763 , n170233 , n170234 , n2766 , n170236 , n170237 , n2769 , 
 n2770 , n2771 , n170241 , n2773 , n170243 , n170244 , n2776 , n170246 , n170247 , n2779 , 
 n170249 , n2781 , n2782 , n170252 , n170253 , n2785 , n170255 , n170256 , n2788 , n170258 , 
 n170259 , n2791 , n170261 , n170262 , n2794 , n170264 , n170265 , n2797 , n170267 , n2799 , 
 n2800 , n170270 , n170271 , n2803 , n170273 , n170274 , n2806 , n170276 , n170277 , n2809 , 
 n2810 , n170280 , n170281 , n2813 , n170283 , n170284 , n2816 , n170286 , n170287 , n2819 , 
 n170289 , n2821 , n2822 , n2823 , n170293 , n170294 , n2826 , n170296 , n170297 , n2829 , 
 n170299 , n170300 , n2832 , n170302 , n170303 , n2835 , n170305 , n2837 , n2838 , n2839 , 
 n2840 , n2841 , n2842 , n2843 , n170313 , n2845 , n2846 , n2847 , n170317 , n2849 , 
 n2850 , n2851 , n170321 , n170322 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
 n170329 , n2861 , n170331 , n170332 , n2864 , n2865 , n2866 , n2867 , n170337 , n2869 , 
 n170339 , n2871 , n170341 , n2873 , n2874 , n170344 , n170345 , n2877 , n2878 , n170348 , 
 n170349 , n170350 , n2882 , n2883 , n170353 , n2885 , n2886 , n170356 , n170357 , n2889 , 
 n170359 , n170360 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n170367 , n170368 , 
 n2900 , n2901 , n170371 , n2903 , n2904 , n170374 , n170375 , n2907 , n170377 , n2909 , 
 n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n170385 , n2917 , n170387 , n170388 , 
 n2920 , n170390 , n170391 , n170392 , n170393 , n2925 , n170395 , n170396 , n2928 , n170398 , 
 n2930 , n170400 , n2932 , n2933 , n2934 , n2935 , n170405 , n2937 , n170407 , n170408 , 
 n2940 , n170410 , n170411 , n2943 , n170413 , n170414 , n170415 , n2947 , n170417 , n2949 , 
 n170419 , n170420 , n2952 , n2953 , n170423 , n2955 , n170425 , n2957 , n170427 , n170428 , 
 n2960 , n170430 , n170431 , n2963 , n2964 , n2965 , n2966 , n2967 , n170437 , n170438 , 
 n2970 , n170440 , n170441 , n2973 , n2974 , n2975 , n2976 , n170446 , n2978 , n2979 , 
 n2980 , n2981 , n2982 , n170452 , n170453 , n2985 , n170455 , n170456 , n2988 , n2989 , 
 n2990 , n2991 , n170461 , n170462 , n2994 , n2995 , n2996 , n2997 , n170467 , n170468 , 
 n3000 , n3001 , n3002 , n3003 , n170473 , n170474 , n3006 , n3007 , n3008 , n3009 , 
 n3010 , n170480 , n170481 , n3013 , n170483 , n170484 , n3016 , n3017 , n3018 , n3019 , 
 n170489 , n170490 , n3022 , n170492 , n3024 , n3025 , n170495 , n170496 , n3028 , n170498 , 
 n3030 , n3031 , n170501 , n3033 , n170503 , n3035 , n170505 , n170506 , n3038 , n170508 , 
 n170509 , n3041 , n170511 , n3043 , n170513 , n3045 , n3046 , n170516 , n3048 , n170518 , 
 n3050 , n170520 , n170521 , n3053 , n170523 , n170524 , n3056 , n170526 , n170527 , n3059 , 
 n3060 , n170530 , n170531 , n3063 , n3064 , n170534 , n170535 , n170536 , n3068 , n170538 , 
 n3070 , n3071 , n170541 , n3073 , n170543 , n3075 , n170545 , n170546 , n3078 , n170548 , 
 n170549 , n3081 , n170551 , n170552 , n3084 , n170554 , n3086 , n170556 , n3088 , n3089 , 
 n170559 , n170560 , n3092 , n170562 , n170563 , n3095 , n170565 , n170566 , n170567 , n170568 , 
 n3100 , n170570 , n170571 , n3103 , n170573 , n170574 , n3106 , n170576 , n170577 , n3109 , 
 n170579 , n3111 , n3112 , n170582 , n170583 , n170584 , n3116 , n170586 , n170587 , n3119 , 
 n170589 , n170590 , n3122 , n170592 , n3124 , n170594 , n3126 , n170596 , n3128 , n3129 , 
 n170599 , n170600 , n170601 , n3133 , n170603 , n170604 , n3136 , n170606 , n170607 , n3139 , 
 n170609 , n3141 , n170611 , n3143 , n170613 , n170614 , n3146 , n170616 , n170617 , n3149 , 
 n3150 , n3151 , n3152 , n3153 , n170623 , n3155 , n170625 , n170626 , n3158 , n3159 , 
 n3160 , n170630 , n170631 , n3163 , n170633 , n3165 , n170635 , n3167 , n3168 , n170638 , 
 n170639 , n3171 , n170641 , n170642 , n170643 , n3175 , n170645 , n170646 , n3178 , n170648 , 
 n170649 , n170650 , n3182 , n170652 , n3184 , n3185 , n170655 , n170656 , n170657 , n3189 , 
 n170659 , n170660 , n3192 , n170662 , n170663 , n3195 , n170665 , n170666 , n3198 , n3199 , 
 n170669 , n170670 , n3202 , n170672 , n3204 , n3205 , n170675 , n3207 , n170677 , n3209 , 
 n3210 , n170680 , n3212 , n170682 , n170683 , n170684 , n3216 , n170686 , n3218 , n3219 , 
 n3220 , n170690 , n170691 , n170692 , n3224 , n170694 , n170695 , n3227 , n170697 , n170698 , 
 n3230 , n170700 , n170701 , n3233 , n170703 , n3235 , n3236 , n170706 , n3238 , n170708 , 
 n170709 , n170710 , n170711 , n3243 , n170713 , n170714 , n3246 , n170716 , n170717 , n3249 , 
 n170719 , n3251 , n170721 , n3253 , n170723 , n3255 , n3256 , n170726 , n170727 , n170728 , 
 n3260 , n170730 , n170731 , n3263 , n170733 , n170734 , n3266 , n170736 , n3268 , n170738 , 
 n3270 , n3271 , n3272 , n3273 , n3274 , n170744 , n170745 , n3277 , n170747 , n170748 , 
 n3280 , n3281 , n3282 , n3283 , n170753 , n170754 , n3286 , n3287 , n3288 , n3289 , 
 n3290 , n170760 , n170761 , n3293 , n170763 , n170764 , n170765 , n170766 , n3298 , n170768 , 
 n170769 , n170770 , n3302 , n170772 , n3304 , n170774 , n3306 , n170776 , n3308 , n170778 , 
 n3310 , n170780 , n3312 , n3313 , n170783 , n170784 , n3316 , n170786 , n170787 , n170788 , 
 n3320 , n170790 , n170791 , n3323 , n170793 , n170794 , n3326 , n3327 , n170797 , n170798 , 
 n3330 , n3331 , n170801 , n170802 , n3334 , n3335 , n3336 , n3337 , n170807 , n170808 , 
 n3340 , n3341 , n3342 , n3343 , n170813 , n170814 , n3346 , n170816 , n170817 , n3349 , 
 n170819 , n3351 , n3352 , n170822 , n3354 , n170824 , n3356 , n3357 , n3358 , n170828 , 
 n170829 , n3361 , n170831 , n3363 , n170833 , n3365 , n3366 , n3367 , n3368 , n3369 , 
 n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
 n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
 n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
 n170869 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n170876 , n3408 , n3409 , 
 n3410 , n3411 , n170881 , n170882 , n3414 , n3415 , n3416 , n3417 , n170887 , n170888 , 
 n3420 , n170890 , n3422 , n170892 , n3424 , n3425 , n170895 , n170896 , n170897 , n3429 , 
 n170899 , n170900 , n3432 , n170902 , n170903 , n3435 , n170905 , n170906 , n3438 , n170908 , 
 n3440 , n3441 , n170911 , n170912 , n170913 , n3445 , n170915 , n170916 , n3448 , n170918 , 
 n170919 , n3451 , n170921 , n3453 , n170923 , n3455 , n170925 , n3457 , n3458 , n170928 , 
 n3460 , n170930 , n3462 , n170932 , n170933 , n3465 , n170935 , n3467 , n170937 , n170938 , 
 n3470 , n170940 , n3472 , n3473 , n170943 , n170944 , n170945 , n3477 , n170947 , n170948 , 
 n3480 , n170950 , n170951 , n3483 , n170953 , n170954 , n170955 , n170956 , n3488 , n170958 , 
 n170959 , n3491 , n170961 , n170962 , n3494 , n170964 , n3496 , n3497 , n170967 , n3499 , 
 n3500 , n170970 , n3502 , n170972 , n170973 , n170974 , n170975 , n3507 , n170977 , n170978 , 
 n3510 , n170980 , n170981 , n3513 , n170983 , n170984 , n3516 , n170986 , n3518 , n170988 , 
 n3520 , n170990 , n170991 , n3523 , n3524 , n170994 , n170995 , n170996 , n3528 , n170998 , 
 n170999 , n3531 , n171001 , n171002 , n3534 , n171004 , n171005 , n3537 , n171007 , n171008 , 
 n3540 , n3541 , n171011 , n3543 , n171013 , n3545 , n3546 , n171016 , n171017 , n171018 , 
 n3550 , n171020 , n171021 , n3553 , n171023 , n3555 , n171025 , n3557 , n171027 , n3559 , 
 n171029 , n171030 , n3562 , n3563 , n171033 , n171034 , n171035 , n3567 , n171037 , n171038 , 
 n3570 , n171040 , n171041 , n3573 , n171043 , n3575 , n171045 , n3577 , n171047 , n3579 , 
 n171049 , n171050 , n3582 , n3583 , n171053 , n3585 , n171055 , n171056 , n171057 , n171058 , 
 n3590 , n171060 , n171061 , n3593 , n171063 , n171064 , n3596 , n171066 , n3598 , n171068 , 
 n3600 , n171070 , n171071 , n3603 , n171073 , n171074 , n3606 , n3607 , n3608 , n3609 , 
 n3610 , n171080 , n171081 , n3613 , n171083 , n171084 , n3616 , n3617 , n3618 , n3619 , 
 n3620 , n171090 , n171091 , n3623 , n171093 , n171094 , n3626 , n3627 , n3628 , n171098 , 
 n171099 , n3631 , n3632 , n3633 , n3634 , n171104 , n171105 , n3637 , n3638 , n3639 , 
 n3640 , n3641 , n171111 , n171112 , n3644 , n3645 , n3646 , n3647 , n171117 , n171118 , 
 n3650 , n3651 , n3652 , n3653 , n3654 , n171124 , n171125 , n3657 , n171127 , n171128 , 
 n171129 , n171130 , n3662 , n171132 , n171133 , n171134 , n3666 , n171136 , n3668 , n3669 , 
 n171139 , n171140 , n3672 , n171142 , n171143 , n3675 , n171145 , n171146 , n3678 , n171148 , 
 n3680 , n3681 , n3682 , n3683 , n171153 , n3685 , n3686 , n171156 , n171157 , n171158 , 
 n3690 , n171160 , n171161 , n3693 , n171163 , n171164 , n3696 , n171166 , n171167 , n3699 , 
 n171169 , n171170 , n171171 , n3703 , n171173 , n3705 , n3706 , n171176 , n171177 , n3709 , 
 n171179 , n3711 , n171181 , n171182 , n3714 , n171184 , n171185 , n3717 , n3718 , n3719 , 
 n3720 , n3721 , n171191 , n171192 , n3724 , n171194 , n171195 , n3727 , n171197 , n171198 , 
 n3730 , n3731 , n3732 , n3733 , n3734 , n171204 , n171205 , n3737 , n171207 , n171208 , 
 n171209 , n3741 , n171211 , n3743 , n3744 , n171214 , n171215 , n171216 , n3748 , n171218 , 
 n171219 , n3751 , n171221 , n171222 , n3754 , n171224 , n171225 , n171226 , n3758 , n3759 , 
 n3760 , n3761 , n3762 , n3763 , n3764 , n171234 , n3766 , n3767 , n171237 , n171238 , 
 n171239 , n3771 , n171241 , n171242 , n3774 , n171244 , n171245 , n3777 , n171247 , n171248 , 
 n3780 , n171250 , n171251 , n3783 , n3784 , n171254 , n3786 , n3787 , n171257 , n171258 , 
 n171259 , n3791 , n171261 , n3793 , n3794 , n171264 , n171265 , n171266 , n3798 , n171268 , 
 n171269 , n3801 , n171271 , n171272 , n3804 , n171274 , n171275 , n3807 , n3808 , n171278 , 
 n3810 , n171280 , n171281 , n3813 , n3814 , n171284 , n3816 , n3817 , n3818 , n171288 , 
 n171289 , n3821 , n171291 , n171292 , n171293 , n171294 , n3826 , n171296 , n171297 , n3829 , 
 n171299 , n3831 , n3832 , n3833 , n3834 , n3835 , n171305 , n171306 , n171307 , n3839 , 
 n171309 , n171310 , n3842 , n171312 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
 n3850 , n3851 , n3852 , n171322 , n171323 , n3855 , n171325 , n171326 , n3858 , n171328 , 
 n3860 , n171330 , n171331 , n171332 , n171333 , n3865 , n171335 , n171336 , n3868 , n171338 , 
 n171339 , n3871 , n3872 , n171342 , n3874 , n3875 , n171345 , n3877 , n171347 , n3879 , 
 n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n171355 , n171356 , n3888 , n171358 , 
 n3890 , n3891 , n171361 , n171362 , n171363 , n3895 , n171365 , n171366 , n3898 , n171368 , 
 n171369 , n3901 , n171371 , n171372 , n171373 , n3905 , n171375 , n3907 , n3908 , n171378 , 
 n171379 , n171380 , n3912 , n171382 , n171383 , n3915 , n171385 , n171386 , n3918 , n171388 , 
 n171389 , n3921 , n171391 , n3923 , n171393 , n3925 , n3926 , n171396 , n171397 , n171398 , 
 n3930 , n171400 , n171401 , n3933 , n171403 , n171404 , n3936 , n171406 , n171407 , n3939 , 
 n171409 , n171410 , n3942 , n3943 , n171413 , n3945 , n171415 , n171416 , n3948 , n3949 , 
 n171419 , n171420 , n171421 , n3953 , n171423 , n3955 , n171425 , n3957 , n3958 , n171428 , 
 n3960 , n171430 , n171431 , n3963 , n3964 , n171434 , n171435 , n3967 , n171437 , n3969 , 
 n171439 , n171440 , n3972 , n171442 , n171443 , n3975 , n171445 , n3977 , n3978 , n171448 , 
 n171449 , n3981 , n171451 , n3983 , n171453 , n171454 , n3986 , n171456 , n171457 , n3989 , 
 n171459 , n3991 , n3992 , n3993 , n3994 , n3995 , n171465 , n3997 , n171467 , n3999 , 
 n4000 , n4001 , n4002 , n4003 , n171473 , n171474 , n4006 , n171476 , n171477 , n4009 , 
 n171479 , n4011 , n171481 , n4013 , n4014 , n4015 , n4016 , n171486 , n4018 , n171488 , 
 n171489 , n4021 , n171491 , n4023 , n171493 , n4025 , n4026 , n171496 , n171497 , n171498 , 
 n4030 , n171500 , n171501 , n4033 , n171503 , n171504 , n4036 , n171506 , n171507 , n4039 , 
 n171509 , n4041 , n4042 , n171512 , n171513 , n171514 , n4046 , n171516 , n171517 , n4049 , 
 n171519 , n171520 , n4052 , n171522 , n4054 , n171524 , n4056 , n171526 , n4058 , n171528 , 
 n4060 , n4061 , n171531 , n4063 , n171533 , n4065 , n4066 , n171536 , n4068 , n171538 , 
 n4070 , n171540 , n171541 , n4073 , n171543 , n171544 , n4076 , n4077 , n171547 , n171548 , 
 n171549 , n4081 , n171551 , n171552 , n4084 , n171554 , n171555 , n4087 , n171557 , n171558 , 
 n171559 , n4091 , n171561 , n4093 , n4094 , n171564 , n171565 , n171566 , n4098 , n171568 , 
 n171569 , n4101 , n171571 , n171572 , n4104 , n171574 , n171575 , n4107 , n171577 , n4109 , 
 n171579 , n4111 , n4112 , n171582 , n4114 , n171584 , n4116 , n171586 , n171587 , n4119 , 
 n171589 , n171590 , n4122 , n171592 , n171593 , n4125 , n4126 , n171596 , n171597 , n4129 , 
 n4130 , n171600 , n171601 , n4133 , n4134 , n171604 , n171605 , n4137 , n4138 , n171608 , 
 n171609 , n4141 , n4142 , n4143 , n171613 , n171614 , n4146 , n171616 , n4148 , n171618 , 
 n4150 , n171620 , n4152 , n4153 , n4154 , n4155 , n4156 , n171626 , n171627 , n4159 , 
 n171629 , n171630 , n4162 , n171632 , n171633 , n4165 , n171635 , n171636 , n4168 , n171638 , 
 n171639 , n4171 , n4172 , n171642 , n171643 , n4175 , n171645 , n171646 , n4178 , n171648 , 
 n171649 , n4181 , n171651 , n171652 , n4184 , n171654 , n171655 , n4187 , n171657 , n171658 , 
 n4190 , n171660 , n4192 , n171662 , n171663 , n4195 , n171665 , n171666 , n4198 , n4199 , 
 n4200 , n171670 , n4202 , n171672 , n4204 , n4205 , n171675 , n171676 , n4208 , n4209 , 
 n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
 n4220 , n4221 , n4222 , n171692 , n171693 , n171694 , n4226 , n171696 , n171697 , n4229 , 
 n171699 , n171700 , n4232 , n171702 , n171703 , n171704 , n4236 , n171706 , n171707 , n4239 , 
 n4240 , n171710 , n171711 , n4243 , n171713 , n171714 , n4246 , n171716 , n171717 , n171718 , 
 n171719 , n4251 , n171721 , n171722 , n4254 , n171724 , n4256 , n4257 , n171727 , n171728 , 
 n4260 , n171730 , n171731 , n4263 , n171733 , n171734 , n4266 , n4267 , n4268 , n4269 , 
 n4270 , n4271 , n4272 , n4273 , n171743 , n171744 , n171745 , n4277 , n171747 , n4279 , 
 n171749 , n171750 , n171751 , n4283 , n171753 , n4285 , n171755 , n4287 , n171757 , n171758 , 
 n4290 , n4291 , n4292 , n171762 , n171763 , n4295 , n4296 , n171766 , n171767 , n4299 , 
 n4300 , n4301 , n171771 , n171772 , n4304 , n4305 , n4306 , n171776 , n171777 , n4309 , 
 n4310 , n4311 , n171781 , n171782 , n171783 , n171784 , n4316 , n171786 , n171787 , n4319 , 
 n171789 , n4321 , n4322 , n171792 , n171793 , n4325 , n171795 , n171796 , n4328 , n171798 , 
 n171799 , n171800 , n171801 , n4333 , n171803 , n171804 , n4336 , n4337 , n171807 , n4339 , 
 n4340 , n171810 , n171811 , n4343 , n171813 , n171814 , n4346 , n171816 , n171817 , n4349 , 
 n171819 , n171820 , n4352 , n171822 , n171823 , n4355 , n171825 , n4357 , n4358 , n171828 , 
 n171829 , n4361 , n171831 , n171832 , n4364 , n171834 , n171835 , n4367 , n4368 , n4369 , 
 n171839 , n171840 , n4372 , n4373 , n4374 , n171844 , n171845 , n4377 , n4378 , n4379 , 
 n171849 , n171850 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
 n4390 , n4391 , n4392 , n4393 , n171863 , n4395 , n4396 , n4397 , n4398 , n4399 , 
 n171869 , n171870 , n4402 , n171872 , n4404 , n4405 , n4406 , n171876 , n4408 , n171878 , 
 n4410 , n171880 , n171881 , n4413 , n4414 , n171884 , n171885 , n4417 , n171887 , n171888 , 
 n4420 , n171890 , n4422 , n4423 , n171893 , n171894 , n4426 , n171896 , n4428 , n171898 , 
 n4430 , n171900 , n4432 , n4433 , n171903 , n171904 , n4436 , n171906 , n171907 , n4439 , 
 n171909 , n171910 , n4442 , n171912 , n4444 , n4445 , n171915 , n171916 , n4448 , n171918 , 
 n171919 , n4451 , n171921 , n4453 , n4454 , n171924 , n171925 , n4457 , n171927 , n171928 , 
 n4460 , n171930 , n171931 , n4463 , n171933 , n171934 , n4466 , n171936 , n171937 , n4469 , 
 n171939 , n4471 , n4472 , n171942 , n171943 , n4475 , n171945 , n171946 , n4478 , n171948 , 
 n171949 , n4481 , n4482 , n171952 , n171953 , n4485 , n171955 , n171956 , n4488 , n171958 , 
 n171959 , n4491 , n171961 , n4493 , n4494 , n171964 , n171965 , n4497 , n171967 , n171968 , 
 n4500 , n171970 , n171971 , n4503 , n171973 , n171974 , n4506 , n171976 , n4508 , n171978 , 
 n171979 , n4511 , n171981 , n171982 , n4514 , n171984 , n4516 , n4517 , n171987 , n171988 , 
 n4520 , n171990 , n171991 , n4523 , n171993 , n171994 , n171995 , n171996 , n4528 , n171998 , 
 n171999 , n4531 , n172001 , n4533 , n4534 , n172004 , n172005 , n4537 , n172007 , n172008 , 
 n4540 , n172010 , n172011 , n4543 , n4544 , n4545 , n4546 , n172016 , n172017 , n4549 , 
 n172019 , n4551 , n4552 , n172022 , n4554 , n4555 , n4556 , n172026 , n4558 , n4559 , 
 n4560 , n172030 , n4562 , n172032 , n172033 , n172034 , n172035 , n4567 , n172037 , n172038 , 
 n4570 , n172040 , n172041 , n4573 , n4574 , n4575 , n172045 , n172046 , n4578 , n172048 , 
 n4580 , n4581 , n172051 , n4583 , n172053 , n4585 , n172055 , n4587 , n4588 , n172058 , 
 n172059 , n4591 , n4592 , n172062 , n4594 , n172064 , n4596 , n4597 , n4598 , n4599 , 
 n4600 , n4601 , n4602 , n4603 , n172073 , n4605 , n172075 , n4607 , n4608 , n4609 , 
 n172079 , n4611 , n4612 , n4613 , n4614 , n4615 , n172085 , n4617 , n172087 , n172088 , 
 n4620 , n172090 , n4622 , n172092 , n4624 , n172094 , n4626 , n4627 , n4628 , n4629 , 
 n4630 , n4631 , n4632 , n4633 , n4634 , n172104 , n4636 , n4637 , n4638 , n4639 , 
 n172109 , n172110 , n4642 , n172112 , n172113 , n172114 , n4646 , n172116 , n172117 , n4649 , 
 n172119 , n172120 , n4652 , n172122 , n172123 , n4655 , n172125 , n172126 , n4658 , n172128 , 
 n4660 , n172130 , n4662 , n4663 , n172133 , n172134 , n4666 , n4667 , n172137 , n172138 , 
 n172139 , n4671 , n172141 , n172142 , n4674 , n4675 , n4676 , n172146 , n4678 , n4679 , 
 n4680 , n172150 , n4682 , n172152 , n172153 , n4685 , n4686 , n4687 , n172157 , n4689 , 
 n4690 , n4691 , n4692 , n172162 , n172163 , n172164 , n4696 , n4697 , n172167 , n172168 , 
 n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
 n172179 , n4711 , n4712 , n172182 , n172183 , n4715 , n4716 , n4717 , n4718 , n4719 , 
 n172189 , n172190 , n4722 , n4723 , n4724 , n172194 , n4726 , n4727 , n172197 , n172198 , 
 n4730 , n172200 , n172201 , n172202 , n4734 , n172204 , n4736 , n4737 , n4738 , n4739 , 
 n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n172215 , n4747 , n4748 , n4749 , 
 n4750 , n4751 , n4752 , n4753 , n172223 , n172224 , n4756 , n172226 , n172227 , n4759 , 
 n172229 , n4761 , n4762 , n172232 , n172233 , n4765 , n172235 , n172236 , n4768 , n172238 , 
 n172239 , n172240 , n172241 , n4773 , n172243 , n172244 , n4776 , n172246 , n4778 , n4779 , 
 n172249 , n172250 , n4782 , n172252 , n172253 , n4785 , n172255 , n172256 , n4788 , n4789 , 
 n172259 , n4791 , n172261 , n4793 , n4794 , n4795 , n172265 , n4797 , n172267 , n172268 , 
 n4800 , n4801 , n4802 , n172272 , n172273 , n4805 , n172275 , n172276 , n4808 , n172278 , 
 n4810 , n172280 , n4812 , n4813 , n172283 , n172284 , n4816 , n172286 , n172287 , n4819 , 
 n172289 , n172290 , n4822 , n172292 , n4824 , n172294 , n4826 , n4827 , n172297 , n172298 , 
 n4830 , n172300 , n172301 , n4833 , n172303 , n172304 , n4836 , n172306 , n172307 , n4839 , 
 n172309 , n172310 , n4842 , n172312 , n4844 , n4845 , n172315 , n172316 , n4848 , n172318 , 
 n172319 , n4851 , n172321 , n172322 , n4854 , n4855 , n4856 , n172326 , n4858 , n4859 , 
 n172329 , n4861 , n4862 , n172332 , n4864 , n172334 , n4866 , n172336 , n172337 , n4869 , 
 n172339 , n172340 , n172341 , n172342 , n4874 , n172344 , n172345 , n4877 , n172347 , n4879 , 
 n4880 , n172350 , n172351 , n4883 , n172353 , n172354 , n4886 , n172356 , n172357 , n4889 , 
 n4890 , n172360 , n4892 , n172362 , n4894 , n4895 , n172365 , n172366 , n4898 , n172368 , 
 n172369 , n4901 , n172371 , n172372 , n4904 , n4905 , n4906 , n172376 , n172377 , n172378 , 
 n172379 , n4911 , n172381 , n172382 , n4914 , n172384 , n4916 , n4917 , n172387 , n172388 , 
 n4920 , n172390 , n172391 , n4923 , n172393 , n172394 , n172395 , n172396 , n4928 , n172398 , 
 n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n172405 , n4937 , n4938 , n4939 , 
 n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n172415 , n4947 , n4948 , n4949 , 
 n172419 , n172420 , n4952 , n4953 , n4954 , n172424 , n172425 , n4957 , n4958 , n4959 , 
 n172429 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
 n4970 , n172440 , n4972 , n4973 , n4974 , n172444 , n172445 , n4977 , n4978 , n4979 , 
 n172449 , n172450 , n4982 , n4983 , n172453 , n4985 , n172455 , n4987 , n172457 , n4989 , 
 n4990 , n172460 , n172461 , n4993 , n4994 , n172464 , n172465 , n4997 , n4998 , n172468 , 
 n5000 , n172470 , n172471 , n5003 , n172473 , n5005 , n172475 , n172476 , n5008 , n172478 , 
 n172479 , n5011 , n5012 , n5013 , n172483 , n172484 , n5016 , n172486 , n5018 , n172488 , 
 n5020 , n5021 , n172491 , n172492 , n5024 , n172494 , n172495 , n172496 , n172497 , n5029 , 
 n172499 , n5031 , n5032 , n172502 , n172503 , n172504 , n5036 , n172506 , n172507 , n5039 , 
 n172509 , n5041 , n5042 , n172512 , n172513 , n5045 , n172515 , n172516 , n5048 , n172518 , 
 n172519 , n172520 , n172521 , n5053 , n172523 , n5055 , n172525 , n172526 , n172527 , n172528 , 
 n5060 , n172530 , n172531 , n172532 , n5064 , n172534 , n172535 , n172536 , n172537 , n5069 , 
 n172539 , n172540 , n5072 , n172542 , n5074 , n5075 , n172545 , n172546 , n5078 , n172548 , 
 n172549 , n5081 , n172551 , n172552 , n5084 , n172554 , n172555 , n5087 , n172557 , n172558 , 
 n5090 , n172560 , n172561 , n5093 , n172563 , n5095 , n5096 , n172566 , n172567 , n5099 , 
 n172569 , n172570 , n5102 , n172572 , n172573 , n5105 , n172575 , n5107 , n172577 , n5109 , 
 n5110 , n172580 , n5112 , n172582 , n172583 , n172584 , n5116 , n172586 , n172587 , n5119 , 
 n172589 , n172590 , n5122 , n5123 , n172593 , n5125 , n172595 , n5127 , n5128 , n172598 , 
 n172599 , n5131 , n172601 , n172602 , n5134 , n172604 , n172605 , n5137 , n5138 , n5139 , 
 n172609 , n172610 , n5142 , n5143 , n5144 , n172614 , n172615 , n5147 , n5148 , n172618 , 
 n172619 , n5151 , n5152 , n5153 , n172623 , n172624 , n5156 , n5157 , n172627 , n172628 , 
 n5160 , n5161 , n5162 , n172632 , n172633 , n5165 , n5166 , n5167 , n172637 , n172638 , 
 n5170 , n5171 , n5172 , n172642 , n172643 , n5175 , n5176 , n5177 , n5178 , n5179 , 
 n5180 , n172650 , n172651 , n5183 , n172653 , n172654 , n5186 , n172656 , n5188 , n5189 , 
 n172659 , n172660 , n5192 , n172662 , n172663 , n5195 , n172665 , n5197 , n172667 , n172668 , 
 n5200 , n172670 , n172671 , n5203 , n172673 , n5205 , n5206 , n172676 , n172677 , n5209 , 
 n172679 , n172680 , n5212 , n172682 , n5214 , n5215 , n5216 , n172686 , n172687 , n5219 , 
 n172689 , n172690 , n5222 , n172692 , n5224 , n5225 , n172695 , n172696 , n5228 , n172698 , 
 n172699 , n5231 , n172701 , n172702 , n5234 , n172704 , n5236 , n172706 , n5238 , n5239 , 
 n172709 , n172710 , n5242 , n172712 , n172713 , n5245 , n172715 , n172716 , n5248 , n172718 , 
 n172719 , n5251 , n172721 , n172722 , n5254 , n172724 , n5256 , n5257 , n172727 , n172728 , 
 n5260 , n172730 , n172731 , n5263 , n172733 , n172734 , n5266 , n5267 , n5268 , n172738 , 
 n5270 , n5271 , n5272 , n172742 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
 n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
 n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
 n5300 , n172770 , n5302 , n5303 , n5304 , n5305 , n172775 , n5307 , n5308 , n5309 , 
 n172779 , n172780 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
 n5320 , n5321 , n5322 , n5323 , n172793 , n5325 , n5326 , n5327 , n172797 , n172798 , 
 n5330 , n5331 , n5332 , n172802 , n172803 , n5335 , n5336 , n5337 , n172807 , n172808 , 
 n5340 , n172810 , n172811 , n5343 , n172813 , n172814 , n172815 , n172816 , n172817 , n5349 , 
 n172819 , n172820 , n5352 , n5353 , n172823 , n5355 , n5356 , n172826 , n172827 , n172828 , 
 n5360 , n172830 , n172831 , n5363 , n172833 , n172834 , n5366 , n5367 , n172837 , n5369 , 
 n5370 , n172840 , n172841 , n172842 , n172843 , n5375 , n172845 , n172846 , n5378 , n172848 , 
 n5380 , n5381 , n172851 , n172852 , n5384 , n172854 , n172855 , n5387 , n172857 , n172858 , 
 n172859 , n172860 , n5392 , n172862 , n172863 , n5395 , n172865 , n5397 , n5398 , n172868 , 
 n172869 , n5401 , n172871 , n172872 , n5404 , n172874 , n172875 , n5407 , n5408 , n172878 , 
 n172879 , n5411 , n5412 , n5413 , n172883 , n172884 , n5416 , n172886 , n5418 , n172888 , 
 n5420 , n5421 , n172891 , n172892 , n5424 , n172894 , n172895 , n5427 , n172897 , n172898 , 
 n172899 , n5431 , n172901 , n5433 , n172903 , n172904 , n5436 , n5437 , n5438 , n5439 , 
 n172909 , n172910 , n5442 , n172912 , n5444 , n5445 , n172915 , n5447 , n172917 , n172918 , 
 n172919 , n172920 , n172921 , n5453 , n172923 , n172924 , n5456 , n172926 , n172927 , n5459 , 
 n172929 , n172930 , n5462 , n172932 , n172933 , n5465 , n172935 , n5467 , n5468 , n5469 , 
 n5470 , n172940 , n172941 , n172942 , n5474 , n172944 , n172945 , n5477 , n172947 , n5479 , 
 n5480 , n172950 , n172951 , n5483 , n172953 , n172954 , n5486 , n172956 , n172957 , n5489 , 
 n5490 , n172960 , n5492 , n172962 , n5494 , n5495 , n172965 , n172966 , n5498 , n172968 , 
 n172969 , n5501 , n172971 , n172972 , n5504 , n5505 , n5506 , n172976 , n172977 , n5509 , 
 n172979 , n172980 , n5512 , n172982 , n172983 , n5515 , n172985 , n5517 , n5518 , n172988 , 
 n172989 , n5521 , n172991 , n172992 , n5524 , n172994 , n5526 , n172996 , n5528 , n172998 , 
 n172999 , n5531 , n173001 , n5533 , n5534 , n5535 , n173005 , n173006 , n5538 , n173008 , 
 n5540 , n5541 , n173011 , n5543 , n5544 , n173014 , n173015 , n5547 , n173017 , n173018 , 
 n5550 , n173020 , n5552 , n5553 , n173023 , n173024 , n5556 , n173026 , n173027 , n5559 , 
 n173029 , n173030 , n5562 , n173032 , n173033 , n173034 , n173035 , n5567 , n173037 , n173038 , 
 n5570 , n173040 , n173041 , n5573 , n5574 , n5575 , n173045 , n173046 , n5578 , n5579 , 
 n5580 , n173050 , n173051 , n5583 , n5584 , n5585 , n173055 , n173056 , n5588 , n5589 , 
 n173059 , n173060 , n5592 , n5593 , n5594 , n173064 , n5596 , n5597 , n5598 , n5599 , 
 n5600 , n173070 , n173071 , n173072 , n5604 , n173074 , n173075 , n5607 , n173077 , n5609 , 
 n5610 , n173080 , n173081 , n5613 , n173083 , n173084 , n5616 , n173086 , n173087 , n5619 , 
 n173089 , n173090 , n5622 , n173092 , n173093 , n173094 , n173095 , n5627 , n173097 , n173098 , 
 n5630 , n173100 , n5632 , n5633 , n173103 , n173104 , n5636 , n173106 , n173107 , n5639 , 
 n173109 , n173110 , n5642 , n173112 , n5644 , n173114 , n5646 , n5647 , n173117 , n173118 , 
 n5650 , n173120 , n173121 , n5653 , n173123 , n173124 , n5656 , n173126 , n173127 , n5659 , 
 n173129 , n173130 , n5662 , n173132 , n173133 , n5665 , n173135 , n173136 , n5668 , n5669 , 
 n5670 , n173140 , n173141 , n5673 , n5674 , n5675 , n173145 , n5677 , n5678 , n5679 , 
 n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n173156 , n5688 , n5689 , 
 n5690 , n173160 , n173161 , n5693 , n5694 , n5695 , n173165 , n173166 , n5698 , n5699 , 
 n5700 , n173170 , n173171 , n5703 , n5704 , n5705 , n173175 , n173176 , n5708 , n5709 , 
 n5710 , n173180 , n5712 , n5713 , n5714 , n173184 , n173185 , n5717 , n173187 , n5719 , 
 n173189 , n5721 , n173191 , n173192 , n5724 , n173194 , n173195 , n5727 , n173197 , n173198 , 
 n5730 , n173200 , n173201 , n5733 , n173203 , n5735 , n5736 , n5737 , n5738 , n5739 , 
 n5740 , n5741 , n5742 , n173212 , n5744 , n5745 , n173215 , n173216 , n5748 , n5749 , 
 n173219 , n173220 , n5752 , n173222 , n173223 , n5755 , n173225 , n5757 , n173227 , n173228 , 
 n173229 , n173230 , n5762 , n173232 , n173233 , n173234 , n5766 , n173236 , n173237 , n5769 , 
 n173239 , n5771 , n173241 , n5773 , n5774 , n173244 , n173245 , n5777 , n173247 , n173248 , 
 n5780 , n173250 , n173251 , n5783 , n173253 , n5785 , n173255 , n5787 , n173257 , n5789 , 
 n5790 , n173260 , n173261 , n5793 , n173263 , n173264 , n5796 , n173266 , n5798 , n173268 , 
 n5800 , n173270 , n5802 , n5803 , n173273 , n173274 , n5806 , n173276 , n173277 , n5809 , 
 n173279 , n5811 , n5812 , n173282 , n5814 , n173284 , n5816 , n173286 , n173287 , n5819 , 
 n173289 , n5821 , n173291 , n5823 , n173293 , n173294 , n5826 , n5827 , n173297 , n5829 , 
 n173299 , n173300 , n173301 , n173302 , n5834 , n173304 , n173305 , n5837 , n173307 , n5839 , 
 n5840 , n5841 , n5842 , n5843 , n173313 , n173314 , n5846 , n173316 , n173317 , n5849 , 
 n173319 , n5851 , n5852 , n173322 , n173323 , n5855 , n173325 , n173326 , n5858 , n173328 , 
 n173329 , n173330 , n173331 , n5863 , n173333 , n173334 , n5866 , n173336 , n5868 , n5869 , 
 n173339 , n173340 , n5872 , n173342 , n173343 , n5875 , n173345 , n173346 , n5878 , n5879 , 
 n5880 , n5881 , n173351 , n173352 , n5884 , n173354 , n173355 , n5887 , n173357 , n5889 , 
 n5890 , n173360 , n5892 , n5893 , n5894 , n173364 , n5896 , n5897 , n5898 , n173368 , 
 n5900 , n5901 , n5902 , n173372 , n173373 , n5905 , n5906 , n173376 , n173377 , n5909 , 
 n5910 , n5911 , n173381 , n173382 , n173383 , n173384 , n5916 , n5917 , n173387 , n5919 , 
 n5920 , n173390 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n173398 , 
 n5930 , n173400 , n5932 , n5933 , n173403 , n5935 , n173405 , n5937 , n173407 , n173408 , 
 n5940 , n173410 , n5942 , n5943 , n173413 , n5945 , n173415 , n5947 , n5948 , n173418 , 
 n173419 , n5951 , n173421 , n173422 , n5954 , n173424 , n5956 , n173426 , n173427 , n5959 , 
 n173429 , n173430 , n5962 , n5963 , n5964 , n173434 , n5966 , n5967 , n173437 , n173438 , 
 n5970 , n173440 , n173441 , n5973 , n173443 , n5975 , n5976 , n5977 , n5978 , n5979 , 
 n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
 n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
 n173469 , n6001 , n173471 , n6003 , n6004 , n173474 , n6006 , n6007 , n6008 , n173478 , 
 n173479 , n6011 , n6012 , n6013 , n173483 , n173484 , n6016 , n6017 , n6018 , n173488 , 
 n173489 , n6021 , n6022 , n6023 , n173493 , n173494 , n6026 , n6027 , n6028 , n173498 , 
 n173499 , n6031 , n6032 , n6033 , n173503 , n173504 , n6036 , n173506 , n173507 , n173508 , 
 n6040 , n6041 , n173511 , n6043 , n6044 , n173514 , n6046 , n6047 , n173517 , n173518 , 
 n6050 , n173520 , n173521 , n6053 , n173523 , n173524 , n6056 , n173526 , n6058 , n6059 , 
 n173529 , n173530 , n6062 , n173532 , n173533 , n6065 , n173535 , n173536 , n6068 , n173538 , 
 n173539 , n6071 , n6072 , n6073 , n6074 , n6075 , n173545 , n173546 , n6078 , n173548 , 
 n6080 , n173550 , n173551 , n173552 , n6084 , n173554 , n173555 , n6087 , n173557 , n6089 , 
 n6090 , n173560 , n173561 , n6093 , n173563 , n173564 , n6096 , n173566 , n173567 , n6099 , 
 n173569 , n173570 , n6102 , n173572 , n173573 , n6105 , n173575 , n6107 , n6108 , n173578 , 
 n173579 , n6111 , n173581 , n173582 , n6114 , n173584 , n173585 , n6117 , n6118 , n6119 , 
 n173589 , n173590 , n6122 , n6123 , n6124 , n173594 , n173595 , n6127 , n6128 , n6129 , 
 n173599 , n173600 , n6132 , n6133 , n173603 , n173604 , n6136 , n6137 , n6138 , n173608 , 
 n173609 , n6141 , n6142 , n6143 , n173613 , n173614 , n6146 , n6147 , n6148 , n173618 , 
 n173619 , n6151 , n6152 , n6153 , n173623 , n173624 , n6156 , n6157 , n6158 , n173628 , 
 n173629 , n6161 , n6162 , n6163 , n173633 , n173634 , n6166 , n173636 , n173637 , n6169 , 
 n173639 , n6171 , n6172 , n6173 , n173643 , n6175 , n6176 , n6177 , n6178 , n173648 , 
 n6180 , n6181 , n6182 , n6183 , n173653 , n6185 , n173655 , n173656 , n173657 , n6189 , 
 n173659 , n173660 , n6192 , n173662 , n6194 , n6195 , n6196 , n6197 , n173667 , n173668 , 
 n173669 , n6201 , n6202 , n173672 , n173673 , n173674 , n6206 , n173676 , n173677 , n6209 , 
 n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
 n6220 , n173690 , n6222 , n173692 , n173693 , n6225 , n6226 , n173696 , n173697 , n6229 , 
 n173699 , n173700 , n6232 , n173702 , n6234 , n6235 , n173705 , n173706 , n6238 , n173708 , 
 n173709 , n6241 , n173711 , n173712 , n6244 , n173714 , n173715 , n173716 , n6248 , n173718 , 
 n6250 , n173720 , n173721 , n6253 , n173723 , n173724 , n6256 , n6257 , n173727 , n173728 , 
 n6260 , n173730 , n173731 , n6263 , n173733 , n173734 , n6266 , n173736 , n6268 , n6269 , 
 n173739 , n173740 , n6272 , n173742 , n173743 , n6275 , n173745 , n173746 , n173747 , n173748 , 
 n6280 , n173750 , n173751 , n6283 , n173753 , n6285 , n6286 , n6287 , n173757 , n173758 , 
 n6290 , n173760 , n173761 , n6293 , n173763 , n173764 , n6296 , n173766 , n6298 , n173768 , 
 n6300 , n6301 , n173771 , n6303 , n173773 , n173774 , n6306 , n173776 , n6308 , n173778 , 
 n173779 , n6311 , n6312 , n173782 , n173783 , n6315 , n6316 , n6317 , n173787 , n173788 , 
 n6320 , n6321 , n6322 , n173792 , n173793 , n6325 , n6326 , n6327 , n6328 , n6329 , 
 n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
 n173809 , n6341 , n173811 , n6343 , n6344 , n173814 , n173815 , n6347 , n173817 , n173818 , 
 n6350 , n173820 , n6352 , n173822 , n173823 , n6355 , n173825 , n173826 , n6358 , n173828 , 
 n6360 , n6361 , n173831 , n173832 , n6364 , n173834 , n173835 , n6367 , n173837 , n6369 , 
 n6370 , n6371 , n173841 , n173842 , n6374 , n173844 , n6376 , n173846 , n173847 , n173848 , 
 n6380 , n173850 , n6382 , n6383 , n173853 , n173854 , n6386 , n173856 , n6388 , n6389 , 
 n173859 , n173860 , n6392 , n173862 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
 n173869 , n6401 , n6402 , n6403 , n173873 , n173874 , n6406 , n6407 , n6408 , n6409 , 
 n173879 , n173880 , n6412 , n6413 , n6414 , n173884 , n6416 , n6417 , n173887 , n173888 , 
 n6420 , n6421 , n173891 , n173892 , n6424 , n6425 , n6426 , n173896 , n173897 , n173898 , 
 n173899 , n6431 , n173901 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n173908 , 
 n6440 , n6441 , n173911 , n6443 , n173913 , n6445 , n6446 , n173916 , n173917 , n6449 , 
 n173919 , n173920 , n6452 , n173922 , n173923 , n6455 , n6456 , n173926 , n173927 , n6459 , 
 n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n173935 , n6467 , n173937 , n173938 , 
 n6470 , n173940 , n173941 , n173942 , n173943 , n6475 , n173945 , n173946 , n6478 , n173948 , 
 n6480 , n6481 , n173951 , n173952 , n6484 , n173954 , n173955 , n6487 , n173957 , n6489 , 
 n173959 , n173960 , n6492 , n173962 , n173963 , n6495 , n173965 , n6497 , n6498 , n173968 , 
 n173969 , n6501 , n173971 , n173972 , n6504 , n173974 , n6506 , n6507 , n173977 , n173978 , 
 n6510 , n173980 , n173981 , n173982 , n6514 , n173984 , n173985 , n6517 , n173987 , n6519 , 
 n6520 , n173990 , n173991 , n6523 , n173993 , n173994 , n6526 , n173996 , n173997 , n6529 , 
 n173999 , n6531 , n6532 , n174002 , n6534 , n6535 , n6536 , n6537 , n6538 , n174008 , 
 n174009 , n6541 , n174011 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n174018 , 
 n174019 , n6551 , n174021 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
 n6560 , n174030 , n174031 , n6563 , n174033 , n6565 , n6566 , n6567 , n6568 , n174038 , 
 n6570 , n6571 , n6572 , n174042 , n174043 , n6575 , n6576 , n6577 , n174047 , n174048 , 
 n6580 , n6581 , n6582 , n174052 , n174053 , n6585 , n6586 , n6587 , n174057 , n174058 , 
 n6590 , n6591 , n6592 , n174062 , n174063 , n6595 , n6596 , n6597 , n174067 , n174068 , 
 n6600 , n6601 , n6602 , n174072 , n174073 , n6605 , n6606 , n6607 , n174077 , n174078 , 
 n6610 , n174080 , n174081 , n6613 , n6614 , n174084 , n174085 , n174086 , n6618 , n6619 , 
 n174089 , n174090 , n6622 , n6623 , n174093 , n174094 , n6626 , n174096 , n6628 , n174098 , 
 n6630 , n174100 , n6632 , n6633 , n174103 , n174104 , n6636 , n6637 , n174107 , n174108 , 
 n6640 , n6641 , n174111 , n174112 , n6644 , n6645 , n174115 , n174116 , n6648 , n6649 , 
 n174119 , n174120 , n6652 , n6653 , n6654 , n174124 , n174125 , n6657 , n6658 , n6659 , 
 n174129 , n174130 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n174137 , n6669 , 
 n6670 , n6671 , n174141 , n174142 , n6674 , n6675 , n6676 , n174146 , n174147 , n6679 , 
 n6680 , n6681 , n174151 , n174152 , n6684 , n6685 , n6686 , n174156 , n174157 , n6689 , 
 n6690 , n6691 , n174161 , n174162 , n6694 , n174164 , n174165 , n6697 , n174167 , n174168 , 
 n6700 , n174170 , n174171 , n6703 , n174173 , n174174 , n174175 , n6707 , n174177 , n174178 , 
 n6710 , n174180 , n6712 , n174182 , n6714 , n174184 , n6716 , n6717 , n174187 , n6719 , 
 n174189 , n174190 , n174191 , n6723 , n174193 , n6725 , n6726 , n6727 , n174197 , n6729 , 
 n6730 , n174200 , n174201 , n174202 , n6734 , n6735 , n174205 , n174206 , n6738 , n174208 , 
 n6740 , n6741 , n6742 , n174212 , n174213 , n6745 , n174215 , n6747 , n6748 , n174218 , 
 n174219 , n6751 , n174221 , n6753 , n174223 , n174224 , n6756 , n174226 , n174227 , n6759 , 
 n174229 , n6761 , n6762 , n174232 , n174233 , n6765 , n174235 , n174236 , n6768 , n174238 , 
 n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
 n6780 , n174250 , n174251 , n6783 , n174253 , n174254 , n6786 , n174256 , n6788 , n6789 , 
 n6790 , n174260 , n6792 , n174262 , n174263 , n6795 , n174265 , n174266 , n6798 , n174268 , 
 n174269 , n6801 , n174271 , n174272 , n174273 , n174274 , n174275 , n6807 , n174277 , n174278 , 
 n174279 , n174280 , n174281 , n6813 , n174283 , n174284 , n174285 , n174286 , n174287 , n6819 , 
 n174289 , n174290 , n174291 , n6823 , n174293 , n174294 , n174295 , n174296 , n174297 , n6829 , 
 n174299 , n174300 , n174301 , n174302 , n174303 , n6835 , n174305 , n174306 , n174307 , n174308 , 
 n174309 , n6841 , n174311 , n6843 , n174313 , n174314 , n174315 , n174316 , n174317 , n174318 , 
 n174319 , n174320 , n174321 , n6853 , n174323 , n6855 , n174325 , n6857 , n174327 , n6859 , 
 n174329 , n6861 , n174331 , n174332 , n174333 , n6865 , n174335 , n174336 , n174337 , n6869 , 
 n174339 , n174340 , n174341 , n6873 , n174343 , n174344 , n174345 , n174346 , n174347 , n6879 , 
 n174349 , n174350 , n174351 , n174352 , n174353 , n6885 , n174355 , n174356 , n174357 , n174358 , 
 n174359 , n6891 , n174361 , n174362 , n174363 , n174364 , n174365 , n6897 , n174367 , n174368 , 
 n174369 , n6901 , n174371 , n6903 , n174373 , n6905 , n174375 , n6907 , n174377 , n6909 , 
 n174379 , n6911 , n174381 , n174382 , n174383 , n174384 , n174385 , n174386 , n174387 , n6919 , 
 n174389 , n174390 , n174391 , n6923 , n174393 , n174394 , n174395 , n6927 , n174397 , n174398 , 
 n174399 , n174400 , n6932 , n174402 , n174403 , n6935 , n174405 , n6937 , n174407 , n174408 , 
 n174409 , n6941 , n174411 , n6943 , n6944 , n174414 , n6946 , n6947 , n174417 , n174418 , 
 n174419 , n6954 , n6955 , n6956 , n6957 , n6958 , n174425 , n6960 , n6961 , n6962 , 
 n174429 , n6964 , n6965 , n174432 , n174433 , n174434 , n6969 , n6970 , n6971 , n174438 , 
 n174439 , n6974 , n6975 , n6976 , n174443 , n174444 , n174445 , n6980 , n6981 , n174448 , 
 n174449 , n6984 , n174451 , n174452 , n6987 , n174454 , n174455 , n174456 , n6991 , n174458 , 
 n174459 , n6997 , n174461 , n174462 , n7000 , n174464 , n7002 , n174466 , n7004 , n7005 , 
 n174469 , n174470 , n174471 , n7009 , n174473 , n174474 , n7012 , n174476 , n174477 , n7015 , 
 n174479 , n174480 , n174481 , n174482 , n7020 , n174484 , n174485 , n7023 , n174487 , n7025 , 
 n7026 , n174490 , n174491 , n174492 , n174493 , n174494 , n7032 , n174496 , n174497 , n174498 , 
 n7036 , n174500 , n174501 , n174502 , n174503 , n174504 , n174505 , n7046 , n174507 , n174508 , 
 n174509 , n7050 , n174511 , n7052 , n7053 , n174514 , n7055 , n174516 , n7057 , n174518 , 
 n174519 , n7060 , n174521 , n174522 , n174523 , n7064 , n174525 , n7066 , n7067 , n174528 , 
 n174529 , n174530 , n7071 , n174532 , n7073 , n7074 , n7075 , n174536 , n174537 , n7078 , 
 n174539 , n7080 , n7081 , n174542 , n174543 , n7084 , n174545 , n7086 , n7087 , n7088 , 
 n174549 , n174550 , n7091 , n174552 , n7093 , n7094 , n7095 , n7096 , n174557 , n7098 , 
 n7099 , n7100 , n174561 , n7102 , n174563 , n174564 , n7105 , n7106 , n7107 , n174568 , 
 n7109 , n7110 , n174571 , n174572 , n7116 , n174574 , n174575 , n7119 , n174577 , n174578 , 
 n7122 , n174580 , n174581 , n7125 , n174583 , n174584 , n7128 , n174586 , n174587 , n7131 , 
 n174589 , n7133 , n174591 , n7135 , n7136 , n7137 , n174595 , n7139 , n174597 , n174598 , 
 n7142 , n174600 , n174601 , n7145 , n7146 , n174604 , n174605 , n7149 , n7150 , n174608 , 
 n174609 , n7153 , n7154 , n174612 , n174613 , n7157 , n174615 , n7159 , n7160 , n174618 , 
 n7162 , n174620 , n174621 , n174622 , n174623 , n7167 , n7168 , n174626 , n174627 , n7171 , 
 n174629 , n174630 , n7174 , n174632 , n7176 , n7177 , n174635 , n174636 , n7183 , n174638 , 
 n174639 , n7186 , n174641 , n7188 , n7189 , n7190 , n174645 , n7192 , n174647 , n7194 , 
 n174649 , n7196 , n7197 , n174652 , n7199 , n174654 , n174655 , n7202 , n174657 , n174658 , 
 n7205 , n7206 , n174661 , n174662 , n174663 , n7210 , n174665 , n174666 , n7213 , n7214 , 
 n174669 , n7216 , n7217 , n174672 , n7219 , n7220 , n174675 , n7222 , n174677 , n7224 , 
 n7225 , n174680 , n174681 , n7228 , n174683 , n174684 , n7231 , n174686 , n174687 , n7234 , 
 n174689 , n174690 , n174691 , n7238 , n7239 , n174694 , n174695 , n7242 , n7243 , n174698 , 
 n174699 , n174700 , n7247 , n174702 , n174703 , n7250 , n174705 , n174706 , n7253 , n174708 , 
 n174709 , n7256 , n174711 , n7258 , n7259 , n174714 , n174715 , n7262 , n174717 , n174718 , 
 n7265 , n174720 , n174721 , n7268 , n174723 , n174724 , n7271 , n174726 , n7276 , n7277 , 
 n174729 , n174730 , n7280 , n174732 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , 
 n7288 , n7289 , n7290 , n174742 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , 
 n7298 , n7299 , n7300 , n174752 , n7302 , n7303 , n7304 , n7305 , n174757 , n7307 , 
 n7308 , n7309 , n174761 , n174762 , n7312 , n7313 , n7314 , n174766 , n174767 , n174768 , 
 n174769 , n7319 , n7320 , n7321 , n174773 , n174774 , n174775 , n7325 , n7326 , n174778 , 
 n174779 , n174780 , n7330 , n174782 , n174783 , n7333 , n7334 , n7335 , n7336 , n7337 , 
 n174789 , n174790 , n7340 , n174792 , n174793 , n7343 , n174795 , n7345 , n174797 , n174798 , 
 n7348 , n7349 , n174801 , n174802 , n7352 , n174804 , n174805 , n7355 , n174807 , n7357 , 
 n174809 , n174810 , n174811 , n7364 , n174813 , n174814 , n174815 , n174816 , n174817 , n7370 , 
 n174819 , n174820 , n174821 , n7374 , n174823 , n7376 , n174825 , n174826 , n7379 , n174828 , 
 n174829 , n7382 , n174831 , n174832 , n7385 , n174834 , n174835 , n7388 , n174837 , n174838 , 
 n7391 , n174840 , n7393 , n7394 , n7395 , n174844 , n7397 , n7398 , n174847 , n7400 , 
 n174849 , n7402 , n7403 , n174852 , n174853 , n7406 , n174855 , n174856 , n7409 , n174858 , 
 n174859 , n7412 , n7413 , n174862 , n174863 , n7416 , n174865 , n174866 , n7419 , n174868 , 
 n174869 , n174870 , n174871 , n7424 , n7425 , n174874 , n174875 , n7428 , n174877 , n174878 , 
 n7431 , n174880 , n174881 , n7434 , n174883 , n174884 , n7437 , n174886 , n7439 , n174888 , 
 n7441 , n7442 , n174891 , n174892 , n7445 , n174894 , n174895 , n7448 , n174897 , n7450 , 
 n7451 , n174900 , n174901 , n7454 , n174903 , n174904 , n7457 , n174906 , n7459 , n174908 , 
 n7461 , n174910 , n7463 , n174912 , n174913 , n7466 , n7467 , n174916 , n174917 , n7470 , 
 n174919 , n174920 , n7476 , n174922 , n7478 , n174924 , n7480 , n174926 , n174927 , n7483 , 
 n7484 , n174930 , n174931 , n7487 , n174933 , n174934 , n7490 , n174936 , n7492 , n174938 , 
 n174939 , n7495 , n7496 , n174942 , n174943 , n7499 , n174945 , n174946 , n7502 , n174948 , 
 n174949 , n7505 , n174951 , n7507 , n174953 , n7509 , n174955 , n174956 , n174957 , n174958 , 
 n7514 , n174960 , n174961 , n7517 , n174963 , n7519 , n7520 , n7521 , n7522 , n7523 , 
 n7524 , n7525 , n7526 , n174972 , n7528 , n7529 , n174975 , n174976 , n7532 , n174978 , 
 n174979 , n7535 , n174981 , n174982 , n7538 , n7539 , n174985 , n174986 , n7542 , n174988 , 
 n174989 , n174990 , n7546 , n7547 , n174993 , n7549 , n174995 , n7551 , n7552 , n7553 , 
 n174999 , n7555 , n175001 , n7557 , n7558 , n7559 , n175005 , n7561 , n7562 , n175008 , 
 n175009 , n7565 , n175011 , n175012 , n7568 , n175014 , n7570 , n7571 , n7572 , n7573 , 
 n7574 , n7575 , n7576 , n7577 , n175023 , n7582 , n7583 , n7584 , n175027 , n7586 , 
 n175029 , n7588 , n175031 , n175032 , n7591 , n175034 , n7593 , n7594 , n175037 , n175038 , 
 n175039 , n7598 , n7599 , n175042 , n7601 , n7602 , n175045 , n175046 , n175047 , n7606 , 
 n175049 , n7608 , n7609 , n175052 , n175053 , n7612 , n175055 , n7614 , n175057 , n175058 , 
 n175059 , n175060 , n7619 , n175062 , n175063 , n175064 , n7623 , n175066 , n175067 , n175068 , 
 n175069 , n7628 , n175071 , n175072 , n7631 , n175074 , n7633 , n7634 , n175077 , n175078 , 
 n7637 , n175080 , n175081 , n7640 , n175083 , n175084 , n7643 , n175086 , n175087 , n175088 , 
 n175089 , n175090 , n175091 , n7650 , n175093 , n175094 , n7653 , n175096 , n175097 , n7656 , 
 n175099 , n175100 , n7659 , n175102 , n7661 , n7662 , n7663 , n7664 , n7665 , n175108 , 
 n175109 , n7668 , n175111 , n175112 , n7671 , n7672 , n7673 , n7674 , n7675 , n175118 , 
 n175119 , n7678 , n175121 , n175122 , n7681 , n175124 , n7683 , n7684 , n175127 , n175128 , 
 n7687 , n175130 , n175131 , n7690 , n175133 , n7692 , n7693 , n7694 , n175137 , n175138 , 
 n7697 , n175140 , n175141 , n7700 , n175143 , n7702 , n7703 , n175146 , n175147 , n7706 , 
 n175149 , n175150 , n7709 , n175152 , n175153 , n175154 , n7716 , n7717 , n7718 , n175158 , 
 n175159 , n175160 , n175161 , n7723 , n175163 , n7725 , n175165 , n175166 , n7728 , n175168 , 
 n175169 , n7731 , n175171 , n7733 , n7734 , n175174 , n175175 , n7737 , n175177 , n175178 , 
 n7740 , n175180 , n175181 , n7743 , n175183 , n175184 , n175185 , n175186 , n7748 , n175188 , 
 n175189 , n7751 , n175191 , n7753 , n7754 , n7755 , n175195 , n7757 , n7758 , n7759 , 
 n175199 , n7761 , n7762 , n7763 , n7764 , n175204 , n7766 , n7767 , n175207 , n7769 , 
 n175209 , n7771 , n175211 , n175212 , n7774 , n7775 , n7776 , n175216 , n7778 , n7779 , 
 n7780 , n7781 , n175221 , n175222 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
 n175229 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n175236 , n7798 , n7799 , 
 n7800 , n175240 , n7802 , n7803 , n7804 , n175244 , n175245 , n7807 , n175247 , n175248 , 
 n7810 , n175250 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n175258 , 
 n7820 , n175260 , n7822 , n175262 , n7824 , n7825 , n7826 , n175266 , n7828 , n7829 , 
 n7830 , n7831 , n175271 , n175272 , n7834 , n175274 , n7836 , n7837 , n175277 , n175278 , 
 n7843 , n7844 , n175281 , n175282 , n175283 , n175284 , n7849 , n7850 , n175287 , n7852 , 
 n7853 , n175290 , n175291 , n175292 , n175293 , n7858 , n175295 , n175296 , n7861 , n175298 , 
 n7863 , n7864 , n175301 , n175302 , n7867 , n175304 , n175305 , n7870 , n175307 , n175308 , 
 n7873 , n175310 , n175311 , n7876 , n175313 , n175314 , n7879 , n175316 , n175317 , n175318 , 
 n175319 , n7884 , n175321 , n175322 , n7887 , n175324 , n7889 , n175326 , n175327 , n175328 , 
 n7893 , n175330 , n175331 , n7896 , n175333 , n175334 , n7899 , n175336 , n175337 , n7902 , 
 n175339 , n175340 , n7905 , n175342 , n7907 , n7908 , n175345 , n175346 , n7911 , n175348 , 
 n175349 , n7914 , n175351 , n175352 , n175353 , n7918 , n7919 , n175356 , n175357 , n175358 , 
 n7923 , n7924 , n175361 , n175362 , n7927 , n7928 , n175365 , n7930 , n175367 , n175368 , 
 n7933 , n175370 , n7935 , n7936 , n7937 , n175374 , n175375 , n7940 , n175377 , n7942 , 
 n7943 , n175380 , n175381 , n7946 , n175383 , n7948 , n7949 , n7950 , n175387 , n175388 , 
 n7953 , n175390 , n7955 , n7956 , n7957 , n7958 , n7959 , n175396 , n7961 , n175398 , 
 n7963 , n175400 , n175401 , n7966 , n7967 , n175404 , n175405 , n7970 , n175407 , n175408 , 
 n7973 , n175410 , n7975 , n7976 , n175413 , n7978 , n7979 , n175416 , n7981 , n175418 , 
 n7983 , n7984 , n7985 , n175422 , n7987 , n7988 , n175425 , n175426 , n7991 , n175428 , 
 n175429 , n175430 , n7998 , n7999 , n8000 , n175434 , n175435 , n8003 , n8004 , n175438 , 
 n175439 , n175440 , n8008 , n175442 , n8010 , n175444 , n8012 , n8013 , n175447 , n175448 , 
 n8016 , n175450 , n175451 , n8019 , n175453 , n175454 , n175455 , n8023 , n8024 , n175458 , 
 n8026 , n175460 , n175461 , n8029 , n8030 , n175464 , n175465 , n8033 , n8034 , n8035 , 
 n175469 , n175470 , n8038 , n8039 , n8040 , n175474 , n8042 , n175476 , n175477 , n175478 , 
 n8046 , n8047 , n175481 , n175482 , n175483 , n175484 , n8052 , n175486 , n175487 , n8055 , 
 n175489 , n8057 , n8058 , n175492 , n175493 , n8061 , n175495 , n175496 , n8064 , n175498 , 
 n175499 , n175500 , n175501 , n8069 , n175503 , n8071 , n175505 , n175506 , n175507 , n175508 , 
 n175509 , n175510 , n175511 , n175512 , n8080 , n175514 , n175515 , n8083 , n175517 , n175518 , 
 n8086 , n175520 , n175521 , n8089 , n175523 , n8091 , n175525 , n8093 , n8094 , n175528 , 
 n175529 , n8097 , n175531 , n175532 , n8100 , n175534 , n175535 , n8103 , n175537 , n175538 , 
 n175539 , n175540 , n175541 , n175542 , n175543 , n8111 , n175545 , n8113 , n8114 , n175548 , 
 n175549 , n8117 , n175551 , n175552 , n8120 , n175554 , n175555 , n8123 , n175557 , n175558 , 
 n8126 , n175560 , n175561 , n8129 , n175563 , n175564 , n8132 , n175566 , n175567 , n8135 , 
 n8136 , n175570 , n175571 , n8142 , n8143 , n8144 , n175575 , n8146 , n175577 , n8148 , 
 n175579 , n8150 , n8151 , n175582 , n175583 , n8154 , n175585 , n175586 , n8157 , n175588 , 
 n175589 , n8160 , n175591 , n175592 , n8163 , n175594 , n8165 , n8166 , n175597 , n175598 , 
 n8169 , n175600 , n175601 , n8172 , n175603 , n175604 , n8175 , n8176 , n175607 , n175608 , 
 n8179 , n175610 , n175611 , n8182 , n175613 , n175614 , n8185 , n175616 , n8187 , n8188 , 
 n175619 , n175620 , n8191 , n175622 , n175623 , n8194 , n175625 , n175626 , n8197 , n175628 , 
 n175629 , n8200 , n175631 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
 n8209 , n175640 , n8211 , n175642 , n8213 , n8214 , n175645 , n175646 , n8217 , n175648 , 
 n175649 , n8220 , n175651 , n8222 , n175653 , n175654 , n8225 , n175656 , n175657 , n8228 , 
 n175659 , n8230 , n8231 , n175662 , n8233 , n175664 , n175665 , n175666 , n8237 , n175668 , 
 n175669 , n175670 , n175671 , n8242 , n8243 , n8244 , n175675 , n175676 , n8247 , n175678 , 
 n175679 , n8250 , n175681 , n8252 , n8253 , n175684 , n175685 , n8256 , n175687 , n175688 , 
 n8259 , n175690 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n175697 , n8268 , 
 n8269 , n8270 , n175701 , n175702 , n8273 , n8274 , n8275 , n175706 , n175707 , n8278 , 
 n8279 , n8280 , n175711 , n175712 , n8283 , n8284 , n8285 , n175716 , n175717 , n8288 , 
 n8289 , n8290 , n175721 , n175722 , n8293 , n175724 , n8295 , n8296 , n8297 , n8298 , 
 n175729 , n175730 , n8301 , n8302 , n175733 , n175734 , n8305 , n175736 , n8307 , n8308 , 
 n175739 , n8310 , n8311 , n175742 , n8316 , n8317 , n8318 , n8319 , n8320 , n175748 , 
 n8322 , n175750 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n175757 , n175758 , 
 n8332 , n175760 , n175761 , n8335 , n175763 , n8337 , n175765 , n175766 , n175767 , n8341 , 
 n175769 , n175770 , n8344 , n175772 , n175773 , n175774 , n175775 , n8349 , n175777 , n175778 , 
 n8352 , n175780 , n8354 , n8355 , n175783 , n8357 , n175785 , n8359 , n175787 , n175788 , 
 n8362 , n175790 , n175791 , n8365 , n175793 , n175794 , n8368 , n175796 , n8370 , n175798 , 
 n175799 , n175800 , n175801 , n8375 , n175803 , n175804 , n175805 , n8379 , n175807 , n175808 , 
 n8382 , n175810 , n175811 , n8385 , n175813 , n175814 , n8388 , n175816 , n175817 , n8391 , 
 n175819 , n8393 , n8394 , n175822 , n175823 , n175824 , n175825 , n175826 , n175827 , n8401 , 
 n175829 , n175830 , n8404 , n175832 , n175833 , n175834 , n175835 , n8409 , n175837 , n175838 , 
 n8412 , n175840 , n8414 , n8415 , n175843 , n175844 , n175845 , n175846 , n175847 , n175848 , 
 n8422 , n175850 , n175851 , n8425 , n175853 , n175854 , n8428 , n175856 , n175857 , n8431 , 
 n175859 , n175860 , n8434 , n175862 , n8436 , n8437 , n175865 , n175866 , n175867 , n8441 , 
 n175869 , n175870 , n8444 , n175872 , n175873 , n8447 , n175875 , n175876 , n8450 , n8451 , 
 n8452 , n175880 , n175881 , n8455 , n8456 , n8457 , n175885 , n8459 , n8460 , n8461 , 
 n175889 , n8463 , n8464 , n8465 , n175893 , n175894 , n8468 , n175896 , n8470 , n175898 , 
 n175899 , n175900 , n8474 , n8475 , n175903 , n8477 , n175905 , n175906 , n175907 , n8484 , 
 n175909 , n175910 , n175911 , n8488 , n175913 , n8490 , n8491 , n175916 , n175917 , n175918 , 
 n175919 , n8496 , n175921 , n175922 , n175923 , n8500 , n175925 , n8502 , n8503 , n175928 , 
 n175929 , n8506 , n175931 , n175932 , n8509 , n175934 , n175935 , n8512 , n175937 , n8514 , 
 n175939 , n8516 , n8517 , n175942 , n175943 , n8520 , n175945 , n175946 , n8523 , n175948 , 
 n175949 , n8526 , n8527 , n8528 , n175953 , n175954 , n8531 , n175956 , n8533 , n175958 , 
 n8535 , n8536 , n175961 , n175962 , n8539 , n175964 , n175965 , n8542 , n175967 , n175968 , 
 n175969 , n175970 , n175971 , n175972 , n175973 , n8550 , n175975 , n8552 , n8553 , n175978 , 
 n175979 , n8556 , n175981 , n175982 , n8559 , n175984 , n175985 , n8562 , n175987 , n8564 , 
 n175989 , n8566 , n8567 , n175992 , n175993 , n8570 , n175995 , n175996 , n8573 , n175998 , 
 n175999 , n8576 , n176001 , n8578 , n176003 , n176004 , n8581 , n176006 , n8583 , n176008 , 
 n176009 , n8586 , n176011 , n176012 , n8589 , n8590 , n8591 , n176016 , n176017 , n8594 , 
 n8595 , n8596 , n176021 , n176022 , n8599 , n8600 , n176025 , n176026 , n8603 , n8604 , 
 n8605 , n8606 , n8607 , n176032 , n176033 , n8610 , n176035 , n176036 , n8613 , n8614 , 
 n8615 , n176040 , n176041 , n176042 , n8619 , n8620 , n8621 , n8622 , n176047 , n176048 , 
 n8625 , n8626 , n8627 , n176052 , n176053 , n8630 , n176055 , n176056 , n8633 , n176058 , 
 n176059 , n8636 , n8637 , n8638 , n176063 , n176064 , n8641 , n176066 , n8643 , n8644 , 
 n176069 , n176070 , n8647 , n176072 , n176073 , n8650 , n8651 , n8652 , n176077 , n8654 , 
 n176079 , n176080 , n8657 , n176082 , n8659 , n8660 , n176085 , n8662 , n176087 , n176088 , 
 n176089 , n8666 , n176091 , n176092 , n176093 , n8670 , n176095 , n176096 , n8676 , n176098 , 
 n176099 , n8679 , n176101 , n176102 , n8682 , n176104 , n176105 , n8685 , n176107 , n8687 , 
 n8688 , n176110 , n8690 , n8691 , n176113 , n176114 , n8694 , n176116 , n8696 , n176118 , 
 n8698 , n176120 , n176121 , n8701 , n176123 , n176124 , n8704 , n8705 , n176127 , n8707 , 
 n176129 , n8709 , n176131 , n8711 , n8712 , n8713 , n8714 , n176136 , n8716 , n176138 , 
 n176139 , n8719 , n8720 , n176142 , n8722 , n176144 , n176145 , n176146 , n176147 , n8727 , 
 n176149 , n176150 , n8730 , n176152 , n176153 , n8733 , n176155 , n176156 , n8736 , n176158 , 
 n176159 , n8739 , n176161 , n176162 , n8742 , n176164 , n8744 , n8745 , n176167 , n176168 , 
 n176169 , n8749 , n176171 , n8751 , n176173 , n8753 , n176175 , n8755 , n8756 , n176178 , 
 n8758 , n176180 , n176181 , n176182 , n176183 , n8763 , n176185 , n176186 , n8766 , n176188 , 
 n8768 , n176190 , n176191 , n8771 , n176193 , n8773 , n176195 , n176196 , n8776 , n176198 , 
 n176199 , n8779 , n176201 , n176202 , n8782 , n176204 , n8784 , n8785 , n176207 , n176208 , 
 n176209 , n8789 , n176211 , n176212 , n176213 , n176214 , n8794 , n8795 , n176217 , n176218 , 
 n8798 , n8799 , n176221 , n176222 , n8802 , n8803 , n176225 , n176226 , n8806 , n176228 , 
 n176229 , n8809 , n176231 , n176232 , n8812 , n176234 , n8814 , n8815 , n176237 , n176238 , 
 n8818 , n176240 , n176241 , n8821 , n176243 , n176244 , n8824 , n176246 , n8826 , n176248 , 
 n8828 , n8829 , n176251 , n176252 , n8832 , n176254 , n176255 , n8835 , n176257 , n176258 , 
 n8838 , n176260 , n8840 , n176262 , n8842 , n8843 , n176265 , n176266 , n8846 , n8847 , 
 n176269 , n176270 , n8850 , n8851 , n8852 , n176274 , n176275 , n8855 , n8856 , n8857 , 
 n176279 , n176280 , n8863 , n8864 , n8865 , n176284 , n176285 , n8868 , n8869 , n176288 , 
 n176289 , n8872 , n8873 , n8874 , n176293 , n176294 , n8877 , n8878 , n8879 , n176298 , 
 n176299 , n8882 , n176301 , n176302 , n8885 , n8886 , n176305 , n176306 , n176307 , n8890 , 
 n8891 , n176310 , n176311 , n176312 , n176313 , n8896 , n176315 , n176316 , n176317 , n176318 , 
 n8901 , n176320 , n176321 , n8904 , n176323 , n8906 , n8907 , n176326 , n176327 , n8910 , 
 n176329 , n176330 , n8913 , n176332 , n176333 , n8916 , n176335 , n176336 , n8919 , n176338 , 
 n176339 , n8922 , n176341 , n8924 , n8925 , n176344 , n176345 , n8928 , n176347 , n176348 , 
 n8931 , n176350 , n176351 , n8934 , n8935 , n8936 , n176355 , n176356 , n176357 , n176358 , 
 n8941 , n176360 , n176361 , n8944 , n176363 , n8946 , n8947 , n176366 , n176367 , n8950 , 
 n176369 , n176370 , n8953 , n176372 , n176373 , n176374 , n176375 , n8958 , n176377 , n176378 , 
 n8961 , n176380 , n8963 , n8964 , n176383 , n176384 , n176385 , n176386 , n176387 , n8970 , 
 n176389 , n176390 , n8973 , n176392 , n8975 , n176394 , n8977 , n8978 , n176397 , n176398 , 
 n176399 , n8982 , n176401 , n176402 , n8985 , n176404 , n176405 , n176406 , n8989 , n176408 , 
 n176409 , n8992 , n8993 , n8994 , n176413 , n176414 , n8997 , n8998 , n8999 , n176418 , 
 n176419 , n9002 , n9003 , n9004 , n176423 , n176424 , n9007 , n9008 , n9009 , n176428 , 
 n176429 , n9012 , n9013 , n9014 , n176433 , n176434 , n176435 , n9018 , n9019 , n176438 , 
 n176439 , n9022 , n9023 , n9024 , n176443 , n176444 , n9027 , n176446 , n176447 , n9030 , 
 n176449 , n176450 , n9033 , n9034 , n176453 , n9036 , n176455 , n9038 , n9039 , n176458 , 
 n176459 , n176460 , n176461 , n9044 , n176463 , n176464 , n9047 , n176466 , n9049 , n9050 , 
 n176469 , n176470 , n9053 , n176472 , n176473 , n9056 , n176475 , n176476 , n9059 , n176478 , 
 n176479 , n9062 , n176481 , n9064 , n176483 , n176484 , n176485 , n176486 , n9069 , n176488 , 
 n176489 , n176490 , n9076 , n176492 , n176493 , n9079 , n176495 , n176496 , n9082 , n9083 , 
 n176499 , n176500 , n9086 , n176502 , n176503 , n9089 , n176505 , n176506 , n9092 , n176508 , 
 n9094 , n9095 , n176511 , n176512 , n9098 , n176514 , n176515 , n9101 , n176517 , n9103 , 
 n176519 , n9105 , n176521 , n9107 , n9108 , n176524 , n176525 , n9111 , n176527 , n176528 , 
 n9114 , n176530 , n9116 , n9117 , n9118 , n9119 , n9120 , n176536 , n176537 , n9123 , 
 n176539 , n9125 , n9126 , n9127 , n9128 , n176544 , n9130 , n9131 , n9132 , n176548 , 
 n176549 , n9135 , n9136 , n9137 , n176553 , n176554 , n9140 , n9141 , n9142 , n176558 , 
 n176559 , n9145 , n9146 , n9147 , n176563 , n176564 , n9150 , n9151 , n9152 , n176568 , 
 n9154 , n9155 , n9156 , n9157 , n176573 , n176574 , n176575 , n9161 , n9162 , n176578 , 
 n176579 , n176580 , n176581 , n9167 , n176583 , n176584 , n9170 , n176586 , n9172 , n9173 , 
 n176589 , n176590 , n9176 , n176592 , n176593 , n9179 , n176595 , n176596 , n176597 , n176598 , 
 n9184 , n176600 , n176601 , n176602 , n176603 , n9189 , n176605 , n176606 , n9192 , n176608 , 
 n9194 , n9195 , n176611 , n176612 , n9198 , n176614 , n176615 , n9201 , n176617 , n176618 , 
 n9204 , n9205 , n176621 , n9207 , n176623 , n9209 , n9210 , n176626 , n176627 , n9213 , 
 n176629 , n176630 , n9216 , n176632 , n176633 , n9219 , n9220 , n9221 , n176637 , n176638 , 
 n9224 , n176640 , n9226 , n176642 , n9228 , n9229 , n176645 , n176646 , n9232 , n9233 , 
 n176649 , n176650 , n9236 , n9237 , n9238 , n176654 , n176655 , n9241 , n9242 , n9243 , 
 n176659 , n176660 , n9246 , n9247 , n9248 , n176664 , n176665 , n9251 , n9252 , n9253 , 
 n176669 , n176670 , n9256 , n9257 , n9258 , n176674 , n176675 , n9261 , n176677 , n9263 , 
 n176679 , n9265 , n176681 , n176682 , n9268 , n9269 , n9270 , n176686 , n176687 , n9273 , 
 n176689 , n176690 , n176691 , n176692 , n176693 , n176694 , n176695 , n9284 , n176697 , n9286 , 
 n176699 , n176700 , n176701 , n9290 , n176703 , n176704 , n9293 , n176706 , n176707 , n176708 , 
 n176709 , n9298 , n176711 , n9300 , n176713 , n176714 , n176715 , n176716 , n9305 , n176718 , 
 n176719 , n176720 , n9309 , n176722 , n176723 , n9312 , n176725 , n176726 , n9315 , n176728 , 
 n176729 , n9318 , n176731 , n176732 , n9321 , n176734 , n176735 , n9324 , n176737 , n9326 , 
 n9327 , n176740 , n176741 , n9330 , n176743 , n176744 , n9333 , n176746 , n176747 , n9336 , 
 n176749 , n176750 , n9339 , n9340 , n176753 , n176754 , n9343 , n176756 , n176757 , n9346 , 
 n176759 , n9348 , n9349 , n176762 , n9351 , n176764 , n176765 , n9354 , n176767 , n176768 , 
 n176769 , n9358 , n176771 , n176772 , n9361 , n176774 , n176775 , n9364 , n176777 , n176778 , 
 n176779 , n9368 , n176781 , n9370 , n176783 , n176784 , n9373 , n176786 , n176787 , n9376 , 
 n9377 , n176790 , n9379 , n9380 , n9381 , n176794 , n176795 , n9384 , n9385 , n9386 , 
 n176799 , n176800 , n9389 , n176802 , n176803 , n9392 , n9393 , n9394 , n176807 , n9396 , 
 n176809 , n9398 , n9399 , n176812 , n176813 , n176814 , n176815 , n9404 , n176817 , n176818 , 
 n9407 , n176820 , n176821 , n9410 , n176823 , n176824 , n9413 , n176826 , n176827 , n9416 , 
 n176829 , n9418 , n9419 , n9420 , n9421 , n176834 , n176835 , n9424 , n9425 , n176838 , 
 n9427 , n176840 , n176841 , n9430 , n9431 , n176844 , n176845 , n9434 , n176847 , n176848 , 
 n176849 , n9438 , n9439 , n176852 , n176853 , n176854 , n176855 , n9444 , n176857 , n176858 , 
 n9447 , n176860 , n9449 , n9450 , n176863 , n176864 , n9453 , n176866 , n176867 , n9456 , 
 n176869 , n176870 , n9459 , n176872 , n9461 , n176874 , n9463 , n9464 , n176877 , n176878 , 
 n9467 , n176880 , n176881 , n9470 , n176883 , n176884 , n9473 , n176886 , n176887 , n9476 , 
 n176889 , n176890 , n9479 , n176892 , n9481 , n9482 , n176895 , n176896 , n9485 , n176898 , 
 n176899 , n9488 , n176901 , n176902 , n9491 , n176904 , n176905 , n176906 , n176907 , n9496 , 
 n176909 , n176910 , n9499 , n176912 , n176913 , n9502 , n9503 , n176916 , n176917 , n9506 , 
 n176919 , n176920 , n9509 , n9510 , n9511 , n176924 , n176925 , n9517 , n9518 , n9519 , 
 n176929 , n176930 , n9522 , n9523 , n9524 , n176934 , n176935 , n9527 , n176937 , n176938 , 
 n9530 , n176940 , n176941 , n176942 , n176943 , n9535 , n9536 , n176946 , n9538 , n9539 , 
 n176949 , n176950 , n9542 , n176952 , n176953 , n176954 , n9546 , n176956 , n176957 , n9549 , 
 n176959 , n176960 , n9552 , n176962 , n176963 , n9555 , n176965 , n176966 , n176967 , n176968 , 
 n9560 , n9561 , n176971 , n176972 , n9564 , n176974 , n176975 , n9567 , n176977 , n176978 , 
 n9570 , n9571 , n176981 , n9573 , n176983 , n9575 , n176985 , n176986 , n9578 , n9579 , 
 n176989 , n176990 , n9582 , n176992 , n176993 , n9585 , n176995 , n9587 , n9588 , n176998 , 
 n176999 , n9591 , n177001 , n177002 , n9594 , n177004 , n177005 , n9597 , n177007 , n177008 , 
 n9600 , n177010 , n9602 , n9603 , n9604 , n177014 , n9606 , n9607 , n9608 , n177018 , 
 n9610 , n177020 , n177021 , n9613 , n9614 , n177024 , n177025 , n9617 , n177027 , n177028 , 
 n9620 , n177030 , n177031 , n9623 , n9624 , n9625 , n177035 , n177036 , n9628 , n9629 , 
 n9630 , n177040 , n177041 , n9633 , n9634 , n177044 , n177045 , n9637 , n177047 , n177048 , 
 n9640 , n9641 , n177051 , n177052 , n177053 , n177054 , n9646 , n177056 , n9648 , n177058 , 
 n177059 , n177060 , n177061 , n9653 , n177063 , n177064 , n177065 , n9657 , n177067 , n177068 , 
 n177069 , n177070 , n9662 , n177072 , n177073 , n9665 , n177075 , n9667 , n9668 , n177078 , 
 n177079 , n9671 , n177081 , n177082 , n9674 , n177084 , n177085 , n9677 , n177087 , n177088 , 
 n177089 , n9681 , n177091 , n177092 , n9684 , n177094 , n9686 , n9687 , n177097 , n177098 , 
 n9690 , n177100 , n177101 , n9693 , n177103 , n9695 , n9696 , n9697 , n9698 , n9699 , 
 n9700 , n177110 , n9702 , n177112 , n177113 , n9705 , n9706 , n9707 , n177117 , n9709 , 
 n177119 , n177120 , n9712 , n177122 , n9714 , n9715 , n177125 , n177126 , n9718 , n177128 , 
 n177129 , n9721 , n177131 , n9723 , n177133 , n9725 , n177135 , n177136 , n9728 , n9729 , 
 n177139 , n177140 , n9732 , n177142 , n9734 , n177144 , n177145 , n9737 , n177147 , n177148 , 
 n9743 , n177150 , n177151 , n9746 , n177153 , n9748 , n177155 , n9750 , n177157 , n9752 , 
 n177159 , n177160 , n9755 , n9756 , n9757 , n9758 , n177165 , n9760 , n177167 , n177168 , 
 n177169 , n9764 , n9765 , n177172 , n9767 , n177174 , n177175 , n9770 , n9771 , n177178 , 
 n177179 , n177180 , n177181 , n177182 , n9777 , n177184 , n177185 , n9780 , n177187 , n9782 , 
 n9783 , n177190 , n177191 , n9786 , n177193 , n177194 , n9789 , n177196 , n177197 , n9792 , 
 n177199 , n177200 , n9795 , n177202 , n177203 , n9798 , n177205 , n177206 , n9801 , n177208 , 
 n9803 , n9804 , n177211 , n177212 , n9807 , n177214 , n177215 , n9810 , n177217 , n177218 , 
 n9813 , n9814 , n9815 , n177222 , n177223 , n9818 , n9819 , n9820 , n177227 , n9822 , 
 n9823 , n9824 , n177231 , n177232 , n9827 , n177234 , n177235 , n9830 , n9831 , n177238 , 
 n177239 , n177240 , n177241 , n177242 , n9837 , n177244 , n177245 , n9840 , n177247 , n9842 , 
 n9843 , n177250 , n177251 , n9846 , n177253 , n177254 , n9849 , n177256 , n9851 , n177258 , 
 n177259 , n9854 , n177261 , n177262 , n9857 , n177264 , n9859 , n9860 , n177267 , n9862 , 
 n177269 , n9864 , n177271 , n177272 , n177273 , n9868 , n177275 , n177276 , n9871 , n177278 , 
 n177279 , n9874 , n177281 , n9876 , n9877 , n177284 , n177285 , n9880 , n177287 , n177288 , 
 n9883 , n177290 , n177291 , n9886 , n177293 , n9888 , n177295 , n9890 , n9891 , n9892 , 
 n177299 , n177300 , n9895 , n9896 , n9897 , n177304 , n177305 , n9900 , n177307 , n177308 , 
 n9903 , n177310 , n177311 , n9906 , n177313 , n177314 , n9909 , n177316 , n177317 , n9912 , 
 n177319 , n177320 , n177321 , n177322 , n177323 , n9918 , n177325 , n177326 , n9921 , n177328 , 
 n177329 , n9924 , n9925 , n177332 , n177333 , n9928 , n177335 , n177336 , n9931 , n177338 , 
 n177339 , n177340 , n177341 , n9936 , n177343 , n9938 , n177345 , n177346 , n177347 , n177348 , 
 n9943 , n177350 , n177351 , n177352 , n9947 , n177354 , n177355 , n9950 , n177357 , n177358 , 
 n9953 , n177360 , n177361 , n9956 , n9957 , n9958 , n177365 , n9960 , n9961 , n9962 , 
 n177369 , n177370 , n9965 , n9966 , n177373 , n177374 , n9969 , n177376 , n177377 , n9972 , 
 n9973 , n177380 , n177381 , n177382 , n177383 , n177384 , n9979 , n177386 , n177387 , n9982 , 
 n177389 , n9984 , n9985 , n177392 , n177393 , n9988 , n177395 , n177396 , n9991 , n177398 , 
 n177399 , n9997 , n177401 , n9999 , n177403 , n177404 , n10002 , n10003 , n177407 , n177408 , 
 n10006 , n177410 , n177411 , n10009 , n10010 , n177414 , n177415 , n10013 , n177417 , n177418 , 
 n10016 , n177420 , n10018 , n177422 , n177423 , n10021 , n177425 , n177426 , n10024 , n10025 , 
 n10026 , n177430 , n177431 , n10029 , n177433 , n177434 , n10032 , n177436 , n10034 , n177438 , 
 n177439 , n177440 , n10038 , n177442 , n177443 , n10041 , n177445 , n177446 , n177447 , n177448 , 
 n10046 , n177450 , n177451 , n10049 , n177453 , n177454 , n10052 , n177456 , n177457 , n177458 , 
 n177459 , n177460 , n10058 , n177462 , n177463 , n177464 , n177465 , n10063 , n177467 , n177468 , 
 n10066 , n177470 , n177471 , n177472 , n177473 , n10071 , n177475 , n10073 , n10074 , n177478 , 
 n177479 , n10077 , n177481 , n177482 , n10080 , n177484 , n177485 , n10083 , n177487 , n177488 , 
 n10086 , n177490 , n177491 , n177492 , n177493 , n177494 , n10092 , n177496 , n177497 , n10095 , 
 n177499 , n177500 , n177501 , n10099 , n177503 , n10101 , n177505 , n177506 , n10104 , n177508 , 
 n10106 , n10107 , n10108 , n177512 , n10110 , n177514 , n177515 , n10113 , n177517 , n177518 , 
 n10116 , n177520 , n177521 , n10119 , n177523 , n10121 , n177525 , n10123 , n177527 , n177528 , 
 n10126 , n10127 , n10128 , n10129 , n177533 , n177534 , n10132 , n177536 , n177537 , n10135 , 
 n177539 , n10137 , n10138 , n177542 , n10140 , n177544 , n177545 , n177546 , n10144 , n177548 , 
 n10146 , n177550 , n10148 , n177552 , n177553 , n177554 , n10152 , n177556 , n177557 , n10155 , 
 n177559 , n177560 , n10158 , n177562 , n177563 , n10161 , n177565 , n10163 , n177567 , n177568 , 
 n177569 , n10167 , n177571 , n177572 , n10170 , n177574 , n177575 , n10173 , n177577 , n177578 , 
 n10176 , n177580 , n177581 , n10179 , n10180 , n10181 , n10182 , n177586 , n177587 , n10185 , 
 n177589 , n10187 , n177591 , n10189 , n10190 , n177594 , n177595 , n177596 , n10194 , n177598 , 
 n177599 , n10197 , n177601 , n177602 , n10200 , n177604 , n177605 , n177606 , n177607 , n177608 , 
 n10206 , n177610 , n177611 , n10209 , n177613 , n177614 , n10212 , n177616 , n10214 , n177618 , 
 n10216 , n10217 , n177621 , n177622 , n10220 , n177624 , n177625 , n177626 , n177627 , n10225 , 
 n177629 , n177630 , n10228 , n177632 , n177633 , n10231 , n177635 , n177636 , n10234 , n177638 , 
 n10236 , n10237 , n177641 , n177642 , n177643 , n10244 , n177645 , n177646 , n177647 , n10248 , 
 n177649 , n10250 , n177651 , n177652 , n10253 , n177654 , n177655 , n10256 , n177657 , n10258 , 
 n177659 , n10260 , n177661 , n177662 , n10263 , n177664 , n10265 , n10266 , n177667 , n10268 , 
 n177669 , n177670 , n10271 , n177672 , n177673 , n10274 , n177675 , n10276 , n177677 , n10278 , 
 n177679 , n177680 , n10281 , n177682 , n10283 , n10284 , n177685 , n177686 , n177687 , n177688 , 
 n177689 , n10290 , n177691 , n177692 , n10293 , n177694 , n10295 , n10296 , n10297 , n10298 , 
 n10299 , n177700 , n177701 , n10302 , n177703 , n177704 , n10305 , n177706 , n10307 , n177708 , 
 n177709 , n10310 , n177711 , n177712 , n10313 , n177714 , n10315 , n177716 , n10317 , n177718 , 
 n177719 , n10320 , n177721 , n177722 , n10323 , n177724 , n177725 , n10326 , n177727 , n177728 , 
 n10329 , n177730 , n177731 , n177732 , n10333 , n177734 , n177735 , n10336 , n177737 , n177738 , 
 n10339 , n177740 , n177741 , n177742 , n10343 , n10344 , n177745 , n10346 , n177747 , n177748 , 
 n10349 , n177750 , n177751 , n177752 , n177753 , n10354 , n177755 , n177756 , n10357 , n177758 , 
 n10359 , n10360 , n177761 , n10362 , n177763 , n10364 , n177765 , n177766 , n10367 , n177768 , 
 n177769 , n10370 , n177771 , n177772 , n10373 , n177774 , n177775 , n10376 , n177777 , n10378 , 
 n10379 , n177780 , n177781 , n177782 , n177783 , n177784 , n10385 , n177786 , n177787 , n10388 , 
 n177789 , n177790 , n10391 , n177792 , n177793 , n177794 , n177795 , n10396 , n177797 , n177798 , 
 n10399 , n177800 , n10401 , n10402 , n177803 , n177804 , n10405 , n177806 , n177807 , n10408 , 
 n177809 , n177810 , n177811 , n177812 , n10413 , n177814 , n177815 , n10416 , n177817 , n10418 , 
 n177819 , n177820 , n10421 , n177822 , n177823 , n177824 , n10425 , n177826 , n177827 , n10428 , 
 n177829 , n177830 , n10431 , n177832 , n177833 , n10434 , n177835 , n177836 , n177837 , n177838 , 
 n10439 , n177840 , n177841 , n10442 , n177843 , n10444 , n10445 , n177846 , n177847 , n177848 , 
 n10449 , n177850 , n177851 , n10452 , n177853 , n177854 , n10455 , n177856 , n177857 , n10458 , 
 n177859 , n177860 , n10461 , n177862 , n177863 , n10464 , n177865 , n10466 , n10467 , n177868 , 
 n177869 , n177870 , n10471 , n177872 , n177873 , n10474 , n177875 , n177876 , n10477 , n177878 , 
 n177879 , n10480 , n10481 , n10482 , n177883 , n177884 , n10485 , n10486 , n10487 , n177888 , 
 n177889 , n10490 , n177891 , n177892 , n10493 , n177894 , n177895 , n10496 , n177897 , n10498 , 
 n10499 , n177900 , n177901 , n177902 , n10503 , n177904 , n177905 , n10506 , n177907 , n177908 , 
 n10509 , n177910 , n177911 , n177912 , n10516 , n10517 , n10518 , n10519 , n177917 , n177918 , 
 n10522 , n177920 , n10524 , n10525 , n177923 , n10527 , n10528 , n177926 , n177927 , n10531 , 
 n177929 , n177930 , n10534 , n177932 , n177933 , n10537 , n177935 , n10539 , n10540 , n177938 , 
 n177939 , n177940 , n10544 , n177942 , n177943 , n177944 , n177945 , n177946 , n10550 , n177948 , 
 n177949 , n10553 , n177951 , n177952 , n10556 , n177954 , n177955 , n177956 , n177957 , n10561 , 
 n177959 , n177960 , n10564 , n177962 , n10566 , n10567 , n177965 , n177966 , n177967 , n10571 , 
 n177969 , n177970 , n10574 , n177972 , n177973 , n10577 , n177975 , n177976 , n177977 , n10581 , 
 n177979 , n177980 , n10584 , n177982 , n10586 , n177984 , n177985 , n10589 , n10590 , n177988 , 
 n177989 , n177990 , n10594 , n177992 , n177993 , n10597 , n177995 , n177996 , n10600 , n177998 , 
 n10602 , n178000 , n178001 , n10605 , n178003 , n178004 , n10608 , n178006 , n10610 , n10611 , 
 n178009 , n178010 , n178011 , n10615 , n178013 , n178014 , n10618 , n178016 , n178017 , n10621 , 
 n178019 , n10623 , n178021 , n178022 , n10626 , n178024 , n10628 , n178026 , n10630 , n178028 , 
 n178029 , n10633 , n178031 , n178032 , n10636 , n178034 , n10638 , n10639 , n178037 , n178038 , 
 n178039 , n10643 , n178041 , n178042 , n10646 , n178044 , n178045 , n10649 , n178047 , n178048 , 
 n178049 , n178050 , n10654 , n178052 , n178053 , n10657 , n178055 , n10659 , n10660 , n178058 , 
 n178059 , n178060 , n10664 , n178062 , n178063 , n10667 , n178065 , n178066 , n10670 , n178068 , 
 n178069 , n10673 , n178071 , n178072 , n10676 , n178074 , n178075 , n10679 , n178077 , n10681 , 
 n10682 , n178080 , n10684 , n178082 , n10686 , n178084 , n178085 , n10689 , n178087 , n178088 , 
 n10692 , n10693 , n10694 , n178092 , n178093 , n10697 , n178095 , n178096 , n178097 , n178098 , 
 n10702 , n178100 , n178101 , n10705 , n178103 , n178104 , n10708 , n10709 , n10710 , n178108 , 
 n178109 , n178110 , n178111 , n10715 , n178113 , n178114 , n178115 , n10719 , n178117 , n10721 , 
 n10722 , n178120 , n178121 , n178122 , n10726 , n178124 , n178125 , n10729 , n178127 , n178128 , 
 n10732 , n178130 , n178131 , n10735 , n178133 , n10737 , n178135 , n10739 , n10740 , n178138 , 
 n178139 , n178140 , n10744 , n178142 , n178143 , n10747 , n178145 , n178146 , n10750 , n178148 , 
 n178149 , n10753 , n178151 , n178152 , n10756 , n178154 , n178155 , n10759 , n178157 , n178158 , 
 n178159 , n10763 , n178161 , n178162 , n10766 , n178164 , n10768 , n10769 , n178167 , n10771 , 
 n178169 , n178170 , n10774 , n178172 , n178173 , n10777 , n178175 , n10782 , n10783 , n178178 , 
 n178179 , n10786 , n178181 , n178182 , n10789 , n178184 , n10791 , n178186 , n10793 , n178188 , 
 n10795 , n10796 , n178191 , n178192 , n178193 , n10800 , n178195 , n178196 , n178197 , n178198 , 
 n178199 , n10806 , n178201 , n10808 , n10809 , n178204 , n10811 , n178206 , n10813 , n10814 , 
 n178209 , n10816 , n10817 , n178212 , n178213 , n10820 , n178215 , n178216 , n10823 , n178218 , 
 n10825 , n178220 , n10827 , n10828 , n178223 , n178224 , n10831 , n10832 , n178227 , n178228 , 
 n10835 , n178230 , n10837 , n178232 , n178233 , n10840 , n10841 , n178236 , n178237 , n178238 , 
 n10845 , n178240 , n178241 , n10848 , n178243 , n178244 , n10851 , n178246 , n178247 , n178248 , 
 n178249 , n10856 , n178251 , n178252 , n10859 , n178254 , n10861 , n10862 , n178257 , n178258 , 
 n10865 , n178260 , n178261 , n10868 , n178263 , n178264 , n10871 , n178266 , n178267 , n10874 , 
 n178269 , n178270 , n10877 , n178272 , n10879 , n10880 , n178275 , n178276 , n10883 , n178278 , 
 n178279 , n178280 , n10887 , n178282 , n178283 , n10890 , n178285 , n178286 , n10893 , n10894 , 
 n10895 , n178290 , n178291 , n10898 , n178293 , n178294 , n178295 , n178296 , n10903 , n178298 , 
 n10905 , n178300 , n178301 , n10908 , n178303 , n10910 , n178305 , n178306 , n10913 , n178308 , 
 n178309 , n10916 , n178311 , n178312 , n10919 , n10920 , n10921 , n178316 , n178317 , n10924 , 
 n178319 , n178320 , n178321 , n178322 , n10929 , n10930 , n178325 , n178326 , n178327 , n10934 , 
 n178329 , n178330 , n178331 , n10938 , n178333 , n178334 , n10941 , n178336 , n178337 , n10944 , 
 n178339 , n178340 , n10947 , n178342 , n10949 , n178344 , n10951 , n10952 , n178347 , n10954 , 
 n178349 , n10956 , n178351 , n178352 , n10959 , n178354 , n178355 , n178356 , n10963 , n178358 , 
 n10965 , n178360 , n178361 , n10968 , n10969 , n178364 , n10971 , n178366 , n10973 , n178368 , 
 n178369 , n10976 , n178371 , n178372 , n10979 , n10980 , n178375 , n10982 , n10983 , n178378 , 
 n10985 , n178380 , n10987 , n10988 , n178383 , n10990 , n10991 , n10992 , n178387 , n178388 , 
 n10995 , n178390 , n178391 , n10998 , n178393 , n11000 , n178395 , n11002 , n11003 , n178398 , 
 n178399 , n178400 , n11007 , n178402 , n178403 , n11010 , n178405 , n178406 , n11013 , n178408 , 
 n178409 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n178418 , 
 n11025 , n178420 , n11027 , n178422 , n11029 , n11030 , n178425 , n178426 , n178427 , n11034 , 
 n178429 , n178430 , n11037 , n178432 , n178433 , n11040 , n178435 , n178436 , n11043 , n11044 , 
 n11045 , n178440 , n178441 , n11048 , n11049 , n11050 , n178445 , n11052 , n178447 , n178448 , 
 n11055 , n178450 , n11057 , n178452 , n11059 , n178454 , n11061 , n178456 , n11063 , n11064 , 
 n178459 , n178460 , n178461 , n11068 , n178463 , n178464 , n11071 , n178466 , n178467 , n11077 , 
 n178469 , n11079 , n11080 , n178472 , n11082 , n178474 , n178475 , n178476 , n11086 , n178478 , 
 n178479 , n11089 , n178481 , n11091 , n11092 , n178484 , n178485 , n178486 , n11096 , n178488 , 
 n178489 , n11099 , n178491 , n178492 , n11102 , n178494 , n11104 , n178496 , n11106 , n11107 , 
 n178499 , n178500 , n11110 , n178502 , n11112 , n11113 , n11114 , n11115 , n178507 , n11117 , 
 n178509 , n178510 , n11120 , n178512 , n178513 , n178514 , n11124 , n178516 , n11126 , n11127 , 
 n178519 , n11129 , n178521 , n11131 , n178523 , n178524 , n11134 , n178526 , n178527 , n11137 , 
 n178529 , n11139 , n178531 , n11141 , n11142 , n178534 , n178535 , n178536 , n11146 , n178538 , 
 n178539 , n11149 , n178541 , n178542 , n11152 , n178544 , n178545 , n11155 , n178547 , n178548 , 
 n11158 , n178550 , n178551 , n11161 , n11162 , n11163 , n178555 , n178556 , n11166 , n178558 , 
 n178559 , n11169 , n178561 , n11171 , n11172 , n178564 , n178565 , n178566 , n11176 , n178568 , 
 n178569 , n11179 , n178571 , n178572 , n11182 , n178574 , n178575 , n11185 , n11186 , n11187 , 
 n178579 , n11189 , n178581 , n11191 , n178583 , n11193 , n178585 , n11195 , n178587 , n11197 , 
 n178589 , n11199 , n11200 , n178592 , n11202 , n178594 , n11204 , n178596 , n178597 , n11207 , 
 n178599 , n178600 , n11210 , n11211 , n11212 , n178604 , n178605 , n11215 , n11216 , n178608 , 
 n11218 , n11219 , n178611 , n178612 , n178613 , n178614 , n11224 , n11225 , n11226 , n11227 , 
 n178619 , n11229 , n178621 , n11231 , n178623 , n11233 , n11234 , n178626 , n178627 , n178628 , 
 n11238 , n178630 , n178631 , n11241 , n178633 , n178634 , n11244 , n178636 , n11246 , n178638 , 
 n11248 , n178640 , n11250 , n11251 , n178643 , n178644 , n178645 , n11255 , n178647 , n178648 , 
 n11258 , n178650 , n178651 , n11261 , n178653 , n11263 , n11264 , n11265 , n11266 , n11267 , 
 n11268 , n178660 , n178661 , n178662 , n11272 , n178664 , n178665 , n11275 , n178667 , n11277 , 
 n11278 , n11279 , n178671 , n178672 , n11282 , n178674 , n11284 , n11285 , n178677 , n178678 , 
 n178679 , n11289 , n178681 , n178682 , n11292 , n178684 , n178685 , n11295 , n178687 , n178688 , 
 n178689 , n178690 , n11300 , n178692 , n11302 , n11303 , n178695 , n11305 , n178697 , n11307 , 
 n178699 , n178700 , n11310 , n178702 , n178703 , n11313 , n11314 , n178706 , n178707 , n11317 , 
 n178709 , n11319 , n178711 , n11321 , n11322 , n178714 , n178715 , n178716 , n11326 , n178718 , 
 n178719 , n11329 , n178721 , n178722 , n11332 , n178724 , n178725 , n11335 , n178727 , n178728 , 
 n11338 , n178730 , n178731 , n11341 , n178733 , n11343 , n178735 , n11345 , n11346 , n178738 , 
 n178739 , n178740 , n11350 , n178742 , n178743 , n11353 , n178745 , n178746 , n11356 , n178748 , 
 n178749 , n178750 , n11363 , n178752 , n11365 , n11366 , n178755 , n178756 , n178757 , n11370 , 
 n178759 , n178760 , n11373 , n178762 , n178763 , n11376 , n178765 , n178766 , n11379 , n178768 , 
 n11381 , n178770 , n178771 , n11384 , n178773 , n178774 , n178775 , n11388 , n178777 , n178778 , 
 n11391 , n178780 , n178781 , n11394 , n178783 , n178784 , n11397 , n178786 , n178787 , n11400 , 
 n178789 , n11402 , n178791 , n11404 , n178793 , n178794 , n178795 , n11408 , n178797 , n178798 , 
 n11411 , n11412 , n178801 , n178802 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , 
 n11421 , n11422 , n11423 , n11424 , n11425 , n178814 , n11427 , n11428 , n11429 , n178818 , 
 n178819 , n11432 , n178821 , n178822 , n11435 , n178824 , n178825 , n11438 , n178827 , n11440 , 
 n11441 , n11442 , n178831 , n11444 , n11445 , n11446 , n11447 , n11448 , n178837 , n178838 , 
 n11451 , n11452 , n178841 , n11454 , n178843 , n178844 , n11457 , n11458 , n178847 , n11460 , 
 n11461 , n178850 , n11463 , n178852 , n11465 , n11466 , n178855 , n11468 , n178857 , n178858 , 
 n11471 , n178860 , n178861 , n11474 , n178863 , n178864 , n11477 , n178866 , n178867 , n11480 , 
 n178869 , n178870 , n178871 , n11484 , n178873 , n11486 , n11487 , n178876 , n178877 , n11490 , 
 n178879 , n178880 , n11493 , n178882 , n178883 , n11496 , n178885 , n11498 , n178887 , n11500 , 
 n11501 , n178890 , n178891 , n11504 , n178893 , n178894 , n11507 , n178896 , n178897 , n11510 , 
 n11511 , n11512 , n178901 , n178902 , n11515 , n11516 , n178905 , n11518 , n178907 , n11520 , 
 n178909 , n178910 , n11523 , n178912 , n178913 , n178914 , n178915 , n178916 , n11529 , n11530 , 
 n178919 , n178920 , n11533 , n178922 , n11535 , n178924 , n11537 , n178926 , n178927 , n178928 , 
 n11541 , n178930 , n178931 , n11544 , n178933 , n178934 , n178935 , n11548 , n178937 , n11550 , 
 n11551 , n178940 , n178941 , n11554 , n178943 , n178944 , n11557 , n178946 , n178947 , n11560 , 
 n178949 , n178950 , n178951 , n11564 , n11565 , n178954 , n178955 , n11568 , n178957 , n178958 , 
 n11571 , n178960 , n178961 , n11574 , n178963 , n178964 , n178965 , n11578 , n178967 , n11580 , 
 n178969 , n178970 , n11583 , n178972 , n11585 , n11586 , n178975 , n178976 , n11589 , n178978 , 
 n178979 , n11592 , n178981 , n11594 , n178983 , n11596 , n178985 , n11598 , n11599 , n178988 , 
 n178989 , n11602 , n178991 , n178992 , n11605 , n178994 , n11607 , n11608 , n11609 , n178998 , 
 n11611 , n179000 , n11613 , n11614 , n179003 , n179004 , n11617 , n179006 , n179007 , n11620 , 
 n179009 , n11622 , n11623 , n179012 , n11625 , n179014 , n11627 , n179016 , n11629 , n11630 , 
 n179019 , n11632 , n179021 , n11634 , n179023 , n179024 , n11637 , n179026 , n179027 , n179028 , 
 n11641 , n179030 , n11643 , n11644 , n179033 , n179034 , n11647 , n179036 , n179037 , n11650 , 
 n179039 , n179040 , n11653 , n179042 , n11655 , n179044 , n11657 , n11658 , n179047 , n179048 , 
 n11661 , n179050 , n179051 , n11664 , n179053 , n179054 , n11667 , n11668 , n11669 , n179058 , 
 n179059 , n179060 , n179061 , n179062 , n179063 , n179064 , n11680 , n179066 , n179067 , n11683 , 
 n179069 , n179070 , n11686 , n11687 , n11688 , n179074 , n179075 , n11691 , n179077 , n179078 , 
 n179079 , n179080 , n11696 , n179082 , n179083 , n11699 , n179085 , n179086 , n11702 , n11703 , 
 n11704 , n11705 , n11706 , n179092 , n11708 , n179094 , n11710 , n179096 , n11712 , n179098 , 
 n11714 , n11715 , n11716 , n179102 , n179103 , n179104 , n11720 , n179106 , n179107 , n11723 , 
 n179109 , n11725 , n179111 , n11727 , n179113 , n179114 , n11730 , n179116 , n11732 , n179118 , 
 n179119 , n11735 , n11736 , n179122 , n11738 , n179124 , n11740 , n179126 , n179127 , n11743 , 
 n179129 , n11745 , n11746 , n179132 , n11748 , n179134 , n11750 , n11751 , n179137 , n179138 , 
 n179139 , n11755 , n179141 , n179142 , n11758 , n179144 , n179145 , n11761 , n179147 , n11763 , 
 n11764 , n11765 , n11766 , n179152 , n11768 , n179154 , n11770 , n179156 , n11772 , n179158 , 
 n179159 , n11775 , n179161 , n11777 , n179163 , n179164 , n11780 , n179166 , n11782 , n179168 , 
 n11784 , n179170 , n11786 , n11787 , n179173 , n179174 , n179175 , n11791 , n179177 , n179178 , 
 n11794 , n179180 , n179181 , n11797 , n179183 , n11799 , n11800 , n179186 , n11802 , n179188 , 
 n11804 , n11805 , n179191 , n11807 , n179193 , n179194 , n11810 , n179196 , n11812 , n11813 , 
 n179199 , n179200 , n179201 , n11817 , n179203 , n179204 , n11820 , n179206 , n179207 , n11823 , 
 n179209 , n11825 , n179211 , n179212 , n11828 , n179214 , n11830 , n11831 , n179217 , n179218 , 
 n179219 , n11835 , n179221 , n179222 , n11838 , n179224 , n179225 , n11841 , n179227 , n179228 , 
 n11844 , n11845 , n179231 , n11847 , n179233 , n179234 , n11850 , n11851 , n179237 , n11853 , 
 n179239 , n11855 , n11856 , n11857 , n11858 , n11859 , n179245 , n179246 , n179247 , n11863 , 
 n179249 , n11865 , n11866 , n179252 , n179253 , n179254 , n11870 , n179256 , n179257 , n11873 , 
 n179259 , n179260 , n11876 , n179262 , n179263 , n11879 , n179265 , n11881 , n11882 , n179268 , 
 n11884 , n179270 , n11886 , n179272 , n179273 , n11889 , n179275 , n11891 , n179277 , n11893 , 
 n179279 , n11895 , n11896 , n179282 , n11898 , n179284 , n11900 , n179286 , n179287 , n11903 , 
 n179289 , n11905 , n179291 , n11907 , n11908 , n11909 , n11910 , n11911 , n179297 , n179298 , 
 n11914 , n179300 , n179301 , n11917 , n179303 , n179304 , n11920 , n11921 , n11922 , n179308 , 
 n179309 , n11925 , n11926 , n179312 , n179313 , n11929 , n179315 , n11931 , n179317 , n11933 , 
 n11934 , n179320 , n179321 , n11937 , n179323 , n179324 , n11940 , n179326 , n179327 , n179328 , 
 n11944 , n179330 , n11946 , n11947 , n179333 , n179334 , n11950 , n179336 , n179337 , n11953 , 
 n179339 , n179340 , n11956 , n179342 , n11958 , n179344 , n11960 , n11961 , n179347 , n179348 , 
 n11964 , n179350 , n179351 , n11967 , n179353 , n179354 , n11970 , n11971 , n11972 , n179358 , 
 n179359 , n11975 , n11976 , n179362 , n179363 , n11982 , n11983 , n11984 , n179367 , n11986 , 
 n179369 , n11988 , n179371 , n11990 , n179373 , n11992 , n179375 , n179376 , n11995 , n11996 , 
 n179379 , n11998 , n179381 , n179382 , n12001 , n12002 , n179385 , n179386 , n179387 , n12006 , 
 n179389 , n179390 , n179391 , n12010 , n179393 , n12012 , n12013 , n179396 , n179397 , n12016 , 
 n12017 , n12018 , n12019 , n179402 , n179403 , n12022 , n12023 , n179406 , n179407 , n12026 , 
 n179409 , n12028 , n179411 , n12030 , n12031 , n179414 , n12033 , n12034 , n12035 , n179418 , 
 n179419 , n12038 , n179421 , n179422 , n179423 , n12042 , n179425 , n12044 , n179427 , n179428 , 
 n12047 , n179430 , n179431 , n12050 , n179433 , n179434 , n179435 , n179436 , n12055 , n179438 , 
 n179439 , n12058 , n179441 , n179442 , n12061 , n179444 , n179445 , n12064 , n179447 , n12066 , 
 n179449 , n12068 , n12069 , n179452 , n179453 , n12072 , n12073 , n179456 , n179457 , n179458 , 
 n12077 , n179460 , n179461 , n12080 , n179463 , n179464 , n12083 , n12084 , n179467 , n179468 , 
 n12087 , n12088 , n12089 , n179472 , n179473 , n12092 , n12093 , n12094 , n179477 , n179478 , 
 n12097 , n12098 , n179481 , n12100 , n179483 , n12102 , n179485 , n12104 , n179487 , n12106 , 
 n12107 , n179490 , n179491 , n12110 , n12111 , n179494 , n179495 , n12114 , n12115 , n179498 , 
 n179499 , n12118 , n12119 , n179502 , n179503 , n12122 , n179505 , n179506 , n12125 , n12126 , 
 n12127 , n179510 , n12129 , n179512 , n179513 , n12132 , n179515 , n12134 , n179517 , n179518 , 
 n12137 , n12138 , n179521 , n179522 , n12141 , n12142 , n179525 , n12144 , n179527 , n12146 , 
 n179529 , n12148 , n12149 , n12150 , n12151 , n179534 , n179535 , n12154 , n179537 , n179538 , 
 n179539 , n179540 , n12159 , n179542 , n179543 , n12162 , n179545 , n179546 , n12165 , n12166 , 
 n179549 , n12168 , n179551 , n12170 , n179553 , n179554 , n12173 , n179556 , n12175 , n12176 , 
 n12177 , n12178 , n12179 , n179562 , n179563 , n12182 , n12183 , n12184 , n179567 , n179568 , 
 n12187 , n12188 , n179571 , n179572 , n12191 , n12192 , n12193 , n179576 , n179577 , n12196 , 
 n179579 , n179580 , n12199 , n179582 , n179583 , n12202 , n179585 , n179586 , n12205 , n179588 , 
 n12207 , n179590 , n12209 , n179592 , n12211 , n179594 , n12213 , n12214 , n179597 , n179598 , 
 n12217 , n179600 , n179601 , n12220 , n179603 , n179604 , n12223 , n179606 , n179607 , n12226 , 
 n12227 , n12228 , n12229 , n12230 , n12231 , n179614 , n179615 , n12234 , n179617 , n179618 , 
 n179619 , n179620 , n12239 , n179622 , n179623 , n12242 , n179625 , n179626 , n12245 , n12246 , 
 n12247 , n12248 , n179631 , n179632 , n12251 , n12252 , n12253 , n12254 , n179637 , n179638 , 
 n12257 , n179640 , n12259 , n179642 , n12261 , n179644 , n179645 , n12264 , n12265 , n179648 , 
 n12267 , n179650 , n179651 , n179652 , n179653 , n12272 , n179655 , n179656 , n12275 , n179658 , 
 n179659 , n12278 , n12279 , n12280 , n179663 , n179664 , n12283 , n12284 , n12285 , n179668 , 
 n12287 , n12288 , n12289 , n179672 , n12291 , n12292 , n179675 , n12294 , n179677 , n12296 , 
 n12297 , n179680 , n179681 , n12300 , n12301 , n179684 , n179685 , n12304 , n179687 , n12306 , 
 n12307 , n12308 , n179691 , n12310 , n12311 , n179694 , n12316 , n12317 , n12318 , n12319 , 
 n179699 , n179700 , n12322 , n12323 , n179703 , n179704 , n12326 , n179706 , n179707 , n12329 , 
 n179709 , n179710 , n12332 , n179712 , n12334 , n12335 , n179715 , n179716 , n179717 , n12339 , 
 n179719 , n12341 , n12342 , n179722 , n12344 , n12345 , n179725 , n12347 , n179727 , n179728 , 
 n12350 , n179730 , n12352 , n179732 , n12354 , n12355 , n179735 , n12357 , n179737 , n179738 , 
 n179739 , n12361 , n179741 , n12363 , n179743 , n179744 , n12366 , n179746 , n179747 , n179748 , 
 n12370 , n179750 , n12372 , n12373 , n179753 , n179754 , n12376 , n12377 , n179757 , n12379 , 
 n179759 , n12381 , n12382 , n12383 , n179763 , n179764 , n12386 , n179766 , n179767 , n179768 , 
 n179769 , n12391 , n179771 , n179772 , n12394 , n179774 , n12396 , n12397 , n12398 , n12399 , 
 n12400 , n179780 , n12402 , n12403 , n12404 , n179784 , n12406 , n179786 , n12408 , n179788 , 
 n179789 , n12411 , n179791 , n12413 , n12414 , n179794 , n12416 , n179796 , n179797 , n179798 , 
 n179799 , n12421 , n179801 , n179802 , n12424 , n179804 , n12426 , n179806 , n12428 , n179808 , 
 n12430 , n12431 , n179811 , n179812 , n12434 , n179814 , n179815 , n179816 , n12438 , n179818 , 
 n179819 , n12441 , n179821 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
 n179829 , n12451 , n179831 , n179832 , n12454 , n179834 , n12456 , n12457 , n179837 , n12459 , 
 n179839 , n179840 , n179841 , n179842 , n12464 , n179844 , n179845 , n12467 , n179847 , n12469 , 
 n12470 , n12471 , n12472 , n12473 , n179853 , n12475 , n179855 , n179856 , n12478 , n179858 , 
 n179859 , n12481 , n179861 , n179862 , n179863 , n179864 , n12486 , n179866 , n179867 , n12489 , 
 n179869 , n12491 , n12492 , n12493 , n12494 , n12495 , n179875 , n12497 , n12498 , n179878 , 
 n179879 , n179880 , n12502 , n12503 , n12504 , n179884 , n12506 , n12507 , n12508 , n179888 , 
 n12510 , n12511 , n179891 , n12513 , n179893 , n12515 , n12516 , n179896 , n12518 , n179898 , 
 n179899 , n179900 , n12522 , n179902 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
 n12530 , n179910 , n12532 , n12533 , n179913 , n12535 , n179915 , n179916 , n12538 , n12539 , 
 n12540 , n12541 , n179921 , n12543 , n179923 , n179924 , n12546 , n12547 , n12548 , n12549 , 
 n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n179936 , n179937 , n12559 , 
 n179939 , n179940 , n12562 , n12563 , n179943 , n12565 , n12566 , n179946 , n179947 , n12569 , 
 n179949 , n12571 , n12572 , n12573 , n179953 , n12575 , n179955 , n12577 , n12578 , n12579 , 
 n12580 , n12581 , n179961 , n12583 , n179963 , n12585 , n179965 , n12587 , n179967 , n179968 , 
 n12590 , n12591 , n179971 , n12593 , n179973 , n12595 , n179975 , n179976 , n12598 , n179978 , 
 n12600 , n12601 , n179981 , n12603 , n179983 , n179984 , n12606 , n179986 , n179987 , n12609 , 
 n12610 , n179990 , n179991 , n12613 , n179993 , n179994 , n12616 , n179996 , n12618 , n12619 , 
 n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
 n12630 , n12631 , n180011 , n12633 , n12634 , n180014 , n180015 , n12637 , n180017 , n12642 , 
 n12643 , n12644 , n12645 , n12646 , n180023 , n12648 , n12649 , n180026 , n12651 , n180028 , 
 n180029 , n12654 , n180031 , n180032 , n12657 , n12658 , n180035 , n12660 , n12661 , n180038 , 
 n180039 , n12664 , n12665 , n12666 , n12667 , n12668 , n180045 , n180046 , n180047 , n12672 , 
 n180049 , n180050 , n180051 , n12676 , n180053 , n12678 , n12679 , n180056 , n180057 , n12682 , 
 n12683 , n180060 , n180061 , n12686 , n180063 , n180064 , n12689 , n12690 , n12691 , n12692 , 
 n12693 , n180070 , n180071 , n12696 , n12697 , n12698 , n180075 , n180076 , n12701 , n12702 , 
 n180079 , n12704 , n180081 , n180082 , n12707 , n180084 , n12709 , n180086 , n180087 , n12712 , 
 n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n180096 , n180097 , n180098 , 
 n180099 , n180100 , n180101 , n12726 , n180103 , n180104 , n180105 , n180106 , n180107 , n12732 , 
 n180109 , n180110 , n12735 , n180112 , n180113 , n12738 , n180115 , n12740 , n180117 , n12742 , 
 n12743 , n180120 , n12745 , n12746 , n12747 , n12748 , n180125 , n180126 , n12751 , n180128 , 
 n12753 , n180130 , n12755 , n12756 , n180133 , n12758 , n180135 , n180136 , n180137 , n12762 , 
 n12763 , n180140 , n12765 , n180142 , n180143 , n12768 , n180145 , n180146 , n12771 , n12772 , 
 n12773 , n180150 , n180151 , n12776 , n180153 , n180154 , n12779 , n180156 , n12781 , n12782 , 
 n180159 , n180160 , n12785 , n180162 , n12787 , n12788 , n180165 , n180166 , n180167 , n12792 , 
 n180169 , n180170 , n12795 , n180172 , n180173 , n12798 , n180175 , n180176 , n180177 , n12802 , 
 n180179 , n12804 , n12805 , n180182 , n180183 , n180184 , n12809 , n180186 , n180187 , n12812 , 
 n180189 , n180190 , n12815 , n180192 , n180193 , n12818 , n180195 , n12820 , n180197 , n180198 , 
 n180199 , n180200 , n12825 , n12826 , n180203 , n180204 , n180205 , n12830 , n180207 , n180208 , 
 n12833 , n180210 , n180211 , n12836 , n180213 , n180214 , n12839 , n180216 , n180217 , n12842 , 
 n180219 , n180220 , n12845 , n180222 , n180223 , n180224 , n12849 , n180226 , n12851 , n12852 , 
 n180229 , n180230 , n180231 , n12856 , n180233 , n180234 , n12859 , n180236 , n180237 , n12862 , 
 n180239 , n180240 , n12865 , n180242 , n12867 , n180244 , n12869 , n12870 , n180247 , n180248 , 
 n12873 , n180250 , n180251 , n12876 , n180253 , n12878 , n180255 , n180256 , n12881 , n180258 , 
 n180259 , n12884 , n180261 , n180262 , n12887 , n180264 , n180265 , n12890 , n12891 , n12892 , 
 n12893 , n12894 , n180271 , n180272 , n12897 , n180274 , n180275 , n12900 , n12901 , n12902 , 
 n12903 , n180280 , n180281 , n12906 , n12907 , n12908 , n12909 , n180286 , n180287 , n12912 , 
 n180289 , n12914 , n12915 , n12916 , n12917 , n180294 , n180295 , n12920 , n180297 , n12922 , 
 n12923 , n12924 , n180301 , n12926 , n180303 , n12928 , n12929 , n180306 , n180307 , n180308 , 
 n12933 , n180310 , n180311 , n12936 , n180313 , n180314 , n12939 , n180316 , n12941 , n180318 , 
 n180319 , n12944 , n180321 , n12946 , n12947 , n180324 , n180325 , n180326 , n12951 , n180328 , 
 n180329 , n12954 , n180331 , n180332 , n12957 , n180334 , n12959 , n12960 , n12961 , n180338 , 
 n180339 , n12964 , n180341 , n12966 , n12967 , n12968 , n180345 , n12970 , n180347 , n12972 , 
 n12973 , n180350 , n12975 , n180352 , n12977 , n180354 , n180355 , n12980 , n180357 , n12982 , 
 n180359 , n12984 , n180361 , n12986 , n180363 , n12988 , n12989 , n180366 , n180367 , n180368 , 
 n12996 , n180370 , n180371 , n12999 , n180373 , n180374 , n13002 , n180376 , n180377 , n180378 , 
 n13006 , n180380 , n13008 , n13009 , n180383 , n180384 , n180385 , n13013 , n180387 , n180388 , 
 n13016 , n180390 , n180391 , n13019 , n180393 , n180394 , n13022 , n180396 , n180397 , n13025 , 
 n180399 , n13027 , n180401 , n180402 , n13030 , n180404 , n13032 , n13033 , n180407 , n13035 , 
 n180409 , n180410 , n13038 , n180412 , n13040 , n180414 , n180415 , n13043 , n180417 , n180418 , 
 n13046 , n180420 , n180421 , n180422 , n13050 , n180424 , n13052 , n13053 , n180427 , n180428 , 
 n13056 , n180430 , n13058 , n180432 , n180433 , n13061 , n180435 , n180436 , n13064 , n13065 , 
 n13066 , n13067 , n13068 , n180442 , n180443 , n13071 , n13072 , n13073 , n13074 , n180448 , 
 n180449 , n13077 , n180451 , n180452 , n13080 , n180454 , n180455 , n180456 , n180457 , n13085 , 
 n180459 , n13087 , n180461 , n180462 , n13090 , n180464 , n180465 , n180466 , n13094 , n180468 , 
 n13096 , n13097 , n180471 , n13099 , n180473 , n13101 , n180475 , n180476 , n13104 , n13105 , 
 n180479 , n13107 , n180481 , n180482 , n13110 , n180484 , n180485 , n13113 , n13114 , n13115 , 
 n13116 , n13117 , n180491 , n180492 , n13120 , n180494 , n180495 , n13123 , n180497 , n180498 , 
 n13126 , n180500 , n180501 , n13129 , n180503 , n180504 , n13132 , n13133 , n13134 , n13135 , 
 n180509 , n180510 , n13138 , n180512 , n180513 , n13141 , n13142 , n180516 , n13144 , n13145 , 
 n180519 , n180520 , n13148 , n13149 , n13150 , n13151 , n180525 , n180526 , n13154 , n180528 , 
 n180529 , n13157 , n180531 , n180532 , n13160 , n180534 , n180535 , n13163 , n13164 , n180538 , 
 n13166 , n13167 , n180541 , n13169 , n13170 , n180544 , n13172 , n180546 , n180547 , n180548 , 
 n13176 , n180550 , n180551 , n13179 , n180553 , n180554 , n180555 , n180556 , n13184 , n180558 , 
 n180559 , n13187 , n180561 , n180562 , n13190 , n180564 , n180565 , n13193 , n180567 , n13195 , 
 n13196 , n180570 , n13198 , n180572 , n13200 , n180574 , n180575 , n13203 , n13204 , n180578 , 
 n13206 , n180580 , n180581 , n13209 , n180583 , n180584 , n13212 , n180586 , n13214 , n13215 , 
 n180589 , n13217 , n13218 , n13219 , n13220 , n13221 , n180595 , n180596 , n13224 , n13225 , 
 n13226 , n13227 , n180601 , n180602 , n13230 , n13231 , n13232 , n13233 , n13234 , n180608 , 
 n13236 , n13237 , n13238 , n13239 , n180613 , n13241 , n13242 , n13243 , n13244 , n180618 , 
 n180619 , n180620 , n13248 , n180622 , n13250 , n13251 , n180625 , n180626 , n180627 , n13255 , 
 n180629 , n180630 , n13258 , n180632 , n180633 , n13261 , n180635 , n180636 , n180637 , n13265 , 
 n180639 , n13267 , n13268 , n180642 , n180643 , n180644 , n13272 , n180646 , n180647 , n13275 , 
 n180649 , n180650 , n13278 , n180652 , n180653 , n13281 , n180655 , n180656 , n13284 , n180658 , 
 n180659 , n13287 , n180661 , n13289 , n180663 , n180664 , n180665 , n180666 , n13294 , n180668 , 
 n180669 , n13297 , n180671 , n180672 , n13300 , n13301 , n180675 , n180676 , n13304 , n180678 , 
 n180679 , n13307 , n180681 , n13309 , n180683 , n13311 , n13312 , n180686 , n180687 , n180688 , 
 n13316 , n180690 , n180691 , n13319 , n180693 , n180694 , n13325 , n180696 , n13327 , n180698 , 
 n13329 , n180700 , n13331 , n13332 , n180703 , n180704 , n180705 , n13336 , n180707 , n180708 , 
 n13339 , n180710 , n180711 , n13342 , n180713 , n13344 , n180715 , n13346 , n180717 , n13348 , 
 n13349 , n180720 , n13351 , n180722 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , 
 n13359 , n13360 , n13361 , n13362 , n180733 , n13364 , n180735 , n13366 , n180737 , n13368 , 
 n180739 , n13370 , n13371 , n180742 , n180743 , n180744 , n13375 , n180746 , n180747 , n13378 , 
 n180749 , n180750 , n13381 , n180752 , n180753 , n13384 , n180755 , n180756 , n13387 , n180758 , 
 n13389 , n13390 , n180761 , n13392 , n13393 , n180764 , n180765 , n180766 , n13397 , n180768 , 
 n180769 , n13400 , n180771 , n180772 , n13403 , n180774 , n180775 , n13406 , n13407 , n180778 , 
 n180779 , n13410 , n13411 , n180782 , n180783 , n13414 , n180785 , n13416 , n13417 , n180788 , 
 n180789 , n180790 , n13421 , n180792 , n180793 , n13424 , n180795 , n180796 , n13427 , n180798 , 
 n13429 , n13430 , n180801 , n13432 , n180803 , n13434 , n13435 , n180806 , n13437 , n180808 , 
 n13439 , n13440 , n180811 , n180812 , n180813 , n13444 , n180815 , n180816 , n13447 , n180818 , 
 n180819 , n13450 , n180821 , n180822 , n13453 , n13454 , n13455 , n13456 , n180827 , n13458 , 
 n180829 , n13460 , n180831 , n13462 , n180833 , n13464 , n180835 , n13466 , n180837 , n13468 , 
 n13469 , n180840 , n180841 , n180842 , n13473 , n180844 , n180845 , n13476 , n180847 , n180848 , 
 n13479 , n180850 , n180851 , n13482 , n180853 , n13484 , n13485 , n13486 , n13487 , n13488 , 
 n180859 , n180860 , n180861 , n13492 , n180863 , n180864 , n180865 , n13496 , n180867 , n13498 , 
 n180869 , n13500 , n13501 , n180872 , n180873 , n180874 , n13505 , n180876 , n180877 , n13508 , 
 n180879 , n180880 , n13511 , n180882 , n180883 , n13514 , n180885 , n180886 , n13517 , n13518 , 
 n180889 , n13520 , n180891 , n180892 , n13523 , n13524 , n180895 , n13526 , n13527 , n13528 , 
 n13529 , n13530 , n13531 , n180902 , n180903 , n13534 , n13535 , n13536 , n13537 , n180908 , 
 n180909 , n180910 , n13541 , n180912 , n13543 , n13544 , n13545 , n13546 , n180917 , n13548 , 
 n180919 , n180920 , n180921 , n13552 , n180923 , n13554 , n13555 , n180926 , n180927 , n13558 , 
 n180929 , n13560 , n180931 , n180932 , n13563 , n180934 , n180935 , n13566 , n13567 , n13568 , 
 n13569 , n13570 , n180941 , n180942 , n13573 , n180944 , n180945 , n13576 , n13577 , n13578 , 
 n13579 , n13580 , n180951 , n180952 , n13583 , n180954 , n180955 , n13586 , n13587 , n13588 , 
 n13589 , n13590 , n180961 , n180962 , n13593 , n180964 , n13595 , n180966 , n13597 , n180968 , 
 n180969 , n13600 , n180971 , n180972 , n13603 , n13604 , n180975 , n180976 , n13607 , n180978 , 
 n180979 , n13610 , n180981 , n180982 , n13613 , n180984 , n180985 , n13616 , n180987 , n180988 , 
 n13619 , n180990 , n180991 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , 
 n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , 
 n181009 , n13640 , n13641 , n181012 , n181013 , n13647 , n13648 , n13649 , n13650 , n13651 , 
 n13652 , n13653 , n13654 , n13655 , n13656 , n181024 , n13658 , n13659 , n13660 , n13661 , 
 n181029 , n181030 , n13664 , n181032 , n13666 , n181034 , n181035 , n13669 , n181037 , n181038 , 
 n13672 , n181040 , n13674 , n181042 , n13676 , n181044 , n13678 , n181046 , n181047 , n13681 , 
 n13682 , n181050 , n13684 , n13685 , n181053 , n181054 , n13688 , n181056 , n181057 , n13691 , 
 n181059 , n181060 , n13694 , n181062 , n13696 , n13697 , n13698 , n13699 , n181067 , n13701 , 
 n181069 , n181070 , n13704 , n181072 , n181073 , n13707 , n181075 , n181076 , n13710 , n181078 , 
 n181079 , n13713 , n181081 , n181082 , n13716 , n181084 , n181085 , n13719 , n181087 , n13721 , 
 n13722 , n13723 , n13724 , n181092 , n181093 , n13727 , n181095 , n13729 , n13730 , n181098 , 
 n181099 , n13733 , n181101 , n181102 , n13736 , n181104 , n181105 , n13739 , n181107 , n13741 , 
 n181109 , n13743 , n13744 , n181112 , n181113 , n181114 , n13748 , n181116 , n181117 , n13751 , 
 n181119 , n181120 , n13754 , n181122 , n181123 , n13757 , n181125 , n181126 , n181127 , n13761 , 
 n181129 , n13763 , n13764 , n181132 , n181133 , n181134 , n13768 , n181136 , n181137 , n13771 , 
 n181139 , n181140 , n13774 , n181142 , n181143 , n13777 , n181145 , n181146 , n13780 , n181148 , 
 n13782 , n181150 , n13784 , n13785 , n181153 , n181154 , n181155 , n13789 , n181157 , n181158 , 
 n13792 , n181160 , n181161 , n13795 , n181163 , n181164 , n13798 , n181166 , n13800 , n13801 , 
 n181169 , n181170 , n181171 , n13805 , n181173 , n181174 , n13808 , n181176 , n181177 , n13811 , 
 n181179 , n13813 , n181181 , n13815 , n13816 , n181184 , n181185 , n13819 , n13820 , n181188 , 
 n181189 , n13823 , n181191 , n13825 , n181193 , n13827 , n13828 , n181196 , n181197 , n181198 , 
 n13832 , n181200 , n181201 , n13835 , n181203 , n181204 , n13838 , n181206 , n181207 , n13841 , 
 n181209 , n13843 , n13844 , n181212 , n13846 , n181214 , n13848 , n181216 , n181217 , n13851 , 
 n181219 , n181220 , n13854 , n181222 , n13856 , n181224 , n13858 , n181226 , n13860 , n13861 , 
 n181229 , n13863 , n181231 , n13865 , n181233 , n181234 , n13868 , n181236 , n13870 , n181238 , 
 n13872 , n181240 , n181241 , n13875 , n13876 , n13877 , n13878 , n181246 , n181247 , n13881 , 
 n13882 , n13883 , n13884 , n13885 , n181253 , n181254 , n13888 , n13889 , n13890 , n13891 , 
 n181259 , n181260 , n13894 , n181262 , n13896 , n181264 , n13898 , n13899 , n181267 , n181268 , 
 n181269 , n13903 , n181271 , n181272 , n13906 , n181274 , n181275 , n13909 , n181277 , n181278 , 
 n13912 , n181280 , n181281 , n13915 , n13916 , n13917 , n13918 , n181286 , n181287 , n13921 , 
 n13922 , n13923 , n13924 , n13925 , n181293 , n181294 , n13928 , n181296 , n181297 , n13931 , 
 n181299 , n181300 , n13934 , n181302 , n181303 , n181304 , n13938 , n181306 , n13940 , n13941 , 
 n181309 , n181310 , n13944 , n181312 , n13946 , n181314 , n181315 , n13949 , n181317 , n13951 , 
 n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , 
 n13962 , n181330 , n181331 , n181332 , n13966 , n181334 , n181335 , n13969 , n181337 , n181338 , 
 n181339 , n13976 , n181341 , n13978 , n13979 , n181344 , n181345 , n181346 , n13983 , n181348 , 
 n181349 , n13986 , n181351 , n181352 , n13989 , n181354 , n181355 , n13992 , n181357 , n13994 , 
 n181359 , n13996 , n13997 , n181362 , n181363 , n181364 , n14001 , n181366 , n181367 , n14004 , 
 n181369 , n181370 , n14007 , n181372 , n181373 , n14010 , n181375 , n181376 , n14013 , n181378 , 
 n181379 , n14016 , n14017 , n181382 , n14019 , n14020 , n181385 , n181386 , n181387 , n181388 , 
 n14025 , n14026 , n181391 , n14028 , n181393 , n181394 , n181395 , n181396 , n14033 , n181398 , 
 n181399 , n14036 , n181401 , n181402 , n14039 , n14040 , n14041 , n14042 , n14043 , n181408 , 
 n181409 , n14046 , n181411 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , 
 n14055 , n14056 , n181421 , n14058 , n181423 , n14060 , n14061 , n14062 , n14063 , n14064 , 
 n181429 , n14066 , n181431 , n14068 , n14069 , n14070 , n14071 , n181436 , n14073 , n14074 , 
 n14075 , n14076 , n14077 , n14078 , n181443 , n181444 , n14081 , n181446 , n14083 , n181448 , 
 n14085 , n14086 , n181451 , n14088 , n181453 , n14090 , n181455 , n181456 , n14093 , n181458 , 
 n181459 , n14096 , n181461 , n14098 , n14099 , n181464 , n14101 , n181466 , n14103 , n181468 , 
 n181469 , n14106 , n181471 , n14108 , n181473 , n14110 , n181475 , n14112 , n14113 , n181478 , 
 n181479 , n181480 , n14117 , n181482 , n181483 , n14120 , n181485 , n181486 , n14123 , n181488 , 
 n14125 , n14126 , n181491 , n14128 , n181493 , n14130 , n14131 , n181496 , n181497 , n14134 , 
 n181499 , n181500 , n181501 , n14138 , n181503 , n181504 , n14141 , n181506 , n181507 , n14144 , 
 n181509 , n14146 , n181511 , n181512 , n14149 , n14150 , n181515 , n14152 , n181517 , n14154 , 
 n181519 , n14156 , n181521 , n14158 , n14159 , n181524 , n181525 , n181526 , n14163 , n181528 , 
 n181529 , n14166 , n181531 , n181532 , n14169 , n181534 , n14171 , n14172 , n181537 , n14174 , 
 n181539 , n14176 , n14177 , n181542 , n181543 , n181544 , n14181 , n181546 , n181547 , n14184 , 
 n181549 , n181550 , n14187 , n181552 , n181553 , n14190 , n181555 , n181556 , n181557 , n14194 , 
 n181559 , n14196 , n14197 , n181562 , n181563 , n181564 , n14201 , n181566 , n181567 , n14204 , 
 n181569 , n181570 , n14207 , n181572 , n181573 , n14210 , n14211 , n181576 , n14213 , n181578 , 
 n181579 , n14216 , n14217 , n181582 , n181583 , n181584 , n14221 , n181586 , n14223 , n181588 , 
 n181589 , n14226 , n14227 , n181592 , n14229 , n181594 , n181595 , n181596 , n181597 , n14234 , 
 n181599 , n181600 , n14237 , n181602 , n181603 , n14240 , n181605 , n181606 , n14243 , n181608 , 
 n14245 , n181610 , n14247 , n14248 , n181613 , n181614 , n14251 , n14252 , n181617 , n181618 , 
 n181619 , n181620 , n14257 , n181622 , n181623 , n181624 , n14261 , n181626 , n14263 , n14264 , 
 n14265 , n14266 , n181631 , n14268 , n181633 , n181634 , n14271 , n181636 , n14273 , n181638 , 
 n14275 , n14276 , n14277 , n181642 , n181643 , n181644 , n14281 , n181646 , n181647 , n14284 , 
 n181649 , n181650 , n14287 , n181652 , n181653 , n14290 , n181655 , n181656 , n14293 , n181658 , 
 n14298 , n14299 , n181661 , n14301 , n181663 , n14303 , n181665 , n181666 , n14306 , n14307 , 
 n181669 , n14309 , n181671 , n181672 , n14312 , n181674 , n181675 , n14315 , n181677 , n14317 , 
 n181679 , n14319 , n181681 , n14321 , n14322 , n181684 , n181685 , n181686 , n14326 , n181688 , 
 n181689 , n14329 , n181691 , n181692 , n14332 , n181694 , n181695 , n14335 , n181697 , n181698 , 
 n14338 , n14339 , n181701 , n181702 , n14342 , n14343 , n181705 , n181706 , n14346 , n14347 , 
 n181709 , n181710 , n14350 , n14351 , n181713 , n14353 , n14354 , n14355 , n14356 , n14357 , 
 n181719 , n14359 , n14360 , n14361 , n14362 , n181724 , n14364 , n14365 , n181727 , n14367 , 
 n14368 , n181730 , n181731 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , 
 n14378 , n181740 , n14380 , n14381 , n14382 , n14383 , n14384 , n181746 , n181747 , n14387 , 
 n181749 , n14389 , n181751 , n181752 , n181753 , n14393 , n181755 , n14395 , n181757 , n181758 , 
 n181759 , n181760 , n14400 , n181762 , n181763 , n14403 , n181765 , n181766 , n14406 , n14407 , 
 n14408 , n14409 , n14410 , n181772 , n181773 , n14413 , n181775 , n181776 , n14416 , n14417 , 
 n14418 , n14419 , n14420 , n181782 , n181783 , n14423 , n181785 , n181786 , n14426 , n14427 , 
 n14428 , n14429 , n181791 , n181792 , n14432 , n14433 , n14434 , n14435 , n14436 , n181798 , 
 n181799 , n14439 , n181801 , n181802 , n14442 , n14443 , n14444 , n14445 , n14446 , n181808 , 
 n14448 , n181810 , n181811 , n14451 , n181813 , n181814 , n14454 , n14455 , n14456 , n14457 , 
 n14458 , n181820 , n181821 , n14461 , n14462 , n181824 , n14464 , n181826 , n181827 , n181828 , 
 n14468 , n181830 , n181831 , n14471 , n181833 , n14473 , n14474 , n181836 , n14476 , n14477 , 
 n181839 , n14479 , n14480 , n181842 , n14482 , n181844 , n181845 , n181846 , n14486 , n181848 , 
 n181849 , n14489 , n181851 , n181852 , n181853 , n181854 , n14494 , n181856 , n181857 , n14497 , 
 n181859 , n14499 , n181861 , n181862 , n14502 , n181864 , n14504 , n14505 , n181867 , n181868 , 
 n181869 , n14509 , n181871 , n181872 , n14512 , n181874 , n181875 , n14515 , n181877 , n181878 , 
 n14518 , n14519 , n14520 , n181882 , n181883 , n181884 , n14524 , n181886 , n181887 , n14527 , 
 n181889 , n14529 , n181891 , n14531 , n181893 , n14533 , n181895 , n14535 , n14536 , n14537 , 
 n14538 , n181900 , n181901 , n181902 , n14542 , n181904 , n181905 , n14545 , n181907 , n181908 , 
 n14548 , n181910 , n181911 , n14551 , n181913 , n181914 , n181915 , n14555 , n181917 , n14557 , 
 n14558 , n181920 , n181921 , n181922 , n14562 , n181924 , n181925 , n14565 , n181927 , n181928 , 
 n14568 , n181930 , n181931 , n181932 , n14572 , n181934 , n14574 , n14575 , n181937 , n181938 , 
 n181939 , n14579 , n181941 , n181942 , n14582 , n181944 , n181945 , n14585 , n181947 , n181948 , 
 n14588 , n181950 , n14590 , n181952 , n14592 , n14593 , n181955 , n181956 , n181957 , n14597 , 
 n181959 , n181960 , n14600 , n181962 , n181963 , n14603 , n181965 , n181966 , n14606 , n181968 , 
 n181969 , n14612 , n181971 , n181972 , n14615 , n14616 , n14617 , n14618 , n14619 , n181978 , 
 n181979 , n14622 , n181981 , n181982 , n14625 , n181984 , n181985 , n14628 , n181987 , n14630 , 
 n181989 , n14632 , n181991 , n181992 , n14635 , n14636 , n181995 , n14638 , n181997 , n181998 , 
 n14641 , n182000 , n14643 , n14644 , n182003 , n14646 , n182005 , n182006 , n14649 , n182008 , 
 n182009 , n14652 , n14653 , n14654 , n14655 , n182014 , n14657 , n182016 , n14659 , n14660 , 
 n182019 , n14662 , n182021 , n14664 , n14665 , n182024 , n182025 , n14668 , n182027 , n182028 , 
 n182029 , n14672 , n182031 , n14674 , n14675 , n182034 , n182035 , n182036 , n14679 , n182038 , 
 n182039 , n14682 , n182041 , n182042 , n14685 , n182044 , n182045 , n14688 , n182047 , n14690 , 
 n182049 , n14692 , n14693 , n182052 , n182053 , n14696 , n182055 , n182056 , n14699 , n182058 , 
 n182059 , n14702 , n182061 , n182062 , n14705 , n182064 , n14707 , n14708 , n14709 , n14710 , 
 n14711 , n14712 , n14713 , n14714 , n182073 , n182074 , n182075 , n14718 , n182077 , n182078 , 
 n14721 , n182080 , n14723 , n182082 , n14725 , n182084 , n14727 , n14728 , n182087 , n182088 , 
 n182089 , n14732 , n182091 , n182092 , n14735 , n182094 , n182095 , n14738 , n182097 , n14740 , 
 n182099 , n14742 , n182101 , n14744 , n14745 , n182104 , n182105 , n182106 , n14749 , n182108 , 
 n182109 , n14752 , n182111 , n182112 , n14755 , n182114 , n14757 , n14758 , n14759 , n14760 , 
 n182119 , n14762 , n14763 , n182122 , n14765 , n14766 , n182125 , n182126 , n14769 , n14770 , 
 n182129 , n182130 , n14773 , n14774 , n182133 , n182134 , n14777 , n14778 , n182137 , n182138 , 
 n14781 , n14782 , n14783 , n14784 , n182143 , n182144 , n14787 , n14788 , n14789 , n14790 , 
 n14791 , n182150 , n182151 , n182152 , n182153 , n14796 , n182155 , n182156 , n14799 , n182158 , 
 n14801 , n14802 , n182161 , n182162 , n14805 , n182164 , n182165 , n14808 , n182167 , n182168 , 
 n14811 , n182170 , n182171 , n14814 , n182173 , n14816 , n14817 , n182176 , n182177 , n14820 , 
 n182179 , n14822 , n182181 , n182182 , n14825 , n182184 , n14827 , n14828 , n182187 , n182188 , 
 n14831 , n182190 , n14833 , n182192 , n182193 , n14836 , n182195 , n182196 , n14839 , n14840 , 
 n14841 , n14842 , n14843 , n182202 , n182203 , n14846 , n182205 , n182206 , n14849 , n14850 , 
 n182209 , n14852 , n182211 , n14854 , n14855 , n182214 , n182215 , n14858 , n182217 , n14860 , 
 n14861 , n182220 , n14863 , n182222 , n182223 , n14866 , n182225 , n14868 , n182227 , n14870 , 
 n14871 , n182230 , n14873 , n182232 , n182233 , n182234 , n182235 , n14878 , n182237 , n182238 , 
 n14881 , n182240 , n182241 , n14884 , n182243 , n182244 , n14887 , n182246 , n182247 , n14890 , 
 n14891 , n14892 , n182251 , n182252 , n14895 , n182254 , n182255 , n14898 , n182257 , n14900 , 
 n182259 , n14902 , n14903 , n182262 , n182263 , n182264 , n14907 , n182266 , n182267 , n182268 , 
 n182269 , n182270 , n14916 , n182272 , n182273 , n182274 , n14920 , n182276 , n14922 , n14923 , 
 n182279 , n182280 , n182281 , n14927 , n182283 , n182284 , n14930 , n182286 , n182287 , n14933 , 
 n182289 , n182290 , n14936 , n182292 , n14938 , n182294 , n14940 , n182296 , n182297 , n14943 , 
 n14944 , n182300 , n14946 , n182302 , n182303 , n14949 , n182305 , n182306 , n14952 , n14953 , 
 n14954 , n14955 , n182311 , n182312 , n14958 , n14959 , n14960 , n14961 , n182317 , n182318 , 
 n182319 , n14965 , n182321 , n182322 , n14968 , n182324 , n14970 , n14971 , n14972 , n14973 , 
 n182329 , n182330 , n182331 , n14977 , n182333 , n182334 , n14980 , n182336 , n14982 , n14983 , 
 n14984 , n14985 , n14986 , n182342 , n182343 , n182344 , n14990 , n182346 , n182347 , n14993 , 
 n182349 , n14995 , n14996 , n182352 , n14998 , n182354 , n182355 , n15001 , n182357 , n15003 , 
 n15004 , n182360 , n182361 , n182362 , n15008 , n182364 , n182365 , n15011 , n182367 , n182368 , 
 n15014 , n182370 , n182371 , n182372 , n182373 , n15019 , n182375 , n182376 , n15022 , n15023 , 
 n182379 , n182380 , n15026 , n182382 , n182383 , n15029 , n15030 , n182386 , n182387 , n182388 , 
 n15034 , n182390 , n15036 , n15037 , n182393 , n182394 , n182395 , n15041 , n182397 , n182398 , 
 n15044 , n182400 , n182401 , n15047 , n182403 , n182404 , n15050 , n182406 , n182407 , n15053 , 
 n15054 , n182410 , n15056 , n15057 , n182413 , n182414 , n15060 , n15061 , n15062 , n15063 , 
 n15064 , n182420 , n182421 , n15067 , n15068 , n182424 , n182425 , n15071 , n15072 , n182428 , 
 n182429 , n182430 , n15076 , n182432 , n15078 , n15079 , n182435 , n15081 , n182437 , n15083 , 
 n182439 , n182440 , n15086 , n182442 , n182443 , n15089 , n182445 , n15091 , n15092 , n182448 , 
 n182449 , n182450 , n15096 , n182452 , n182453 , n15099 , n182455 , n182456 , n15102 , n182458 , 
 n15104 , n182460 , n15106 , n182462 , n15108 , n15109 , n182465 , n182466 , n182467 , n15113 , 
 n182469 , n182470 , n15116 , n182472 , n182473 , n15119 , n182475 , n15121 , n182477 , n15123 , 
 n182479 , n182480 , n15126 , n15127 , n182483 , n15129 , n15130 , n182486 , n15132 , n15133 , 
 n15134 , n15135 , n15136 , n182492 , n182493 , n15139 , n182495 , n15141 , n15142 , n15143 , 
 n15144 , n182500 , n15146 , n15147 , n15148 , n15149 , n182505 , n182506 , n15152 , n15153 , 
 n15154 , n15155 , n15156 , n182512 , n182513 , n15159 , n15160 , n15161 , n15162 , n182518 , 
 n182519 , n182520 , n15166 , n15167 , n15168 , n15169 , n182525 , n182526 , n15172 , n15173 , 
 n15174 , n182530 , n182531 , n182532 , n15178 , n182534 , n182535 , n15181 , n182537 , n182538 , 
 n15184 , n182540 , n182541 , n15187 , n15188 , n15189 , n15190 , n15191 , n182547 , n182548 , 
 n15194 , n182550 , n15196 , n182552 , n182553 , n15199 , n182555 , n182556 , n15202 , n182558 , 
 n182559 , n15208 , n15209 , n15210 , n182563 , n182564 , n15213 , n182566 , n182567 , n15216 , 
 n182569 , n182570 , n15219 , n182572 , n182573 , n15222 , n182575 , n182576 , n15225 , n182578 , 
 n182579 , n15228 , n182581 , n182582 , n15231 , n15232 , n182585 , n182586 , n15235 , n15236 , 
 n182589 , n182590 , n15239 , n15240 , n15241 , n182594 , n182595 , n15244 , n15245 , n15246 , 
 n15247 , n182600 , n182601 , n15250 , n182603 , n182604 , n15253 , n182606 , n182607 , n15256 , 
 n182609 , n182610 , n182611 , n182612 , n15261 , n182614 , n182615 , n182616 , n182617 , n15266 , 
 n15267 , n182620 , n15269 , n182622 , n182623 , n15272 , n15273 , n182626 , n182627 , n15276 , 
 n182629 , n182630 , n15279 , n182632 , n182633 , n15282 , n182635 , n182636 , n15285 , n15286 , 
 n15287 , n15288 , n15289 , n182642 , n182643 , n182644 , n15293 , n182646 , n182647 , n15296 , 
 n182649 , n15298 , n182651 , n182652 , n182653 , n182654 , n15303 , n182656 , n182657 , n15306 , 
 n182659 , n182660 , n15309 , n15310 , n15311 , n15312 , n182665 , n182666 , n15315 , n182668 , 
 n182669 , n15318 , n182671 , n182672 , n182673 , n15322 , n182675 , n15324 , n15325 , n182678 , 
 n182679 , n182680 , n15329 , n182682 , n182683 , n15332 , n182685 , n182686 , n15335 , n182688 , 
 n182689 , n15338 , n182691 , n15340 , n182693 , n15342 , n15343 , n182696 , n182697 , n182698 , 
 n182699 , n182700 , n182701 , n15350 , n182703 , n182704 , n15353 , n182706 , n182707 , n15356 , 
 n182709 , n182710 , n15359 , n182712 , n15361 , n15362 , n182715 , n182716 , n182717 , n15366 , 
 n182719 , n182720 , n15369 , n182722 , n182723 , n15372 , n182725 , n182726 , n182727 , n15376 , 
 n182729 , n15378 , n15379 , n182732 , n182733 , n182734 , n15383 , n182736 , n182737 , n15386 , 
 n182739 , n182740 , n15389 , n182742 , n182743 , n15392 , n182745 , n15394 , n182747 , n15396 , 
 n15397 , n182750 , n182751 , n182752 , n15401 , n182754 , n182755 , n15404 , n182757 , n182758 , 
 n15407 , n182760 , n182761 , n15410 , n182763 , n15412 , n182765 , n15414 , n182767 , n15416 , 
 n15417 , n182770 , n182771 , n182772 , n15421 , n182774 , n182775 , n15424 , n182777 , n182778 , 
 n15427 , n182780 , n182781 , n182782 , n15431 , n182784 , n15433 , n15434 , n182787 , n182788 , 
 n182789 , n15438 , n182791 , n182792 , n15441 , n182794 , n182795 , n15444 , n182797 , n182798 , 
 n15447 , n182800 , n15449 , n182802 , n15451 , n15452 , n182805 , n182806 , n15455 , n182808 , 
 n182809 , n15458 , n182811 , n182812 , n15461 , n182814 , n15463 , n182816 , n15465 , n182818 , 
 n182819 , n15468 , n15469 , n15470 , n15471 , n182824 , n182825 , n15474 , n182827 , n15476 , 
 n182829 , n15478 , n15479 , n182832 , n15481 , n182834 , n15483 , n182836 , n182837 , n182838 , 
 n182839 , n15491 , n15492 , n15493 , n182843 , n182844 , n182845 , n15497 , n182847 , n182848 , 
 n15500 , n182850 , n15502 , n15503 , n182853 , n15505 , n182855 , n15507 , n15508 , n182858 , 
 n182859 , n15511 , n182861 , n15513 , n182863 , n182864 , n15516 , n182866 , n15518 , n182868 , 
 n15520 , n15521 , n15522 , n15523 , n182873 , n182874 , n15526 , n15527 , n15528 , n182878 , 
 n182879 , n182880 , n15532 , n182882 , n182883 , n15535 , n182885 , n182886 , n182887 , n182888 , 
 n15540 , n182890 , n15542 , n182892 , n182893 , n182894 , n182895 , n15547 , n182897 , n182898 , 
 n15550 , n182900 , n182901 , n15553 , n15554 , n15555 , n15556 , n15557 , n182907 , n182908 , 
 n15560 , n182910 , n182911 , n15563 , n182913 , n182914 , n15566 , n15567 , n15568 , n15569 , 
 n182919 , n182920 , n15572 , n182922 , n15574 , n182924 , n15576 , n15577 , n182927 , n182928 , 
 n15580 , n182930 , n15582 , n182932 , n182933 , n15585 , n182935 , n182936 , n15588 , n182938 , 
 n182939 , n15591 , n182941 , n182942 , n15594 , n182944 , n15596 , n182946 , n15598 , n182948 , 
 n15600 , n182950 , n182951 , n15603 , n182953 , n15605 , n15606 , n15607 , n15608 , n15609 , 
 n15610 , n182960 , n182961 , n15613 , n15614 , n15615 , n15616 , n15617 , n182967 , n182968 , 
 n15620 , n15621 , n15622 , n15623 , n182973 , n182974 , n15626 , n15627 , n15628 , n15629 , 
 n15630 , n182980 , n182981 , n15633 , n15634 , n15635 , n182985 , n182986 , n182987 , n15639 , 
 n182989 , n182990 , n15642 , n182992 , n15644 , n15645 , n15646 , n15647 , n15648 , n182998 , 
 n182999 , n183000 , n15652 , n183002 , n183003 , n15655 , n183005 , n15657 , n15658 , n183008 , 
 n183009 , n15661 , n183011 , n15663 , n183013 , n183014 , n15666 , n183016 , n15668 , n15669 , 
 n183019 , n15671 , n183021 , n15673 , n183023 , n183024 , n15676 , n183026 , n183027 , n15679 , 
 n15680 , n15681 , n15682 , n15683 , n183033 , n183034 , n15686 , n183036 , n183037 , n15689 , 
 n15690 , n15691 , n15692 , n183042 , n183043 , n15695 , n183045 , n15697 , n183047 , n15699 , 
 n183049 , n15701 , n15702 , n15703 , n15704 , n183054 , n183055 , n15707 , n15708 , n15709 , 
 n15710 , n183060 , n183061 , n15713 , n15714 , n15715 , n15716 , n15717 , n183067 , n183068 , 
 n15720 , n183070 , n183071 , n15723 , n183073 , n183074 , n15726 , n183076 , n183077 , n183078 , 
 n15730 , n183080 , n15732 , n15733 , n183083 , n183084 , n183085 , n15737 , n183087 , n183088 , 
 n15740 , n183090 , n183091 , n15743 , n183093 , n183094 , n15746 , n183096 , n15748 , n183098 , 
 n15750 , n183100 , n183101 , n15753 , n15754 , n183104 , n183105 , n183106 , n15758 , n183108 , 
 n183109 , n15764 , n183111 , n183112 , n15767 , n183114 , n183115 , n15770 , n183117 , n183118 , 
 n15773 , n15774 , n15775 , n183122 , n183123 , n183124 , n15779 , n183126 , n183127 , n15782 , 
 n183129 , n15784 , n183131 , n15786 , n183133 , n183134 , n15789 , n183136 , n15791 , n15792 , 
 n183139 , n15794 , n183141 , n15796 , n183143 , n15798 , n183145 , n15800 , n15801 , n183148 , 
 n183149 , n183150 , n15805 , n183152 , n183153 , n15808 , n183155 , n183156 , n15811 , n183158 , 
 n15813 , n183160 , n15815 , n183162 , n15817 , n183164 , n15819 , n15820 , n183167 , n183168 , 
 n183169 , n15824 , n183171 , n183172 , n15827 , n183174 , n183175 , n15830 , n183177 , n183178 , 
 n183179 , n15834 , n183181 , n15836 , n183183 , n183184 , n15839 , n15840 , n183187 , n183188 , 
 n183189 , n15844 , n183191 , n183192 , n15847 , n183194 , n183195 , n15850 , n183197 , n183198 , 
 n15853 , n183200 , n15855 , n183202 , n15857 , n15858 , n183205 , n183206 , n183207 , n15862 , 
 n183209 , n183210 , n15865 , n183212 , n183213 , n15868 , n183215 , n183216 , n15871 , n183218 , 
 n183219 , n15874 , n183221 , n183222 , n15877 , n183224 , n183225 , n15880 , n183227 , n183228 , 
 n15883 , n183230 , n183231 , n15886 , n183233 , n183234 , n15889 , n15890 , n183237 , n183238 , 
 n183239 , n183240 , n183241 , n15896 , n183243 , n183244 , n15899 , n183246 , n15901 , n183248 , 
 n183249 , n15904 , n183251 , n15906 , n15907 , n15908 , n15909 , n183256 , n183257 , n15912 , 
 n183259 , n15914 , n183261 , n15916 , n15917 , n15918 , n15919 , n183266 , n15921 , n15922 , 
 n15923 , n15924 , n183271 , n183272 , n183273 , n15928 , n183275 , n15930 , n15931 , n183278 , 
 n183279 , n183280 , n15935 , n183282 , n183283 , n15938 , n183285 , n183286 , n15941 , n183288 , 
 n183289 , n183290 , n15945 , n183292 , n15947 , n15948 , n183295 , n183296 , n183297 , n15952 , 
 n183299 , n183300 , n15955 , n183302 , n183303 , n15958 , n183305 , n183306 , n15961 , n183308 , 
 n15963 , n183310 , n183311 , n183312 , n15967 , n183314 , n183315 , n15970 , n183317 , n15972 , 
 n183319 , n183320 , n183321 , n183322 , n15977 , n183324 , n183325 , n15980 , n183327 , n183328 , 
 n15983 , n15984 , n183331 , n183332 , n15987 , n183334 , n183335 , n15990 , n183337 , n183338 , 
 n15993 , n183340 , n183341 , n183342 , n15997 , n183344 , n15999 , n16000 , n183347 , n183348 , 
 n183349 , n16004 , n183351 , n183352 , n16007 , n183354 , n183355 , n16010 , n183357 , n183358 , 
 n16013 , n183360 , n16015 , n183362 , n16017 , n16018 , n183365 , n183366 , n183367 , n183368 , 
 n183369 , n183370 , n16028 , n183372 , n183373 , n16031 , n183375 , n183376 , n16034 , n183378 , 
 n183379 , n16037 , n183381 , n183382 , n16040 , n183384 , n16042 , n16043 , n183387 , n183388 , 
 n16046 , n183390 , n183391 , n16049 , n183393 , n183394 , n16052 , n183396 , n16054 , n16055 , 
 n183399 , n183400 , n16058 , n183402 , n16060 , n183404 , n183405 , n16063 , n183407 , n16065 , 
 n16066 , n16067 , n16068 , n16069 , n183413 , n16071 , n183415 , n16073 , n16074 , n16075 , 
 n16076 , n16077 , n183421 , n183422 , n16080 , n16081 , n183425 , n183426 , n16084 , n16085 , 
 n183429 , n16087 , n183431 , n16089 , n16090 , n16091 , n16092 , n183436 , n183437 , n16095 , 
 n183439 , n16097 , n16098 , n183442 , n183443 , n183444 , n16102 , n183446 , n183447 , n16105 , 
 n183449 , n183450 , n16108 , n183452 , n183453 , n183454 , n16112 , n183456 , n16114 , n16115 , 
 n183459 , n183460 , n183461 , n16119 , n183463 , n183464 , n16122 , n183466 , n183467 , n16125 , 
 n183469 , n183470 , n16128 , n183472 , n16130 , n183474 , n16132 , n16133 , n183477 , n183478 , 
 n183479 , n16137 , n183481 , n183482 , n16140 , n183484 , n183485 , n16143 , n183487 , n183488 , 
 n16146 , n183490 , n183491 , n16149 , n16150 , n183494 , n16152 , n16153 , n183497 , n183498 , 
 n16156 , n183500 , n183501 , n16159 , n16160 , n16161 , n16162 , n183506 , n183507 , n16165 , 
 n16166 , n16167 , n16168 , n16169 , n183513 , n183514 , n16172 , n183516 , n183517 , n16175 , 
 n16176 , n16177 , n16178 , n16179 , n183523 , n183524 , n16182 , n183526 , n16184 , n183528 , 
 n16186 , n183530 , n183531 , n16189 , n183533 , n183534 , n16192 , n183536 , n183537 , n16195 , 
 n183539 , n183540 , n16198 , n183542 , n183543 , n16201 , n183545 , n16203 , n16204 , n183548 , 
 n16206 , n183550 , n183551 , n16209 , n183553 , n183554 , n16212 , n183556 , n16214 , n16215 , 
 n16216 , n183560 , n16218 , n183562 , n16220 , n16221 , n183565 , n16223 , n183567 , n16225 , 
 n16226 , n183570 , n16228 , n183572 , n16230 , n183574 , n183575 , n183576 , n16234 , n183578 , 
 n183579 , n16237 , n183581 , n183582 , n16240 , n16241 , n183585 , n183586 , n16244 , n183588 , 
 n183589 , n16247 , n183591 , n183592 , n183593 , n16251 , n183595 , n16253 , n16254 , n183598 , 
 n16256 , n183600 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , 
 n16266 , n16267 , n16268 , n16269 , n183613 , n183614 , n16272 , n183616 , n183617 , n16275 , 
 n183619 , n16280 , n16281 , n16282 , n16283 , n183624 , n16285 , n16286 , n183627 , n16288 , 
 n183629 , n183630 , n183631 , n16292 , n183633 , n183634 , n16295 , n183636 , n16297 , n16298 , 
 n16299 , n16300 , n16301 , n16302 , n16303 , n183644 , n183645 , n183646 , n16307 , n183648 , 
 n183649 , n16310 , n183651 , n183652 , n183653 , n16314 , n183655 , n183656 , n183657 , n16318 , 
 n183659 , n183660 , n16321 , n183662 , n183663 , n16324 , n183665 , n16326 , n16327 , n16328 , 
 n16329 , n183670 , n16331 , n183672 , n183673 , n16334 , n183675 , n183676 , n16337 , n183678 , 
 n16339 , n183680 , n16341 , n183682 , n183683 , n16344 , n183685 , n183686 , n16347 , n183688 , 
 n183689 , n16350 , n183691 , n183692 , n16353 , n16354 , n183695 , n183696 , n16357 , n183698 , 
 n183699 , n16360 , n183701 , n183702 , n16363 , n183704 , n183705 , n16366 , n16367 , n183708 , 
 n183709 , n16370 , n183711 , n183712 , n16373 , n183714 , n16375 , n183716 , n16377 , n183718 , 
 n183719 , n16380 , n183721 , n183722 , n16383 , n183724 , n183725 , n183726 , n183727 , n16388 , 
 n183729 , n183730 , n16391 , n183732 , n16393 , n183734 , n16395 , n16396 , n183737 , n183738 , 
 n183739 , n183740 , n183741 , n16402 , n183743 , n16404 , n16405 , n183746 , n16407 , n16408 , 
 n16409 , n16410 , n183751 , n183752 , n16413 , n16414 , n16415 , n16416 , n16417 , n183758 , 
 n183759 , n16420 , n16421 , n16422 , n16423 , n183764 , n183765 , n16426 , n183767 , n183768 , 
 n16429 , n183770 , n183771 , n183772 , n16433 , n183774 , n16435 , n16436 , n183777 , n183778 , 
 n183779 , n16440 , n183781 , n183782 , n16443 , n183784 , n183785 , n16446 , n183787 , n183788 , 
 n16449 , n183790 , n16451 , n183792 , n16453 , n16454 , n16455 , n183796 , n183797 , n183798 , 
 n16459 , n183800 , n183801 , n16462 , n183803 , n183804 , n16465 , n183806 , n183807 , n16468 , 
 n183809 , n183810 , n16471 , n183812 , n183813 , n16474 , n183815 , n183816 , n183817 , n16478 , 
 n183819 , n16480 , n16481 , n183822 , n183823 , n183824 , n16485 , n183826 , n183827 , n16488 , 
 n183829 , n183830 , n16491 , n183832 , n183833 , n183834 , n16495 , n183836 , n16497 , n16498 , 
 n183839 , n183840 , n183841 , n16502 , n183843 , n183844 , n16505 , n183846 , n183847 , n16508 , 
 n183849 , n183850 , n16511 , n183852 , n16513 , n183854 , n16515 , n16516 , n183857 , n183858 , 
 n183859 , n16523 , n183861 , n183862 , n16526 , n183864 , n183865 , n16529 , n183867 , n183868 , 
 n16532 , n183870 , n183871 , n183872 , n16536 , n183874 , n16538 , n16539 , n183877 , n183878 , 
 n183879 , n16543 , n183881 , n183882 , n16546 , n183884 , n183885 , n16549 , n183887 , n183888 , 
 n183889 , n183890 , n16554 , n183892 , n16556 , n183894 , n183895 , n16559 , n183897 , n16561 , 
 n183899 , n16563 , n16564 , n183902 , n16566 , n183904 , n183905 , n183906 , n183907 , n16571 , 
 n183909 , n183910 , n16574 , n183912 , n183913 , n16577 , n183915 , n183916 , n16580 , n183918 , 
 n183919 , n16583 , n183921 , n183922 , n16586 , n183924 , n16588 , n16589 , n183927 , n183928 , 
 n183929 , n16593 , n183931 , n183932 , n16596 , n183934 , n183935 , n16599 , n183937 , n183938 , 
 n16602 , n16603 , n16604 , n16605 , n16606 , n183944 , n183945 , n16609 , n183947 , n183948 , 
 n16612 , n183950 , n183951 , n16615 , n16616 , n16617 , n16618 , n183956 , n183957 , n16621 , 
 n183959 , n183960 , n16624 , n183962 , n183963 , n16627 , n183965 , n16629 , n183967 , n183968 , 
 n183969 , n183970 , n16634 , n183972 , n183973 , n183974 , n183975 , n183976 , n16640 , n183978 , 
 n183979 , n16643 , n16644 , n16645 , n16646 , n16647 , n183985 , n183986 , n16650 , n183988 , 
 n183989 , n16653 , n16654 , n16655 , n16656 , n183994 , n183995 , n16659 , n183997 , n183998 , 
 n16662 , n184000 , n184001 , n16665 , n184003 , n184004 , n16668 , n184006 , n184007 , n16671 , 
 n184009 , n184010 , n16674 , n16675 , n184013 , n16677 , n184015 , n184016 , n16680 , n16681 , 
 n184019 , n16683 , n184021 , n16685 , n184023 , n184024 , n184025 , n16689 , n16690 , n16691 , 
 n184029 , n16693 , n184031 , n184032 , n16696 , n184034 , n184035 , n16699 , n184037 , n16701 , 
 n16702 , n184040 , n16704 , n184042 , n184043 , n16707 , n16708 , n16709 , n184047 , n16711 , 
 n16712 , n184050 , n16714 , n184052 , n16716 , n16717 , n16718 , n184056 , n16720 , n184058 , 
 n184059 , n16723 , n184061 , n184062 , n16726 , n184064 , n184065 , n16729 , n184067 , n184068 , 
 n16732 , n184070 , n184071 , n16735 , n184073 , n184074 , n16738 , n184076 , n184077 , n16741 , 
 n16742 , n184080 , n16744 , n184082 , n184083 , n16747 , n16748 , n184086 , n16750 , n184088 , 
 n184089 , n16756 , n184091 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n184099 , n16766 , n184101 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n184110 , n16777 , n184112 , n16779 , n16780 , n184115 , n16782 , n184117 , n184118 , 
 n16785 , n184120 , n16787 , n16788 , n16789 , n184124 , n184125 , n16792 , n184127 , n16794 , 
 n184129 , n16796 , n184131 , n184132 , n16799 , n184134 , n184135 , n16802 , n184137 , n16804 , 
 n16805 , n16806 , n184141 , n16808 , n184143 , n184144 , n184145 , n184146 , n16813 , n184148 , 
 n184149 , n16816 , n184151 , n16818 , n16819 , n184154 , n184155 , n184156 , n16823 , n184158 , 
 n184159 , n16826 , n184161 , n184162 , n16829 , n184164 , n184165 , n184166 , n184167 , n16834 , 
 n184169 , n184170 , n16837 , n184172 , n184173 , n184174 , n184175 , n16842 , n184177 , n184178 , 
 n16845 , n184180 , n16847 , n16848 , n184183 , n16850 , n184185 , n16852 , n184187 , n184188 , 
 n16855 , n184190 , n184191 , n16858 , n184193 , n184194 , n184195 , n184196 , n16863 , n184198 , 
 n184199 , n16866 , n184201 , n16868 , n16869 , n184204 , n184205 , n16872 , n184207 , n184208 , 
 n16875 , n184210 , n184211 , n16878 , n184213 , n184214 , n16881 , n184216 , n184217 , n16884 , 
 n184219 , n16886 , n16887 , n184222 , n184223 , n184224 , n16891 , n184226 , n184227 , n16894 , 
 n184229 , n184230 , n16897 , n184232 , n184233 , n16900 , n184235 , n16902 , n184237 , n184238 , 
 n184239 , n16906 , n184241 , n184242 , n16909 , n184244 , n16911 , n184246 , n184247 , n16914 , 
 n184249 , n184250 , n16917 , n184252 , n184253 , n184254 , n16921 , n184256 , n184257 , n16924 , 
 n184259 , n16926 , n184261 , n16928 , n16929 , n184264 , n184265 , n16932 , n16933 , n184268 , 
 n184269 , n16936 , n184271 , n184272 , n16939 , n184274 , n16941 , n16942 , n184277 , n184278 , 
 n16945 , n184280 , n184281 , n16948 , n184283 , n184284 , n16951 , n184286 , n184287 , n184288 , 
 n16955 , n184290 , n16957 , n184292 , n184293 , n16960 , n184295 , n184296 , n16963 , n184298 , 
 n184299 , n16966 , n16967 , n16968 , n184303 , n184304 , n16971 , n184306 , n184307 , n184308 , 
 n184309 , n184310 , n16980 , n184312 , n16982 , n16983 , n184315 , n16985 , n184317 , n16987 , 
 n184319 , n184320 , n16990 , n184322 , n184323 , n16993 , n184325 , n16995 , n16996 , n184328 , 
 n184329 , n184330 , n17000 , n184332 , n184333 , n17003 , n184335 , n184336 , n17006 , n184338 , 
 n17008 , n184340 , n184341 , n17011 , n17012 , n184344 , n17014 , n17015 , n184347 , n184348 , 
 n17018 , n184350 , n184351 , n184352 , n17022 , n184354 , n17024 , n17025 , n184357 , n184358 , 
 n17028 , n184360 , n184361 , n17031 , n184363 , n184364 , n184365 , n17035 , n184367 , n184368 , 
 n17038 , n184370 , n17040 , n17041 , n184373 , n184374 , n17044 , n184376 , n184377 , n17047 , 
 n184379 , n17049 , n17050 , n184382 , n184383 , n17053 , n184385 , n184386 , n17056 , n184388 , 
 n17058 , n17059 , n184391 , n184392 , n17062 , n184394 , n184395 , n17065 , n184397 , n17067 , 
 n17068 , n17069 , n17070 , n184402 , n184403 , n17073 , n184405 , n184406 , n17076 , n184408 , 
 n17078 , n17079 , n184411 , n184412 , n17082 , n184414 , n184415 , n17085 , n184417 , n184418 , 
 n184419 , n184420 , n17090 , n184422 , n184423 , n17093 , n184425 , n17095 , n17096 , n184428 , 
 n184429 , n17099 , n184431 , n184432 , n17102 , n184434 , n184435 , n17105 , n17106 , n184438 , 
 n17108 , n184440 , n17110 , n17111 , n184443 , n184444 , n184445 , n17115 , n184447 , n184448 , 
 n17118 , n184450 , n184451 , n17121 , n184453 , n184454 , n17124 , n17125 , n17126 , n184458 , 
 n17128 , n17129 , n184461 , n184462 , n17132 , n184464 , n184465 , n184466 , n184467 , n17137 , 
 n184469 , n184470 , n17140 , n184472 , n17142 , n17143 , n184475 , n184476 , n17146 , n184478 , 
 n184479 , n17149 , n184481 , n184482 , n17152 , n17153 , n184485 , n17155 , n184487 , n17157 , 
 n17158 , n184490 , n184491 , n184492 , n17162 , n184494 , n184495 , n17165 , n184497 , n184498 , 
 n17168 , n184500 , n184501 , n17171 , n17172 , n17173 , n184505 , n17175 , n17176 , n17177 , 
 n17178 , n17179 , n17180 , n17181 , n184513 , n17183 , n17184 , n17185 , n17186 , n17187 , 
 n184519 , n17192 , n184521 , n184522 , n17195 , n184524 , n184525 , n184526 , n17199 , n184528 , 
 n17201 , n17202 , n184531 , n184532 , n184533 , n17206 , n184535 , n184536 , n17209 , n184538 , 
 n184539 , n17212 , n184541 , n184542 , n17215 , n184544 , n17217 , n184546 , n17219 , n17220 , 
 n184549 , n184550 , n184551 , n17224 , n184553 , n184554 , n17227 , n184556 , n184557 , n17230 , 
 n184559 , n184560 , n17233 , n17234 , n17235 , n184564 , n17237 , n17238 , n17239 , n17240 , 
 n17241 , n17242 , n184571 , n184572 , n17245 , n184574 , n17247 , n17248 , n184577 , n184578 , 
 n184579 , n17252 , n184581 , n184582 , n17255 , n184584 , n184585 , n17258 , n184587 , n184588 , 
 n17261 , n184590 , n17263 , n184592 , n17265 , n17266 , n184595 , n17268 , n184597 , n17270 , 
 n184599 , n184600 , n17273 , n184602 , n184603 , n17276 , n184605 , n17278 , n184607 , n17280 , 
 n17281 , n17282 , n184611 , n184612 , n17285 , n17286 , n184615 , n184616 , n17289 , n184618 , 
 n184619 , n184620 , n17293 , n17294 , n184623 , n17296 , n184625 , n17298 , n184627 , n184628 , 
 n17301 , n184630 , n184631 , n184632 , n17305 , n184634 , n17307 , n17308 , n184637 , n184638 , 
 n17311 , n184640 , n184641 , n17314 , n184643 , n184644 , n17317 , n17318 , n17319 , n17320 , 
 n17321 , n17322 , n184651 , n17324 , n17325 , n184654 , n184655 , n17328 , n184657 , n17330 , 
 n184659 , n17332 , n17333 , n184662 , n184663 , n17336 , n184665 , n184666 , n17339 , n184668 , 
 n184669 , n17342 , n184671 , n184672 , n17345 , n184674 , n184675 , n17348 , n184677 , n184678 , 
 n17351 , n184680 , n184681 , n184682 , n17355 , n184684 , n17357 , n17358 , n184687 , n184688 , 
 n17361 , n184690 , n184691 , n17364 , n184693 , n184694 , n17367 , n184696 , n17369 , n184698 , 
 n17371 , n17372 , n184701 , n184702 , n17375 , n184704 , n184705 , n17378 , n184707 , n184708 , 
 n17381 , n17382 , n17383 , n184712 , n184713 , n17386 , n17387 , n17388 , n184717 , n184718 , 
 n17394 , n17395 , n17396 , n184722 , n184723 , n17399 , n184725 , n184726 , n17402 , n17403 , 
 n17404 , n184730 , n184731 , n17407 , n17408 , n184734 , n184735 , n17411 , n17412 , n184738 , 
 n184739 , n17415 , n17416 , n184742 , n17418 , n17419 , n184745 , n184746 , n17422 , n17423 , 
 n17424 , n184750 , n184751 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , 
 n184759 , n17435 , n17436 , n17437 , n184763 , n184764 , n17440 , n17441 , n17442 , n184768 , 
 n184769 , n17445 , n184771 , n184772 , n184773 , n17449 , n184775 , n17451 , n17452 , n184778 , 
 n184779 , n17455 , n184781 , n184782 , n17458 , n184784 , n184785 , n184786 , n17462 , n184788 , 
 n17464 , n17465 , n184791 , n184792 , n17468 , n184794 , n184795 , n17471 , n184797 , n184798 , 
 n17474 , n184800 , n17476 , n184802 , n184803 , n17479 , n17480 , n17481 , n184807 , n184808 , 
 n17484 , n17485 , n184811 , n184812 , n17488 , n184814 , n17490 , n17491 , n17492 , n184818 , 
 n184819 , n17495 , n17496 , n17497 , n17498 , n184824 , n184825 , n17501 , n17502 , n17503 , 
 n17504 , n17505 , n184831 , n184832 , n17508 , n17509 , n17510 , n184836 , n184837 , n17513 , 
 n17514 , n17515 , n184841 , n184842 , n17518 , n17519 , n184845 , n184846 , n17522 , n17523 , 
 n17524 , n184850 , n184851 , n17527 , n17528 , n184854 , n17530 , n17531 , n17532 , n184858 , 
 n184859 , n17535 , n17536 , n17537 , n184863 , n184864 , n17540 , n17541 , n184867 , n184868 , 
 n17544 , n17545 , n17546 , n17547 , n17548 , n184874 , n184875 , n17551 , n17552 , n17553 , 
 n17554 , n184880 , n184881 , n17557 , n17558 , n17559 , n184885 , n184886 , n17562 , n17563 , 
 n17564 , n184890 , n184891 , n17567 , n17568 , n17569 , n184895 , n184896 , n17572 , n17573 , 
 n17574 , n184900 , n184901 , n17577 , n184903 , n184904 , n17580 , n184906 , n184907 , n17583 , 
 n184909 , n184910 , n184911 , n17590 , n17591 , n184914 , n184915 , n17594 , n17595 , n17596 , 
 n17597 , n184920 , n184921 , n17600 , n17601 , n184924 , n184925 , n17604 , n17605 , n17606 , 
 n17607 , n17608 , n184931 , n184932 , n17611 , n17612 , n17613 , n184936 , n184937 , n17616 , 
 n17617 , n17618 , n184941 , n184942 , n17621 , n17622 , n17623 , n184946 , n184947 , n17626 , 
 n184949 , n184950 , n17629 , n184952 , n184953 , n17632 , n184955 , n184956 , n17635 , n17636 , 
 n184959 , n184960 , n17639 , n17640 , n184963 , n184964 , n17643 , n17644 , n184967 , n184968 , 
 n17647 , n17648 , n17649 , n17650 , n17651 , n184974 , n184975 , n17654 , n17655 , n17656 , 
 n184979 , n184980 , n17659 , n184982 , n184983 , n17662 , n17663 , n184986 , n184987 , n17666 , 
 n184989 , n184990 , n17669 , n184992 , n184993 , n17672 , n184995 , n184996 , n17675 , n17676 , 
 n184999 , n17678 , n185001 , n17680 , n17681 , n185004 , n17683 , n185006 , n17685 , n185008 , 
 n185009 , n17688 , n185011 , n185012 , n185013 , n185014 , n17693 , n185016 , n185017 , n185018 , 
 n17697 , n185020 , n17699 , n185022 , n185023 , n17702 , n17703 , n185026 , n17705 , n185028 , 
 n17707 , n185030 , n185031 , n17710 , n185033 , n185034 , n17713 , n185036 , n185037 , n17716 , 
 n185039 , n185040 , n17719 , n185042 , n185043 , n17722 , n185045 , n185046 , n17725 , n185048 , 
 n185049 , n17728 , n185051 , n185052 , n17731 , n17732 , n17733 , n17734 , n17735 , n185058 , 
 n185059 , n17738 , n17739 , n17740 , n17741 , n185064 , n185065 , n17744 , n17745 , n17746 , 
 n17747 , n185070 , n185071 , n17750 , n185073 , n17752 , n185075 , n17754 , n17755 , n185078 , 
 n185079 , n17758 , n185081 , n185082 , n17761 , n185084 , n185085 , n17764 , n185087 , n185088 , 
 n185089 , n185090 , n17772 , n185092 , n17774 , n185094 , n185095 , n185096 , n185097 , n17779 , 
 n185099 , n185100 , n17782 , n185102 , n185103 , n17785 , n17786 , n17787 , n17788 , n17789 , 
 n185109 , n185110 , n17792 , n185112 , n185113 , n17795 , n17796 , n17797 , n17798 , n17799 , 
 n17800 , n185120 , n17802 , n185122 , n185123 , n17805 , n185125 , n17807 , n185127 , n185128 , 
 n185129 , n185130 , n17812 , n185132 , n185133 , n17815 , n185135 , n185136 , n185137 , n17819 , 
 n185139 , n17821 , n17822 , n185142 , n185143 , n185144 , n17826 , n185146 , n185147 , n17829 , 
 n185149 , n185150 , n17832 , n185152 , n185153 , n185154 , n17836 , n185156 , n17838 , n17839 , 
 n185159 , n17841 , n185161 , n17843 , n185163 , n185164 , n17846 , n185166 , n185167 , n17849 , 
 n185169 , n17851 , n185171 , n17853 , n17854 , n185174 , n185175 , n185176 , n17858 , n185178 , 
 n185179 , n17861 , n185181 , n185182 , n17864 , n185184 , n185185 , n17867 , n185187 , n185188 , 
 n17870 , n17871 , n185191 , n185192 , n17874 , n185194 , n17876 , n17877 , n185197 , n17879 , 
 n185199 , n17881 , n185201 , n185202 , n17884 , n185204 , n17886 , n185206 , n17888 , n185208 , 
 n17890 , n17891 , n185211 , n185212 , n185213 , n17895 , n185215 , n185216 , n17898 , n185218 , 
 n185219 , n17901 , n185221 , n17903 , n185223 , n17905 , n185225 , n185226 , n17908 , n185228 , 
 n185229 , n17911 , n185231 , n185232 , n17914 , n185234 , n185235 , n17917 , n185237 , n185238 , 
 n17920 , n185240 , n185241 , n17923 , n185243 , n17925 , n17926 , n17927 , n17928 , n185248 , 
 n185249 , n17931 , n185251 , n17933 , n17934 , n185254 , n185255 , n185256 , n17938 , n185258 , 
 n185259 , n17944 , n185261 , n185262 , n17947 , n185264 , n185265 , n185266 , n17951 , n185268 , 
 n17953 , n17954 , n185271 , n17956 , n185273 , n185274 , n17959 , n185276 , n17961 , n185278 , 
 n17963 , n17964 , n185281 , n185282 , n185283 , n17968 , n185285 , n185286 , n17971 , n185288 , 
 n185289 , n17974 , n185291 , n185292 , n17977 , n185294 , n185295 , n17980 , n185297 , n17982 , 
 n185299 , n17984 , n17985 , n185302 , n185303 , n185304 , n17989 , n185306 , n185307 , n17992 , 
 n185309 , n185310 , n17995 , n185312 , n185313 , n185314 , n17999 , n185316 , n18001 , n18002 , 
 n185319 , n185320 , n185321 , n18006 , n185323 , n185324 , n18009 , n185326 , n185327 , n18012 , 
 n185329 , n185330 , n18015 , n185332 , n18017 , n185334 , n18019 , n18020 , n185337 , n185338 , 
 n185339 , n18024 , n185341 , n185342 , n18027 , n185344 , n185345 , n18030 , n185347 , n185348 , 
 n18033 , n185350 , n185351 , n18036 , n185353 , n185354 , n18039 , n185356 , n185357 , n185358 , 
 n18043 , n18044 , n18045 , n18046 , n18047 , n185364 , n185365 , n18050 , n185367 , n185368 , 
 n18053 , n18054 , n18055 , n18056 , n185373 , n185374 , n18059 , n18060 , n18061 , n18062 , 
 n18063 , n185380 , n185381 , n18066 , n185383 , n185384 , n18069 , n18070 , n18071 , n18072 , 
 n18073 , n185390 , n185391 , n18076 , n185393 , n185394 , n18079 , n18080 , n18081 , n18082 , 
 n185399 , n185400 , n18085 , n185402 , n18087 , n185404 , n18089 , n185406 , n185407 , n18092 , 
 n185409 , n185410 , n18095 , n185412 , n185413 , n18098 , n185415 , n185416 , n18101 , n185418 , 
 n18106 , n185420 , n185421 , n18109 , n185423 , n185424 , n185425 , n185426 , n185427 , n18115 , 
 n185429 , n185430 , n18118 , n185432 , n185433 , n185434 , n185435 , n18123 , n185437 , n185438 , 
 n18126 , n185440 , n185441 , n18129 , n185443 , n185444 , n18132 , n185446 , n185447 , n185448 , 
 n18136 , n185450 , n185451 , n18139 , n185453 , n185454 , n18142 , n185456 , n18144 , n185458 , 
 n185459 , n18147 , n185461 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , 
 n185469 , n18157 , n18158 , n185472 , n185473 , n185474 , n18162 , n185476 , n185477 , n18165 , 
 n185479 , n185480 , n18168 , n185482 , n185483 , n18171 , n185485 , n185486 , n18174 , n185488 , 
 n185489 , n18177 , n185491 , n185492 , n18180 , n185494 , n185495 , n18183 , n18184 , n185498 , 
 n18186 , n185500 , n18188 , n185502 , n185503 , n185504 , n18192 , n185506 , n185507 , n18195 , 
 n185509 , n185510 , n18198 , n18199 , n185513 , n185514 , n18202 , n185516 , n185517 , n18205 , 
 n185519 , n185520 , n18208 , n185522 , n185523 , n18211 , n185525 , n185526 , n18214 , n185528 , 
 n18216 , n18217 , n185531 , n185532 , n18220 , n18221 , n18222 , n18223 , n185537 , n185538 , 
 n18226 , n18227 , n18228 , n18229 , n185543 , n185544 , n18232 , n185546 , n18234 , n185548 , 
 n18236 , n18237 , n185551 , n185552 , n185553 , n18241 , n185555 , n185556 , n18244 , n185558 , 
 n185559 , n18247 , n185561 , n185562 , n18250 , n185564 , n18252 , n18253 , n185567 , n185568 , 
 n185569 , n185570 , n185571 , n18262 , n185573 , n18264 , n185575 , n18266 , n185577 , n18268 , 
 n18269 , n185580 , n185581 , n185582 , n18273 , n185584 , n185585 , n18276 , n185587 , n185588 , 
 n18279 , n185590 , n18281 , n185592 , n18283 , n185594 , n185595 , n18286 , n185597 , n185598 , 
 n185599 , n18290 , n185601 , n18292 , n18293 , n185604 , n185605 , n185606 , n18297 , n185608 , 
 n185609 , n18300 , n185611 , n185612 , n18303 , n185614 , n185615 , n18306 , n185617 , n18308 , 
 n185619 , n18310 , n18311 , n185622 , n18313 , n185624 , n18315 , n185626 , n185627 , n18318 , 
 n185629 , n185630 , n18321 , n185632 , n185633 , n18324 , n185635 , n185636 , n18327 , n18328 , 
 n185639 , n18330 , n185641 , n185642 , n18333 , n18334 , n18335 , n18336 , n18337 , n185648 , 
 n185649 , n18340 , n185651 , n185652 , n18343 , n18344 , n18345 , n18346 , n18347 , n185658 , 
 n185659 , n18350 , n185661 , n185662 , n18353 , n18354 , n18355 , n18356 , n185667 , n185668 , 
 n18359 , n185670 , n185671 , n18362 , n185673 , n185674 , n18365 , n185676 , n185677 , n185678 , 
 n18369 , n185680 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n185688 , 
 n185689 , n18380 , n185691 , n185692 , n18383 , n185694 , n18385 , n18386 , n185697 , n18388 , 
 n185699 , n185700 , n18391 , n185702 , n18393 , n18394 , n185705 , n18396 , n185707 , n185708 , 
 n18402 , n185710 , n185711 , n18405 , n185713 , n185714 , n18408 , n185716 , n185717 , n185718 , 
 n185719 , n18413 , n185721 , n185722 , n18416 , n185724 , n185725 , n18419 , n18420 , n185728 , 
 n18422 , n18423 , n185731 , n18425 , n185733 , n18427 , n18428 , n18429 , n185737 , n18431 , 
 n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n185746 , n18440 , n185748 , 
 n185749 , n18443 , n185751 , n185752 , n185753 , n185754 , n18448 , n185756 , n185757 , n18451 , 
 n18452 , n185760 , n18454 , n185762 , n185763 , n18457 , n18458 , n185766 , n18460 , n185768 , 
 n18462 , n185770 , n18464 , n18465 , n185773 , n185774 , n185775 , n185776 , n18470 , n185778 , 
 n18472 , n185780 , n185781 , n18475 , n18476 , n185784 , n18478 , n18479 , n185787 , n18481 , 
 n185789 , n18483 , n185791 , n185792 , n18486 , n185794 , n185795 , n185796 , n18490 , n185798 , 
 n185799 , n185800 , n18494 , n185802 , n185803 , n18497 , n185805 , n185806 , n18500 , n185808 , 
 n185809 , n18503 , n185811 , n18505 , n18506 , n18507 , n185815 , n18509 , n185817 , n18511 , 
 n185819 , n185820 , n18514 , n18515 , n185823 , n18517 , n185825 , n18519 , n185827 , n185828 , 
 n18522 , n18523 , n185831 , n18525 , n185833 , n185834 , n18528 , n185836 , n185837 , n18531 , 
 n185839 , n18536 , n185841 , n18538 , n185843 , n185844 , n18541 , n185846 , n18543 , n185848 , 
 n18545 , n18546 , n18547 , n185852 , n18549 , n185854 , n185855 , n185856 , n18553 , n185858 , 
 n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n185866 , n18563 , n185868 , 
 n185869 , n18566 , n185871 , n18568 , n18569 , n185874 , n18571 , n185876 , n18573 , n185878 , 
 n185879 , n18576 , n185881 , n185882 , n185883 , n185884 , n18581 , n185886 , n185887 , n18584 , 
 n185889 , n185890 , n18587 , n185892 , n185893 , n18590 , n185895 , n185896 , n185897 , n18594 , 
 n185899 , n18596 , n185901 , n185902 , n18599 , n185904 , n18601 , n185906 , n185907 , n18604 , 
 n18605 , n185910 , n18607 , n185912 , n185913 , n18610 , n18611 , n185916 , n18613 , n185918 , 
 n18615 , n185920 , n18617 , n185922 , n185923 , n18620 , n185925 , n18622 , n18623 , n185928 , 
 n185929 , n18626 , n185931 , n18628 , n185933 , n185934 , n18631 , n185936 , n185937 , n185938 , 
 n185939 , n18636 , n185941 , n185942 , n18639 , n185944 , n185945 , n18642 , n18643 , n185948 , 
 n18645 , n18646 , n185951 , n18648 , n185953 , n18650 , n185955 , n18652 , n18653 , n185958 , 
 n18658 , n185960 , n185961 , n18661 , n185963 , n185964 , n18664 , n185966 , n185967 , n18667 , 
 n185969 , n185970 , n18670 , n185972 , n185973 , n18673 , n18674 , n185976 , n18676 , n18677 , 
 n185979 , n18679 , n185981 , n18681 , n185983 , n185984 , n185985 , n18685 , n185987 , n185988 , 
 n18688 , n185990 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n185997 , n18697 , 
 n185999 , n186000 , n18700 , n186002 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , 
 n18708 , n18709 , n18710 , n18711 , n186013 , n186014 , n18714 , n186016 , n18716 , n18717 , 
 n186019 , n186020 , n18720 , n186022 , n186023 , n18723 , n186025 , n186026 , n18726 , n186028 , 
 n186029 , n18729 , n186031 , n186032 , n18732 , n186034 , n186035 , n18735 , n186037 , n18737 , 
 n18738 , n186040 , n18740 , n186042 , n186043 , n18743 , n186045 , n186046 , n18746 , n186048 , 
 n186049 , n18749 , n18750 , n186052 , n18752 , n186054 , n186055 , n18755 , n18756 , n18757 , 
 n18758 , n18759 , n186061 , n18761 , n186063 , n186064 , n18764 , n186066 , n186067 , n18767 , 
 n186069 , n186070 , n186071 , n18774 , n186073 , n18776 , n186075 , n186076 , n186077 , n18780 , 
 n186079 , n186080 , n18783 , n186082 , n18785 , n18786 , n18787 , n186086 , n18789 , n186088 , 
 n18791 , n18792 , n186091 , n18794 , n186093 , n186094 , n186095 , n18798 , n186097 , n186098 , 
 n18801 , n186100 , n186101 , n186102 , n18805 , n186104 , n18807 , n18808 , n18809 , n18810 , 
 n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , 
 n186119 , n186120 , n18823 , n186122 , n18825 , n18826 , n186125 , n186126 , n18829 , n186128 , 
 n18831 , n186130 , n186131 , n18834 , n186133 , n186134 , n18837 , n186136 , n186137 , n18840 , 
 n18841 , n186140 , n18843 , n18844 , n186143 , n18846 , n186145 , n186146 , n18849 , n186148 , 
 n186149 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , 
 n18861 , n18862 , n186161 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n186168 , 
 n18874 , n18875 , n186171 , n186172 , n18878 , n186174 , n186175 , n18881 , n186177 , n186178 , 
 n186179 , n186180 , n18886 , n186182 , n186183 , n18889 , n18890 , n18891 , n186187 , n186188 , 
 n186189 , n18895 , n186191 , n186192 , n18898 , n186194 , n186195 , n18901 , n186197 , n186198 , 
 n18904 , n18905 , n18906 , n18907 , n186203 , n18909 , n186205 , n186206 , n18912 , n186208 , 
 n186209 , n186210 , n186211 , n18917 , n186213 , n186214 , n18920 , n186216 , n186217 , n18923 , 
 n186219 , n186220 , n18926 , n186222 , n186223 , n18929 , n186225 , n186226 , n18932 , n18933 , 
 n18934 , n18935 , n18936 , n18937 , n18938 , n186234 , n186235 , n18941 , n186237 , n18943 , 
 n186239 , n18945 , n186241 , n186242 , n18948 , n18949 , n186245 , n186246 , n18952 , n186248 , 
 n186249 , n18955 , n186251 , n186252 , n18958 , n186254 , n186255 , n186256 , n186257 , n18963 , 
 n186259 , n186260 , n18969 , n186262 , n186263 , n18972 , n186265 , n186266 , n186267 , n186268 , 
 n18977 , n186270 , n186271 , n18980 , n186273 , n18982 , n186275 , n18984 , n186277 , n186278 , 
 n18987 , n186280 , n18989 , n186282 , n18991 , n18992 , n186285 , n18994 , n186287 , n186288 , 
 n18997 , n18998 , n18999 , n186292 , n19001 , n186294 , n186295 , n19004 , n186297 , n186298 , 
 n186299 , n186300 , n19009 , n186302 , n186303 , n19012 , n186305 , n186306 , n19015 , n186308 , 
 n186309 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , 
 n19027 , n19028 , n19029 , n19030 , n19031 , n186324 , n19033 , n186326 , n186327 , n186328 , 
 n186329 , n19038 , n186331 , n186332 , n19041 , n186334 , n186335 , n19044 , n186337 , n186338 , 
 n19050 , n186340 , n186341 , n19053 , n186343 , n186344 , n186345 , n186346 , n19058 , n186348 , 
 n186349 , n19061 , n186351 , n186352 , n19064 , n19065 , n186355 , n186356 , n19068 , n19069 , 
 n19070 , n186360 , n186361 , n19073 , n19074 , n19075 , n186365 , n186366 , n186367 , n186368 , 
 n19080 , n186370 , n19082 , n186372 , n186373 , n186374 , n186375 , n186376 , n19088 , n19089 , 
 n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n186388 , 
 n19100 , n19101 , n19102 , n19103 , n186393 , n19105 , n186395 , n186396 , n186397 , n186398 , 
 n19110 , n186400 , n186401 , n19113 , n186403 , n186404 , n19116 , n186406 , n19118 , n19119 , 
 n186409 , n186410 , n19125 , n186412 , n186413 , n19128 , n19129 , n19130 , n19131 , n19132 , 
 n186419 , n19134 , n186421 , n19136 , n186423 , n19138 , n186425 , n19140 , n186427 , n19142 , 
 n186429 , n186430 , n19145 , n186432 , n186433 , n19148 , n186435 , n186436 , n19151 , n19152 , 
 n186439 , n19154 , n186441 , n186442 , n19157 , n186444 , n186445 , n186446 , n186447 , n19162 , 
 n186449 , n186450 , n19165 , n186452 , n186453 , n19168 , n186455 , n19170 , n186457 , n186458 , 
 n19173 , n186460 , n186461 , n19176 , n19177 , n186464 , n19179 , n19180 , n186467 , n186468 , 
 n19186 , n186470 , n186471 , n19189 , n186473 , n19191 , n186475 , n186476 , n19194 , n186478 , 
 n186479 , n19197 , n186481 , n19199 , n19200 , n19201 , n186485 , n186486 , n19204 , n186488 , 
 n186489 , n19207 , n186491 , n186492 , n19210 , n186494 , n19212 , n19213 , n186497 , n186498 , 
 n19216 , n186500 , n186501 , n19219 , n186503 , n19221 , n19222 , n186506 , n186507 , n19225 , 
 n186509 , n186510 , n19228 , n186512 , n19230 , n19231 , n186515 , n186516 , n19234 , n186518 , 
 n186519 , n19240 , n186521 , n186522 , n19243 , n186524 , n186525 , n186526 , n19247 , n186528 , 
 n186529 , n19250 , n19251 , n186532 , n19253 , n186534 , n186535 , n186536 , n19257 , n186538 , 
 n186539 , n19260 , n186541 , n19262 , n19263 , n19264 , n19265 , n186546 , n186547 , n186548 , 
 n19269 , n186550 , n186551 , n19272 , n186553 , n186554 , n19275 , n186556 , n19277 , n186558 , 
 n186559 , n186560 , n186561 , n186562 , n186563 , n186564 , n186565 , n186566 , n186567 , n186568 , 
 n186569 , n186570 , n186571 , n186572 , n186573 , n186574 , n186575 , n186576 , n186577 , n186578 , 
 n186579 , n186580 , n186581 , n186582 , n186583 , n186584 , n186585 , n186586 , n186587 , n186588 , 
 n186589 , n186590 , n186591 , n186592 , n186593 , n186594 , n186595 , n186596 , n186597 , n186598 , 
 n186599 , n186600 , n186601 , n186602 , n186603 , n186604 , n186605 , n186606 , n186607 , n186608 , 
 n186609 , n186610 , n186611 , n186612 , n186613 , n186614 , n186615 , n186616 , n186617 , n186618 , 
 n186619 , n186620 , n186621 , n186622 , n186623 , n186624 , n186625 , n186626 , n186627 , n186628 , 
 n186629 , n186630 , n186631 , n186632 , n186633 , n186634 , n186635 , n186636 , n186637 , n186638 , 
 n186639 , n186640 , n186641 , n186642 , n186643 , n186644 , n186645 , n186646 , n186647 , n186648 , 
 n186649 , n186650 , n186651 , n186652 , n186653 , n186654 , n186655 , n186656 , n186657 , n186658 , 
 n186659 , n186660 , n186661 , n186662 , n186663 , n186664 , n186665 , n186666 , n186667 , n186668 , 
 n186669 , n186670 , n186671 , n186672 , n186673 , n186674 , n186675 , n186676 , n186677 , n186678 , 
 n186679 , n186680 , n186681 , n186682 , n186683 , n186684 , n186685 , n186686 , n186687 , n19411 , 
 n186689 , n186690 , n186691 , n19415 , n186693 , n186694 , n19418 , n186696 , n186697 , n19421 , 
 n186699 , n186700 , n19424 , n19425 , n19426 , n186704 , n186705 , n19429 , n186707 , n186708 , 
 n19432 , n186710 , n186711 , n186712 , n186713 , n19437 , n186715 , n186716 , n186717 , n19441 , 
 n186719 , n19443 , n19444 , n186722 , n19446 , n186724 , n19448 , n186726 , n186727 , n19451 , 
 n186729 , n186730 , n19454 , n186732 , n19456 , n186734 , n19458 , n19459 , n186737 , n19461 , 
 n186739 , n19463 , n186741 , n186742 , n19466 , n186744 , n186745 , n19469 , n186747 , n186748 , 
 n186749 , n19473 , n186751 , n19475 , n19476 , n186754 , n186755 , n186756 , n19480 , n186758 , 
 n186759 , n19483 , n186761 , n186762 , n19486 , n186764 , n186765 , n186766 , n19490 , n186768 , 
 n19492 , n19493 , n19494 , n186772 , n186773 , n186774 , n19498 , n186776 , n186777 , n19501 , 
 n186779 , n186780 , n19504 , n186782 , n186783 , n19507 , n186785 , n19509 , n186787 , n19511 , 
 n186789 , n186790 , n19514 , n19515 , n186793 , n186794 , n19518 , n186796 , n186797 , n19521 , 
 n186799 , n186800 , n19524 , n186802 , n186803 , n19527 , n186805 , n186806 , n19530 , n186808 , 
 n19532 , n186810 , n19534 , n19535 , n186813 , n19537 , n186815 , n19539 , n186817 , n186818 , 
 n19542 , n186820 , n186821 , n186822 , n19546 , n186824 , n19548 , n19549 , n186827 , n19551 , 
 n186829 , n19553 , n186831 , n186832 , n19556 , n186834 , n186835 , n19559 , n186837 , n19561 , 
 n186839 , n19563 , n19564 , n186842 , n19566 , n186844 , n19568 , n186846 , n186847 , n19571 , 
 n186849 , n186850 , n19574 , n186852 , n186853 , n19577 , n186855 , n186856 , n19580 , n19581 , 
 n186859 , n186860 , n19584 , n19585 , n186863 , n186864 , n19588 , n19589 , n19590 , n186868 , 
 n186869 , n19593 , n19594 , n19595 , n186873 , n186874 , n19598 , n186876 , n19600 , n19601 , 
 n19602 , n186880 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , 
 n19612 , n19613 , n186891 , n19615 , n186893 , n186894 , n19618 , n19619 , n186897 , n19621 , 
 n186899 , n186900 , n186901 , n186902 , n19626 , n186904 , n186905 , n19629 , n186907 , n19631 , 
 n19632 , n186910 , n186911 , n19635 , n186913 , n186914 , n19638 , n186916 , n186917 , n19641 , 
 n19642 , n186920 , n19644 , n186922 , n19646 , n186924 , n186925 , n19649 , n19650 , n186928 , 
 n186929 , n19653 , n186931 , n186932 , n19656 , n186934 , n186935 , n19659 , n19660 , n19661 , 
 n186939 , n186940 , n19664 , n186942 , n186943 , n19667 , n19668 , n19669 , n186947 , n19671 , 
 n186949 , n19673 , n19674 , n186952 , n186953 , n19677 , n186955 , n186956 , n19680 , n186958 , 
 n186959 , n19683 , n186961 , n186962 , n19686 , n186964 , n186965 , n19689 , n186967 , n19691 , 
 n19692 , n186970 , n186971 , n19695 , n186973 , n186974 , n19698 , n186976 , n186977 , n19701 , 
 n19702 , n186980 , n19704 , n186982 , n186983 , n19707 , n186985 , n19709 , n186987 , n186988 , 
 n19712 , n19713 , n186991 , n186992 , n19716 , n186994 , n186995 , n19719 , n186997 , n19721 , 
 n19722 , n187000 , n187001 , n19725 , n187003 , n187004 , n19728 , n187006 , n187007 , n19731 , 
 n187009 , n187010 , n19734 , n187012 , n187013 , n19737 , n187015 , n187016 , n187017 , n19741 , 
 n187019 , n19743 , n187021 , n187022 , n19746 , n187024 , n187025 , n19749 , n19750 , n19751 , 
 n19752 , n19753 , n19754 , n187032 , n19756 , n19757 , n19758 , n19759 , n187037 , n187038 , 
 n19762 , n187040 , n19764 , n19765 , n19766 , n187044 , n19768 , n187046 , n19770 , n187048 , 
 n19772 , n19773 , n19774 , n187052 , n187053 , n19777 , n187055 , n19779 , n19780 , n187058 , 
 n187059 , n19783 , n187061 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , 
 n19792 , n187070 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , 
 n19802 , n19803 , n19804 , n187082 , n19806 , n19807 , n19808 , n187086 , n187087 , n19811 , 
 n187089 , n187090 , n19814 , n19815 , n19816 , n187094 , n187095 , n187096 , n187097 , n187098 , 
 n19822 , n187100 , n187101 , n19825 , n187103 , n187104 , n19828 , n19829 , n187107 , n187108 , 
 n19832 , n187110 , n187111 , n19835 , n187113 , n19837 , n187115 , n19839 , n19840 , n187118 , 
 n187119 , n19843 , n187121 , n187122 , n19846 , n187124 , n187125 , n19849 , n187127 , n187128 , 
 n19852 , n187130 , n187131 , n19855 , n187133 , n19857 , n19858 , n187136 , n187137 , n19861 , 
 n187139 , n187140 , n19864 , n187142 , n187143 , n19867 , n19868 , n19869 , n187147 , n187148 , 
 n19872 , n19873 , n187151 , n19875 , n187153 , n187154 , n19878 , n187156 , n187157 , n19881 , 
 n187159 , n19883 , n19884 , n187162 , n187163 , n19887 , n187165 , n187166 , n19890 , n187168 , 
 n187169 , n19893 , n187171 , n19895 , n187173 , n19897 , n19898 , n187176 , n187177 , n19901 , 
 n187179 , n187180 , n19904 , n187182 , n187183 , n19907 , n19908 , n187186 , n19910 , n187188 , 
 n19912 , n19913 , n187191 , n187192 , n19916 , n187194 , n187195 , n19919 , n187197 , n187198 , 
 n19922 , n19923 , n19924 , n187202 , n187203 , n187204 , n187205 , n19929 , n187207 , n187208 , 
 n19932 , n187210 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , 
 n19942 , n19943 , n187221 , n187222 , n19946 , n187224 , n187225 , n19949 , n187227 , n187228 , 
 n187229 , n187230 , n19954 , n187232 , n187233 , n19957 , n187235 , n19959 , n19960 , n187238 , 
 n187239 , n19963 , n187241 , n187242 , n19966 , n187244 , n187245 , n19969 , n187247 , n187248 , 
 n19972 , n187250 , n187251 , n19975 , n187253 , n19977 , n19978 , n187256 , n187257 , n19981 , 
 n187259 , n187260 , n19984 , n187262 , n187263 , n19987 , n19988 , n19989 , n187267 , n187268 , 
 n19992 , n187270 , n187271 , n19995 , n187273 , n187274 , n187275 , n187276 , n20000 , n187278 , 
 n187279 , n20003 , n187281 , n20005 , n20006 , n187284 , n187285 , n20009 , n187287 , n187288 , 
 n20012 , n187290 , n187291 , n20015 , n187293 , n187294 , n20018 , n187296 , n187297 , n20021 , 
 n187299 , n20023 , n20024 , n187302 , n187303 , n20027 , n187305 , n187306 , n20030 , n187308 , 
 n187309 , n20033 , n20034 , n20035 , n187313 , n187314 , n20038 , n20039 , n20040 , n187318 , 
 n187319 , n20043 , n20044 , n20045 , n187323 , n187324 , n20048 , n20049 , n20050 , n20051 , 
 n20052 , n187330 , n20054 , n187332 , n20056 , n187334 , n20058 , n187336 , n20060 , n20061 , 
 n187339 , n187340 , n20064 , n20065 , n187343 , n187344 , n20068 , n20069 , n187347 , n187348 , 
 n20072 , n20073 , n187351 , n20075 , n20076 , n20077 , n187355 , n20079 , n20080 , n20081 , 
 n20082 , n20083 , n20084 , n20085 , n20086 , n187364 , n20088 , n187366 , n20090 , n187368 , 
 n20092 , n20093 , n187371 , n187372 , n20096 , n20097 , n187375 , n187376 , n187377 , n20101 , 
 n20102 , n187380 , n20104 , n20105 , n187383 , n187384 , n20108 , n187386 , n187387 , n20111 , 
 n187389 , n187390 , n187391 , n187392 , n20116 , n187394 , n187395 , n20119 , n187397 , n187398 , 
 n20122 , n20123 , n20124 , n187402 , n187403 , n20127 , n187405 , n20129 , n187407 , n187408 , 
 n187409 , n20133 , n187411 , n187412 , n20136 , n187414 , n20138 , n20139 , n187417 , n187418 , 
 n187419 , n20143 , n187421 , n187422 , n20146 , n187424 , n187425 , n20149 , n187427 , n187428 , 
 n20152 , n187430 , n187431 , n20155 , n187433 , n187434 , n20158 , n20159 , n20160 , n20161 , 
 n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n187447 , n20171 , 
 n187449 , n187450 , n20174 , n187452 , n187453 , n20177 , n20178 , n20179 , n20180 , n20181 , 
 n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n187467 , n20191 , 
 n187469 , n187470 , n20194 , n20195 , n20196 , n20197 , n187475 , n20199 , n187477 , n187478 , 
 n20202 , n187480 , n20204 , n187482 , n187483 , n20207 , n187485 , n187486 , n20210 , n20211 , 
 n20212 , n187490 , n187491 , n20215 , n20216 , n20217 , n187495 , n187496 , n20220 , n20221 , 
 n20222 , n187500 , n187501 , n20225 , n187503 , n187504 , n187505 , n20229 , n187507 , n20231 , 
 n20232 , n187510 , n20234 , n187512 , n20236 , n187514 , n20238 , n20239 , n20240 , n20241 , 
 n20242 , n20243 , n20244 , n20245 , n20246 , n187524 , n20248 , n187526 , n20250 , n187528 , 
 n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n187538 , 
 n187539 , n20263 , n187541 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , 
 n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n187557 , n20281 , 
 n187559 , n20283 , n187561 , n20285 , n187563 , n20287 , n20288 , n20289 , n20290 , n20291 , 
 n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , 
 n20302 , n187580 , n20304 , n20305 , n187583 , n187584 , n20308 , n187586 , n187587 , n20311 , 
 n187589 , n20313 , n20314 , n20315 , n187593 , n187594 , n20318 , n187596 , n20320 , n20321 , 
 n187599 , n20323 , n187601 , n187602 , n20326 , n187604 , n20328 , n187606 , n187607 , n20331 , 
 n187609 , n187610 , n20334 , n20335 , n187613 , n20337 , n20338 , n20339 , n20340 , n187618 , 
 n20342 , n187620 , n187621 , n20345 , n187623 , n187624 , n20348 , n187626 , n187627 , n20351 , 
 n187629 , n187630 , n20354 , n187632 , n20356 , n20357 , n20358 , n187636 , n187637 , n187638 , 
 n20362 , n187640 , n187641 , n20365 , n187643 , n187644 , n20368 , n187646 , n187647 , n20371 , 
 n187649 , n187650 , n20374 , n20375 , n187653 , n187654 , n20378 , n187656 , n187657 , n20381 , 
 n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , 
 n187669 , n20393 , n20394 , n20395 , n20396 , n187674 , n20398 , n187676 , n20400 , n187678 , 
 n187679 , n20403 , n187681 , n187682 , n20406 , n187684 , n187685 , n187686 , n187687 , n20411 , 
 n187689 , n187690 , n20414 , n187692 , n20416 , n20417 , n20418 , n20419 , n20420 , n187698 , 
 n20422 , n20423 , n187701 , n20425 , n187703 , n187704 , n20428 , n187706 , n20430 , n20431 , 
 n20432 , n187710 , n20434 , n20435 , n20436 , n20437 , n187715 , n20439 , n20440 , n20441 , 
 n187719 , n187720 , n20444 , n187722 , n187723 , n20447 , n187725 , n187726 , n20450 , n187728 , 
 n20452 , n187730 , n187731 , n20455 , n187733 , n20457 , n20458 , n20459 , n20460 , n20461 , 
 n20462 , n20463 , n187741 , n20465 , n20466 , n187744 , n20468 , n187746 , n20470 , n187748 , 
 n187749 , n20473 , n187751 , n187752 , n20476 , n187754 , n20478 , n187756 , n20480 , n20481 , 
 n187759 , n187760 , n187761 , n20485 , n187763 , n187764 , n20488 , n187766 , n187767 , n20491 , 
 n187769 , n187770 , n20494 , n187772 , n187773 , n187774 , n187775 , n20499 , n187777 , n187778 , 
 n20502 , n187780 , n187781 , n187782 , n20506 , n187784 , n20508 , n20509 , n187787 , n20511 , 
 n187789 , n20513 , n187791 , n187792 , n20516 , n187794 , n187795 , n20519 , n187797 , n20521 , 
 n20522 , n187800 , n187801 , n187802 , n20526 , n187804 , n187805 , n20529 , n187807 , n187808 , 
 n20532 , n187810 , n20534 , n187812 , n20536 , n187814 , n20538 , n20539 , n20540 , n20541 , 
 n20542 , n187820 , n20544 , n187822 , n20546 , n20547 , n20548 , n187826 , n20550 , n187828 , 
 n20552 , n20553 , n20554 , n187832 , n20556 , n20557 , n20558 , n187836 , n187837 , n187838 , 
 n20562 , n187840 , n187841 , n20565 , n187843 , n187844 , n20568 , n187846 , n20570 , n187848 , 
 n187849 , n20573 , n187851 , n187852 , n20576 , n187854 , n20578 , n187856 , n20580 , n187858 , 
 n20582 , n187860 , n20584 , n20585 , n187863 , n20587 , n187865 , n187866 , n20590 , n187868 , 
 n20592 , n187870 , n187871 , n20595 , n187873 , n20597 , n187875 , n20599 , n187877 , n20601 , 
 n20602 , n187880 , n20604 , n187882 , n20606 , n187884 , n187885 , n20609 , n187887 , n20611 , 
 n20612 , n20613 , n20614 , n20615 , n20616 , n187894 , n20618 , n187896 , n187897 , n20621 , 
 n187899 , n187900 , n20624 , n187902 , n187903 , n187904 , n20628 , n187906 , n187907 , n20631 , 
 n20632 , n20633 , n20634 , n20635 , n187913 , n187914 , n20638 , n187916 , n20640 , n20641 , 
 n187919 , n20643 , n187921 , n187922 , n20646 , n187924 , n187925 , n20649 , n187927 , n187928 , 
 n20652 , n187930 , n20654 , n187932 , n20656 , n20657 , n187935 , n20659 , n187937 , n20661 , 
 n187939 , n187940 , n20664 , n187942 , n187943 , n20667 , n20668 , n187946 , n20670 , n20671 , 
 n20672 , n20673 , n20674 , n20675 , n187953 , n20677 , n20678 , n20679 , n20680 , n20681 , 
 n20682 , n20683 , n187961 , n20685 , n187963 , n187964 , n187965 , n187966 , n20690 , n187968 , 
 n187969 , n187970 , n187971 , n20695 , n187973 , n187974 , n20698 , n187976 , n187977 , n20701 , 
 n187979 , n187980 , n20704 , n187982 , n20706 , n187984 , n20708 , n187986 , n187987 , n20711 , 
 n187989 , n20713 , n187991 , n187992 , n20716 , n187994 , n20718 , n187996 , n187997 , n20721 , 
 n187999 , n188000 , n20724 , n20725 , n20726 , n20727 , n188005 , n20729 , n20730 , n188008 , 
 n20732 , n188010 , n188011 , n188012 , n20736 , n188014 , n188015 , n20739 , n188017 , n20741 , 
 n188019 , n188020 , n20744 , n188022 , n188023 , n20747 , n188025 , n20749 , n20750 , n188028 , 
 n188029 , n20753 , n188031 , n188032 , n20756 , n188034 , n188035 , n20759 , n188037 , n20761 , 
 n20762 , n188040 , n188041 , n20765 , n188043 , n188044 , n20768 , n20769 , n188047 , n20771 , 
 n20772 , n188050 , n188051 , n20775 , n188053 , n188054 , n20778 , n188056 , n20780 , n20781 , 
 n188059 , n188060 , n20784 , n188062 , n20786 , n20787 , n20788 , n20789 , n188067 , n20791 , 
 n188069 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n188078 , 
 n188079 , n188080 , n20804 , n188082 , n188083 , n20807 , n188085 , n20809 , n20810 , n20811 , 
 n20812 , n188090 , n188091 , n20815 , n188093 , n20817 , n20818 , n20819 , n188097 , n188098 , 
 n188099 , n20823 , n188101 , n188102 , n20826 , n188104 , n20828 , n20829 , n188107 , n188108 , 
 n188109 , n20833 , n188111 , n188112 , n20836 , n188114 , n20838 , n20839 , n20840 , n20841 , 
 n20842 , n20843 , n188121 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , 
 n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , 
 n20862 , n20863 , n188141 , n20865 , n188143 , n188144 , n20868 , n188146 , n188147 , n188148 , 
 n188149 , n20873 , n188151 , n188152 , n20876 , n20877 , n188155 , n20879 , n20880 , n188158 , 
 n188159 , n188160 , n20884 , n188162 , n188163 , n20887 , n188165 , n188166 , n20890 , n188168 , 
 n20892 , n188170 , n20894 , n188172 , n20896 , n20897 , n188175 , n188176 , n20900 , n188178 , 
 n20902 , n20903 , n188181 , n20905 , n188183 , n20907 , n188185 , n20909 , n20910 , n20911 , 
 n20912 , n188190 , n188191 , n188192 , n20916 , n188194 , n188195 , n20919 , n188197 , n20921 , 
 n20922 , n188200 , n20924 , n188202 , n20926 , n20927 , n20928 , n20929 , n188207 , n20931 , 
 n188209 , n20933 , n188211 , n20935 , n188213 , n188214 , n20938 , n188216 , n188217 , n20941 , 
 n20942 , n188220 , n188221 , n188222 , n20946 , n188224 , n188225 , n20949 , n188227 , n188228 , 
 n20952 , n188230 , n20954 , n188232 , n20956 , n188234 , n20958 , n20959 , n188237 , n20961 , 
 n188239 , n188240 , n20964 , n188242 , n188243 , n188244 , n20968 , n188246 , n20970 , n20971 , 
 n20972 , n188250 , n20974 , n188252 , n20976 , n20977 , n188255 , n20979 , n188257 , n188258 , 
 n20982 , n20983 , n188261 , n20985 , n20986 , n188264 , n20988 , n20989 , n20990 , n20991 , 
 n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n188277 , n188278 , 
 n188279 , n21003 , n188281 , n188282 , n21006 , n188284 , n21008 , n21009 , n21010 , n21011 , 
 n21012 , n188290 , n188291 , n188292 , n21016 , n188294 , n188295 , n21019 , n188297 , n21021 , 
 n21022 , n188300 , n21024 , n188302 , n188303 , n21027 , n188305 , n21029 , n21030 , n21031 , 
 n188309 , n188310 , n21034 , n188312 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , 
 n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , 
 n21052 , n21053 , n21054 , n21055 , n188333 , n21057 , n188335 , n21059 , n21060 , n188338 , 
 n21062 , n188340 , n21064 , n188342 , n188343 , n21067 , n188345 , n21069 , n21070 , n21071 , 
 n21072 , n21073 , n21074 , n21075 , n21076 , n188354 , n21078 , n188356 , n21080 , n188358 , 
 n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n188368 , 
 n21092 , n188370 , n21094 , n21095 , n21096 , n188374 , n21098 , n188376 , n21100 , n21101 , 
 n188379 , n188380 , n188381 , n21105 , n188383 , n188384 , n21108 , n188386 , n188387 , n21111 , 
 n188389 , n188390 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n188397 , n21121 , 
 n21122 , n188400 , n188401 , n21125 , n21126 , n188404 , n188405 , n188406 , n21130 , n188408 , 
 n21132 , n21133 , n188411 , n188412 , n188413 , n21137 , n188415 , n188416 , n21140 , n188418 , 
 n188419 , n21143 , n188421 , n188422 , n21146 , n188424 , n188425 , n21149 , n21150 , n188428 , 
 n21152 , n21153 , n188431 , n188432 , n21156 , n188434 , n21158 , n21159 , n21160 , n21161 , 
 n21162 , n21163 , n21164 , n188442 , n21166 , n188444 , n21168 , n21169 , n188447 , n21171 , 
 n188449 , n188450 , n188451 , n188452 , n21176 , n188454 , n188455 , n21179 , n188457 , n21181 , 
 n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n188466 , n21190 , n188468 , 
 n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , 
 n21202 , n21203 , n21204 , n21205 , n188483 , n21207 , n188485 , n21209 , n21210 , n188488 , 
 n21212 , n21213 , n188491 , n21215 , n188493 , n188494 , n21218 , n21219 , n188497 , n188498 , 
 n21222 , n188500 , n188501 , n21225 , n21226 , n21227 , n21228 , n188506 , n21230 , n188508 , 
 n21232 , n21233 , n188511 , n188512 , n21236 , n188514 , n188515 , n21239 , n188517 , n188518 , 
 n188519 , n21243 , n188521 , n188522 , n21246 , n21247 , n188525 , n21249 , n21250 , n188528 , 
 n188529 , n21253 , n188531 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , 
 n188539 , n188540 , n21264 , n21265 , n188543 , n21267 , n21268 , n188546 , n188547 , n188548 , 
 n188549 , n21273 , n188551 , n188552 , n21276 , n188554 , n21278 , n21279 , n188557 , n21281 , 
 n188559 , n188560 , n188561 , n21285 , n188563 , n188564 , n21288 , n188566 , n188567 , n188568 , 
 n188569 , n21293 , n188571 , n188572 , n21296 , n188574 , n21298 , n21299 , n188577 , n188578 , 
 n21302 , n188580 , n188581 , n21305 , n188583 , n188584 , n21308 , n188586 , n188587 , n21311 , 
 n188589 , n21313 , n188591 , n188592 , n188593 , n188594 , n21318 , n188596 , n188597 , n188598 , 
 n21322 , n188600 , n188601 , n21325 , n188603 , n21327 , n21328 , n21329 , n21330 , n188608 , 
 n21332 , n21333 , n188611 , n188612 , n21336 , n188614 , n188615 , n21339 , n188617 , n188618 , 
 n21342 , n188620 , n188621 , n21345 , n188623 , n188624 , n21348 , n188626 , n188627 , n21351 , 
 n188629 , n188630 , n21354 , n188632 , n21356 , n21357 , n188635 , n188636 , n188637 , n21361 , 
 n188639 , n188640 , n21364 , n188642 , n188643 , n21367 , n188645 , n188646 , n21370 , n188648 , 
 n188649 , n21373 , n188651 , n188652 , n21376 , n188654 , n188655 , n21379 , n188657 , n21381 , 
 n21382 , n188660 , n188661 , n188662 , n21386 , n188664 , n188665 , n21389 , n188667 , n188668 , 
 n21392 , n188670 , n188671 , n21395 , n188673 , n188674 , n21398 , n21399 , n21400 , n188678 , 
 n21402 , n188680 , n21404 , n21405 , n188683 , n188684 , n188685 , n21409 , n188687 , n188688 , 
 n21412 , n188690 , n188691 , n21415 , n188693 , n188694 , n21418 , n188696 , n188697 , n188698 , 
 n188699 , n21423 , n188701 , n188702 , n21426 , n188704 , n188705 , n188706 , n188707 , n21431 , 
 n188709 , n21433 , n21434 , n21435 , n188713 , n188714 , n188715 , n21439 , n188717 , n188718 , 
 n21442 , n188720 , n21444 , n188722 , n188723 , n21447 , n188725 , n21449 , n21450 , n21451 , 
 n188729 , n188730 , n188731 , n21455 , n188733 , n188734 , n21458 , n188736 , n21460 , n21461 , 
 n188739 , n188740 , n21464 , n188742 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , 
 n188749 , n21473 , n188751 , n21475 , n21476 , n188754 , n188755 , n188756 , n21480 , n188758 , 
 n188759 , n21483 , n188761 , n21485 , n21486 , n21487 , n21488 , n188766 , n21490 , n188768 , 
 n188769 , n21493 , n188771 , n188772 , n21496 , n188774 , n21498 , n21499 , n188777 , n188778 , 
 n188779 , n21503 , n188781 , n188782 , n21506 , n188784 , n188785 , n21509 , n188787 , n21511 , 
 n21512 , n188790 , n188791 , n21515 , n188793 , n21517 , n21518 , n21519 , n21520 , n21521 , 
 n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n188805 , n21529 , n188807 , n21531 , 
 n21532 , n21533 , n21534 , n188812 , n188813 , n21537 , n188815 , n188816 , n21540 , n188818 , 
 n21542 , n21543 , n188821 , n21545 , n188823 , n188824 , n188825 , n188826 , n21550 , n188828 , 
 n188829 , n21553 , n188831 , n188832 , n21556 , n188834 , n21558 , n21559 , n188837 , n21561 , 
 n188839 , n188840 , n188841 , n188842 , n21566 , n188844 , n188845 , n21569 , n188847 , n188848 , 
 n21572 , n21573 , n21574 , n188852 , n21576 , n21577 , n21578 , n188856 , n188857 , n21581 , 
 n188859 , n188860 , n21584 , n21585 , n21586 , n21587 , n21588 , n188866 , n21590 , n21591 , 
 n188869 , n188870 , n21594 , n21595 , n188873 , n188874 , n188875 , n21599 , n188877 , n21601 , 
 n21602 , n188880 , n188881 , n21605 , n21606 , n188884 , n21608 , n21609 , n21610 , n21611 , 
 n188889 , n21613 , n21614 , n21615 , n188893 , n188894 , n21618 , n21619 , n188897 , n21621 , 
 n21622 , n188900 , n21624 , n188902 , n21626 , n188904 , n21628 , n188906 , n21630 , n21631 , 
 n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , 
 n21642 , n21643 , n21644 , n188922 , n21646 , n188924 , n21648 , n21649 , n21650 , n21651 , 
 n21652 , n21653 , n21654 , n21655 , n21656 , n188934 , n21658 , n21659 , n21660 , n188938 , 
 n188939 , n21663 , n188941 , n188942 , n21666 , n21667 , n21668 , n21669 , n21670 , n188948 , 
 n21672 , n21673 , n188951 , n188952 , n188953 , n21677 , n188955 , n21679 , n21680 , n188958 , 
 n188959 , n21683 , n188961 , n188962 , n21686 , n188964 , n188965 , n21689 , n188967 , n21691 , 
 n188969 , n21693 , n21694 , n188972 , n188973 , n21697 , n188975 , n188976 , n21700 , n188978 , 
 n188979 , n21703 , n21704 , n188982 , n21706 , n188984 , n188985 , n21709 , n21710 , n188988 , 
 n21712 , n21713 , n188991 , n188992 , n21716 , n188994 , n188995 , n21719 , n188997 , n21721 , 
 n21722 , n189000 , n189001 , n21725 , n189003 , n189004 , n21728 , n189006 , n189007 , n21731 , 
 n189009 , n189010 , n21734 , n189012 , n189013 , n21737 , n21738 , n21739 , n21740 , n189018 , 
 n189019 , n21743 , n189021 , n21745 , n21746 , n21747 , n21748 , n189026 , n189027 , n21751 , 
 n189029 , n21753 , n21754 , n189032 , n21756 , n189034 , n189035 , n21759 , n189037 , n189038 , 
 n189039 , n21763 , n189041 , n21765 , n21766 , n21767 , n21768 , n21769 , n189047 , n21771 , 
 n21772 , n21773 , n189051 , n21775 , n189053 , n189054 , n21778 , n189056 , n21780 , n21781 , 
 n21782 , n189060 , n189061 , n21785 , n189063 , n21787 , n21788 , n21789 , n189067 , n189068 , 
 n21792 , n189070 , n21794 , n21795 , n21796 , n21797 , n21798 , n189076 , n189077 , n21801 , 
 n189079 , n21803 , n21804 , n21805 , n21806 , n189084 , n189085 , n21809 , n189087 , n189088 , 
 n21812 , n189090 , n21814 , n21815 , n189093 , n189094 , n21818 , n189096 , n189097 , n21821 , 
 n189099 , n21823 , n189101 , n21825 , n189103 , n21827 , n189105 , n189106 , n189107 , n189108 , 
 n21832 , n189110 , n189111 , n21835 , n189113 , n21837 , n21838 , n189116 , n189117 , n21841 , 
 n189119 , n189120 , n21844 , n189122 , n189123 , n21847 , n189125 , n21849 , n21850 , n189128 , 
 n21852 , n21853 , n189131 , n189132 , n21856 , n189134 , n189135 , n21859 , n189137 , n189138 , 
 n21862 , n21863 , n189141 , n189142 , n21866 , n189144 , n189145 , n21869 , n189147 , n189148 , 
 n21872 , n189150 , n21874 , n21875 , n189153 , n189154 , n21878 , n189156 , n189157 , n21881 , 
 n189159 , n189160 , n21884 , n189162 , n189163 , n21887 , n189165 , n189166 , n21890 , n189168 , 
 n21892 , n189170 , n21894 , n21895 , n189173 , n189174 , n21898 , n189176 , n189177 , n21901 , 
 n189179 , n189180 , n21904 , n189182 , n21906 , n189184 , n21908 , n21909 , n189187 , n189188 , 
 n21912 , n189190 , n189191 , n21915 , n189193 , n189194 , n21918 , n21919 , n21920 , n189198 , 
 n21922 , n189200 , n21924 , n21925 , n189203 , n189204 , n21928 , n189206 , n189207 , n21931 , 
 n189209 , n21933 , n189211 , n21935 , n189213 , n189214 , n21938 , n189216 , n189217 , n189218 , 
 n189219 , n21943 , n189221 , n189222 , n21946 , n189224 , n21948 , n189226 , n21950 , n189228 , 
 n189229 , n21953 , n21954 , n21955 , n189233 , n21957 , n189235 , n21959 , n189237 , n189238 , 
 n189239 , n21963 , n189241 , n189242 , n21966 , n189244 , n21968 , n21969 , n189247 , n189248 , 
 n189249 , n21973 , n189251 , n189252 , n21976 , n189254 , n189255 , n21979 , n189257 , n189258 , 
 n21982 , n189260 , n21984 , n21985 , n189263 , n189264 , n21988 , n189266 , n189267 , n21991 , 
 n189269 , n189270 , n21994 , n21995 , n21996 , n189274 , n189275 , n21999 , n189277 , n189278 , 
 n22002 , n189280 , n189281 , n22005 , n189283 , n22007 , n22008 , n22009 , n189287 , n189288 , 
 n22012 , n189290 , n189291 , n22015 , n189293 , n189294 , n22018 , n22019 , n22020 , n22021 , 
 n22022 , n189300 , n22024 , n189302 , n22026 , n22027 , n189305 , n189306 , n22030 , n189308 , 
 n189309 , n22033 , n189311 , n189312 , n22036 , n22037 , n189315 , n22039 , n189317 , n189318 , 
 n22042 , n189320 , n22044 , n189322 , n189323 , n22047 , n22048 , n189326 , n189327 , n22051 , 
 n189329 , n189330 , n22054 , n189332 , n22056 , n22057 , n189335 , n189336 , n22060 , n189338 , 
 n189339 , n22063 , n189341 , n189342 , n22066 , n189344 , n189345 , n22069 , n189347 , n189348 , 
 n22072 , n22073 , n22074 , n189352 , n22076 , n22077 , n22078 , n189356 , n22080 , n22081 , 
 n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , 
 n22092 , n22093 , n22094 , n22095 , n22096 , n189374 , n22098 , n22099 , n22100 , n22101 , 
 n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n189387 , n22111 , 
 n22112 , n22113 , n22114 , n189392 , n22116 , n189394 , n189395 , n189396 , n22120 , n22121 , 
 n189399 , n22123 , n189401 , n189402 , n22126 , n189404 , n22128 , n22129 , n189407 , n22131 , 
 n22132 , n22133 , n189411 , n189412 , n22136 , n189414 , n189415 , n189416 , n189417 , n22141 , 
 n189419 , n189420 , n22144 , n189422 , n189423 , n22147 , n22148 , n22149 , n189427 , n189428 , 
 n22152 , n189430 , n189431 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n189438 , 
 n189439 , n189440 , n189441 , n22165 , n189443 , n189444 , n189445 , n22169 , n189447 , n22171 , 
 n22172 , n189450 , n22174 , n189452 , n22176 , n189454 , n189455 , n22179 , n189457 , n189458 , 
 n22182 , n22183 , n22184 , n22185 , n22186 , n189464 , n189465 , n189466 , n22190 , n189468 , 
 n189469 , n22193 , n189471 , n22195 , n189473 , n22197 , n189475 , n189476 , n189477 , n22201 , 
 n189479 , n22203 , n22204 , n189482 , n22206 , n189484 , n189485 , n189486 , n22210 , n189488 , 
 n22212 , n22213 , n189491 , n189492 , n189493 , n22217 , n189495 , n189496 , n22220 , n189498 , 
 n189499 , n22223 , n189501 , n189502 , n22226 , n189504 , n22228 , n189506 , n22230 , n22231 , 
 n189509 , n189510 , n189511 , n22235 , n189513 , n189514 , n22238 , n189516 , n189517 , n22241 , 
 n189519 , n189520 , n22244 , n189522 , n189523 , n22247 , n22248 , n189526 , n22250 , n189528 , 
 n22252 , n22253 , n189531 , n22255 , n189533 , n189534 , n22258 , n22259 , n189537 , n22261 , 
 n189539 , n189540 , n22264 , n189542 , n189543 , n189544 , n22268 , n189546 , n189547 , n22271 , 
 n189549 , n189550 , n22274 , n22275 , n189553 , n189554 , n189555 , n22279 , n189557 , n189558 , 
 n22282 , n189560 , n189561 , n22285 , n189563 , n189564 , n22288 , n22289 , n22290 , n189568 , 
 n22292 , n189570 , n22294 , n189572 , n22296 , n189574 , n22298 , n189576 , n22300 , n189578 , 
 n22302 , n22303 , n22304 , n189582 , n22306 , n189584 , n22308 , n189586 , n189587 , n22311 , 
 n189589 , n189590 , n22314 , n189592 , n189593 , n22317 , n22318 , n22319 , n22320 , n189598 , 
 n189599 , n189600 , n22324 , n189602 , n189603 , n22327 , n189605 , n22329 , n22330 , n22331 , 
 n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n189616 , n189617 , n189618 , 
 n22342 , n189620 , n189621 , n22345 , n189623 , n22347 , n22348 , n22349 , n189627 , n22351 , 
 n189629 , n22353 , n22354 , n189632 , n22356 , n189634 , n22358 , n189636 , n189637 , n22361 , 
 n189639 , n22363 , n189641 , n22365 , n22366 , n189644 , n189645 , n22369 , n22370 , n189648 , 
 n189649 , n22373 , n22374 , n22375 , n189653 , n189654 , n189655 , n22379 , n189657 , n189658 , 
 n22382 , n189660 , n22384 , n189662 , n22386 , n189664 , n22388 , n189666 , n22390 , n22391 , 
 n189669 , n189670 , n189671 , n22395 , n189673 , n189674 , n22398 , n189676 , n189677 , n22401 , 
 n189679 , n189680 , n22404 , n189682 , n189683 , n22407 , n22408 , n189686 , n22410 , n189688 , 
 n22412 , n189690 , n189691 , n22415 , n189693 , n189694 , n189695 , n22419 , n189697 , n22421 , 
 n22422 , n189700 , n189701 , n22425 , n189703 , n189704 , n189705 , n22429 , n189707 , n189708 , 
 n22432 , n189710 , n189711 , n22435 , n189713 , n189714 , n22438 , n22439 , n189717 , n22441 , 
 n22442 , n189720 , n189721 , n22445 , n22446 , n189724 , n22448 , n189726 , n189727 , n22451 , 
 n22452 , n189730 , n189731 , n22455 , n22456 , n22457 , n22458 , n22459 , n189737 , n189738 , 
 n189739 , n189740 , n22464 , n189742 , n22466 , n22467 , n189745 , n189746 , n189747 , n22471 , 
 n189749 , n189750 , n22474 , n189752 , n189753 , n22477 , n189755 , n189756 , n22480 , n22481 , 
 n22482 , n22483 , n22484 , n189762 , n22486 , n189764 , n189765 , n22489 , n22490 , n22491 , 
 n22492 , n22493 , n189771 , n189772 , n22496 , n189774 , n189775 , n22499 , n189777 , n189778 , 
 n22502 , n189780 , n189781 , n22505 , n22506 , n189784 , n22508 , n22509 , n189787 , n189788 , 
 n22512 , n189790 , n22514 , n22515 , n189793 , n22517 , n22518 , n189796 , n189797 , n22521 , 
 n189799 , n22523 , n189801 , n189802 , n22526 , n189804 , n22528 , n189806 , n189807 , n22531 , 
 n189809 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , 
 n22542 , n22543 , n189821 , n22545 , n189823 , n189824 , n22548 , n189826 , n189827 , n189828 , 
 n22552 , n189830 , n22554 , n189832 , n189833 , n22557 , n189835 , n22559 , n189837 , n22561 , 
 n189839 , n189840 , n189841 , n22565 , n189843 , n22567 , n22568 , n189846 , n189847 , n22571 , 
 n22572 , n189850 , n189851 , n22575 , n189853 , n189854 , n22578 , n22579 , n189857 , n189858 , 
 n22582 , n22583 , n22584 , n22585 , n189863 , n22587 , n189865 , n22589 , n22590 , n22591 , 
 n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , 
 n22602 , n22603 , n22604 , n22605 , n22606 , n189884 , n22608 , n189886 , n22610 , n22611 , 
 n189889 , n189890 , n22614 , n189892 , n189893 , n22617 , n189895 , n22619 , n189897 , n189898 , 
 n22622 , n189900 , n189901 , n22625 , n189903 , n22627 , n22628 , n189906 , n189907 , n22631 , 
 n189909 , n189910 , n22634 , n189912 , n22636 , n22637 , n189915 , n189916 , n22640 , n189918 , 
 n189919 , n22643 , n189921 , n189922 , n22646 , n189924 , n22648 , n22649 , n189927 , n189928 , 
 n22652 , n189930 , n189931 , n22655 , n189933 , n189934 , n22658 , n189936 , n22660 , n189938 , 
 n189939 , n22663 , n189941 , n189942 , n22666 , n189944 , n22668 , n22669 , n189947 , n189948 , 
 n22672 , n189950 , n189951 , n22675 , n189953 , n22677 , n189955 , n189956 , n22680 , n189958 , 
 n22682 , n22683 , n189961 , n189962 , n22686 , n189964 , n189965 , n189966 , n22690 , n189968 , 
 n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , 
 n189979 , n189980 , n22704 , n189982 , n189983 , n22707 , n189985 , n22709 , n22710 , n189988 , 
 n189989 , n22713 , n189991 , n189992 , n22716 , n189994 , n22718 , n189996 , n189997 , n22721 , 
 n189999 , n190000 , n22724 , n190002 , n22726 , n22727 , n190005 , n190006 , n22730 , n190008 , 
 n190009 , n22733 , n190011 , n22735 , n22736 , n190014 , n190015 , n22739 , n190017 , n190018 , 
 n22742 , n190020 , n190021 , n22745 , n190023 , n22747 , n22748 , n190026 , n190027 , n22751 , 
 n190029 , n190030 , n22754 , n190032 , n190033 , n22757 , n190035 , n22759 , n22760 , n22761 , 
 n22762 , n22763 , n22764 , n22765 , n190043 , n22767 , n22768 , n190046 , n22770 , n22771 , 
 n22772 , n190050 , n22774 , n22775 , n22776 , n190054 , n190055 , n22779 , n22780 , n190058 , 
 n22782 , n22783 , n22784 , n190062 , n190063 , n190064 , n190065 , n22789 , n190067 , n22791 , 
 n190069 , n190070 , n190071 , n190072 , n22796 , n190074 , n190075 , n190076 , n22800 , n190078 , 
 n190079 , n190080 , n190081 , n22805 , n190083 , n190084 , n22808 , n22809 , n190087 , n22811 , 
 n22812 , n190090 , n190091 , n22815 , n190093 , n190094 , n22818 , n190096 , n190097 , n22821 , 
 n190099 , n190100 , n190101 , n190102 , n22826 , n190104 , n190105 , n22829 , n190107 , n22831 , 
 n22832 , n190110 , n190111 , n22835 , n190113 , n190114 , n22838 , n190116 , n190117 , n22841 , 
 n190119 , n190120 , n22844 , n190122 , n22846 , n22847 , n22848 , n190126 , n22850 , n190128 , 
 n190129 , n190130 , n22854 , n190132 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , 
 n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , 
 n190149 , n190150 , n22874 , n190152 , n190153 , n190154 , n22878 , n190156 , n22880 , n22881 , 
 n22882 , n22883 , n190161 , n22885 , n22886 , n22887 , n190165 , n190166 , n22890 , n22891 , 
 n190169 , n190170 , n22894 , n190172 , n190173 , n22897 , n190175 , n190176 , n190177 , n22901 , 
 n190179 , n190180 , n22904 , n22905 , n22906 , n190184 , n190185 , n22909 , n22910 , n22911 , 
 n22912 , n22913 , n190191 , n22915 , n22916 , n22917 , n22918 , n190196 , n190197 , n190198 , 
 n22922 , n190200 , n190201 , n22925 , n190203 , n190204 , n190205 , n22929 , n190207 , n22931 , 
 n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n190217 , n190218 , 
 n22942 , n190220 , n190221 , n22945 , n190223 , n22947 , n22948 , n22949 , n190227 , n190228 , 
 n22952 , n190230 , n190231 , n22955 , n190233 , n190234 , n22958 , n22959 , n190237 , n190238 , 
 n22962 , n22963 , n190241 , n22965 , n190243 , n22967 , n22968 , n190246 , n22970 , n190248 , 
 n190249 , n190250 , n22974 , n190252 , n190253 , n22977 , n190255 , n22979 , n22980 , n22981 , 
 n190259 , n190260 , n22984 , n190262 , n22986 , n190264 , n22988 , n190266 , n190267 , n22991 , 
 n190269 , n22993 , n22994 , n22995 , n190273 , n22997 , n190275 , n22999 , n23000 , n190278 , 
 n190279 , n23003 , n23004 , n190282 , n23006 , n23007 , n190285 , n23009 , n23010 , n190288 , 
 n23012 , n190290 , n190291 , n23015 , n190293 , n190294 , n23018 , n190296 , n23020 , n23021 , 
 n190299 , n190300 , n23024 , n23025 , n190303 , n190304 , n23028 , n190306 , n190307 , n23031 , 
 n23032 , n23033 , n190311 , n190312 , n23036 , n23037 , n23038 , n190316 , n190317 , n23041 , 
 n23042 , n23043 , n190321 , n190322 , n23046 , n190324 , n23048 , n190326 , n190327 , n23051 , 
 n190329 , n190330 , n23054 , n190332 , n23056 , n190334 , n190335 , n23059 , n190337 , n190338 , 
 n23062 , n23063 , n190341 , n190342 , n190343 , n23067 , n190345 , n190346 , n23070 , n190348 , 
 n190349 , n23073 , n190351 , n190352 , n190353 , n23077 , n190355 , n190356 , n23080 , n190358 , 
 n23082 , n23083 , n190361 , n190362 , n23086 , n190364 , n190365 , n190366 , n23090 , n190368 , 
 n190369 , n23093 , n190371 , n23095 , n190373 , n190374 , n23098 , n190376 , n190377 , n23101 , 
 n190379 , n23103 , n23104 , n190382 , n190383 , n190384 , n23108 , n190386 , n190387 , n23111 , 
 n190389 , n190390 , n23114 , n190392 , n23116 , n190394 , n190395 , n190396 , n23120 , n190398 , 
 n190399 , n23123 , n190401 , n23125 , n23126 , n23127 , n190405 , n190406 , n23130 , n190408 , 
 n190409 , n23133 , n190411 , n190412 , n190413 , n190414 , n23138 , n190416 , n190417 , n23141 , 
 n190419 , n190420 , n23144 , n23145 , n190423 , n190424 , n23148 , n190426 , n190427 , n23151 , 
 n190429 , n23153 , n23154 , n23155 , n23156 , n23157 , n190435 , n23159 , n190437 , n190438 , 
 n23162 , n23163 , n190441 , n23165 , n190443 , n23167 , n23168 , n190446 , n190447 , n23171 , 
 n190449 , n190450 , n23174 , n190452 , n23176 , n190454 , n190455 , n23179 , n23180 , n190458 , 
 n190459 , n190460 , n23184 , n190462 , n190463 , n23187 , n190465 , n190466 , n23190 , n190468 , 
 n190469 , n23193 , n190471 , n190472 , n23196 , n190474 , n190475 , n23199 , n190477 , n190478 , 
 n23202 , n190480 , n190481 , n23205 , n190483 , n23207 , n190485 , n190486 , n23210 , n23211 , 
 n190489 , n23213 , n190491 , n190492 , n190493 , n190494 , n23218 , n190496 , n190497 , n23221 , 
 n190499 , n190500 , n23224 , n190502 , n190503 , n23227 , n190505 , n190506 , n23230 , n190508 , 
 n23232 , n190510 , n190511 , n190512 , n190513 , n23237 , n190515 , n190516 , n190517 , n23241 , 
 n190519 , n190520 , n23244 , n23245 , n190523 , n190524 , n23248 , n23249 , n190527 , n190528 , 
 n23252 , n23253 , n23254 , n190532 , n190533 , n23257 , n190535 , n23259 , n190537 , n23261 , 
 n190539 , n190540 , n190541 , n23265 , n190543 , n190544 , n23268 , n190546 , n23270 , n190548 , 
 n190549 , n23273 , n190551 , n190552 , n190553 , n190554 , n23278 , n190556 , n190557 , n23281 , 
 n190559 , n23283 , n23284 , n190562 , n190563 , n190564 , n23288 , n190566 , n190567 , n23291 , 
 n190569 , n190570 , n23294 , n190572 , n190573 , n23297 , n190575 , n23299 , n190577 , n23301 , 
 n23302 , n190580 , n190581 , n190582 , n23306 , n190584 , n190585 , n23309 , n190587 , n190588 , 
 n23312 , n190590 , n190591 , n23315 , n190593 , n190594 , n23318 , n190596 , n23320 , n23321 , 
 n190599 , n23323 , n23324 , n190602 , n190603 , n23327 , n190605 , n190606 , n23330 , n190608 , 
 n190609 , n190610 , n23334 , n190612 , n23336 , n23337 , n190615 , n190616 , n23340 , n190618 , 
 n190619 , n23343 , n190621 , n190622 , n23346 , n23347 , n190625 , n23349 , n190627 , n23351 , 
 n23352 , n23353 , n190631 , n190632 , n23356 , n190634 , n190635 , n23359 , n190637 , n190638 , 
 n23362 , n23363 , n23364 , n190642 , n190643 , n23367 , n190645 , n190646 , n23370 , n190648 , 
 n23372 , n190650 , n190651 , n23375 , n190653 , n190654 , n190655 , n23379 , n190657 , n23381 , 
 n23382 , n190660 , n190661 , n190662 , n23386 , n190664 , n190665 , n23389 , n190667 , n190668 , 
 n23392 , n190670 , n190671 , n23395 , n190673 , n23397 , n190675 , n23399 , n23400 , n190678 , 
 n190679 , n23403 , n190681 , n190682 , n23406 , n190684 , n190685 , n23409 , n190687 , n190688 , 
 n23412 , n190690 , n190691 , n23415 , n23416 , n23417 , n23418 , n190696 , n190697 , n23421 , 
 n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n190707 , n23431 , 
 n23432 , n23433 , n190711 , n23435 , n23436 , n23437 , n23438 , n190716 , n23440 , n23441 , 
 n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n190727 , n23451 , 
 n190729 , n23453 , n23454 , n190732 , n190733 , n190734 , n23458 , n190736 , n190737 , n23461 , 
 n190739 , n190740 , n23464 , n190742 , n190743 , n190744 , n23468 , n190746 , n23470 , n23471 , 
 n190749 , n190750 , n23474 , n190752 , n190753 , n190754 , n23478 , n190756 , n190757 , n23481 , 
 n190759 , n190760 , n190761 , n23485 , n190763 , n23487 , n23488 , n23489 , n23490 , n23491 , 
 n23492 , n23493 , n190771 , n23495 , n190773 , n190774 , n23498 , n23499 , n190777 , n23501 , 
 n190779 , n190780 , n23504 , n23505 , n190783 , n190784 , n23508 , n190786 , n23510 , n190788 , 
 n190789 , n23513 , n190791 , n23515 , n190793 , n190794 , n23518 , n190796 , n23520 , n23521 , 
 n190799 , n190800 , n23524 , n190802 , n23526 , n190804 , n190805 , n23529 , n190807 , n190808 , 
 n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n190816 , n23540 , n23541 , 
 n23542 , n190820 , n190821 , n190822 , n23546 , n190824 , n190825 , n23549 , n190827 , n23551 , 
 n190829 , n23553 , n190831 , n23555 , n190833 , n23557 , n23558 , n190836 , n190837 , n190838 , 
 n23562 , n190840 , n190841 , n23565 , n190843 , n190844 , n23568 , n190846 , n190847 , n23571 , 
 n23572 , n23573 , n190851 , n190852 , n23576 , n190854 , n23578 , n23579 , n23580 , n23581 , 
 n190859 , n23583 , n190861 , n23585 , n190863 , n23587 , n23588 , n23589 , n23590 , n190868 , 
 n23592 , n190870 , n23594 , n190872 , n23596 , n23597 , n23598 , n190876 , n190877 , n23601 , 
 n190879 , n23603 , n23604 , n190882 , n190883 , n23607 , n190885 , n23609 , n23610 , n23611 , 
 n23612 , n23613 , n23614 , n190892 , n23616 , n190894 , n23618 , n23619 , n23620 , n23621 , 
 n190899 , n23623 , n190901 , n190902 , n190903 , n23627 , n190905 , n23629 , n23630 , n23631 , 
 n23632 , n190910 , n23634 , n190912 , n190913 , n23637 , n190915 , n23639 , n190917 , n23641 , 
 n23642 , n190920 , n23644 , n190922 , n23646 , n190924 , n190925 , n23649 , n190927 , n190928 , 
 n23652 , n23653 , n23654 , n190932 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , 
 n190939 , n23663 , n190941 , n23665 , n23666 , n190944 , n190945 , n190946 , n23670 , n190948 , 
 n190949 , n23673 , n190951 , n190952 , n23676 , n190954 , n190955 , n23679 , n190957 , n23681 , 
 n23682 , n190960 , n190961 , n190962 , n23686 , n190964 , n190965 , n23689 , n190967 , n190968 , 
 n23692 , n190970 , n23694 , n23695 , n23696 , n23697 , n23698 , n190976 , n190977 , n190978 , 
 n23702 , n190980 , n190981 , n23705 , n190983 , n23707 , n23708 , n23709 , n23710 , n23711 , 
 n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , 
 n190999 , n191000 , n23724 , n23725 , n23726 , n23727 , n191005 , n191006 , n23730 , n191008 , 
 n23732 , n191010 , n23734 , n23735 , n191013 , n23737 , n191015 , n191016 , n191017 , n191018 , 
 n23742 , n191020 , n191021 , n23745 , n191023 , n191024 , n23748 , n191026 , n191027 , n23751 , 
 n23752 , n23753 , n23754 , n191032 , n191033 , n23757 , n23758 , n191036 , n191037 , n23761 , 
 n23762 , n191040 , n23764 , n191042 , n191043 , n23767 , n23768 , n191046 , n191047 , n23771 , 
 n23772 , n23773 , n191051 , n23775 , n23776 , n23777 , n191055 , n23779 , n191057 , n23781 , 
 n23782 , n191060 , n23784 , n191062 , n191063 , n191064 , n23788 , n191066 , n23790 , n191068 , 
 n191069 , n23793 , n191071 , n191072 , n23796 , n23797 , n191075 , n23799 , n23800 , n191078 , 
 n191079 , n23803 , n23804 , n23805 , n191083 , n191084 , n23808 , n191086 , n191087 , n23811 , 
 n23812 , n23813 , n23814 , n23815 , n191093 , n191094 , n23818 , n23819 , n23820 , n191098 , 
 n23822 , n23823 , n23824 , n23825 , n191103 , n191104 , n191105 , n191106 , n23830 , n191108 , 
 n191109 , n191110 , n23834 , n191112 , n23836 , n23837 , n191115 , n191116 , n191117 , n23841 , 
 n191119 , n191120 , n23844 , n191122 , n191123 , n23847 , n191125 , n191126 , n23850 , n191128 , 
 n23852 , n191130 , n23854 , n23855 , n191133 , n191134 , n191135 , n23859 , n191137 , n191138 , 
 n23862 , n191140 , n191141 , n23865 , n191143 , n191144 , n23868 , n191146 , n191147 , n23871 , 
 n191149 , n23873 , n23874 , n23875 , n23876 , n191154 , n191155 , n191156 , n23880 , n191158 , 
 n191159 , n23883 , n191161 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , 
 n23892 , n23893 , n191171 , n191172 , n191173 , n23897 , n191175 , n191176 , n23900 , n191178 , 
 n23902 , n23903 , n23904 , n191182 , n23906 , n191184 , n23908 , n23909 , n191187 , n191188 , 
 n191189 , n23913 , n191191 , n191192 , n23916 , n191194 , n191195 , n23919 , n191197 , n191198 , 
 n23922 , n191200 , n191201 , n23925 , n191203 , n191204 , n23928 , n23929 , n191207 , n191208 , 
 n191209 , n23933 , n191211 , n191212 , n23936 , n191214 , n191215 , n23939 , n191217 , n23941 , 
 n191219 , n191220 , n23944 , n191222 , n23946 , n23947 , n191225 , n23949 , n191227 , n191228 , 
 n191229 , n191230 , n23954 , n191232 , n191233 , n23957 , n191235 , n191236 , n23960 , n191238 , 
 n191239 , n23963 , n191241 , n23965 , n191243 , n23967 , n23968 , n23969 , n23970 , n23971 , 
 n191249 , n191250 , n191251 , n23975 , n191253 , n23977 , n23978 , n191256 , n191257 , n191258 , 
 n23982 , n191260 , n191261 , n23985 , n191263 , n191264 , n23988 , n191266 , n191267 , n23991 , 
 n191269 , n23993 , n23994 , n191272 , n191273 , n191274 , n23998 , n191276 , n191277 , n24001 , 
 n191279 , n191280 , n24004 , n191282 , n24006 , n191284 , n24008 , n191286 , n24010 , n24011 , 
 n191289 , n191290 , n191291 , n24015 , n191293 , n191294 , n24018 , n191296 , n191297 , n24021 , 
 n191299 , n24023 , n191301 , n24025 , n24026 , n24027 , n24028 , n24029 , n191307 , n191308 , 
 n24032 , n191310 , n191311 , n24035 , n191313 , n24037 , n24038 , n24039 , n191317 , n191318 , 
 n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n191327 , n24051 , 
 n24052 , n24053 , n191331 , n191332 , n24056 , n24057 , n24058 , n191336 , n24060 , n24061 , 
 n24062 , n24063 , n24064 , n24065 , n191343 , n24067 , n24068 , n24069 , n24070 , n24071 , 
 n191349 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n191357 , n191358 , 
 n24082 , n191360 , n24084 , n191362 , n191363 , n191364 , n191365 , n24089 , n191367 , n24091 , 
 n24092 , n191370 , n24094 , n191372 , n191373 , n24097 , n191375 , n191376 , n24100 , n191378 , 
 n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n191386 , n24110 , n24111 , 
 n24112 , n24113 , n24114 , n24115 , n191393 , n24117 , n24118 , n191396 , n191397 , n24121 , 
 n24122 , n191400 , n191401 , n24125 , n24126 , n191404 , n191405 , n191406 , n191407 , n24131 , 
 n191409 , n191410 , n24134 , n191412 , n24136 , n24137 , n191415 , n191416 , n24140 , n191418 , 
 n191419 , n24143 , n191421 , n24145 , n191423 , n191424 , n24148 , n191426 , n24150 , n24151 , 
 n191429 , n191430 , n24154 , n191432 , n191433 , n191434 , n24158 , n191436 , n191437 , n24161 , 
 n191439 , n24163 , n24164 , n191442 , n191443 , n24167 , n191445 , n191446 , n24170 , n191448 , 
 n191449 , n24173 , n191451 , n24175 , n24176 , n24177 , n191455 , n24179 , n191457 , n191458 , 
 n24182 , n191460 , n191461 , n24185 , n191463 , n24187 , n24188 , n24189 , n191467 , n24191 , 
 n191469 , n191470 , n191471 , n191472 , n24196 , n191474 , n191475 , n24199 , n191477 , n24201 , 
 n24202 , n191480 , n191481 , n24205 , n191483 , n191484 , n24208 , n191486 , n191487 , n24211 , 
 n191489 , n191490 , n24214 , n191492 , n191493 , n24217 , n191495 , n24219 , n24220 , n191498 , 
 n191499 , n24223 , n191501 , n191502 , n24226 , n191504 , n191505 , n24229 , n24230 , n24231 , 
 n191509 , n191510 , n24234 , n191512 , n191513 , n24237 , n24238 , n191516 , n191517 , n24241 , 
 n191519 , n191520 , n24244 , n191522 , n24246 , n24247 , n191525 , n191526 , n24250 , n191528 , 
 n191529 , n24253 , n191531 , n24255 , n191533 , n191534 , n24258 , n191536 , n24260 , n24261 , 
 n24262 , n191540 , n191541 , n24265 , n191543 , n24267 , n24268 , n24269 , n191547 , n191548 , 
 n24272 , n191550 , n191551 , n191552 , n191553 , n24277 , n191555 , n191556 , n24280 , n191558 , 
 n191559 , n24283 , n24284 , n191562 , n24286 , n24287 , n24288 , n191566 , n24290 , n191568 , 
 n191569 , n191570 , n191571 , n24295 , n191573 , n191574 , n24298 , n191576 , n191577 , n24301 , 
 n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , 
 n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n191597 , n191598 , 
 n24322 , n191600 , n24324 , n191602 , n191603 , n24327 , n191605 , n191606 , n191607 , n24331 , 
 n191609 , n24333 , n24334 , n24335 , n191613 , n24337 , n24338 , n24339 , n191617 , n191618 , 
 n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n191627 , n24351 , 
 n191629 , n24353 , n24354 , n191632 , n191633 , n191634 , n24358 , n191636 , n24360 , n24361 , 
 n24362 , n191640 , n191641 , n24365 , n191643 , n24367 , n24368 , n191646 , n191647 , n24371 , 
 n191649 , n191650 , n24374 , n191652 , n24376 , n24377 , n191655 , n191656 , n24380 , n191658 , 
 n191659 , n24383 , n191661 , n24385 , n24386 , n24387 , n191665 , n191666 , n24390 , n191668 , 
 n191669 , n24393 , n191671 , n24395 , n24396 , n191674 , n191675 , n24399 , n191677 , n191678 , 
 n24402 , n191680 , n24404 , n24405 , n191683 , n191684 , n24408 , n191686 , n191687 , n24411 , 
 n191689 , n24413 , n24414 , n191692 , n191693 , n24417 , n191695 , n191696 , n24420 , n191698 , 
 n191699 , n24423 , n191701 , n191702 , n24426 , n191704 , n191705 , n24429 , n191707 , n24431 , 
 n24432 , n191710 , n191711 , n24435 , n191713 , n191714 , n24438 , n191716 , n191717 , n24441 , 
 n24442 , n24443 , n191721 , n191722 , n24446 , n191724 , n24448 , n24449 , n24450 , n191728 , 
 n191729 , n24453 , n191731 , n24455 , n24456 , n191734 , n24458 , n191736 , n24460 , n24461 , 
 n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n191745 , n24469 , n24470 , n24471 , 
 n191749 , n24473 , n24474 , n24475 , n191753 , n191754 , n24478 , n24479 , n24480 , n191758 , 
 n191759 , n24483 , n24484 , n191762 , n191763 , n24487 , n24488 , n191766 , n191767 , n24491 , 
 n24492 , n24493 , n191771 , n24495 , n24496 , n191774 , n191775 , n191776 , n24500 , n191778 , 
 n24502 , n24503 , n24504 , n191782 , n191783 , n24507 , n191785 , n24509 , n191787 , n191788 , 
 n191789 , n24513 , n191791 , n24515 , n191793 , n191794 , n191795 , n24519 , n191797 , n24521 , 
 n191799 , n24523 , n191801 , n24525 , n24526 , n24527 , n24528 , n191806 , n191807 , n24531 , 
 n191809 , n24533 , n24534 , n191812 , n24536 , n191814 , n24538 , n191816 , n191817 , n24541 , 
 n191819 , n191820 , n24544 , n191822 , n24546 , n24547 , n191825 , n191826 , n24550 , n191828 , 
 n191829 , n24553 , n191831 , n191832 , n24556 , n191834 , n24558 , n24559 , n191837 , n191838 , 
 n24562 , n191840 , n191841 , n24565 , n191843 , n24567 , n24568 , n191846 , n191847 , n24571 , 
 n191849 , n191850 , n24574 , n191852 , n24576 , n191854 , n191855 , n24579 , n191857 , n24581 , 
 n24582 , n191860 , n191861 , n24585 , n191863 , n191864 , n24588 , n191866 , n24590 , n24591 , 
 n191869 , n191870 , n24594 , n191872 , n191873 , n24597 , n191875 , n24599 , n191877 , n191878 , 
 n24602 , n191880 , n191881 , n24605 , n191883 , n24607 , n24608 , n191886 , n191887 , n24611 , 
 n191889 , n191890 , n24614 , n191892 , n24616 , n24617 , n191895 , n191896 , n24620 , n191898 , 
 n191899 , n191900 , n191901 , n24625 , n191903 , n191904 , n24628 , n191906 , n191907 , n24631 , 
 n24632 , n191910 , n24634 , n24635 , n24636 , n24637 , n24638 , n191916 , n24640 , n191918 , 
 n191919 , n24643 , n191921 , n191922 , n191923 , n24647 , n191925 , n24649 , n191927 , n191928 , 
 n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , 
 n24662 , n191940 , n24664 , n24665 , n191943 , n191944 , n24668 , n191946 , n24670 , n191948 , 
 n191949 , n24673 , n191951 , n191952 , n191953 , n24677 , n191955 , n24679 , n191957 , n191958 , 
 n24682 , n191960 , n191961 , n24685 , n191963 , n191964 , n24688 , n24689 , n24690 , n191968 , 
 n191969 , n24693 , n24694 , n24695 , n24696 , n191974 , n24698 , n191976 , n24700 , n191978 , 
 n24702 , n24703 , n24704 , n24705 , n24706 , n191984 , n24708 , n191986 , n191987 , n24711 , 
 n191989 , n24713 , n191991 , n191992 , n24716 , n24717 , n191995 , n191996 , n24720 , n191998 , 
 n191999 , n24723 , n192001 , n24725 , n24726 , n192004 , n192005 , n24729 , n192007 , n192008 , 
 n24732 , n192010 , n192011 , n192012 , n192013 , n24737 , n192015 , n192016 , n24740 , n192018 , 
 n24742 , n24743 , n192021 , n192022 , n24746 , n192024 , n192025 , n24749 , n192027 , n192028 , 
 n24752 , n24753 , n192031 , n24755 , n192033 , n24757 , n24758 , n192036 , n192037 , n24761 , 
 n192039 , n192040 , n24764 , n192042 , n192043 , n24767 , n24768 , n24769 , n192047 , n192048 , 
 n192049 , n192050 , n24774 , n192052 , n192053 , n24777 , n192055 , n24779 , n24780 , n192058 , 
 n192059 , n24783 , n192061 , n192062 , n24786 , n192064 , n192065 , n24789 , n192067 , n192068 , 
 n24792 , n192070 , n192071 , n24795 , n192073 , n24797 , n24798 , n192076 , n192077 , n24801 , 
 n192079 , n192080 , n24804 , n192082 , n192083 , n24807 , n24808 , n192086 , n192087 , n24811 , 
 n192089 , n192090 , n24814 , n192092 , n192093 , n24817 , n192095 , n24819 , n24820 , n192098 , 
 n192099 , n24823 , n192101 , n192102 , n24826 , n192104 , n192105 , n24829 , n192107 , n192108 , 
 n24832 , n192110 , n192111 , n24835 , n24836 , n24837 , n192115 , n192116 , n24840 , n24841 , 
 n24842 , n192120 , n192121 , n24845 , n192123 , n192124 , n192125 , n24849 , n192127 , n24851 , 
 n192129 , n192130 , n24854 , n192132 , n192133 , n24857 , n192135 , n192136 , n24860 , n24861 , 
 n24862 , n192140 , n192141 , n24865 , n24866 , n24867 , n192145 , n192146 , n24870 , n24871 , 
 n24872 , n192150 , n24874 , n24875 , n192153 , n192154 , n24878 , n24879 , n24880 , n192158 , 
 n192159 , n24883 , n192161 , n192162 , n24886 , n192164 , n24888 , n192166 , n192167 , n24891 , 
 n192169 , n192170 , n24894 , n192172 , n24896 , n24897 , n192175 , n192176 , n192177 , n24901 , 
 n192179 , n192180 , n24904 , n192182 , n192183 , n24907 , n192185 , n192186 , n192187 , n24911 , 
 n192189 , n192190 , n24914 , n192192 , n24916 , n24917 , n192195 , n192196 , n192197 , n24921 , 
 n192199 , n192200 , n24924 , n192202 , n192203 , n24927 , n192205 , n24929 , n192207 , n192208 , 
 n24932 , n192210 , n192211 , n24935 , n192213 , n24937 , n24938 , n192216 , n192217 , n192218 , 
 n24942 , n192220 , n192221 , n24945 , n192223 , n192224 , n24948 , n192226 , n24950 , n24951 , 
 n24952 , n24953 , n24954 , n192232 , n192233 , n24957 , n192235 , n192236 , n24960 , n192238 , 
 n24962 , n24963 , n192241 , n192242 , n192243 , n24967 , n192245 , n192246 , n24970 , n192248 , 
 n192249 , n24973 , n192251 , n192252 , n192253 , n192254 , n24978 , n192256 , n192257 , n24981 , 
 n192259 , n24983 , n24984 , n192262 , n192263 , n192264 , n24988 , n192266 , n192267 , n24991 , 
 n192269 , n192270 , n24994 , n192272 , n192273 , n24997 , n192275 , n192276 , n25000 , n192278 , 
 n192279 , n25003 , n192281 , n25005 , n25006 , n192284 , n192285 , n192286 , n25010 , n192288 , 
 n192289 , n25013 , n192291 , n192292 , n25016 , n192294 , n192295 , n25019 , n192297 , n25021 , 
 n25022 , n25023 , n25024 , n192302 , n25026 , n192304 , n25028 , n25029 , n25030 , n192308 , 
 n192309 , n25033 , n192311 , n25035 , n25036 , n25037 , n192315 , n192316 , n192317 , n25041 , 
 n192319 , n192320 , n25044 , n192322 , n25046 , n25047 , n192325 , n192326 , n25050 , n192328 , 
 n25052 , n192330 , n25054 , n192332 , n25056 , n25057 , n192335 , n192336 , n192337 , n25061 , 
 n192339 , n192340 , n25064 , n192342 , n25066 , n25067 , n25068 , n192346 , n192347 , n25071 , 
 n192349 , n192350 , n192351 , n192352 , n25076 , n192354 , n192355 , n25079 , n192357 , n25081 , 
 n25082 , n192360 , n192361 , n192362 , n25086 , n192364 , n192365 , n25089 , n192367 , n192368 , 
 n25092 , n192370 , n192371 , n25095 , n192373 , n192374 , n25098 , n192376 , n192377 , n25101 , 
 n192379 , n25103 , n25104 , n192382 , n192383 , n192384 , n25108 , n192386 , n192387 , n25111 , 
 n192389 , n192390 , n25114 , n192392 , n192393 , n25117 , n192395 , n192396 , n25120 , n192398 , 
 n25122 , n192400 , n25124 , n25125 , n192403 , n192404 , n192405 , n25129 , n192407 , n192408 , 
 n25132 , n192410 , n192411 , n25135 , n192413 , n192414 , n192415 , n192416 , n25140 , n192418 , 
 n192419 , n25143 , n192421 , n25145 , n25146 , n192424 , n192425 , n25149 , n192427 , n192428 , 
 n25152 , n192430 , n192431 , n25155 , n192433 , n192434 , n25158 , n192436 , n192437 , n25161 , 
 n192439 , n25163 , n25164 , n192442 , n192443 , n25167 , n192445 , n192446 , n25170 , n192448 , 
 n25172 , n192450 , n192451 , n25175 , n192453 , n192454 , n25178 , n192456 , n25180 , n25181 , 
 n192459 , n192460 , n25184 , n192462 , n192463 , n25187 , n192465 , n25189 , n25190 , n192468 , 
 n192469 , n25193 , n192471 , n192472 , n192473 , n25197 , n192475 , n192476 , n25200 , n192478 , 
 n25202 , n25203 , n192481 , n192482 , n25206 , n192484 , n192485 , n25209 , n192487 , n192488 , 
 n25212 , n192490 , n25214 , n25215 , n192493 , n25217 , n192495 , n192496 , n25220 , n192498 , 
 n25222 , n192500 , n25224 , n25225 , n192503 , n25227 , n192505 , n192506 , n25230 , n192508 , 
 n192509 , n192510 , n192511 , n25235 , n192513 , n192514 , n25238 , n192516 , n25240 , n25241 , 
 n192519 , n192520 , n25244 , n192522 , n192523 , n25247 , n192525 , n192526 , n25250 , n192528 , 
 n192529 , n25253 , n192531 , n192532 , n25256 , n192534 , n25258 , n25259 , n192537 , n192538 , 
 n192539 , n25263 , n192541 , n192542 , n25266 , n192544 , n192545 , n25269 , n192547 , n192548 , 
 n25272 , n25273 , n192551 , n25275 , n192553 , n192554 , n25278 , n192556 , n25280 , n192558 , 
 n192559 , n25283 , n25284 , n192562 , n192563 , n25287 , n192565 , n192566 , n25290 , n192568 , 
 n25292 , n25293 , n192571 , n25295 , n192573 , n192574 , n192575 , n25299 , n192577 , n192578 , 
 n25302 , n192580 , n192581 , n25305 , n192583 , n192584 , n25308 , n192586 , n192587 , n25311 , 
 n192589 , n192590 , n25314 , n192592 , n192593 , n25317 , n25318 , n192596 , n25320 , n25321 , 
 n192599 , n192600 , n192601 , n25325 , n192603 , n192604 , n25328 , n192606 , n192607 , n25331 , 
 n192609 , n192610 , n192611 , n192612 , n25336 , n192614 , n192615 , n25339 , n192617 , n25341 , 
 n25342 , n192620 , n25344 , n192622 , n25346 , n192624 , n192625 , n25349 , n192627 , n192628 , 
 n25352 , n192630 , n192631 , n25355 , n192633 , n192634 , n25358 , n192636 , n25360 , n25361 , 
 n192639 , n192640 , n192641 , n25365 , n192643 , n192644 , n25368 , n192646 , n192647 , n25371 , 
 n192649 , n192650 , n25374 , n25375 , n25376 , n192654 , n192655 , n25379 , n25380 , n25381 , 
 n192659 , n192660 , n25384 , n192662 , n25386 , n192664 , n192665 , n25389 , n192667 , n192668 , 
 n192669 , n192670 , n25394 , n192672 , n192673 , n25397 , n192675 , n25399 , n25400 , n192678 , 
 n192679 , n192680 , n25404 , n192682 , n192683 , n25407 , n192685 , n192686 , n25410 , n192688 , 
 n192689 , n25413 , n192691 , n25415 , n192693 , n25417 , n25418 , n192696 , n192697 , n192698 , 
 n25422 , n192700 , n192701 , n25425 , n192703 , n192704 , n25428 , n192706 , n192707 , n25431 , 
 n25432 , n25433 , n192711 , n192712 , n192713 , n25437 , n192715 , n25439 , n25440 , n192718 , 
 n192719 , n25443 , n192721 , n192722 , n25446 , n192724 , n192725 , n192726 , n25450 , n192728 , 
 n25452 , n25453 , n192731 , n192732 , n25456 , n192734 , n192735 , n25459 , n192737 , n192738 , 
 n25462 , n192740 , n25464 , n192742 , n25466 , n25467 , n192745 , n192746 , n25470 , n192748 , 
 n192749 , n25473 , n192751 , n192752 , n25476 , n192754 , n192755 , n192756 , n192757 , n25481 , 
 n192759 , n192760 , n25484 , n192762 , n192763 , n192764 , n192765 , n25489 , n192767 , n192768 , 
 n25492 , n25493 , n192771 , n192772 , n25496 , n192774 , n192775 , n25499 , n192777 , n25501 , 
 n192779 , n25503 , n25504 , n192782 , n192783 , n25507 , n192785 , n192786 , n192787 , n25511 , 
 n192789 , n192790 , n25514 , n192792 , n192793 , n25517 , n25518 , n25519 , n192797 , n25521 , 
 n192799 , n25523 , n25524 , n192802 , n25526 , n192804 , n25528 , n25529 , n192807 , n192808 , 
 n25532 , n192810 , n192811 , n25535 , n192813 , n192814 , n25538 , n192816 , n192817 , n25541 , 
 n192819 , n192820 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n192827 , n25551 , 
 n192829 , n192830 , n25554 , n192832 , n25556 , n192834 , n25558 , n25559 , n192837 , n192838 , 
 n192839 , n25563 , n192841 , n192842 , n25566 , n192844 , n192845 , n25569 , n192847 , n192848 , 
 n25572 , n192850 , n192851 , n25575 , n25576 , n192854 , n25578 , n192856 , n25580 , n25581 , 
 n192859 , n192860 , n192861 , n25585 , n192863 , n192864 , n25588 , n192866 , n192867 , n25591 , 
 n192869 , n192870 , n25594 , n192872 , n192873 , n192874 , n192875 , n25599 , n192877 , n192878 , 
 n25602 , n192880 , n192881 , n25605 , n25606 , n25607 , n192885 , n192886 , n25610 , n25611 , 
 n25612 , n192890 , n192891 , n25615 , n25616 , n25617 , n192895 , n25619 , n192897 , n192898 , 
 n25622 , n192900 , n25624 , n25625 , n192903 , n192904 , n25628 , n192906 , n192907 , n25631 , 
 n192909 , n192910 , n25634 , n192912 , n25636 , n192914 , n25638 , n25639 , n192917 , n192918 , 
 n25642 , n192920 , n192921 , n25645 , n192923 , n192924 , n25648 , n192926 , n192927 , n25651 , 
 n25652 , n192930 , n25654 , n192932 , n25656 , n192934 , n192935 , n25659 , n192937 , n192938 , 
 n192939 , n192940 , n25664 , n192942 , n192943 , n25667 , n192945 , n25669 , n25670 , n192948 , 
 n192949 , n192950 , n25674 , n192952 , n192953 , n25677 , n192955 , n192956 , n25680 , n192958 , 
 n192959 , n25683 , n192961 , n192962 , n25686 , n25687 , n192965 , n25689 , n25690 , n192968 , 
 n192969 , n25693 , n192971 , n25695 , n25696 , n25697 , n192975 , n25699 , n25700 , n192978 , 
 n192979 , n25703 , n25704 , n25705 , n192983 , n25707 , n192985 , n25709 , n192987 , n192988 , 
 n192989 , n25713 , n192991 , n192992 , n192993 , n25717 , n192995 , n25719 , n25720 , n192998 , 
 n192999 , n25723 , n193001 , n193002 , n25726 , n193004 , n193005 , n25729 , n193007 , n25731 , 
 n193009 , n25733 , n25734 , n193012 , n193013 , n25737 , n193015 , n193016 , n25740 , n193018 , 
 n193019 , n25743 , n25744 , n25745 , n193023 , n193024 , n25748 , n25749 , n193027 , n193028 , 
 n25752 , n25753 , n25754 , n193032 , n25756 , n193034 , n25758 , n25759 , n25760 , n193038 , 
 n193039 , n25763 , n193041 , n25765 , n25766 , n193044 , n193045 , n193046 , n25770 , n193048 , 
 n193049 , n25773 , n193051 , n193052 , n25776 , n193054 , n193055 , n25779 , n193057 , n25781 , 
 n193059 , n25783 , n25784 , n193062 , n193063 , n193064 , n25788 , n193066 , n193067 , n25791 , 
 n193069 , n193070 , n25794 , n193072 , n193073 , n25797 , n193075 , n193076 , n25800 , n25801 , 
 n25802 , n193080 , n193081 , n25805 , n193083 , n25807 , n193085 , n25809 , n25810 , n193088 , 
 n25812 , n193090 , n193091 , n193092 , n193093 , n25817 , n193095 , n193096 , n25820 , n193098 , 
 n193099 , n193100 , n193101 , n25825 , n193103 , n193104 , n193105 , n25829 , n193107 , n25831 , 
 n25832 , n193110 , n193111 , n25835 , n193113 , n193114 , n25838 , n193116 , n193117 , n25841 , 
 n193119 , n25843 , n193121 , n25845 , n25846 , n193124 , n193125 , n25849 , n193127 , n193128 , 
 n25852 , n193130 , n193131 , n25855 , n193133 , n193134 , n25858 , n25859 , n25860 , n25861 , 
 n25862 , n193140 , n193141 , n25865 , n193143 , n193144 , n25868 , n193146 , n193147 , n25871 , 
 n25872 , n193150 , n193151 , n25875 , n25876 , n25877 , n25878 , n193156 , n193157 , n25881 , 
 n25882 , n193160 , n193161 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , 
 n25892 , n25893 , n193171 , n25895 , n25896 , n25897 , n193175 , n193176 , n25900 , n25901 , 
 n25902 , n25903 , n193181 , n25905 , n25906 , n25907 , n193185 , n193186 , n25910 , n25911 , 
 n193189 , n193190 , n25914 , n193192 , n193193 , n25917 , n193195 , n193196 , n25920 , n25921 , 
 n193199 , n25923 , n25924 , n193202 , n193203 , n25927 , n25928 , n193206 , n25930 , n193208 , 
 n25932 , n193210 , n25934 , n25935 , n193213 , n193214 , n25938 , n193216 , n193217 , n25941 , 
 n193219 , n193220 , n193221 , n25945 , n193223 , n193224 , n25948 , n193226 , n193227 , n25951 , 
 n193229 , n25953 , n193231 , n193232 , n193233 , n193234 , n25958 , n193236 , n193237 , n25961 , 
 n193239 , n193240 , n25964 , n193242 , n193243 , n25967 , n25968 , n25969 , n193247 , n193248 , 
 n25972 , n25973 , n25974 , n25975 , n193253 , n193254 , n25978 , n25979 , n25980 , n25981 , 
 n25982 , n25983 , n25984 , n25985 , n193263 , n25987 , n25988 , n25989 , n25990 , n25991 , 
 n25992 , n25993 , n25994 , n25995 , n25996 , n193274 , n25998 , n25999 , n193277 , n193278 , 
 n26002 , n193280 , n26004 , n193282 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , 
 n26012 , n193290 , n26014 , n193292 , n193293 , n26017 , n26018 , n26019 , n193297 , n193298 , 
 n26022 , n26023 , n26024 , n26025 , n26026 , n193304 , n193305 , n26029 , n26030 , n26031 , 
 n26032 , n193310 , n193311 , n26035 , n26036 , n26037 , n193315 , n193316 , n26040 , n193318 , 
 n193319 , n26043 , n26044 , n26045 , n193323 , n193324 , n26048 , n26049 , n26050 , n193328 , 
 n193329 , n26053 , n26054 , n26055 , n26056 , n26057 , n193335 , n193336 , n26060 , n26061 , 
 n26062 , n26063 , n193341 , n193342 , n193343 , n26067 , n193345 , n26069 , n26070 , n193348 , 
 n193349 , n26073 , n193351 , n193352 , n26076 , n193354 , n193355 , n26079 , n193357 , n26081 , 
 n26082 , n193360 , n193361 , n26085 , n193363 , n193364 , n26088 , n193366 , n26090 , n193368 , 
 n26092 , n193370 , n26094 , n26095 , n193373 , n193374 , n26098 , n193376 , n193377 , n26101 , 
 n193379 , n26103 , n193381 , n26105 , n193383 , n26107 , n26108 , n193386 , n26110 , n193388 , 
 n193389 , n193390 , n26114 , n193392 , n26116 , n193394 , n26118 , n26119 , n26120 , n26121 , 
 n193399 , n193400 , n26124 , n193402 , n26126 , n193404 , n26128 , n26129 , n193407 , n193408 , 
 n26132 , n193410 , n193411 , n26135 , n193413 , n193414 , n26138 , n193416 , n26140 , n26141 , 
 n193419 , n193420 , n26144 , n193422 , n193423 , n26147 , n193425 , n26149 , n193427 , n26151 , 
 n193429 , n26153 , n26154 , n193432 , n193433 , n26157 , n193435 , n193436 , n26160 , n193438 , 
 n26162 , n26163 , n26164 , n193442 , n26166 , n193444 , n193445 , n26169 , n26170 , n193448 , 
 n193449 , n26173 , n193451 , n193452 , n26176 , n26177 , n26178 , n26179 , n26180 , n193458 , 
 n26182 , n26183 , n26184 , n193462 , n26186 , n26187 , n26188 , n193466 , n193467 , n26191 , 
 n193469 , n193470 , n26194 , n26195 , n26196 , n193474 , n26198 , n26199 , n193477 , n26201 , 
 n26202 , n26203 , n26204 , n26205 , n193483 , n26207 , n26208 , n26209 , n193487 , n26211 , 
 n193489 , n193490 , n26214 , n193492 , n26216 , n26217 , n26218 , n26219 , n26220 , n193498 , 
 n193499 , n26223 , n26224 , n26225 , n26226 , n193504 , n193505 , n26229 , n193507 , n26231 , 
 n26232 , n26233 , n26234 , n193512 , n193513 , n26237 , n26238 , n26239 , n26240 , n26241 , 
 n193519 , n193520 , n26244 , n193522 , n193523 , n26247 , n193525 , n193526 , n26250 , n26251 , 
 n26252 , n26253 , n193531 , n193532 , n193533 , n193534 , n26258 , n193536 , n193537 , n193538 , 
 n26262 , n193540 , n26264 , n26265 , n193543 , n193544 , n193545 , n26269 , n193547 , n193548 , 
 n26272 , n193550 , n193551 , n26275 , n193553 , n193554 , n26278 , n193556 , n26280 , n193558 , 
 n26282 , n26283 , n193561 , n193562 , n193563 , n26287 , n193565 , n193566 , n26290 , n193568 , 
 n193569 , n26293 , n193571 , n193572 , n26296 , n193574 , n193575 , n193576 , n26300 , n193578 , 
 n26302 , n26303 , n193581 , n193582 , n193583 , n26307 , n193585 , n193586 , n26310 , n193588 , 
 n193589 , n26313 , n193591 , n193592 , n193593 , n26317 , n193595 , n26319 , n26320 , n193598 , 
 n193599 , n193600 , n26324 , n193602 , n193603 , n26327 , n193605 , n193606 , n26330 , n193608 , 
 n193609 , n26333 , n193611 , n26335 , n193613 , n26337 , n26338 , n193616 , n193617 , n193618 , 
 n26342 , n193620 , n193621 , n26345 , n193623 , n193624 , n26348 , n193626 , n193627 , n26351 , 
 n193629 , n193630 , n26354 , n193632 , n26356 , n193634 , n26358 , n26359 , n193637 , n26361 , 
 n193639 , n26363 , n193641 , n193642 , n26366 , n193644 , n193645 , n26369 , n193647 , n26371 , 
 n26372 , n193650 , n26374 , n193652 , n26376 , n193654 , n193655 , n26379 , n193657 , n26381 , 
 n193659 , n193660 , n26384 , n193662 , n26386 , n193664 , n26388 , n193666 , n26390 , n193668 , 
 n193669 , n26393 , n26394 , n26395 , n26396 , n26397 , n193675 , n193676 , n26400 , n193678 , 
 n193679 , n26403 , n26404 , n26405 , n26406 , n26407 , n193685 , n193686 , n26410 , n193688 , 
 n26412 , n26413 , n26414 , n26415 , n26416 , n193694 , n26418 , n193696 , n193697 , n26421 , 
 n193699 , n26423 , n26424 , n26425 , n193703 , n193704 , n26428 , n193706 , n26430 , n26431 , 
 n193709 , n193710 , n26434 , n193712 , n193713 , n26437 , n193715 , n26439 , n26440 , n193718 , 
 n193719 , n193720 , n26444 , n193722 , n193723 , n26447 , n193725 , n193726 , n26450 , n193728 , 
 n26452 , n193730 , n193731 , n26455 , n193733 , n193734 , n26458 , n193736 , n26460 , n26461 , 
 n193739 , n193740 , n193741 , n26465 , n193743 , n193744 , n26468 , n193746 , n193747 , n26471 , 
 n193749 , n26473 , n193751 , n193752 , n26476 , n193754 , n193755 , n26479 , n193757 , n26481 , 
 n26482 , n193760 , n193761 , n193762 , n26486 , n193764 , n193765 , n26489 , n193767 , n193768 , 
 n26492 , n193770 , n26494 , n193772 , n193773 , n26497 , n193775 , n26499 , n26500 , n193778 , 
 n193779 , n26503 , n193781 , n193782 , n193783 , n26507 , n193785 , n26509 , n26510 , n26511 , 
 n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n193797 , n193798 , 
 n26522 , n193800 , n193801 , n26525 , n193803 , n26527 , n26528 , n193806 , n193807 , n193808 , 
 n26532 , n193810 , n193811 , n26535 , n193813 , n193814 , n26538 , n193816 , n193817 , n193818 , 
 n26542 , n193820 , n193821 , n26545 , n193823 , n26547 , n26548 , n193826 , n193827 , n193828 , 
 n26552 , n193830 , n193831 , n26555 , n193833 , n193834 , n26558 , n193836 , n26560 , n193838 , 
 n193839 , n26563 , n193841 , n193842 , n26566 , n26567 , n193845 , n26569 , n26570 , n26571 , 
 n193849 , n193850 , n193851 , n26575 , n193853 , n193854 , n26578 , n193856 , n193857 , n26581 , 
 n193859 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , 
 n26592 , n26593 , n26594 , n26595 , n193873 , n193874 , n193875 , n26599 , n193877 , n193878 , 
 n26602 , n193880 , n26604 , n26605 , n193883 , n193884 , n26608 , n193886 , n193887 , n193888 , 
 n26612 , n193890 , n193891 , n26615 , n193893 , n193894 , n193895 , n193896 , n26620 , n193898 , 
 n26622 , n193900 , n193901 , n193902 , n26626 , n193904 , n26628 , n193906 , n26630 , n193908 , 
 n193909 , n26633 , n193911 , n26635 , n193913 , n26637 , n26638 , n193916 , n193917 , n193918 , 
 n26642 , n193920 , n193921 , n26645 , n193923 , n193924 , n26648 , n193926 , n193927 , n26651 , 
 n26652 , n193930 , n26654 , n193932 , n26656 , n26657 , n193935 , n193936 , n193937 , n26661 , 
 n193939 , n193940 , n26664 , n193942 , n193943 , n26667 , n193945 , n193946 , n26670 , n26671 , 
 n26672 , n193950 , n193951 , n193952 , n26676 , n193954 , n26678 , n26679 , n193957 , n193958 , 
 n26682 , n193960 , n193961 , n26685 , n193963 , n193964 , n193965 , n193966 , n26690 , n193968 , 
 n26692 , n193970 , n193971 , n193972 , n193973 , n26697 , n193975 , n193976 , n193977 , n26701 , 
 n193979 , n193980 , n193981 , n193982 , n26706 , n193984 , n193985 , n26709 , n193987 , n26711 , 
 n26712 , n193990 , n193991 , n26715 , n193993 , n193994 , n26718 , n193996 , n193997 , n26721 , 
 n193999 , n194000 , n26724 , n194002 , n194003 , n26727 , n194005 , n194006 , n194007 , n26731 , 
 n194009 , n26733 , n26734 , n194012 , n194013 , n26737 , n194015 , n194016 , n26740 , n194018 , 
 n194019 , n26743 , n194021 , n194022 , n26746 , n194024 , n194025 , n26749 , n194027 , n26751 , 
 n26752 , n194030 , n194031 , n194032 , n26756 , n194034 , n194035 , n26759 , n194037 , n194038 , 
 n26762 , n194040 , n194041 , n26765 , n26766 , n26767 , n194045 , n194046 , n26770 , n194048 , 
 n194049 , n26773 , n26774 , n26775 , n194053 , n194054 , n194055 , n194056 , n26780 , n194058 , 
 n194059 , n26783 , n194061 , n26785 , n26786 , n194064 , n194065 , n194066 , n26790 , n194068 , 
 n194069 , n26793 , n194071 , n194072 , n26796 , n194074 , n194075 , n26799 , n194077 , n194078 , 
 n26802 , n194080 , n194081 , n26805 , n194083 , n26807 , n26808 , n194086 , n194087 , n194088 , 
 n26812 , n194090 , n194091 , n26815 , n194093 , n194094 , n26818 , n194096 , n194097 , n26821 , 
 n26822 , n194100 , n194101 , n26825 , n26826 , n194104 , n26828 , n194106 , n26830 , n26831 , 
 n194109 , n194110 , n26834 , n194112 , n194113 , n26837 , n194115 , n194116 , n26840 , n194118 , 
 n194119 , n26843 , n194121 , n194122 , n26846 , n26847 , n194125 , n26849 , n194127 , n26851 , 
 n26852 , n194130 , n194131 , n26855 , n194133 , n194134 , n26858 , n194136 , n194137 , n194138 , 
 n194139 , n26863 , n194141 , n194142 , n26866 , n194144 , n26868 , n26869 , n194147 , n26871 , 
 n194149 , n26873 , n194151 , n194152 , n26876 , n194154 , n194155 , n26879 , n26880 , n194158 , 
 n26882 , n194160 , n26884 , n26885 , n194163 , n194164 , n26888 , n194166 , n194167 , n26891 , 
 n194169 , n194170 , n26894 , n26895 , n26896 , n194174 , n194175 , n26899 , n26900 , n26901 , 
 n194179 , n194180 , n26904 , n26905 , n26906 , n194184 , n194185 , n26909 , n26910 , n26911 , 
 n26912 , n26913 , n194191 , n194192 , n26916 , n194194 , n194195 , n194196 , n194197 , n26921 , 
 n194199 , n194200 , n26924 , n194202 , n26926 , n26927 , n194205 , n194206 , n26930 , n194208 , 
 n194209 , n26933 , n194211 , n26935 , n26936 , n26937 , n194215 , n194216 , n26940 , n194218 , 
 n26942 , n26943 , n194221 , n194222 , n26946 , n194224 , n194225 , n26949 , n194227 , n26951 , 
 n26952 , n194230 , n194231 , n26955 , n194233 , n194234 , n26958 , n194236 , n26960 , n194238 , 
 n26962 , n194240 , n26964 , n194242 , n194243 , n26967 , n194245 , n194246 , n26970 , n194248 , 
 n194249 , n26973 , n194251 , n26975 , n26976 , n194254 , n194255 , n26979 , n194257 , n194258 , 
 n26982 , n194260 , n194261 , n26985 , n194263 , n26987 , n194265 , n26989 , n26990 , n194268 , 
 n194269 , n26993 , n194271 , n194272 , n26996 , n194274 , n194275 , n26999 , n194277 , n27001 , 
 n194279 , n27003 , n27004 , n194282 , n194283 , n27007 , n194285 , n194286 , n27010 , n194288 , 
 n194289 , n27013 , n194291 , n194292 , n194293 , n194294 , n27018 , n194296 , n194297 , n27021 , 
 n194299 , n194300 , n27024 , n194302 , n194303 , n27027 , n194305 , n27029 , n194307 , n27031 , 
 n27032 , n194310 , n194311 , n27035 , n194313 , n194314 , n27038 , n194316 , n27040 , n194318 , 
 n27042 , n194320 , n27044 , n27045 , n194323 , n194324 , n27048 , n194326 , n194327 , n27051 , 
 n194329 , n27053 , n27054 , n27055 , n194333 , n194334 , n27058 , n194336 , n27060 , n27061 , 
 n27062 , n27063 , n194341 , n194342 , n27066 , n194344 , n27068 , n194346 , n27070 , n27071 , 
 n194349 , n27073 , n27074 , n27075 , n194353 , n27077 , n27078 , n27079 , n194357 , n194358 , 
 n27082 , n194360 , n194361 , n27085 , n194363 , n27087 , n27088 , n27089 , n194367 , n194368 , 
 n27092 , n27093 , n194371 , n194372 , n27096 , n27097 , n27098 , n194376 , n27100 , n194378 , 
 n194379 , n27103 , n194381 , n194382 , n194383 , n194384 , n27108 , n194386 , n194387 , n27111 , 
 n27112 , n27113 , n27114 , n194392 , n194393 , n27117 , n194395 , n27119 , n194397 , n27121 , 
 n194399 , n194400 , n27124 , n194402 , n194403 , n27127 , n194405 , n27129 , n27130 , n194408 , 
 n194409 , n27133 , n194411 , n194412 , n27136 , n194414 , n194415 , n27139 , n27140 , n27141 , 
 n194419 , n194420 , n27144 , n194422 , n194423 , n27147 , n194425 , n194426 , n27150 , n194428 , 
 n27152 , n27153 , n194431 , n194432 , n27156 , n194434 , n194435 , n27159 , n194437 , n194438 , 
 n194439 , n194440 , n27164 , n194442 , n194443 , n27167 , n194445 , n27169 , n27170 , n194448 , 
 n194449 , n27173 , n194451 , n194452 , n27176 , n194454 , n194455 , n27179 , n27180 , n194458 , 
 n27182 , n194460 , n27184 , n27185 , n194463 , n194464 , n27188 , n194466 , n194467 , n27191 , 
 n194469 , n194470 , n27194 , n27195 , n27196 , n194474 , n194475 , n27199 , n27200 , n27201 , 
 n194479 , n194480 , n27204 , n27205 , n27206 , n194484 , n194485 , n27209 , n27210 , n27211 , 
 n194489 , n194490 , n27214 , n194492 , n27216 , n194494 , n27218 , n194496 , n27220 , n27221 , 
 n194499 , n27223 , n194501 , n27225 , n194503 , n194504 , n27228 , n194506 , n27230 , n194508 , 
 n27232 , n194510 , n27234 , n27235 , n194513 , n194514 , n27238 , n194516 , n194517 , n27241 , 
 n194519 , n27243 , n194521 , n194522 , n194523 , n27247 , n194525 , n27249 , n194527 , n194528 , 
 n194529 , n194530 , n27254 , n194532 , n194533 , n194534 , n27258 , n194536 , n194537 , n27261 , 
 n194539 , n27263 , n194541 , n27265 , n27266 , n194544 , n194545 , n27269 , n194547 , n194548 , 
 n27272 , n194550 , n194551 , n27275 , n27276 , n194554 , n194555 , n27279 , n27280 , n194558 , 
 n194559 , n27283 , n194561 , n194562 , n27286 , n27287 , n27288 , n27289 , n194567 , n194568 , 
 n194569 , n194570 , n27294 , n194572 , n27296 , n194574 , n194575 , n194576 , n194577 , n27301 , 
 n194579 , n194580 , n27304 , n194582 , n194583 , n27307 , n194585 , n27309 , n194587 , n27311 , 
 n27312 , n194590 , n194591 , n27315 , n194593 , n194594 , n27318 , n194596 , n194597 , n194598 , 
 n27322 , n194600 , n27324 , n27325 , n194603 , n194604 , n27328 , n194606 , n194607 , n27331 , 
 n194609 , n194610 , n27334 , n194612 , n27336 , n194614 , n27338 , n27339 , n194617 , n194618 , 
 n27342 , n194620 , n194621 , n27345 , n194623 , n194624 , n27348 , n194626 , n194627 , n27351 , 
 n194629 , n194630 , n27354 , n27355 , n27356 , n27357 , n27358 , n194636 , n194637 , n27361 , 
 n194639 , n27363 , n194641 , n194642 , n27366 , n194644 , n27368 , n27369 , n27370 , n194648 , 
 n194649 , n194650 , n27374 , n194652 , n194653 , n27377 , n194655 , n27379 , n194657 , n194658 , 
 n27382 , n194660 , n27384 , n27385 , n27386 , n194664 , n194665 , n194666 , n27390 , n194668 , 
 n194669 , n27393 , n194671 , n27395 , n27396 , n194674 , n194675 , n27399 , n194677 , n27401 , 
 n27402 , n27403 , n27404 , n194682 , n194683 , n27407 , n194685 , n27409 , n27410 , n27411 , 
 n27412 , n194690 , n194691 , n27415 , n194693 , n27417 , n27418 , n194696 , n194697 , n27421 , 
 n27422 , n194700 , n194701 , n27425 , n194703 , n27427 , n27428 , n194706 , n27430 , n194708 , 
 n27432 , n27433 , n194711 , n194712 , n27436 , n194714 , n194715 , n27439 , n194717 , n194718 , 
 n27442 , n194720 , n27444 , n27445 , n194723 , n194724 , n27448 , n194726 , n194727 , n27451 , 
 n194729 , n27453 , n194731 , n194732 , n27456 , n194734 , n194735 , n27459 , n194737 , n27461 , 
 n27462 , n194740 , n194741 , n27465 , n194743 , n194744 , n27468 , n194746 , n194747 , n194748 , 
 n194749 , n27473 , n194751 , n27475 , n194753 , n194754 , n194755 , n194756 , n27480 , n194758 , 
 n194759 , n194760 , n27484 , n194762 , n194763 , n27487 , n194765 , n194766 , n27490 , n194768 , 
 n194769 , n27493 , n194771 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , 
 n194779 , n194780 , n27504 , n194782 , n27506 , n194784 , n194785 , n194786 , n194787 , n27511 , 
 n194789 , n194790 , n194791 , n27515 , n194793 , n194794 , n194795 , n194796 , n27520 , n194798 , 
 n194799 , n27523 , n194801 , n27525 , n27526 , n194804 , n194805 , n27529 , n194807 , n194808 , 
 n194809 , n27533 , n194811 , n194812 , n27536 , n194814 , n194815 , n27539 , n194817 , n27541 , 
 n27542 , n27543 , n27544 , n27545 , n194823 , n27547 , n27548 , n27549 , n194827 , n194828 , 
 n27552 , n27553 , n194831 , n194832 , n27556 , n27557 , n194835 , n194836 , n27560 , n194838 , 
 n194839 , n27563 , n194841 , n27565 , n27566 , n27567 , n194845 , n194846 , n27570 , n194848 , 
 n27572 , n194850 , n27574 , n27575 , n27576 , n194854 , n194855 , n27579 , n27580 , n194858 , 
 n27582 , n27583 , n194861 , n27585 , n27586 , n194864 , n194865 , n27589 , n27590 , n194868 , 
 n194869 , n27593 , n27594 , n194872 , n194873 , n27597 , n194875 , n27599 , n194877 , n27601 , 
 n27602 , n27603 , n194881 , n194882 , n27606 , n194884 , n194885 , n27609 , n194887 , n194888 , 
 n194889 , n27613 , n194891 , n27615 , n194893 , n194894 , n27618 , n27619 , n27620 , n27621 , 
 n27622 , n194900 , n194901 , n27625 , n27626 , n27627 , n194905 , n194906 , n27630 , n194908 , 
 n194909 , n27633 , n194911 , n27635 , n194913 , n194914 , n27638 , n194916 , n27640 , n194918 , 
 n194919 , n194920 , n194921 , n27645 , n194923 , n194924 , n194925 , n27649 , n194927 , n194928 , 
 n27652 , n27653 , n194931 , n27655 , n194933 , n27657 , n27658 , n27659 , n194937 , n194938 , 
 n27662 , n194940 , n194941 , n27665 , n194943 , n194944 , n27668 , n194946 , n194947 , n27671 , 
 n194949 , n194950 , n27674 , n194952 , n194953 , n27677 , n194955 , n27679 , n27680 , n194958 , 
 n27682 , n194960 , n27684 , n194962 , n194963 , n27687 , n194965 , n194966 , n27690 , n194968 , 
 n194969 , n27693 , n194971 , n27695 , n194973 , n27697 , n194975 , n194976 , n27700 , n194978 , 
 n194979 , n194980 , n194981 , n27705 , n194983 , n194984 , n27708 , n194986 , n27710 , n27711 , 
 n194989 , n194990 , n194991 , n27715 , n194993 , n194994 , n27718 , n194996 , n194997 , n27721 , 
 n194999 , n27723 , n27724 , n195002 , n27726 , n27727 , n195005 , n27729 , n27730 , n195008 , 
 n195009 , n195010 , n27734 , n195012 , n27736 , n27737 , n195015 , n195016 , n27740 , n27741 , 
 n195019 , n195020 , n195021 , n195022 , n27746 , n195024 , n195025 , n27749 , n195027 , n27751 , 
 n27752 , n195030 , n195031 , n27755 , n195033 , n195034 , n27758 , n195036 , n195037 , n195038 , 
 n195039 , n27763 , n195041 , n195042 , n27766 , n195044 , n27768 , n195046 , n195047 , n195048 , 
 n195049 , n27773 , n195051 , n195052 , n27776 , n195054 , n195055 , n195056 , n27780 , n195058 , 
 n195059 , n27783 , n195061 , n195062 , n27786 , n27787 , n195065 , n195066 , n27790 , n27791 , 
 n27792 , n195070 , n195071 , n27795 , n27796 , n195074 , n27798 , n195076 , n27800 , n27801 , 
 n195079 , n27803 , n195081 , n27805 , n195083 , n195084 , n27808 , n195086 , n195087 , n195088 , 
 n195089 , n27813 , n195091 , n195092 , n27816 , n195094 , n27818 , n27819 , n195097 , n195098 , 
 n195099 , n27823 , n195101 , n195102 , n27826 , n195104 , n195105 , n27829 , n195107 , n195108 , 
 n27832 , n195110 , n195111 , n27835 , n195113 , n195114 , n27838 , n195116 , n27840 , n27841 , 
 n195119 , n195120 , n195121 , n27845 , n195123 , n195124 , n27848 , n195126 , n195127 , n27851 , 
 n195129 , n195130 , n27854 , n27855 , n27856 , n195134 , n195135 , n27859 , n27860 , n27861 , 
 n195139 , n195140 , n27864 , n27865 , n27866 , n27867 , n195145 , n195146 , n27870 , n195148 , 
 n27872 , n27873 , n195151 , n27875 , n195153 , n27877 , n27878 , n195156 , n195157 , n195158 , 
 n27882 , n195160 , n195161 , n27885 , n195163 , n195164 , n27888 , n195166 , n27890 , n195168 , 
 n27892 , n195170 , n27894 , n27895 , n195173 , n195174 , n195175 , n27899 , n195177 , n195178 , 
 n27902 , n195180 , n195181 , n27905 , n195183 , n27907 , n195185 , n195186 , n195187 , n27911 , 
 n195189 , n195190 , n27914 , n195192 , n27916 , n27917 , n195195 , n195196 , n195197 , n27921 , 
 n195199 , n195200 , n27924 , n195202 , n195203 , n27927 , n195205 , n27929 , n195207 , n195208 , 
 n27932 , n195210 , n195211 , n27935 , n195213 , n27937 , n27938 , n195216 , n195217 , n195218 , 
 n27942 , n195220 , n195221 , n27945 , n195223 , n195224 , n27948 , n195226 , n27950 , n27951 , 
 n27952 , n195230 , n195231 , n27955 , n195233 , n195234 , n27958 , n195236 , n27960 , n27961 , 
 n195239 , n195240 , n195241 , n27965 , n195243 , n195244 , n27968 , n195246 , n195247 , n27971 , 
 n195249 , n27973 , n27974 , n195252 , n27976 , n27977 , n27978 , n27979 , n195257 , n195258 , 
 n195259 , n27983 , n195261 , n195262 , n27986 , n195264 , n27988 , n195266 , n195267 , n195268 , 
 n27992 , n195270 , n27994 , n27995 , n27996 , n195274 , n195275 , n27999 , n195277 , n28001 , 
 n195279 , n28003 , n195281 , n195282 , n195283 , n28007 , n195285 , n28009 , n28010 , n195288 , 
 n195289 , n28013 , n195291 , n195292 , n28016 , n195294 , n195295 , n28019 , n195297 , n195298 , 
 n28022 , n195300 , n195301 , n195302 , n195303 , n28027 , n195305 , n195306 , n28030 , n195308 , 
 n195309 , n28033 , n28034 , n28035 , n195313 , n195314 , n195315 , n195316 , n28040 , n195318 , 
 n195319 , n195320 , n28044 , n195322 , n28046 , n28047 , n195325 , n195326 , n28050 , n195328 , 
 n195329 , n195330 , n28054 , n195332 , n195333 , n28057 , n195335 , n195336 , n28060 , n195338 , 
 n28062 , n195340 , n28064 , n28065 , n195343 , n195344 , n195345 , n28069 , n195347 , n195348 , 
 n28072 , n195350 , n195351 , n28075 , n195353 , n195354 , n28078 , n195356 , n195357 , n195358 , 
 n28082 , n195360 , n28084 , n28085 , n195363 , n195364 , n195365 , n28089 , n195367 , n195368 , 
 n28092 , n195370 , n195371 , n28095 , n195373 , n195374 , n195375 , n195376 , n28100 , n195378 , 
 n195379 , n28103 , n195381 , n28105 , n28106 , n195384 , n195385 , n195386 , n28110 , n195388 , 
 n195389 , n28113 , n195391 , n195392 , n28116 , n195394 , n195395 , n28119 , n28120 , n195398 , 
 n28122 , n195400 , n28124 , n28125 , n195403 , n195404 , n195405 , n28129 , n195407 , n195408 , 
 n28132 , n195410 , n195411 , n28135 , n195413 , n195414 , n28138 , n195416 , n195417 , n28141 , 
 n195419 , n28143 , n195421 , n28145 , n28146 , n195424 , n195425 , n195426 , n28150 , n195428 , 
 n195429 , n28153 , n195431 , n195432 , n28156 , n195434 , n195435 , n28159 , n195437 , n28161 , 
 n195439 , n28163 , n28164 , n195442 , n195443 , n195444 , n28168 , n195446 , n195447 , n28171 , 
 n195449 , n195450 , n28174 , n195452 , n195453 , n28177 , n195455 , n195456 , n28180 , n28181 , 
 n195459 , n195460 , n28184 , n28185 , n195463 , n195464 , n195465 , n195466 , n28190 , n195468 , 
 n195469 , n28193 , n195471 , n28195 , n28196 , n195474 , n195475 , n195476 , n28200 , n195478 , 
 n195479 , n28203 , n195481 , n195482 , n28206 , n195484 , n195485 , n28209 , n28210 , n195488 , 
 n28212 , n195490 , n195491 , n28215 , n28216 , n195494 , n195495 , n28219 , n195497 , n28221 , 
 n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , 
 n195509 , n28233 , n28234 , n28235 , n28236 , n195514 , n28238 , n195516 , n195517 , n195518 , 
 n28242 , n195520 , n28244 , n28245 , n195523 , n195524 , n28248 , n195526 , n195527 , n28251 , 
 n195529 , n28253 , n195531 , n28255 , n195533 , n28257 , n28258 , n195536 , n195537 , n28261 , 
 n195539 , n195540 , n28264 , n195542 , n28266 , n28267 , n195545 , n195546 , n28270 , n195548 , 
 n195549 , n28273 , n195551 , n195552 , n28276 , n195554 , n28278 , n28279 , n195557 , n195558 , 
 n28282 , n195560 , n195561 , n28285 , n195563 , n195564 , n28288 , n195566 , n28290 , n195568 , 
 n28292 , n195570 , n195571 , n28295 , n28296 , n195574 , n28298 , n28299 , n195577 , n28301 , 
 n28302 , n28303 , n28304 , n195582 , n28306 , n28307 , n195585 , n28309 , n195587 , n28311 , 
 n195589 , n28313 , n195591 , n28315 , n28316 , n28317 , n28318 , n28319 , n195597 , n195598 , 
 n195599 , n28323 , n195601 , n28325 , n195603 , n28327 , n195605 , n195606 , n195607 , n28331 , 
 n195609 , n28333 , n28334 , n195612 , n195613 , n195614 , n28338 , n195616 , n195617 , n28341 , 
 n195619 , n195620 , n28344 , n195622 , n195623 , n28347 , n195625 , n28349 , n28350 , n28351 , 
 n195629 , n195630 , n28354 , n195632 , n28356 , n28357 , n28358 , n195636 , n195637 , n28361 , 
 n195639 , n195640 , n28364 , n195642 , n28366 , n28367 , n195645 , n28369 , n195647 , n28371 , 
 n195649 , n195650 , n28374 , n195652 , n28376 , n28377 , n195655 , n28379 , n195657 , n28381 , 
 n195659 , n28383 , n28384 , n195662 , n195663 , n28387 , n195665 , n195666 , n195667 , n28391 , 
 n195669 , n195670 , n28394 , n195672 , n195673 , n28397 , n195675 , n195676 , n28400 , n195678 , 
 n28402 , n28403 , n195681 , n195682 , n195683 , n28407 , n195685 , n195686 , n28410 , n195688 , 
 n195689 , n28413 , n195691 , n28415 , n195693 , n28417 , n195695 , n28419 , n28420 , n195698 , 
 n195699 , n195700 , n28424 , n195702 , n195703 , n28427 , n195705 , n195706 , n28430 , n195708 , 
 n28432 , n195710 , n28434 , n195712 , n195713 , n28437 , n195715 , n28439 , n195717 , n28441 , 
 n28442 , n195720 , n195721 , n28445 , n195723 , n28447 , n195725 , n195726 , n28450 , n195728 , 
 n195729 , n195730 , n28454 , n195732 , n28456 , n28457 , n195735 , n195736 , n195737 , n28461 , 
 n195739 , n195740 , n28464 , n195742 , n195743 , n28467 , n195745 , n195746 , n195747 , n195748 , 
 n28472 , n195750 , n28474 , n195752 , n195753 , n195754 , n195755 , n28479 , n195757 , n195758 , 
 n195759 , n28483 , n195761 , n195762 , n195763 , n28487 , n195765 , n28489 , n28490 , n195768 , 
 n195769 , n195770 , n28494 , n195772 , n195773 , n28497 , n195775 , n195776 , n28500 , n195778 , 
 n195779 , n28503 , n195781 , n195782 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , 
 n28512 , n28513 , n28514 , n195792 , n28516 , n195794 , n195795 , n28519 , n28520 , n28521 , 
 n28522 , n28523 , n195801 , n195802 , n28526 , n28527 , n28528 , n28529 , n195807 , n195808 , 
 n28532 , n195810 , n28534 , n195812 , n28536 , n28537 , n195815 , n195816 , n28540 , n195818 , 
 n195819 , n195820 , n28544 , n195822 , n195823 , n28547 , n195825 , n195826 , n195827 , n28551 , 
 n195829 , n28553 , n28554 , n195832 , n195833 , n195834 , n28558 , n195836 , n195837 , n28561 , 
 n195839 , n195840 , n28564 , n195842 , n195843 , n28567 , n195845 , n28569 , n195847 , n28571 , 
 n28572 , n195850 , n195851 , n195852 , n28576 , n195854 , n195855 , n28579 , n195857 , n195858 , 
 n28582 , n195860 , n195861 , n28585 , n195863 , n195864 , n28588 , n195866 , n195867 , n28591 , 
 n195869 , n195870 , n28594 , n195872 , n195873 , n28597 , n28598 , n28599 , n195877 , n28601 , 
 n195879 , n195880 , n28604 , n195882 , n28606 , n195884 , n195885 , n195886 , n195887 , n28611 , 
 n195889 , n195890 , n195891 , n28615 , n195893 , n195894 , n195895 , n28619 , n195897 , n28621 , 
 n28622 , n195900 , n195901 , n28625 , n195903 , n195904 , n28628 , n195906 , n195907 , n28631 , 
 n195909 , n195910 , n28634 , n28635 , n195913 , n28637 , n195915 , n28639 , n28640 , n195918 , 
 n195919 , n28643 , n195921 , n195922 , n28646 , n195924 , n28648 , n195926 , n28650 , n195928 , 
 n195929 , n28653 , n195931 , n28655 , n195933 , n28657 , n28658 , n195936 , n28660 , n195938 , 
 n28662 , n195940 , n195941 , n28665 , n195943 , n195944 , n28668 , n195946 , n28670 , n195948 , 
 n28672 , n28673 , n195951 , n195952 , n28676 , n195954 , n195955 , n28679 , n195957 , n195958 , 
 n28682 , n28683 , n195961 , n195962 , n28686 , n195964 , n195965 , n28689 , n195967 , n195968 , 
 n28692 , n195970 , n28694 , n28695 , n195973 , n195974 , n28698 , n195976 , n195977 , n28701 , 
 n195979 , n195980 , n28704 , n195982 , n195983 , n28707 , n195985 , n195986 , n28710 , n28711 , 
 n195989 , n195990 , n28714 , n195992 , n195993 , n28717 , n195995 , n195996 , n28720 , n28721 , 
 n195999 , n196000 , n28724 , n196002 , n196003 , n28727 , n196005 , n196006 , n196007 , n28731 , 
 n196009 , n196010 , n28734 , n28735 , n28736 , n196014 , n196015 , n196016 , n28740 , n196018 , 
 n28742 , n28743 , n196021 , n196022 , n28746 , n196024 , n196025 , n28749 , n196027 , n196028 , 
 n28752 , n196030 , n196031 , n28755 , n196033 , n28757 , n196035 , n28759 , n28760 , n196038 , 
 n196039 , n28763 , n196041 , n196042 , n28766 , n196044 , n196045 , n28769 , n196047 , n196048 , 
 n196049 , n196050 , n28774 , n196052 , n196053 , n28777 , n196055 , n196056 , n28780 , n28781 , 
 n196059 , n196060 , n28784 , n196062 , n196063 , n28787 , n196065 , n196066 , n28790 , n196068 , 
 n28792 , n28793 , n196071 , n196072 , n28796 , n28797 , n196075 , n196076 , n28800 , n28801 , 
 n28802 , n196080 , n196081 , n28805 , n196083 , n196084 , n28808 , n196086 , n196087 , n28811 , 
 n28812 , n28813 , n196091 , n196092 , n196093 , n28817 , n196095 , n28819 , n28820 , n196098 , 
 n196099 , n28823 , n196101 , n196102 , n28826 , n196104 , n28828 , n196106 , n28830 , n196108 , 
 n28832 , n196110 , n28834 , n28835 , n196113 , n196114 , n28838 , n196116 , n196117 , n28841 , 
 n196119 , n196120 , n28844 , n196122 , n196123 , n28847 , n28848 , n196126 , n28850 , n196128 , 
 n28852 , n28853 , n196131 , n196132 , n28856 , n196134 , n196135 , n28859 , n196137 , n196138 , 
 n28862 , n196140 , n196141 , n196142 , n28866 , n196144 , n28868 , n196146 , n196147 , n28871 , 
 n196149 , n196150 , n28874 , n196152 , n28876 , n196154 , n196155 , n28879 , n28880 , n196158 , 
 n28882 , n28883 , n196161 , n196162 , n28886 , n28887 , n196165 , n196166 , n28890 , n28891 , 
 n28892 , n196170 , n196171 , n28895 , n28896 , n196174 , n196175 , n28899 , n28900 , n28901 , 
 n196179 , n28903 , n196181 , n196182 , n28906 , n196184 , n196185 , n28909 , n196187 , n28911 , 
 n196189 , n28913 , n28914 , n196192 , n196193 , n28917 , n28918 , n196196 , n196197 , n28921 , 
 n196199 , n28923 , n28924 , n196202 , n196203 , n28927 , n28928 , n196206 , n196207 , n28931 , 
 n196209 , n28933 , n28934 , n28935 , n196213 , n196214 , n28938 , n28939 , n28940 , n28941 , 
 n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n196227 , n28951 , 
 n196229 , n28953 , n28954 , n196232 , n196233 , n28957 , n196235 , n28959 , n196237 , n196238 , 
 n28962 , n196240 , n28964 , n28965 , n28966 , n196244 , n28968 , n28969 , n196247 , n196248 , 
 n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n196257 , n28981 , 
 n28982 , n28983 , n196261 , n28985 , n28986 , n28987 , n28988 , n196266 , n28990 , n196268 , 
 n196269 , n196270 , n28994 , n28995 , n196273 , n28997 , n196275 , n196276 , n29000 , n196278 , 
 n196279 , n29003 , n29004 , n29005 , n196283 , n196284 , n29008 , n29009 , n196287 , n29011 , 
 n196289 , n29013 , n29014 , n29015 , n29016 , n196294 , n29018 , n29019 , n29020 , n196298 , 
 n29022 , n196300 , n29024 , n196302 , n29026 , n29027 , n196305 , n196306 , n29030 , n196308 , 
 n196309 , n196310 , n29034 , n196312 , n196313 , n29037 , n196315 , n29039 , n29040 , n29041 , 
 n196319 , n29043 , n196321 , n29045 , n29046 , n196324 , n196325 , n196326 , n29050 , n196328 , 
 n196329 , n29053 , n196331 , n196332 , n29056 , n196334 , n196335 , n196336 , n196337 , n29061 , 
 n196339 , n196340 , n29064 , n196342 , n29066 , n29067 , n196345 , n196346 , n196347 , n29071 , 
 n196349 , n196350 , n29074 , n196352 , n196353 , n29077 , n196355 , n196356 , n29080 , n196358 , 
 n196359 , n29083 , n196361 , n196362 , n29086 , n196364 , n29088 , n29089 , n196367 , n196368 , 
 n196369 , n29093 , n196371 , n196372 , n29096 , n196374 , n196375 , n29099 , n196377 , n196378 , 
 n29102 , n29103 , n29104 , n196382 , n196383 , n29107 , n196385 , n29109 , n196387 , n29111 , 
 n29112 , n196390 , n196391 , n196392 , n29116 , n196394 , n196395 , n29119 , n196397 , n196398 , 
 n29122 , n196400 , n196401 , n196402 , n29126 , n196404 , n29128 , n196406 , n196407 , n29131 , 
 n29132 , n196410 , n29134 , n196412 , n196413 , n29137 , n196415 , n196416 , n29140 , n196418 , 
 n196419 , n29143 , n196421 , n29145 , n29146 , n196424 , n196425 , n196426 , n29150 , n196428 , 
 n196429 , n29153 , n196431 , n196432 , n29156 , n196434 , n196435 , n29159 , n29160 , n29161 , 
 n196439 , n196440 , n29164 , n196442 , n29166 , n196444 , n29168 , n196446 , n196447 , n29171 , 
 n196449 , n196450 , n29174 , n29175 , n196453 , n196454 , n196455 , n29179 , n196457 , n196458 , 
 n29182 , n196460 , n196461 , n29185 , n196463 , n196464 , n29188 , n196466 , n29190 , n29191 , 
 n196469 , n196470 , n29194 , n196472 , n196473 , n29197 , n196475 , n29199 , n196477 , n196478 , 
 n29202 , n196480 , n29204 , n29205 , n196483 , n196484 , n196485 , n29209 , n196487 , n196488 , 
 n29212 , n196490 , n196491 , n29215 , n196493 , n196494 , n29218 , n196496 , n196497 , n29221 , 
 n196499 , n196500 , n29224 , n196502 , n196503 , n196504 , n29228 , n196506 , n29230 , n29231 , 
 n196509 , n196510 , n196511 , n29235 , n196513 , n196514 , n29238 , n196516 , n196517 , n29241 , 
 n196519 , n196520 , n29244 , n196522 , n29246 , n196524 , n29248 , n29249 , n196527 , n196528 , 
 n196529 , n29253 , n196531 , n196532 , n29256 , n196534 , n196535 , n29259 , n196537 , n196538 , 
 n29262 , n196540 , n196541 , n29265 , n196543 , n196544 , n196545 , n196546 , n29270 , n196548 , 
 n196549 , n196550 , n196551 , n29275 , n196553 , n196554 , n29278 , n196556 , n29280 , n29281 , 
 n196559 , n196560 , n29284 , n196562 , n196563 , n29287 , n196565 , n196566 , n29290 , n29291 , 
 n196569 , n29293 , n196571 , n29295 , n29296 , n196574 , n196575 , n29299 , n196577 , n196578 , 
 n29302 , n196580 , n196581 , n29305 , n196583 , n29307 , n196585 , n29309 , n29310 , n196588 , 
 n196589 , n29313 , n196591 , n196592 , n29316 , n196594 , n196595 , n29319 , n196597 , n196598 , 
 n196599 , n196600 , n29324 , n196602 , n196603 , n29327 , n196605 , n196606 , n29330 , n196608 , 
 n29332 , n29333 , n196611 , n196612 , n29336 , n196614 , n196615 , n29339 , n196617 , n196618 , 
 n29342 , n196620 , n196621 , n29345 , n196623 , n196624 , n29348 , n29349 , n29350 , n196628 , 
 n196629 , n29353 , n196631 , n196632 , n29356 , n196634 , n196635 , n29359 , n196637 , n196638 , 
 n29362 , n196640 , n29364 , n29365 , n196643 , n196644 , n29368 , n196646 , n196647 , n29371 , 
 n196649 , n196650 , n29374 , n196652 , n196653 , n29377 , n196655 , n196656 , n29380 , n196658 , 
 n29382 , n29383 , n196661 , n196662 , n29386 , n196664 , n196665 , n29389 , n196667 , n196668 , 
 n29392 , n29393 , n29394 , n196672 , n196673 , n29397 , n29398 , n196676 , n196677 , n29401 , 
 n29402 , n29403 , n196681 , n196682 , n29406 , n29407 , n29408 , n196686 , n196687 , n29411 , 
 n196689 , n196690 , n29414 , n29415 , n29416 , n196694 , n196695 , n196696 , n29420 , n196698 , 
 n196699 , n196700 , n196701 , n29425 , n196703 , n196704 , n29428 , n196706 , n29430 , n29431 , 
 n196709 , n196710 , n29434 , n196712 , n196713 , n29437 , n196715 , n196716 , n29440 , n196718 , 
 n196719 , n29443 , n196721 , n196722 , n29446 , n196724 , n196725 , n29449 , n196727 , n29451 , 
 n29452 , n196730 , n196731 , n29455 , n196733 , n196734 , n29458 , n196736 , n196737 , n29461 , 
 n196739 , n196740 , n196741 , n196742 , n29466 , n196744 , n196745 , n29469 , n196747 , n196748 , 
 n29472 , n196750 , n196751 , n29475 , n196753 , n196754 , n29478 , n196756 , n29480 , n29481 , 
 n196759 , n196760 , n29484 , n196762 , n196763 , n29487 , n196765 , n196766 , n29490 , n29491 , 
 n196769 , n29493 , n196771 , n196772 , n29496 , n196774 , n196775 , n29499 , n196777 , n29501 , 
 n29502 , n196780 , n196781 , n29505 , n196783 , n196784 , n29508 , n196786 , n196787 , n29511 , 
 n29512 , n29513 , n196791 , n196792 , n29516 , n29517 , n29518 , n196796 , n196797 , n29521 , 
 n196799 , n196800 , n29524 , n196802 , n196803 , n29527 , n196805 , n29529 , n29530 , n196808 , 
 n196809 , n29533 , n196811 , n196812 , n29536 , n196814 , n196815 , n196816 , n196817 , n29541 , 
 n196819 , n196820 , n29544 , n196822 , n29546 , n29547 , n196825 , n196826 , n29550 , n196828 , 
 n196829 , n29553 , n196831 , n196832 , n29556 , n196834 , n29558 , n196836 , n29560 , n29561 , 
 n196839 , n196840 , n29564 , n196842 , n196843 , n29567 , n196845 , n196846 , n29570 , n196848 , 
 n196849 , n196850 , n196851 , n29575 , n196853 , n196854 , n29578 , n196856 , n196857 , n29581 , 
 n29582 , n196860 , n196861 , n29585 , n29586 , n196864 , n196865 , n29589 , n196867 , n196868 , 
 n29592 , n29593 , n29594 , n196872 , n196873 , n29597 , n29598 , n29599 , n196877 , n196878 , 
 n29602 , n196880 , n29604 , n29605 , n196883 , n196884 , n196885 , n29609 , n196887 , n29611 , 
 n29612 , n196890 , n29614 , n196892 , n29616 , n196894 , n196895 , n29619 , n29620 , n196898 , 
 n29622 , n196900 , n196901 , n29625 , n196903 , n196904 , n29628 , n29629 , n29630 , n29631 , 
 n29632 , n196910 , n196911 , n29635 , n196913 , n196914 , n29638 , n29639 , n29640 , n29641 , 
 n196919 , n196920 , n29644 , n29645 , n29646 , n29647 , n29648 , n196926 , n196927 , n29651 , 
 n196929 , n196930 , n196931 , n29655 , n196933 , n29657 , n196935 , n196936 , n29660 , n29661 , 
 n196939 , n29663 , n196941 , n196942 , n196943 , n196944 , n29668 , n196946 , n196947 , n29671 , 
 n196949 , n196950 , n196951 , n29675 , n196953 , n29677 , n29678 , n196956 , n196957 , n196958 , 
 n29682 , n196960 , n196961 , n29685 , n196963 , n196964 , n29688 , n196966 , n196967 , n196968 , 
 n29692 , n196970 , n29694 , n29695 , n196973 , n196974 , n196975 , n29699 , n196977 , n196978 , 
 n29702 , n196980 , n196981 , n29705 , n196983 , n196984 , n29708 , n196986 , n29710 , n196988 , 
 n29712 , n29713 , n196991 , n196992 , n196993 , n29717 , n196995 , n196996 , n29720 , n196998 , 
 n196999 , n29723 , n197001 , n197002 , n29726 , n197004 , n197005 , n29729 , n197007 , n29731 , 
 n197009 , n29733 , n29734 , n197012 , n197013 , n197014 , n29738 , n197016 , n197017 , n29741 , 
 n197019 , n197020 , n29744 , n197022 , n29746 , n29747 , n29748 , n197026 , n197027 , n197028 , 
 n29752 , n197030 , n197031 , n29755 , n197033 , n29757 , n29758 , n197036 , n29760 , n197038 , 
 n29762 , n29763 , n197041 , n197042 , n197043 , n29767 , n197045 , n197046 , n29770 , n197048 , 
 n197049 , n29773 , n197051 , n29775 , n197053 , n29777 , n197055 , n197056 , n29780 , n197058 , 
 n197059 , n29783 , n197061 , n29785 , n29786 , n197064 , n197065 , n29789 , n197067 , n197068 , 
 n197069 , n29793 , n197071 , n197072 , n29796 , n197074 , n197075 , n29799 , n197077 , n29801 , 
 n197079 , n29803 , n29804 , n197082 , n197083 , n197084 , n29808 , n197086 , n197087 , n29811 , 
 n197089 , n197090 , n29814 , n197092 , n197093 , n29817 , n197095 , n197096 , n197097 , n29821 , 
 n197099 , n29823 , n29824 , n197102 , n197103 , n29827 , n197105 , n197106 , n197107 , n29831 , 
 n197109 , n197110 , n29834 , n197112 , n197113 , n197114 , n29838 , n197116 , n29840 , n29841 , 
 n197119 , n197120 , n197121 , n29845 , n197123 , n197124 , n29848 , n197126 , n197127 , n29851 , 
 n197129 , n197130 , n29854 , n197132 , n29856 , n197134 , n29858 , n29859 , n197137 , n197138 , 
 n197139 , n29863 , n197141 , n197142 , n29866 , n197144 , n197145 , n29869 , n197147 , n197148 , 
 n29872 , n197150 , n197151 , n29875 , n29876 , n29877 , n29878 , n29879 , n197157 , n197158 , 
 n29882 , n197160 , n197161 , n29885 , n29886 , n29887 , n29888 , n29889 , n197167 , n197168 , 
 n29892 , n197170 , n197171 , n29895 , n29896 , n29897 , n29898 , n29899 , n197177 , n197178 , 
 n29902 , n29903 , n29904 , n197182 , n29906 , n29907 , n29908 , n29909 , n197187 , n197188 , 
 n29912 , n197190 , n29914 , n197192 , n197193 , n197194 , n197195 , n29919 , n197197 , n29921 , 
 n29922 , n29923 , n197201 , n197202 , n29926 , n197204 , n197205 , n29929 , n197207 , n197208 , 
 n197209 , n197210 , n29934 , n197212 , n29936 , n197214 , n197215 , n197216 , n197217 , n29941 , 
 n197219 , n29943 , n29944 , n29945 , n197223 , n197224 , n29948 , n197226 , n197227 , n197228 , 
 n29952 , n29953 , n197231 , n29955 , n29956 , n197234 , n29958 , n197236 , n29960 , n197238 , 
 n197239 , n29963 , n197241 , n197242 , n197243 , n29967 , n29968 , n197246 , n29970 , n197248 , 
 n197249 , n29973 , n29974 , n197252 , n197253 , n29977 , n29978 , n29979 , n29980 , n197258 , 
 n197259 , n29983 , n197261 , n197262 , n29986 , n197264 , n197265 , n197266 , n29990 , n197268 , 
 n29992 , n197270 , n197271 , n29995 , n197273 , n197274 , n29998 , n197276 , n197277 , n30001 , 
 n197279 , n197280 , n30004 , n197282 , n197283 , n197284 , n30008 , n197286 , n197287 , n30011 , 
 n197289 , n197290 , n30014 , n197292 , n197293 , n197294 , n30018 , n197296 , n197297 , n30021 , 
 n197299 , n197300 , n30024 , n197302 , n197303 , n30027 , n197305 , n30029 , n30030 , n30031 , 
 n197309 , n197310 , n30034 , n197312 , n197313 , n30037 , n30038 , n30039 , n30040 , n197318 , 
 n197319 , n30043 , n197321 , n197322 , n30046 , n197324 , n30048 , n197326 , n30050 , n197328 , 
 n30052 , n197330 , n30054 , n30055 , n30056 , n197334 , n30058 , n30059 , n197337 , n197338 , 
 n197339 , n30063 , n197341 , n30065 , n30066 , n197344 , n197345 , n30069 , n197347 , n30071 , 
 n197349 , n197350 , n30074 , n197352 , n197353 , n30077 , n197355 , n197356 , n30080 , n197358 , 
 n197359 , n30083 , n197361 , n197362 , n197363 , n197364 , n197365 , n30089 , n197367 , n197368 , 
 n197369 , n197370 , n30094 , n197372 , n197373 , n30097 , n197375 , n197376 , n30100 , n197378 , 
 n197379 , n30103 , n197381 , n197382 , n197383 , n30107 , n197385 , n197386 , n197387 , n30111 , 
 n197389 , n197390 , n30114 , n197392 , n197393 , n30117 , n30118 , n197396 , n197397 , n30121 , 
 n197399 , n197400 , n30124 , n197402 , n197403 , n30127 , n197405 , n197406 , n30130 , n197408 , 
 n197409 , n30133 , n197411 , n197412 , n30136 , n197414 , n197415 , n30139 , n197417 , n30141 , 
 n197419 , n197420 , n197421 , n197422 , n30146 , n197424 , n30148 , n30149 , n30150 , n197428 , 
 n197429 , n30153 , n197431 , n197432 , n30156 , n197434 , n197435 , n30159 , n30160 , n197438 , 
 n197439 , n197440 , n197441 , n30165 , n197443 , n30167 , n30168 , n30169 , n197447 , n197448 , 
 n30172 , n197450 , n197451 , n197452 , n197453 , n30177 , n197455 , n30179 , n197457 , n30181 , 
 n30182 , n30183 , n30184 , n30185 , n197463 , n30187 , n30188 , n30189 , n30190 , n197468 , 
 n197469 , n30193 , n30194 , n30195 , n30196 , n197474 , n197475 , n30199 , n197477 , n30201 , 
 n197479 , n30203 , n197481 , n197482 , n30206 , n30207 , n197485 , n197486 , n197487 , n30211 , 
 n197489 , n197490 , n30214 , n197492 , n197493 , n30217 , n197495 , n197496 , n30220 , n197498 , 
 n197499 , n30223 , n197501 , n197502 , n197503 , n30227 , n197505 , n197506 , n30230 , n197508 , 
 n197509 , n30233 , n30234 , n197512 , n30236 , n197514 , n197515 , n30239 , n197517 , n197518 , 
 n30242 , n30243 , n197521 , n197522 , n30246 , n197524 , n197525 , n30249 , n197527 , n197528 , 
 n30252 , n197530 , n197531 , n30255 , n197533 , n197534 , n30258 , n197536 , n197537 , n197538 , 
 n30262 , n197540 , n30264 , n197542 , n197543 , n30267 , n30268 , n30269 , n30270 , n197548 , 
 n197549 , n30273 , n197551 , n197552 , n30276 , n197554 , n197555 , n197556 , n197557 , n30281 , 
 n197559 , n197560 , n30284 , n197562 , n197563 , n30287 , n197565 , n30289 , n30290 , n30291 , 
 n30292 , n30293 , n30294 , n30295 , n197573 , n30297 , n197575 , n30299 , n197577 , n197578 , 
 n30302 , n30303 , n197581 , n30305 , n197583 , n30307 , n30308 , n197586 , n30310 , n197588 , 
 n197589 , n30313 , n197591 , n197592 , n30316 , n197594 , n197595 , n197596 , n30320 , n197598 , 
 n30322 , n197600 , n197601 , n30325 , n30326 , n197604 , n30328 , n197606 , n197607 , n30331 , 
 n30332 , n197610 , n30334 , n197612 , n197613 , n30337 , n197615 , n197616 , n30340 , n197618 , 
 n30342 , n197620 , n197621 , n30345 , n197623 , n197624 , n30348 , n197626 , n30350 , n197628 , 
 n197629 , n30353 , n30354 , n197632 , n30356 , n197634 , n30358 , n30359 , n197637 , n30361 , 
 n197639 , n197640 , n30364 , n197642 , n197643 , n30367 , n197645 , n197646 , n30370 , n30371 , 
 n197649 , n30373 , n30374 , n197652 , n30376 , n197654 , n197655 , n30379 , n30380 , n197658 , 
 n30382 , n30383 , n30384 , n30385 , n30386 , n197664 , n30388 , n197666 , n30390 , n30391 , 
 n197669 , n30393 , n197671 , n197672 , n197673 , n30397 , n30398 , n197676 , n30400 , n30401 , 
 n197679 , n197680 , n30404 , n197682 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , 
 n30412 , n197690 , n30414 , n197692 , n197693 , n197694 , n197695 , n30419 , n197697 , n197698 , 
 n197699 , n30423 , n197701 , n197702 , n30426 , n197704 , n197705 , n30429 , n197707 , n197708 , 
 n30432 , n197710 , n197711 , n30435 , n197713 , n197714 , n30438 , n197716 , n30440 , n197718 , 
 n30442 , n197720 , n197721 , n30445 , n30446 , n197724 , n197725 , n30449 , n30450 , n197728 , 
 n30452 , n30453 , n197731 , n30455 , n197733 , n30457 , n197735 , n197736 , n30460 , n197738 , 
 n197739 , n197740 , n30464 , n197742 , n197743 , n30467 , n197745 , n30469 , n197747 , n197748 , 
 n30472 , n30473 , n197751 , n30475 , n197753 , n197754 , n197755 , n197756 , n30480 , n197758 , 
 n197759 , n30483 , n197761 , n197762 , n30486 , n197764 , n197765 , n30489 , n30490 , n197768 , 
 n197769 , n30493 , n30494 , n197772 , n30496 , n30497 , n30498 , n197776 , n30500 , n197778 , 
 n30502 , n30503 , n197781 , n30505 , n197783 , n197784 , n30508 , n197786 , n197787 , n197788 , 
 n197789 , n30513 , n197791 , n197792 , n30516 , n197794 , n197795 , n30519 , n30520 , n197798 , 
 n30522 , n30523 , n197801 , n30525 , n30526 , n197804 , n30528 , n197806 , n30530 , n30531 , 
 n197809 , n30533 , n197811 , n197812 , n30536 , n197814 , n197815 , n197816 , n30540 , n197818 , 
 n30542 , n30543 , n197821 , n30545 , n197823 , n197824 , n30548 , n197826 , n197827 , n30551 , 
 n30552 , n197830 , n30554 , n30555 , n197833 , n30557 , n30558 , n30559 , n197837 , n30561 , 
 n197839 , n30563 , n30564 , n197842 , n30566 , n197844 , n197845 , n197846 , n30570 , n197848 , 
 n30572 , n197850 , n197851 , n30575 , n197853 , n197854 , n30578 , n30579 , n197857 , n30581 , 
 n30582 , n197860 , n30584 , n30585 , n197863 , n30587 , n197865 , n30589 , n30590 , n197868 , 
 n30592 , n197870 , n197871 , n197872 , n197873 , n30597 , n197875 , n197876 , n30600 , n197878 , 
 n197879 , n30603 , n30604 , n197882 , n30606 , n30607 , n197885 , n30609 , n30610 , n30611 , 
 n197889 , n197890 , n30614 , n197892 , n197893 , n197894 , n30618 , n197896 , n197897 , n30621 , 
 n30622 , n197900 , n30624 , n30625 , n197903 , n30627 , n30628 , n197906 , n197907 , n30631 , 
 n197909 , n197910 , n197911 , n30635 , n197913 , n30637 , n197915 , n197916 , n30640 , n197918 , 
 n30642 , n30643 , n30644 , n197922 , n30646 , n197924 , n30648 , n197926 , n30650 , n30651 , 
 n30652 , n197930 , n197931 , n30655 , n197933 , n30657 , n30658 , n197936 , n30660 , n197938 , 
 n197939 , n30663 , n197941 , n30665 , n30666 , n30667 , n197945 , n30669 , n197947 , n30671 , 
 n197949 , n197950 , n30674 , n197952 , n30676 , n30677 , n197955 , n197956 , n30680 , n197958 , 
 n30682 , n197960 , n197961 , n30685 , n197963 , n197964 , n197965 , n30689 , n197967 , n30691 , 
 n197969 , n197970 , n30694 , n30695 , n197973 , n30697 , n197975 , n197976 , n30700 , n30701 , 
 n197979 , n30703 , n30704 , n197982 , n197983 , n30707 , n197985 , n30709 , n197987 , n30711 , 
 n197989 , n197990 , n30714 , n197992 , n30716 , n30717 , n30718 , n197996 , n30720 , n30721 , 
 n197999 , n198000 , n30724 , n198002 , n30726 , n30727 , n30728 , n198006 , n30730 , n30731 , 
 n198009 , n30733 , n30734 , n198012 , n198013 , n30737 , n198015 , n30739 , n198017 , n198018 , 
 n30742 , n30743 , n30744 , n30745 , n198023 , n198024 , n30748 , n198026 , n198027 , n30751 , 
 n198029 , n30753 , n198031 , n30755 , n198033 , n198034 , n30758 , n198036 , n30760 , n30761 , 
 n30762 , n198040 , n198041 , n30765 , n30766 , n30767 , n198045 , n198046 , n30770 , n198048 , 
 n198049 , n30773 , n198051 , n198052 , n198053 , n30777 , n30778 , n30779 , n30780 , n198058 , 
 n198059 , n198060 , n198061 , n30785 , n198063 , n30787 , n198065 , n198066 , n30790 , n198068 , 
 n198069 , n30793 , n198071 , n198072 , n30796 , n30797 , n198075 , n198076 , n30800 , n30801 , 
 n30802 , n30803 , n198081 , n198082 , n30806 , n198084 , n198085 , n30809 , n198087 , n198088 , 
 n30812 , n198090 , n198091 , n30815 , n198093 , n30817 , n30818 , n198096 , n198097 , n30821 , 
 n198099 , n198100 , n198101 , n30825 , n198103 , n198104 , n30828 , n198106 , n198107 , n30831 , 
 n198109 , n198110 , n30834 , n198112 , n198113 , n30837 , n198115 , n198116 , n198117 , n30841 , 
 n198119 , n198120 , n30844 , n30845 , n198123 , n198124 , n198125 , n30849 , n198127 , n198128 , 
 n30852 , n198130 , n30854 , n198132 , n30856 , n198134 , n198135 , n30859 , n198137 , n198138 , 
 n30862 , n198140 , n198141 , n30865 , n198143 , n198144 , n30868 , n198146 , n198147 , n30871 , 
 n30872 , n198150 , n198151 , n30875 , n198153 , n198154 , n198155 , n30879 , n198157 , n30881 , 
 n198159 , n30883 , n198161 , n198162 , n198163 , n30887 , n198165 , n198166 , n30890 , n198168 , 
 n30892 , n30893 , n30894 , n30895 , n198173 , n30897 , n198175 , n198176 , n198177 , n30901 , 
 n198179 , n198180 , n30904 , n198182 , n198183 , n30907 , n198185 , n30909 , n198187 , n30911 , 
 n198189 , n198190 , n30914 , n30915 , n30916 , n30917 , n198195 , n198196 , n30920 , n198198 , 
 n198199 , n30923 , n198201 , n30925 , n198203 , n198204 , n30928 , n198206 , n198207 , n30931 , 
 n198209 , n198210 , n30934 , n198212 , n198213 , n30937 , n198215 , n198216 , n198217 , n198218 , 
 n30942 , n198220 , n198221 , n30945 , n198223 , n198224 , n30948 , n198226 , n198227 , n30951 , 
 n30952 , n198230 , n30954 , n198232 , n198233 , n30957 , n30958 , n198236 , n30960 , n30961 , 
 n30962 , n30963 , n198241 , n30965 , n198243 , n198244 , n198245 , n30969 , n198247 , n198248 , 
 n30972 , n198250 , n30974 , n198252 , n198253 , n30977 , n198255 , n198256 , n30980 , n30981 , 
 n198259 , n30983 , n198261 , n198262 , n198263 , n30987 , n30988 , n198266 , n30990 , n30991 , 
 n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n198276 , n198277 , n198278 , 
 n31002 , n198280 , n198281 , n31005 , n198283 , n198284 , n31008 , n198286 , n198287 , n31011 , 
 n198289 , n198290 , n31014 , n198292 , n198293 , n31017 , n198295 , n31019 , n198297 , n198298 , 
 n31022 , n198300 , n31024 , n31025 , n198303 , n31027 , n198305 , n31029 , n31030 , n198308 , 
 n198309 , n31033 , n198311 , n198312 , n31036 , n198314 , n198315 , n31039 , n198317 , n31041 , 
 n198319 , n31043 , n31044 , n198322 , n198323 , n31047 , n198325 , n198326 , n31050 , n198328 , 
 n31052 , n198330 , n198331 , n198332 , n31056 , n198334 , n198335 , n31059 , n198337 , n31061 , 
 n198339 , n31063 , n31064 , n31065 , n31066 , n198344 , n31068 , n198346 , n198347 , n31071 , 
 n198349 , n198350 , n198351 , n31075 , n198353 , n31077 , n31078 , n31079 , n198357 , n198358 , 
 n198359 , n31083 , n198361 , n31085 , n31086 , n198364 , n198365 , n31089 , n198367 , n198368 , 
 n31092 , n198370 , n198371 , n31095 , n198373 , n31097 , n31098 , n31099 , n198377 , n198378 , 
 n31102 , n198380 , n31104 , n198382 , n198383 , n198384 , n31108 , n198386 , n198387 , n31111 , 
 n198389 , n31113 , n198391 , n31115 , n198393 , n31117 , n31118 , n198396 , n198397 , n31121 , 
 n198399 , n198400 , n31124 , n198402 , n31126 , n31127 , n31128 , n31129 , n31130 , n198408 , 
 n31132 , n198410 , n31134 , n31135 , n31136 , n31137 , n198415 , n31139 , n198417 , n198418 , 
 n31142 , n198420 , n31144 , n198422 , n31146 , n31147 , n31148 , n31149 , n198427 , n31151 , 
 n198429 , n31153 , n198431 , n31155 , n31156 , n198434 , n198435 , n31159 , n198437 , n198438 , 
 n31162 , n198440 , n198441 , n31165 , n198443 , n198444 , n31168 , n198446 , n198447 , n198448 , 
 n31172 , n198450 , n31174 , n31175 , n198453 , n31177 , n198455 , n31179 , n31180 , n31181 , 
 n198459 , n198460 , n31184 , n198462 , n31186 , n198464 , n198465 , n31189 , n198467 , n31191 , 
 n198469 , n198470 , n31194 , n198472 , n198473 , n198474 , n31198 , n198476 , n31200 , n31201 , 
 n198479 , n31203 , n198481 , n31205 , n31206 , n31207 , n198485 , n31209 , n198487 , n198488 , 
 n31212 , n198490 , n31214 , n31215 , n31216 , n198494 , n31218 , n198496 , n198497 , n31221 , 
 n198499 , n31223 , n198501 , n198502 , n198503 , n198504 , n31228 , n198506 , n31230 , n31231 , 
 n31232 , n198510 , n198511 , n31235 , n198513 , n198514 , n31238 , n31239 , n198517 , n198518 , 
 n198519 , n198520 , n31244 , n198522 , n31246 , n31247 , n31248 , n198526 , n198527 , n31251 , 
 n198529 , n198530 , n31254 , n198532 , n198533 , n31257 , n198535 , n198536 , n31260 , n198538 , 
 n198539 , n198540 , n31264 , n198542 , n31266 , n31267 , n31268 , n198546 , n198547 , n31271 , 
 n198549 , n198550 , n31274 , n198552 , n31276 , n198554 , n198555 , n31279 , n198557 , n198558 , 
 n31282 , n198560 , n198561 , n198562 , n198563 , n31287 , n198565 , n31289 , n31290 , n31291 , 
 n198569 , n198570 , n31294 , n31295 , n31296 , n198574 , n198575 , n31299 , n198577 , n198578 , 
 n31302 , n198580 , n198581 , n31305 , n198583 , n198584 , n31308 , n198586 , n198587 , n31311 , 
 n198589 , n198590 , n31314 , n198592 , n31316 , n31317 , n31318 , n198596 , n198597 , n198598 , 
 n198599 , n31323 , n198601 , n31325 , n31326 , n31327 , n198605 , n198606 , n31330 , n198608 , 
 n198609 , n31333 , n31334 , n198612 , n198613 , n31337 , n31338 , n31339 , n31340 , n198618 , 
 n198619 , n31343 , n198621 , n198622 , n31346 , n198624 , n198625 , n31349 , n198627 , n198628 , 
 n31352 , n198630 , n198631 , n198632 , n31356 , n198634 , n31358 , n31359 , n31360 , n198638 , 
 n198639 , n31363 , n31364 , n198642 , n198643 , n31367 , n198645 , n198646 , n198647 , n198648 , 
 n31372 , n198650 , n31374 , n31375 , n31376 , n198654 , n198655 , n31379 , n31380 , n198658 , 
 n198659 , n31383 , n198661 , n198662 , n31386 , n198664 , n198665 , n198666 , n198667 , n31391 , 
 n198669 , n31393 , n31394 , n31395 , n198673 , n31397 , n31398 , n31399 , n31400 , n198678 , 
 n198679 , n31403 , n198681 , n31405 , n31406 , n31407 , n31408 , n198686 , n198687 , n31411 , 
 n198689 , n31413 , n31414 , n31415 , n31416 , n198694 , n198695 , n31419 , n198697 , n31421 , 
 n31422 , n31423 , n198701 , n31425 , n198703 , n198704 , n31428 , n198706 , n31430 , n198708 , 
 n198709 , n31433 , n198711 , n31435 , n31436 , n31437 , n198715 , n198716 , n31440 , n31441 , 
 n198719 , n198720 , n31444 , n198722 , n31446 , n31447 , n198725 , n31449 , n31450 , n31451 , 
 n31452 , n198730 , n31454 , n31455 , n198733 , n31457 , n198735 , n31459 , n198737 , n31461 , 
 n198739 , n198740 , n31464 , n198742 , n198743 , n31467 , n198745 , n31469 , n31470 , n198748 , 
 n31472 , n198750 , n198751 , n31475 , n198753 , n198754 , n31478 , n31479 , n198757 , n198758 , 
 n31482 , n198760 , n198761 , n31485 , n198763 , n198764 , n31488 , n198766 , n198767 , n31491 , 
 n198769 , n31493 , n198771 , n198772 , n31496 , n198774 , n198775 , n31499 , n198777 , n198778 , 
 n31502 , n31503 , n198781 , n31505 , n31506 , n198784 , n31508 , n198786 , n31510 , n198788 , 
 n198789 , n31513 , n198791 , n198792 , n31516 , n31517 , n198795 , n31519 , n198797 , n198798 , 
 n198799 , n198800 , n31524 , n198802 , n198803 , n31527 , n198805 , n198806 , n31530 , n198808 , 
 n198809 , n31533 , n198811 , n198812 , n31536 , n198814 , n198815 , n31539 , n198817 , n198818 , 
 n198819 , n198820 , n31544 , n198822 , n198823 , n31547 , n198825 , n198826 , n31550 , n198828 , 
 n31552 , n198830 , n198831 , n31555 , n31556 , n198834 , n31558 , n198836 , n198837 , n198838 , 
 n31562 , n198840 , n198841 , n31565 , n198843 , n198844 , n31568 , n198846 , n198847 , n198848 , 
 n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , 
 n198859 , n31583 , n198861 , n198862 , n31586 , n198864 , n198865 , n31589 , n198867 , n198868 , 
 n31592 , n198870 , n198871 , n31595 , n198873 , n198874 , n31598 , n198876 , n198877 , n198878 , 
 n31602 , n198880 , n198881 , n198882 , n31606 , n198884 , n198885 , n198886 , n31610 , n198888 , 
 n198889 , n31613 , n198891 , n198892 , n31616 , n198894 , n31618 , n31619 , n198897 , n31621 , 
 n198899 , n31623 , n198901 , n198902 , n31626 , n198904 , n198905 , n31629 , n198907 , n198908 , 
 n31632 , n198910 , n198911 , n31635 , n31636 , n198914 , n198915 , n31639 , n198917 , n198918 , 
 n31642 , n198920 , n198921 , n31645 , n198923 , n31647 , n31648 , n198926 , n198927 , n31651 , 
 n198929 , n31653 , n31654 , n31655 , n198933 , n31657 , n198935 , n31659 , n31660 , n31661 , 
 n31662 , n31663 , n31664 , n31665 , n198943 , n31667 , n31668 , n198946 , n31670 , n198948 , 
 n198949 , n31673 , n198951 , n198952 , n198953 , n198954 , n31678 , n198956 , n198957 , n31681 , 
 n198959 , n198960 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n198967 , n31691 , 
 n31692 , n198970 , n198971 , n198972 , n31696 , n198974 , n198975 , n31699 , n198977 , n198978 , 
 n31702 , n198980 , n198981 , n31705 , n198983 , n198984 , n198985 , n198986 , n31710 , n198988 , 
 n198989 , n31713 , n198991 , n31715 , n198993 , n198994 , n198995 , n31719 , n198997 , n198998 , 
 n31722 , n199000 , n199001 , n31725 , n199003 , n31727 , n199005 , n199006 , n31730 , n199008 , 
 n199009 , n31733 , n199011 , n31735 , n31736 , n199014 , n31738 , n199016 , n31740 , n199018 , 
 n199019 , n31743 , n199021 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n199028 , 
 n31752 , n199030 , n31754 , n199032 , n31756 , n31757 , n199035 , n31759 , n31760 , n31761 , 
 n199039 , n31763 , n199041 , n199042 , n31766 , n199044 , n199045 , n31769 , n31770 , n199048 , 
 n199049 , n31773 , n199051 , n199052 , n31776 , n199054 , n199055 , n199056 , n31780 , n199058 , 
 n199059 , n31783 , n199061 , n199062 , n31786 , n199064 , n31788 , n31789 , n31790 , n31791 , 
 n31792 , n199070 , n31794 , n199072 , n199073 , n31797 , n31798 , n31799 , n199077 , n31801 , 
 n199079 , n199080 , n31804 , n199082 , n199083 , n31807 , n199085 , n199086 , n31810 , n199088 , 
 n199089 , n31813 , n199091 , n199092 , n31816 , n199094 , n199095 , n31819 , n31820 , n31821 , 
 n199099 , n199100 , n31824 , n199102 , n31826 , n31827 , n199105 , n31829 , n199107 , n31831 , 
 n199109 , n31833 , n199111 , n199112 , n31836 , n199114 , n199115 , n31839 , n31840 , n199118 , 
 n31842 , n31843 , n199121 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , 
 n31852 , n199130 , n31854 , n199132 , n31856 , n31857 , n199135 , n31859 , n199137 , n199138 , 
 n31862 , n199140 , n31864 , n199142 , n199143 , n199144 , n31868 , n199146 , n31870 , n31871 , 
 n199149 , n31873 , n31874 , n31875 , n199153 , n31877 , n31878 , n199156 , n31880 , n199158 , 
 n31882 , n199160 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n199167 , n31891 , 
 n199169 , n199170 , n31894 , n199172 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , 
 n31902 , n199180 , n31904 , n199182 , n31906 , n199184 , n31908 , n31909 , n199187 , n31911 , 
 n199189 , n199190 , n31914 , n31915 , n199193 , n31917 , n199195 , n199196 , n31920 , n199198 , 
 n199199 , n199200 , n31924 , n199202 , n199203 , n199204 , n31928 , n199206 , n199207 , n31931 , 
 n199209 , n199210 , n31934 , n199212 , n199213 , n31937 , n31938 , n199216 , n31940 , n31941 , 
 n199219 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n199227 , n199228 , 
 n199229 , n31953 , n199231 , n199232 , n31956 , n199234 , n199235 , n31959 , n31960 , n199238 , 
 n31962 , n31963 , n199241 , n31965 , n31966 , n199244 , n31968 , n199246 , n31970 , n31971 , 
 n199249 , n31973 , n199251 , n199252 , n199253 , n199254 , n31978 , n199256 , n199257 , n31981 , 
 n199259 , n199260 , n31984 , n31985 , n199263 , n31987 , n31988 , n199266 , n31990 , n31991 , 
 n199269 , n31993 , n199271 , n199272 , n199273 , n31997 , n199275 , n199276 , n32000 , n199278 , 
 n199279 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , 
 n32012 , n32013 , n32014 , n32015 , n199293 , n32017 , n199295 , n199296 , n32020 , n199298 , 
 n199299 , n32023 , n32024 , n32025 , n199303 , n32027 , n199305 , n32029 , n199307 , n32031 , 
 n199309 , n199310 , n32034 , n32035 , n199313 , n32037 , n32038 , n199316 , n32040 , n32041 , 
 n199319 , n32043 , n199321 , n32045 , n32046 , n199324 , n32048 , n199326 , n199327 , n199328 , 
 n199329 , n32053 , n199331 , n199332 , n32056 , n199334 , n199335 , n32059 , n199337 , n199338 , 
 n32062 , n32063 , n199341 , n32065 , n32066 , n199344 , n32068 , n32069 , n199347 , n199348 , 
 n32072 , n199350 , n199351 , n199352 , n32076 , n199354 , n199355 , n32079 , n32080 , n199358 , 
 n32082 , n199360 , n199361 , n32085 , n32086 , n199364 , n32088 , n32089 , n32090 , n32091 , 
 n32092 , n32093 , n32094 , n32095 , n199373 , n199374 , n32098 , n199376 , n32100 , n199378 , 
 n199379 , n32103 , n199381 , n199382 , n32106 , n32107 , n199385 , n32109 , n32110 , n199388 , 
 n32112 , n32113 , n199391 , n32115 , n199393 , n32117 , n32118 , n199396 , n32120 , n199398 , 
 n199399 , n32123 , n199401 , n32125 , n32126 , n32127 , n199405 , n199406 , n32130 , n199408 , 
 n199409 , n32133 , n199411 , n199412 , n199413 , n32137 , n199415 , n199416 , n199417 , n32141 , 
 n199419 , n199420 , n199421 , n32145 , n199423 , n32147 , n32148 , n32149 , n32150 , n32151 , 
 n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n199435 , n199436 , n32160 , n199438 , 
 n199439 , n199440 , n32164 , n199442 , n199443 , n32167 , n199445 , n199446 , n32170 , n199448 , 
 n32172 , n32173 , n32174 , n32175 , n199453 , n199454 , n32178 , n199456 , n199457 , n32181 , 
 n199459 , n199460 , n199461 , n32185 , n199463 , n199464 , n32188 , n199466 , n32190 , n32191 , 
 n199469 , n32193 , n32194 , n199472 , n32196 , n32197 , n199475 , n32199 , n199477 , n32201 , 
 n199479 , n199480 , n32204 , n32205 , n199483 , n32207 , n199485 , n199486 , n32210 , n199488 , 
 n199489 , n32213 , n199491 , n199492 , n32216 , n199494 , n199495 , n32219 , n199497 , n199498 , 
 n199499 , n32223 , n199501 , n32225 , n199503 , n199504 , n32228 , n199506 , n199507 , n32231 , 
 n32232 , n199510 , n32234 , n32235 , n199513 , n32237 , n32238 , n32239 , n199517 , n199518 , 
 n199519 , n199520 , n32244 , n199522 , n199523 , n32247 , n199525 , n32249 , n32250 , n199528 , 
 n199529 , n32253 , n199531 , n199532 , n32256 , n199534 , n199535 , n32259 , n199537 , n199538 , 
 n32262 , n199540 , n199541 , n32265 , n199543 , n32267 , n32268 , n199546 , n199547 , n32271 , 
 n199549 , n199550 , n32274 , n199552 , n199553 , n32277 , n199555 , n199556 , n32280 , n199558 , 
 n199559 , n32283 , n199561 , n32285 , n32286 , n199564 , n199565 , n32289 , n199567 , n199568 , 
 n32292 , n199570 , n199571 , n32295 , n32296 , n199574 , n199575 , n32299 , n199577 , n199578 , 
 n32302 , n199580 , n199581 , n32305 , n199583 , n32307 , n32308 , n199586 , n199587 , n32311 , 
 n199589 , n199590 , n32314 , n199592 , n199593 , n32317 , n199595 , n199596 , n32320 , n199598 , 
 n199599 , n32323 , n32324 , n32325 , n199603 , n199604 , n32328 , n32329 , n199607 , n199608 , 
 n32332 , n199610 , n199611 , n32335 , n199613 , n199614 , n199615 , n199616 , n32340 , n199618 , 
 n199619 , n32343 , n199621 , n32345 , n32346 , n199624 , n199625 , n32349 , n199627 , n199628 , 
 n32352 , n199630 , n199631 , n32355 , n199633 , n199634 , n32358 , n199636 , n199637 , n32361 , 
 n199639 , n32363 , n32364 , n199642 , n199643 , n32367 , n199645 , n199646 , n32370 , n199648 , 
 n199649 , n32373 , n32374 , n32375 , n199653 , n199654 , n199655 , n199656 , n32380 , n199658 , 
 n199659 , n32383 , n199661 , n32385 , n32386 , n199664 , n199665 , n32389 , n199667 , n199668 , 
 n32392 , n199670 , n199671 , n199672 , n199673 , n32397 , n199675 , n199676 , n32400 , n199678 , 
 n32402 , n32403 , n199681 , n199682 , n32406 , n199684 , n199685 , n32409 , n199687 , n199688 , 
 n32412 , n199690 , n199691 , n32415 , n199693 , n199694 , n32418 , n199696 , n32420 , n32421 , 
 n199699 , n199700 , n32424 , n199702 , n199703 , n32427 , n199705 , n199706 , n32430 , n32431 , 
 n32432 , n199710 , n199711 , n32435 , n199713 , n199714 , n32438 , n199716 , n32440 , n199718 , 
 n199719 , n32443 , n199721 , n32445 , n199723 , n32447 , n32448 , n199726 , n199727 , n32451 , 
 n199729 , n199730 , n32454 , n199732 , n199733 , n32457 , n199735 , n199736 , n32460 , n199738 , 
 n199739 , n32463 , n199741 , n32465 , n32466 , n199744 , n199745 , n32469 , n199747 , n199748 , 
 n32472 , n199750 , n199751 , n32475 , n32476 , n32477 , n199755 , n199756 , n32480 , n32481 , 
 n32482 , n199760 , n199761 , n32485 , n32486 , n32487 , n199765 , n32489 , n32490 , n199768 , 
 n32492 , n32493 , n32494 , n199772 , n199773 , n32497 , n32498 , n199776 , n199777 , n32501 , 
 n32502 , n32503 , n199781 , n199782 , n32506 , n199784 , n199785 , n199786 , n199787 , n32511 , 
 n199789 , n199790 , n32514 , n199792 , n199793 , n32517 , n32518 , n199796 , n199797 , n32521 , 
 n32522 , n32523 , n199801 , n32525 , n32526 , n32527 , n199805 , n32529 , n32530 , n32531 , 
 n32532 , n32533 , n32534 , n199812 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , 
 n32542 , n32543 , n32544 , n32545 , n199823 , n32547 , n32548 , n32549 , n32550 , n32551 , 
 n32552 , n32553 , n32554 , n199832 , n32556 , n32557 , n32558 , n32559 , n32560 , n199838 , 
 n199839 , n32563 , n32564 , n32565 , n32566 , n199844 , n199845 , n32569 , n32570 , n32571 , 
 n32572 , n199850 , n199851 , n32575 , n199853 , n32577 , n199855 , n32579 , n32580 , n199858 , 
 n199859 , n32583 , n199861 , n199862 , n32586 , n199864 , n199865 , n199866 , n32590 , n199868 , 
 n32592 , n32593 , n199871 , n199872 , n32596 , n199874 , n199875 , n32599 , n199877 , n199878 , 
 n32602 , n199880 , n32604 , n199882 , n32606 , n32607 , n199885 , n199886 , n32610 , n199888 , 
 n199889 , n32613 , n199891 , n199892 , n32616 , n199894 , n199895 , n32619 , n199897 , n199898 , 
 n32622 , n32623 , n32624 , n32625 , n199903 , n199904 , n32628 , n199906 , n199907 , n32631 , 
 n199909 , n199910 , n199911 , n32635 , n199913 , n32637 , n32638 , n199916 , n199917 , n32641 , 
 n199919 , n199920 , n32644 , n199922 , n199923 , n32647 , n199925 , n32649 , n199927 , n32651 , 
 n32652 , n199930 , n199931 , n32655 , n199933 , n199934 , n32658 , n199936 , n199937 , n32661 , 
 n199939 , n199940 , n199941 , n32665 , n199943 , n199944 , n199945 , n32669 , n199947 , n32671 , 
 n32672 , n199950 , n199951 , n32675 , n199953 , n199954 , n32678 , n199956 , n199957 , n32681 , 
 n199959 , n199960 , n32684 , n199962 , n32686 , n199964 , n199965 , n199966 , n199967 , n32691 , 
 n199969 , n199970 , n32694 , n199972 , n199973 , n32697 , n199975 , n199976 , n32700 , n32701 , 
 n32702 , n32703 , n32704 , n199982 , n199983 , n32707 , n199985 , n199986 , n32710 , n199988 , 
 n199989 , n32713 , n32714 , n32715 , n32716 , n32717 , n199995 , n199996 , n32720 , n199998 , 
 n32722 , n32723 , n200001 , n200002 , n32726 , n200004 , n200005 , n200006 , n32730 , n200008 , 
 n200009 , n32733 , n200011 , n200012 , n32736 , n32737 , n200015 , n32739 , n32740 , n200018 , 
 n200019 , n32743 , n32744 , n32745 , n32746 , n32747 , n200025 , n200026 , n32750 , n200028 , 
 n200029 , n32753 , n32754 , n32755 , n32756 , n200034 , n200035 , n32759 , n32760 , n32761 , 
 n32762 , n200040 , n200041 , n32765 , n32766 , n32767 , n32768 , n200046 , n200047 , n32771 , 
 n32772 , n32773 , n200051 , n200052 , n32776 , n200054 , n200055 , n32779 , n32780 , n32781 , 
 n32782 , n32783 , n200061 , n200062 , n32786 , n200064 , n200065 , n32789 , n32790 , n32791 , 
 n32792 , n32793 , n200071 , n200072 , n32796 , n200074 , n32798 , n32799 , n32800 , n32801 , 
 n32802 , n200080 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , 
 n32812 , n200090 , n200091 , n32815 , n32816 , n200094 , n200095 , n32819 , n32820 , n32821 , 
 n32822 , n200100 , n200101 , n32825 , n32826 , n32827 , n200105 , n200106 , n32830 , n200108 , 
 n200109 , n32833 , n32834 , n32835 , n32836 , n32837 , n200115 , n200116 , n32840 , n32841 , 
 n32842 , n200120 , n32844 , n32845 , n200123 , n200124 , n32848 , n32849 , n200127 , n200128 , 
 n32852 , n32853 , n32854 , n32855 , n32856 , n200134 , n200135 , n32859 , n200137 , n32861 , 
 n32862 , n32863 , n200141 , n32865 , n32866 , n32867 , n32868 , n200146 , n32870 , n32871 , 
 n32872 , n32873 , n32874 , n32875 , n200153 , n200154 , n32878 , n200156 , n200157 , n32881 , 
 n32882 , n32883 , n200161 , n32885 , n32886 , n200164 , n32888 , n200166 , n32890 , n32891 , 
 n200169 , n200170 , n32894 , n200172 , n200173 , n32897 , n200175 , n200176 , n200177 , n32901 , 
 n200179 , n32903 , n32904 , n200182 , n200183 , n32907 , n200185 , n200186 , n32910 , n200188 , 
 n200189 , n32913 , n200191 , n32915 , n200193 , n32917 , n32918 , n32919 , n200197 , n200198 , 
 n32922 , n200200 , n200201 , n32925 , n200203 , n200204 , n32928 , n32929 , n32930 , n200208 , 
 n200209 , n32933 , n200211 , n200212 , n32936 , n32937 , n200215 , n32939 , n200217 , n200218 , 
 n200219 , n32943 , n200221 , n32945 , n32946 , n200224 , n200225 , n32949 , n200227 , n200228 , 
 n32952 , n200230 , n200231 , n200232 , n32956 , n200234 , n32958 , n32959 , n200237 , n200238 , 
 n32962 , n200240 , n200241 , n32965 , n200243 , n200244 , n32968 , n200246 , n32970 , n200248 , 
 n32972 , n32973 , n200251 , n200252 , n32976 , n200254 , n200255 , n32979 , n200257 , n200258 , 
 n32982 , n200260 , n200261 , n32985 , n32986 , n32987 , n200265 , n200266 , n32990 , n32991 , 
 n200269 , n200270 , n32994 , n32995 , n32996 , n200274 , n200275 , n32999 , n33000 , n33001 , 
 n200279 , n200280 , n33004 , n33005 , n200283 , n200284 , n33008 , n200286 , n200287 , n33011 , 
 n200289 , n200290 , n33014 , n33015 , n33016 , n33017 , n200295 , n200296 , n33020 , n33021 , 
 n33022 , n200300 , n200301 , n33025 , n200303 , n200304 , n33028 , n200306 , n33030 , n33031 , 
 n200309 , n200310 , n33034 , n200312 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , 
 n33042 , n33043 , n200321 , n33045 , n200323 , n200324 , n33048 , n33049 , n33050 , n33051 , 
 n33052 , n200330 , n200331 , n33055 , n200333 , n200334 , n33058 , n33059 , n33060 , n33061 , 
 n33062 , n33063 , n200341 , n33065 , n33066 , n33067 , n200345 , n200346 , n33070 , n33071 , 
 n33072 , n33073 , n200351 , n200352 , n200353 , n200354 , n200355 , n33079 , n200357 , n200358 , 
 n200359 , n33083 , n200361 , n33085 , n33086 , n200364 , n200365 , n33089 , n200367 , n200368 , 
 n33092 , n200370 , n200371 , n33095 , n200373 , n33097 , n200375 , n33099 , n33100 , n200378 , 
 n200379 , n33103 , n200381 , n200382 , n33106 , n200384 , n200385 , n33109 , n33110 , n33111 , 
 n200389 , n200390 , n33114 , n200392 , n33116 , n200394 , n33118 , n33119 , n200397 , n200398 , 
 n33122 , n200400 , n200401 , n33125 , n200403 , n200404 , n200405 , n33129 , n200407 , n33131 , 
 n33132 , n200410 , n200411 , n33135 , n200413 , n200414 , n33138 , n200416 , n200417 , n33141 , 
 n200419 , n33143 , n200421 , n33145 , n33146 , n200424 , n200425 , n33149 , n200427 , n200428 , 
 n33152 , n200430 , n200431 , n33155 , n33156 , n33157 , n200435 , n200436 , n33160 , n200438 , 
 n200439 , n33163 , n33164 , n33165 , n200443 , n200444 , n33168 , n33169 , n33170 , n33171 , 
 n200449 , n200450 , n33174 , n33175 , n33176 , n200454 , n200455 , n33179 , n33180 , n33181 , 
 n200459 , n200460 , n33184 , n200462 , n200463 , n33187 , n33188 , n33189 , n200467 , n200468 , 
 n33192 , n33193 , n200471 , n200472 , n33196 , n33197 , n200475 , n200476 , n33200 , n33201 , 
 n33202 , n33203 , n33204 , n200482 , n200483 , n33207 , n200485 , n200486 , n33210 , n33211 , 
 n33212 , n33213 , n33214 , n200492 , n200493 , n33217 , n33218 , n33219 , n200497 , n200498 , 
 n33222 , n33223 , n33224 , n200502 , n200503 , n33227 , n33228 , n33229 , n33230 , n33231 , 
 n200509 , n200510 , n33234 , n33235 , n200513 , n200514 , n33238 , n33239 , n33240 , n33241 , 
 n200519 , n200520 , n33244 , n33245 , n33246 , n200524 , n200525 , n33249 , n200527 , n200528 , 
 n33252 , n33253 , n33254 , n200532 , n200533 , n33257 , n200535 , n200536 , n33260 , n33261 , 
 n33262 , n200540 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n200547 , n200548 , 
 n33272 , n200550 , n200551 , n200552 , n200553 , n33277 , n200555 , n200556 , n33280 , n200558 , 
 n200559 , n33283 , n200561 , n200562 , n33286 , n200564 , n200565 , n33289 , n200567 , n33291 , 
 n200569 , n33293 , n200571 , n33295 , n33296 , n200574 , n200575 , n33299 , n200577 , n200578 , 
 n33302 , n200580 , n200581 , n200582 , n33306 , n33307 , n200585 , n33309 , n200587 , n200588 , 
 n33312 , n33313 , n200591 , n200592 , n33316 , n33317 , n200595 , n200596 , n33320 , n33321 , 
 n33322 , n33323 , n200601 , n200602 , n33326 , n33327 , n33328 , n33329 , n33330 , n200608 , 
 n33332 , n33333 , n33334 , n200612 , n200613 , n33337 , n33338 , n33339 , n200617 , n200618 , 
 n33342 , n33343 , n33344 , n200622 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , 
 n200629 , n200630 , n33354 , n33355 , n33356 , n33357 , n200635 , n200636 , n33360 , n33361 , 
 n33362 , n200640 , n200641 , n33365 , n33366 , n33367 , n33368 , n200646 , n200647 , n33371 , 
 n33372 , n33373 , n200651 , n200652 , n33376 , n200654 , n200655 , n33379 , n200657 , n33381 , 
 n33382 , n33383 , n33384 , n33385 , n200663 , n33387 , n33388 , n33389 , n33390 , n33391 , 
 n33392 , n33393 , n200671 , n33395 , n200673 , n33397 , n200675 , n33399 , n33400 , n200678 , 
 n200679 , n33403 , n33404 , n200682 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , 
 n33412 , n33413 , n200691 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , 
 n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , 
 n200709 , n33433 , n33434 , n33435 , n200713 , n200714 , n33438 , n33439 , n33440 , n33441 , 
 n200719 , n200720 , n33444 , n33445 , n33446 , n200724 , n200725 , n33449 , n33450 , n33451 , 
 n200729 , n33453 , n33454 , n33455 , n33456 , n33457 , n200735 , n33459 , n33460 , n33461 , 
 n33462 , n33463 , n33464 , n33465 , n200743 , n33467 , n33468 , n200746 , n200747 , n33471 , 
 n33472 , n33473 , n33474 , n33475 , n200753 , n33477 , n33478 , n200756 , n200757 , n33481 , 
 n33482 , n33483 , n33484 , n33485 , n200763 , n200764 , n33488 , n33489 , n33490 , n200768 , 
 n200769 , n33493 , n33494 , n200772 , n200773 , n33497 , n33498 , n33499 , n200777 , n200778 , 
 n33502 , n33503 , n33504 , n200782 , n200783 , n33507 , n200785 , n33509 , n33510 , n33511 , 
 n200789 , n200790 , n33514 , n33515 , n33516 , n33517 , n200795 , n33519 , n33520 , n33521 , 
 n200799 , n200800 , n33524 , n33525 , n33526 , n200804 , n200805 , n33529 , n33530 , n33531 , 
 n33532 , n200810 , n200811 , n33535 , n33536 , n200814 , n200815 , n33539 , n33540 , n33541 , 
 n200819 , n200820 , n33544 , n33545 , n33546 , n200824 , n200825 , n33549 , n33550 , n33551 , 
 n200829 , n200830 , n33554 , n33555 , n33556 , n200834 , n33558 , n33559 , n33560 , n33561 , 
 n33562 , n33563 , n33564 , n33565 , n200843 , n33567 , n33568 , n33569 , n33570 , n33571 , 
 n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , 
 n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , 
 n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , 
 n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n200885 , n200886 , n33610 , n33611 , 
 n33612 , n33613 , n200891 , n200892 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , 
 n33622 , n33623 , n33624 , n33625 , n33626 , n200904 , n33628 , n33629 , n33630 , n200908 , 
 n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , 
 n33642 , n33643 , n33644 , n33645 , n200923 , n33647 , n33648 , n33649 , n33650 , n200928 , 
 n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n200935 , n33659 , n33660 , n200938 , 
 n200939 , n33663 , n33664 , n200942 , n200943 , n33667 , n33668 , n33669 , n33670 , n200948 , 
 n200949 , n33673 , n33674 , n33675 , n200953 , n200954 , n33678 , n200956 , n33680 , n33681 , 
 n33682 , n33683 , n33684 , n200962 , n200963 , n33687 , n33688 , n200966 , n200967 , n33691 , 
 n33692 , n200970 , n200971 , n33695 , n33696 , n33697 , n200975 , n33699 , n33700 , n33701 , 
 n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n200987 , n200988 , 
 n33712 , n200990 , n200991 , n33715 , n200993 , n33717 , n33718 , n200996 , n200997 , n33721 , 
 n200999 , n201000 , n33724 , n201002 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , 
 n33732 , n33733 , n33734 , n201012 , n33736 , n201014 , n201015 , n33739 , n201017 , n33741 , 
 n33742 , n201020 , n201021 , n33745 , n201023 , n201024 , n33748 , n201026 , n33750 , n201028 , 
 n33752 , n33753 , n201031 , n201032 , n33756 , n201034 , n201035 , n33759 , n201037 , n201038 , 
 n33762 , n33763 , n201041 , n33765 , n201043 , n33767 , n33768 , n201046 , n201047 , n33771 , 
 n201049 , n201050 , n33774 , n201052 , n201053 , n33777 , n33778 , n33779 , n201057 , n201058 , 
 n33782 , n201060 , n33784 , n33785 , n201063 , n201064 , n33788 , n201066 , n201067 , n33791 , 
 n201069 , n33793 , n33794 , n201072 , n201073 , n33797 , n201075 , n201076 , n33800 , n201078 , 
 n201079 , n201080 , n33804 , n201082 , n201083 , n33807 , n201085 , n33809 , n33810 , n201088 , 
 n201089 , n33813 , n201091 , n201092 , n33816 , n201094 , n33818 , n201096 , n201097 , n33821 , 
 n201099 , n201100 , n33824 , n201102 , n33826 , n33827 , n201105 , n201106 , n33830 , n201108 , 
 n201109 , n33833 , n201111 , n33835 , n201113 , n201114 , n33838 , n201116 , n33840 , n33841 , 
 n33842 , n201120 , n33844 , n201122 , n33846 , n33847 , n201125 , n201126 , n33850 , n201128 , 
 n201129 , n33853 , n201131 , n201132 , n201133 , n201134 , n33858 , n201136 , n201137 , n33861 , 
 n201139 , n33863 , n33864 , n201142 , n201143 , n33867 , n201145 , n201146 , n33870 , n201148 , 
 n201149 , n33873 , n201151 , n201152 , n33876 , n201154 , n201155 , n33879 , n201157 , n33881 , 
 n33882 , n201160 , n201161 , n33885 , n201163 , n201164 , n33888 , n201166 , n201167 , n33891 , 
 n33892 , n33893 , n201171 , n33895 , n33896 , n33897 , n201175 , n201176 , n33900 , n201178 , 
 n201179 , n33903 , n201181 , n33905 , n33906 , n201184 , n201185 , n33909 , n201187 , n201188 , 
 n33912 , n201190 , n201191 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n201198 , 
 n33922 , n201200 , n201201 , n33925 , n201203 , n33927 , n33928 , n33929 , n33930 , n33931 , 
 n201209 , n33933 , n33934 , n33935 , n201213 , n201214 , n33938 , n201216 , n33940 , n33941 , 
 n33942 , n33943 , n33944 , n201222 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , 
 n201229 , n33953 , n33954 , n33955 , n201233 , n33957 , n201235 , n33959 , n33960 , n201238 , 
 n201239 , n33963 , n201241 , n201242 , n33966 , n201244 , n33968 , n33969 , n33970 , n33971 , 
 n33972 , n33973 , n33974 , n33975 , n33976 , n201254 , n33978 , n33979 , n33980 , n201258 , 
 n33982 , n201260 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , 
 n201269 , n33993 , n33994 , n33995 , n201273 , n201274 , n33998 , n33999 , n34000 , n201278 , 
 n201279 , n34003 , n34004 , n34005 , n201283 , n201284 , n34008 , n34009 , n34010 , n201288 , 
 n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n201295 , n34019 , n34020 , n34021 , 
 n34022 , n201300 , n201301 , n34025 , n201303 , n34027 , n201305 , n34029 , n34030 , n34031 , 
 n34032 , n201310 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n201318 , 
 n34042 , n34043 , n34044 , n34045 , n201323 , n34047 , n34048 , n34049 , n201327 , n201328 , 
 n34052 , n34053 , n34054 , n201332 , n34056 , n34057 , n34058 , n34059 , n201337 , n34061 , 
 n34062 , n34063 , n34064 , n34065 , n201343 , n34067 , n34068 , n34069 , n34070 , n34071 , 
 n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , 
 n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , 
 n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , 
 n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , 
 n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , 
 n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n201406 , n201407 , n34131 , 
 n201409 , n201410 , n34134 , n201412 , n34136 , n34137 , n201415 , n201416 , n34140 , n201418 , 
 n201419 , n34143 , n201421 , n34145 , n201423 , n201424 , n34148 , n201426 , n201427 , n34151 , 
 n201429 , n34153 , n34154 , n201432 , n201433 , n34157 , n201435 , n201436 , n34160 , n201438 , 
 n34162 , n34163 , n34164 , n201442 , n201443 , n34167 , n201445 , n34169 , n201447 , n201448 , 
 n201449 , n201450 , n34174 , n201452 , n201453 , n201454 , n34178 , n201456 , n34180 , n201458 , 
 n201459 , n34183 , n201461 , n201462 , n34186 , n201464 , n34188 , n34189 , n201467 , n201468 , 
 n34192 , n201470 , n201471 , n34195 , n201473 , n34197 , n34198 , n34199 , n34200 , n34201 , 
 n34202 , n34203 , n201481 , n201482 , n34206 , n201484 , n34208 , n34209 , n34210 , n34211 , 
 n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n201498 , 
 n34222 , n34223 , n34224 , n201502 , n201503 , n34227 , n34228 , n34229 , n201507 , n34231 , 
 n201509 , n34233 , n34234 , n201512 , n34236 , n34237 , n34238 , n201516 , n34240 , n34241 , 
 n34242 , n201520 , n201521 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n201528 , 
 n201529 , n34253 , n34254 , n34255 , n201533 , n34257 , n34258 , n201536 , n201537 , n34261 , 
 n34262 , n201540 , n201541 , n34265 , n34266 , n201544 , n201545 , n34269 , n34270 , n201548 , 
 n201549 , n34273 , n34274 , n201552 , n201553 , n201554 , n201555 , n34279 , n201557 , n201558 , 
 n34282 , n201560 , n34284 , n34285 , n201563 , n201564 , n201565 , n34289 , n201567 , n201568 , 
 n34292 , n201570 , n201571 , n34295 , n201573 , n201574 , n201575 , n34299 , n201577 , n34301 , 
 n34302 , n201580 , n201581 , n201582 , n34306 , n201584 , n201585 , n34309 , n201587 , n201588 , 
 n34312 , n201590 , n201591 , n34315 , n201593 , n201594 , n34318 , n201596 , n34320 , n201598 , 
 n201599 , n201600 , n201601 , n34325 , n201603 , n201604 , n201605 , n34329 , n201607 , n201608 , 
 n34332 , n201610 , n201611 , n34335 , n201613 , n34337 , n201615 , n34339 , n34340 , n201618 , 
 n201619 , n201620 , n34344 , n201622 , n201623 , n34347 , n201625 , n201626 , n34350 , n201628 , 
 n201629 , n201630 , n34354 , n201632 , n34356 , n34357 , n201635 , n201636 , n201637 , n34361 , 
 n201639 , n201640 , n34364 , n201642 , n201643 , n34367 , n201645 , n201646 , n34370 , n34371 , 
 n201649 , n201650 , n34374 , n201652 , n34376 , n34377 , n201655 , n34379 , n201657 , n34381 , 
 n34382 , n201660 , n34384 , n34385 , n34386 , n201664 , n201665 , n34389 , n34390 , n34391 , 
 n201669 , n201670 , n201671 , n201672 , n34396 , n201674 , n201675 , n34399 , n201677 , n201678 , 
 n34402 , n201680 , n201681 , n34405 , n201683 , n34407 , n34408 , n201686 , n201687 , n201688 , 
 n34412 , n201690 , n201691 , n34415 , n201693 , n201694 , n34418 , n201696 , n201697 , n34421 , 
 n34422 , n201700 , n201701 , n34425 , n201703 , n34427 , n201705 , n34429 , n34430 , n201708 , 
 n201709 , n34433 , n201711 , n201712 , n34436 , n201714 , n201715 , n34439 , n201717 , n201718 , 
 n34442 , n201720 , n201721 , n201722 , n201723 , n34447 , n201725 , n201726 , n34450 , n201728 , 
 n34452 , n34453 , n201731 , n201732 , n201733 , n34457 , n201735 , n201736 , n34460 , n201738 , 
 n201739 , n34463 , n201741 , n201742 , n34466 , n201744 , n201745 , n34469 , n201747 , n201748 , 
 n34472 , n201750 , n34474 , n34475 , n201753 , n201754 , n201755 , n34479 , n201757 , n201758 , 
 n34482 , n201760 , n201761 , n34485 , n201763 , n201764 , n34488 , n34489 , n201767 , n201768 , 
 n34492 , n201770 , n201771 , n34495 , n201773 , n201774 , n34498 , n201776 , n34500 , n34501 , 
 n201779 , n201780 , n201781 , n34505 , n201783 , n201784 , n34508 , n201786 , n201787 , n34511 , 
 n201789 , n201790 , n34514 , n201792 , n201793 , n34517 , n201795 , n201796 , n34520 , n201798 , 
 n34522 , n201800 , n34524 , n34525 , n201803 , n201804 , n34528 , n201806 , n201807 , n34531 , 
 n201809 , n201810 , n201811 , n201812 , n34536 , n201814 , n201815 , n34539 , n201817 , n34541 , 
 n34542 , n201820 , n201821 , n34545 , n201823 , n201824 , n34548 , n201826 , n201827 , n34551 , 
 n201829 , n34553 , n201831 , n34555 , n34556 , n201834 , n201835 , n34559 , n201837 , n201838 , 
 n34562 , n201840 , n201841 , n34565 , n201843 , n201844 , n34568 , n201846 , n201847 , n34571 , 
 n201849 , n201850 , n201851 , n34575 , n201853 , n201854 , n34578 , n34579 , n201857 , n34581 , 
 n201859 , n201860 , n34584 , n34585 , n201863 , n201864 , n201865 , n34589 , n34590 , n201868 , 
 n34592 , n201870 , n201871 , n34595 , n34596 , n201874 , n201875 , n34599 , n34600 , n34601 , 
 n34602 , n201880 , n201881 , n201882 , n34606 , n201884 , n201885 , n34609 , n201887 , n34611 , 
 n201889 , n201890 , n34614 , n201892 , n34616 , n34617 , n34618 , n201896 , n201897 , n201898 , 
 n34622 , n201900 , n201901 , n34625 , n201903 , n34627 , n34628 , n201906 , n201907 , n34631 , 
 n201909 , n34633 , n34634 , n34635 , n201913 , n201914 , n201915 , n34639 , n201917 , n201918 , 
 n34642 , n201920 , n34644 , n34645 , n201923 , n34647 , n34648 , n201926 , n201927 , n34651 , 
 n201929 , n201930 , n34654 , n201932 , n201933 , n34657 , n201935 , n34659 , n34660 , n201938 , 
 n201939 , n34663 , n201941 , n201942 , n201943 , n34667 , n201945 , n201946 , n34670 , n201948 , 
 n201949 , n201950 , n34674 , n201952 , n34676 , n34677 , n201955 , n201956 , n201957 , n34681 , 
 n201959 , n201960 , n34684 , n201962 , n201963 , n34687 , n201965 , n201966 , n34690 , n201968 , 
 n34692 , n201970 , n34694 , n34695 , n201973 , n34697 , n201975 , n34699 , n201977 , n201978 , 
 n34702 , n201980 , n201981 , n34705 , n201983 , n201984 , n34708 , n201986 , n201987 , n34711 , 
 n201989 , n201990 , n34714 , n34715 , n34716 , n201994 , n201995 , n34719 , n34720 , n34721 , 
 n201999 , n202000 , n34724 , n202002 , n34726 , n34727 , n34728 , n34729 , n202007 , n202008 , 
 n34732 , n202010 , n34734 , n34735 , n34736 , n34737 , n34738 , n202016 , n202017 , n34741 , 
 n202019 , n34743 , n34744 , n34745 , n34746 , n34747 , n202025 , n34749 , n34750 , n202028 , 
 n34752 , n34753 , n34754 , n34755 , n202033 , n202034 , n34758 , n202036 , n34760 , n34761 , 
 n34762 , n202040 , n34764 , n202042 , n34766 , n34767 , n202045 , n202046 , n34770 , n202048 , 
 n202049 , n34773 , n202051 , n34775 , n34776 , n34777 , n202055 , n34779 , n202057 , n34781 , 
 n34782 , n202060 , n202061 , n34785 , n202063 , n202064 , n34788 , n202066 , n34790 , n34791 , 
 n34792 , n202070 , n34794 , n34795 , n34796 , n202074 , n202075 , n34799 , n34800 , n34801 , 
 n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , 
 n34812 , n34813 , n34814 , n202092 , n34816 , n202094 , n34818 , n202096 , n202097 , n34821 , 
 n34822 , n202100 , n34824 , n202102 , n34826 , n202104 , n202105 , n34829 , n34830 , n202108 , 
 n34832 , n202110 , n34834 , n34835 , n202113 , n202114 , n34838 , n202116 , n202117 , n34841 , 
 n202119 , n202120 , n202121 , n34845 , n202123 , n34847 , n34848 , n202126 , n202127 , n34851 , 
 n202129 , n202130 , n34854 , n202132 , n202133 , n34857 , n202135 , n34859 , n202137 , n34861 , 
 n34862 , n202140 , n202141 , n34865 , n202143 , n202144 , n34868 , n202146 , n202147 , n34871 , 
 n202149 , n202150 , n202151 , n34875 , n202153 , n34877 , n34878 , n202156 , n202157 , n34881 , 
 n202159 , n202160 , n34884 , n202162 , n202163 , n34887 , n202165 , n34889 , n34890 , n202168 , 
 n202169 , n34893 , n202171 , n202172 , n34896 , n202174 , n34898 , n202176 , n34900 , n202178 , 
 n34902 , n34903 , n202181 , n202182 , n34906 , n202184 , n202185 , n34909 , n202187 , n34911 , 
 n202189 , n34913 , n202191 , n34915 , n202193 , n34917 , n34918 , n202196 , n202197 , n34921 , 
 n202199 , n202200 , n34924 , n202202 , n202203 , n34927 , n202205 , n34929 , n34930 , n202208 , 
 n202209 , n34933 , n202211 , n202212 , n34936 , n202214 , n34938 , n202216 , n202217 , n34941 , 
 n202219 , n202220 , n34944 , n34945 , n202223 , n34947 , n202225 , n34949 , n202227 , n202228 , 
 n34952 , n202230 , n202231 , n34955 , n202233 , n202234 , n34958 , n202236 , n34960 , n202238 , 
 n34962 , n202240 , n202241 , n34965 , n34966 , n202244 , n34968 , n202246 , n202247 , n34971 , 
 n34972 , n34973 , n34974 , n34975 , n202253 , n34977 , n202255 , n202256 , n34980 , n34981 , 
 n34982 , n34983 , n202261 , n202262 , n34986 , n34987 , n34988 , n34989 , n34990 , n202268 , 
 n202269 , n34993 , n202271 , n202272 , n34996 , n34997 , n34998 , n202276 , n202277 , n35001 , 
 n35002 , n35003 , n35004 , n35005 , n202283 , n202284 , n202285 , n35009 , n202287 , n35011 , 
 n35012 , n202290 , n202291 , n35015 , n202293 , n35017 , n202295 , n202296 , n35020 , n202298 , 
 n35022 , n35023 , n35024 , n35025 , n35026 , n202304 , n202305 , n35029 , n202307 , n35031 , 
 n35032 , n35033 , n35034 , n35035 , n202313 , n202314 , n35038 , n202316 , n35040 , n35041 , 
 n35042 , n35043 , n202321 , n202322 , n35046 , n202324 , n35048 , n202326 , n35050 , n35051 , 
 n202329 , n35053 , n35054 , n35055 , n35056 , n35057 , n202335 , n35059 , n35060 , n35061 , 
 n35062 , n35063 , n202341 , n35065 , n35066 , n202344 , n35068 , n35069 , n35070 , n35071 , 
 n35072 , n202350 , n202351 , n35075 , n202353 , n202354 , n35078 , n35079 , n202357 , n35081 , 
 n35082 , n202360 , n202361 , n35085 , n202363 , n202364 , n35088 , n35089 , n35090 , n202368 , 
 n202369 , n202370 , n35094 , n202372 , n35096 , n202374 , n202375 , n35099 , n35100 , n202378 , 
 n202379 , n35103 , n35104 , n202382 , n202383 , n202384 , n35108 , n35109 , n202387 , n35111 , 
 n35112 , n202390 , n202391 , n35115 , n202393 , n202394 , n35118 , n35119 , n35120 , n202398 , 
 n35122 , n202400 , n202401 , n202402 , n202403 , n35127 , n202405 , n202406 , n35130 , n202408 , 
 n202409 , n35133 , n202411 , n202412 , n35136 , n35137 , n35138 , n202416 , n35140 , n35141 , 
 n35142 , n35143 , n35144 , n202422 , n202423 , n35147 , n202425 , n35149 , n35150 , n202428 , 
 n202429 , n35153 , n35154 , n202432 , n202433 , n202434 , n35158 , n35159 , n35160 , n202438 , 
 n35162 , n35163 , n202441 , n202442 , n35166 , n35167 , n35168 , n35169 , n35170 , n202448 , 
 n202449 , n35173 , n202451 , n202452 , n35176 , n35177 , n35178 , n35179 , n202457 , n202458 , 
 n35182 , n35183 , n35184 , n202462 , n202463 , n35187 , n202465 , n35189 , n202467 , n202468 , 
 n35192 , n35193 , n35194 , n35195 , n202473 , n35197 , n202475 , n202476 , n202477 , n35201 , 
 n202479 , n202480 , n35204 , n202482 , n202483 , n35207 , n35208 , n35209 , n35210 , n202488 , 
 n202489 , n35213 , n202491 , n35215 , n202493 , n202494 , n35218 , n202496 , n35220 , n202498 , 
 n35222 , n202500 , n202501 , n35225 , n202503 , n35227 , n35228 , n35229 , n35230 , n35231 , 
 n35232 , n202510 , n202511 , n35235 , n35236 , n35237 , n35238 , n202516 , n202517 , n35241 , 
 n35242 , n35243 , n202521 , n202522 , n202523 , n35247 , n202525 , n35249 , n35250 , n202528 , 
 n202529 , n35253 , n35254 , n202532 , n202533 , n202534 , n35258 , n35259 , n202537 , n35261 , 
 n35262 , n202540 , n202541 , n35265 , n35266 , n35267 , n202545 , n202546 , n35270 , n202548 , 
 n202549 , n35273 , n202551 , n35275 , n35276 , n35277 , n35278 , n35279 , n202557 , n35281 , 
 n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n202566 , n35290 , n35291 , 
 n202569 , n202570 , n35294 , n35295 , n202573 , n202574 , n35298 , n35299 , n35300 , n35301 , 
 n35302 , n202580 , n202581 , n35305 , n202583 , n35307 , n35308 , n35309 , n202587 , n35311 , 
 n35312 , n35313 , n35314 , n202592 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , 
 n202599 , n35323 , n35324 , n202602 , n202603 , n35327 , n202605 , n35329 , n35330 , n202608 , 
 n202609 , n35333 , n202611 , n202612 , n35336 , n202614 , n202615 , n202616 , n35340 , n202618 , 
 n35342 , n35343 , n202621 , n202622 , n35346 , n202624 , n202625 , n35349 , n202627 , n202628 , 
 n35352 , n202630 , n35354 , n202632 , n35356 , n35357 , n202635 , n202636 , n35360 , n35361 , 
 n202639 , n202640 , n35364 , n35365 , n35366 , n202644 , n202645 , n35369 , n35370 , n202648 , 
 n202649 , n35373 , n35374 , n35375 , n35376 , n35377 , n202655 , n202656 , n35380 , n35381 , 
 n35382 , n35383 , n202661 , n202662 , n35386 , n35387 , n35388 , n35389 , n35390 , n202668 , 
 n202669 , n35393 , n35394 , n35395 , n202673 , n202674 , n35398 , n35399 , n35400 , n202678 , 
 n202679 , n35403 , n35404 , n202682 , n202683 , n35407 , n202685 , n202686 , n35410 , n202688 , 
 n35412 , n202690 , n202691 , n202692 , n202693 , n35417 , n202695 , n202696 , n35420 , n202698 , 
 n202699 , n35423 , n35424 , n202702 , n35426 , n35427 , n35428 , n202706 , n202707 , n35431 , 
 n35432 , n35433 , n202711 , n202712 , n35436 , n202714 , n202715 , n35439 , n35440 , n35441 , 
 n202719 , n202720 , n35444 , n202722 , n202723 , n35447 , n35448 , n35449 , n35450 , n202728 , 
 n35452 , n202730 , n202731 , n202732 , n202733 , n35457 , n202735 , n202736 , n35460 , n202738 , 
 n202739 , n35463 , n35464 , n35465 , n202743 , n202744 , n35468 , n35469 , n35470 , n202748 , 
 n202749 , n35473 , n35474 , n35475 , n202753 , n35477 , n35478 , n35479 , n202757 , n35481 , 
 n35482 , n35483 , n35484 , n35485 , n35486 , n202764 , n35488 , n35489 , n202767 , n202768 , 
 n35492 , n35493 , n35494 , n35495 , n35496 , n202774 , n202775 , n35499 , n35500 , n35501 , 
 n202779 , n202780 , n35504 , n35505 , n202783 , n202784 , n35508 , n35509 , n35510 , n202788 , 
 n202789 , n35513 , n35514 , n35515 , n35516 , n202794 , n202795 , n35519 , n35520 , n35521 , 
 n202799 , n202800 , n35524 , n35525 , n35526 , n202804 , n202805 , n35529 , n35530 , n35531 , 
 n202809 , n35533 , n35534 , n35535 , n202813 , n35537 , n35538 , n35539 , n35540 , n35541 , 
 n35542 , n35543 , n35544 , n35545 , n202823 , n35547 , n35548 , n35549 , n35550 , n202828 , 
 n35552 , n35553 , n202831 , n35555 , n35556 , n35557 , n202835 , n35559 , n35560 , n35561 , 
 n202839 , n35563 , n35564 , n35565 , n202843 , n202844 , n35568 , n35569 , n35570 , n202848 , 
 n35572 , n35573 , n35574 , n202852 , n35576 , n35577 , n35578 , n35579 , n202857 , n35581 , 
 n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n202865 , n35589 , n35590 , n35591 , 
 n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , 
 n35602 , n202880 , n35604 , n35605 , n35606 , n35607 , n35608 , n202886 , n35610 , n35611 , 
 n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , 
 n202899 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n202908 , 
 n35632 , n35633 , n35634 , n35635 , n202913 , n202914 , n35638 , n35639 , n35640 , n35641 , 
 n35642 , n202920 , n202921 , n35645 , n35646 , n202924 , n35648 , n35649 , n35650 , n35651 , 
 n35652 , n35653 , n202931 , n35655 , n202933 , n202934 , n35658 , n35659 , n35660 , n202938 , 
 n35662 , n35663 , n202941 , n202942 , n35666 , n35667 , n35668 , n35669 , n202947 , n202948 , 
 n35672 , n35673 , n35674 , n202952 , n202953 , n35677 , n202955 , n35679 , n35680 , n35681 , 
 n202959 , n35683 , n35684 , n35685 , n35686 , n202964 , n35688 , n35689 , n35690 , n35691 , 
 n35692 , n35693 , n35694 , n202972 , n35696 , n35697 , n35698 , n35699 , n202977 , n35701 , 
 n35702 , n35703 , n35704 , n202982 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , 
 n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , 
 n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , 
 n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , 
 n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , 
 n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , 
 n203039 , n203040 , n35764 , n35765 , n35766 , n35767 , n203045 , n203046 , n35770 , n35771 , 
 n35772 , n203050 , n203051 , n35775 , n203053 , n35777 , n35778 , n35779 , n35780 , n35781 , 
 n203059 , n35783 , n35784 , n35785 , n35786 , n203064 , n203065 , n35789 , n35790 , n35791 , 
 n35792 , n203070 , n203071 , n35795 , n35796 , n35797 , n203075 , n203076 , n35800 , n35801 , 
 n35802 , n203080 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n203088 , 
 n35812 , n35813 , n35814 , n35815 , n203093 , n35817 , n35818 , n35819 , n35820 , n35821 , 
 n35822 , n35823 , n35824 , n203102 , n35826 , n35827 , n35828 , n203106 , n203107 , n35831 , 
 n203109 , n203110 , n203111 , n35835 , n203113 , n35837 , n35838 , n203116 , n203117 , n35841 , 
 n203119 , n203120 , n203121 , n35845 , n203123 , n203124 , n35848 , n203126 , n203127 , n35851 , 
 n203129 , n203130 , n35854 , n203132 , n203133 , n35857 , n203135 , n35859 , n35860 , n203138 , 
 n203139 , n203140 , n35864 , n203142 , n203143 , n35867 , n203145 , n203146 , n35870 , n203148 , 
 n203149 , n35873 , n203151 , n35875 , n203153 , n35877 , n35878 , n35879 , n203157 , n35881 , 
 n203159 , n35883 , n35884 , n203162 , n203163 , n203164 , n35888 , n203166 , n203167 , n35891 , 
 n203169 , n203170 , n35894 , n203172 , n203173 , n203174 , n203175 , n35899 , n203177 , n203178 , 
 n35902 , n203180 , n35904 , n35905 , n203183 , n203184 , n203185 , n35909 , n203187 , n203188 , 
 n35912 , n203190 , n203191 , n35915 , n203193 , n203194 , n35918 , n35919 , n35920 , n35921 , 
 n203199 , n203200 , n35924 , n203202 , n203203 , n203204 , n35928 , n203206 , n35930 , n203208 , 
 n203209 , n35933 , n203211 , n35935 , n203213 , n203214 , n203215 , n35939 , n203217 , n35941 , 
 n35942 , n35943 , n35944 , n35945 , n35946 , n203224 , n35948 , n203226 , n35950 , n35951 , 
 n35952 , n35953 , n35954 , n203232 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , 
 n35962 , n35963 , n203241 , n203242 , n35966 , n203244 , n203245 , n35969 , n203247 , n35971 , 
 n35972 , n203250 , n203251 , n35975 , n203253 , n203254 , n35978 , n203256 , n35980 , n203258 , 
 n35982 , n203260 , n35984 , n35985 , n203263 , n203264 , n35988 , n203266 , n203267 , n35991 , 
 n203269 , n203270 , n203271 , n35995 , n203273 , n35997 , n203275 , n203276 , n36000 , n203278 , 
 n203279 , n203280 , n36004 , n203282 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , 
 n36012 , n36013 , n36014 , n36015 , n36016 , n203294 , n203295 , n36019 , n203297 , n203298 , 
 n36022 , n203300 , n203301 , n36025 , n203303 , n36027 , n203305 , n36029 , n36030 , n203308 , 
 n203309 , n36033 , n203311 , n203312 , n36036 , n203314 , n203315 , n36039 , n36040 , n203318 , 
 n36042 , n203320 , n203321 , n36045 , n203323 , n36047 , n36048 , n203326 , n36050 , n203328 , 
 n36052 , n36053 , n203331 , n203332 , n36056 , n203334 , n203335 , n36059 , n203337 , n203338 , 
 n36062 , n203340 , n203341 , n36065 , n203343 , n203344 , n36068 , n203346 , n203347 , n36071 , 
 n36072 , n203350 , n36074 , n36075 , n203353 , n203354 , n36078 , n36079 , n203357 , n203358 , 
 n36082 , n36083 , n203361 , n36085 , n36086 , n36087 , n36088 , n203366 , n36090 , n203368 , 
 n36092 , n36093 , n203371 , n203372 , n36096 , n203374 , n203375 , n36099 , n203377 , n203378 , 
 n36102 , n203380 , n36104 , n36105 , n203383 , n36107 , n36108 , n36109 , n203387 , n36111 , 
 n203389 , n203390 , n36114 , n36115 , n36116 , n36117 , n203395 , n36119 , n203397 , n36121 , 
 n36122 , n36123 , n36124 , n36125 , n36126 , n203404 , n36128 , n203406 , n203407 , n36131 , 
 n203409 , n36133 , n36134 , n203412 , n203413 , n36137 , n203415 , n203416 , n36140 , n203418 , 
 n36142 , n36143 , n36144 , n36145 , n36146 , n203424 , n36148 , n36149 , n36150 , n36151 , 
 n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n203436 , n203437 , n36161 , 
 n203439 , n36163 , n203441 , n203442 , n203443 , n203444 , n36168 , n203446 , n203447 , n36171 , 
 n203449 , n203450 , n36174 , n36175 , n203453 , n203454 , n36178 , n36179 , n36180 , n203458 , 
 n203459 , n36183 , n36184 , n36185 , n203463 , n36187 , n36188 , n36189 , n36190 , n36191 , 
 n203469 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n203477 , n36201 , 
 n203479 , n36203 , n203481 , n203482 , n36206 , n203484 , n36208 , n36209 , n203487 , n36211 , 
 n203489 , n36213 , n203491 , n203492 , n36216 , n203494 , n36218 , n36219 , n36220 , n36221 , 
 n36222 , n36223 , n36224 , n203502 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , 
 n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , 
 n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , 
 n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , 
 n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , 
 n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , 
 n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , 
 n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , 
 n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , 
 n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , 
 n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , 
 n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , 
 n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , 
 n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n203636 , n36360 , n36361 , 
 n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , 
 n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , 
 n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , 
 n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , 
 n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , 
 n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , 
 n36422 , n36423 , n36424 , n36425 , n36426 , n203704 , n36428 , n36429 , n36430 , n36431 , 
 n203709 , n203710 , n36434 , n36435 , n36436 , n36437 , n203715 , n203716 , n203717 , n36441 , 
 n203719 , n36443 , n36444 , n203722 , n36446 , n203724 , n36448 , n203726 , n203727 , n36451 , 
 n203729 , n203730 , n36454 , n203732 , n36456 , n203734 , n36458 , n36459 , n36460 , n203738 , 
 n36462 , n203740 , n36464 , n203742 , n36466 , n36467 , n203745 , n203746 , n203747 , n36471 , 
 n203749 , n203750 , n36474 , n203752 , n203753 , n36477 , n203755 , n203756 , n36480 , n203758 , 
 n203759 , n36483 , n203761 , n203762 , n203763 , n36487 , n203765 , n36489 , n203767 , n203768 , 
 n203769 , n203770 , n36494 , n203772 , n203773 , n36497 , n203775 , n203776 , n36500 , n36501 , 
 n203779 , n203780 , n203781 , n36505 , n203783 , n36507 , n36508 , n203786 , n203787 , n203788 , 
 n36512 , n203790 , n203791 , n36515 , n203793 , n203794 , n36518 , n203796 , n203797 , n36521 , 
 n203799 , n36523 , n203801 , n36525 , n36526 , n203804 , n203805 , n203806 , n36530 , n203808 , 
 n203809 , n36533 , n203811 , n203812 , n36536 , n203814 , n203815 , n36539 , n203817 , n203818 , 
 n36542 , n203820 , n203821 , n36545 , n203823 , n203824 , n36548 , n36549 , n36550 , n36551 , 
 n36552 , n203830 , n203831 , n36555 , n203833 , n36557 , n36558 , n36559 , n36560 , n36561 , 
 n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , 
 n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , 
 n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , 
 n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , 
 n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , 
 n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , 
 n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , 
 n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , 
 n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , 
 n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , 
 n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , 
 n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , 
 n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , 
 n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , 
 n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , 
 n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , 
 n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , 
 n204009 , n36733 , n204011 , n36735 , n36736 , n204014 , n204015 , n204016 , n36740 , n204018 , 
 n204019 , n36743 , n204021 , n204022 , n36746 , n204024 , n204025 , n204026 , n36750 , n204028 , 
 n36752 , n36753 , n204031 , n204032 , n36756 , n204034 , n204035 , n36759 , n204037 , n36761 , 
 n204039 , n204040 , n36764 , n204042 , n204043 , n36767 , n204045 , n204046 , n36770 , n36771 , 
 n36772 , n36773 , n36774 , n204052 , n204053 , n36777 , n36778 , n36779 , n204057 , n204058 , 
 n36782 , n204060 , n204061 , n204062 , n36786 , n204064 , n36788 , n36789 , n204067 , n204068 , 
 n204069 , n36793 , n204071 , n204072 , n36796 , n204074 , n204075 , n36799 , n204077 , n204078 , 
 n36802 , n204080 , n36804 , n204082 , n36806 , n36807 , n204085 , n204086 , n36810 , n204088 , 
 n204089 , n36813 , n204091 , n204092 , n36816 , n204094 , n204095 , n36819 , n36820 , n36821 , 
 n36822 , n204100 , n204101 , n36825 , n36826 , n36827 , n204105 , n204106 , n36830 , n36831 , 
 n36832 , n204110 , n204111 , n36835 , n36836 , n36837 , n36838 , n36839 , n204117 , n204118 , 
 n36842 , n204120 , n204121 , n204122 , n36846 , n204124 , n36848 , n36849 , n204127 , n204128 , 
 n36852 , n204130 , n204131 , n36855 , n204133 , n36857 , n204135 , n204136 , n36860 , n204138 , 
 n204139 , n36863 , n204141 , n36865 , n204143 , n204144 , n36868 , n204146 , n36870 , n204148 , 
 n36872 , n36873 , n204151 , n204152 , n204153 , n36877 , n204155 , n204156 , n36880 , n204158 , 
 n204159 , n36883 , n204161 , n204162 , n204163 , n204164 , n36888 , n204166 , n36890 , n204168 , 
 n204169 , n36893 , n204171 , n36895 , n204173 , n204174 , n204175 , n36899 , n204177 , n204178 , 
 n204179 , n36903 , n204181 , n204182 , n36906 , n36907 , n204185 , n36909 , n36910 , n204188 , 
 n204189 , n36913 , n36914 , n204192 , n204193 , n36917 , n204195 , n204196 , n36920 , n204198 , 
 n204199 , n36923 , n204201 , n36925 , n36926 , n36927 , n36928 , n204206 , n204207 , n36931 , 
 n36932 , n204210 , n204211 , n36935 , n36936 , n36937 , n36938 , n36939 , n204217 , n204218 , 
 n36942 , n36943 , n36944 , n204222 , n36946 , n36947 , n36948 , n36949 , n36950 , n204228 , 
 n36952 , n36953 , n204231 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , 
 n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , 
 n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , 
 n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , 
 n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , 
 n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , 
 n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , 
 n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , 
 n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , 
 n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , 
 n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , 
 n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , 
 n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , 
 n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , 
 n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , 
 n37102 , n37103 , n37104 , n204382 , n204383 , n37107 , n37108 , n37109 , n37110 , n204388 , 
 n204389 , n37113 , n204391 , n37115 , n204393 , n204394 , n37118 , n204396 , n37120 , n37121 , 
 n204399 , n204400 , n37124 , n204402 , n204403 , n37127 , n204405 , n204406 , n37130 , n204408 , 
 n204409 , n37133 , n37134 , n37135 , n37136 , n204414 , n204415 , n37139 , n37140 , n204418 , 
 n204419 , n204420 , n37144 , n204422 , n37146 , n37147 , n204425 , n204426 , n37150 , n204428 , 
 n204429 , n37153 , n204431 , n37155 , n204433 , n204434 , n37158 , n204436 , n204437 , n37161 , 
 n204439 , n204440 , n37164 , n204442 , n204443 , n204444 , n37168 , n204446 , n204447 , n37171 , 
 n37172 , n204450 , n37174 , n37175 , n204453 , n204454 , n37178 , n37179 , n204457 , n204458 , 
 n37182 , n204460 , n204461 , n37185 , n204463 , n204464 , n37188 , n37189 , n37190 , n204468 , 
 n37192 , n204470 , n204471 , n204472 , n37196 , n204474 , n37198 , n37199 , n204477 , n37201 , 
 n204479 , n204480 , n37204 , n204482 , n204483 , n37207 , n204485 , n204486 , n204487 , n37211 , 
 n204489 , n204490 , n37214 , n37215 , n204493 , n204494 , n37218 , n204496 , n204497 , n204498 , 
 n204499 , n204500 , n37224 , n204502 , n204503 , n204504 , n37228 , n204506 , n204507 , n37231 , 
 n37232 , n204510 , n204511 , n37235 , n37236 , n37237 , n37238 , n37239 , n204517 , n204518 , 
 n37242 , n204520 , n204521 , n37245 , n37246 , n37247 , n37248 , n37249 , n204527 , n204528 , 
 n37252 , n204530 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n204537 , n37261 , 
 n37262 , n204540 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n204548 , 
 n37272 , n37273 , n37274 , n37275 , n204553 , n204554 , n204555 , n204556 , n37280 , n204558 , 
 n204559 , n204560 , n37284 , n204562 , n37286 , n204564 , n204565 , n204566 , n204567 , n37291 , 
 n204569 , n204570 , n37294 , n204572 , n204573 , n37297 , n204575 , n204576 , n37300 , n204578 , 
 n204579 , n204580 , n37304 , n37305 , n204583 , n37307 , n37308 , n204586 , n204587 , n37311 , 
 n37312 , n204590 , n204591 , n37315 , n204593 , n204594 , n37318 , n37319 , n37320 , n37321 , 
 n37322 , n204600 , n204601 , n37325 , n204603 , n37327 , n37328 , n37329 , n37330 , n37331 , 
 n204609 , n204610 , n37334 , n204612 , n204613 , n37337 , n37338 , n37339 , n37340 , n204618 , 
 n204619 , n37343 , n204621 , n204622 , n37346 , n204624 , n37348 , n204626 , n204627 , n204628 , 
 n204629 , n37353 , n204631 , n204632 , n37356 , n204634 , n204635 , n37359 , n204637 , n204638 , 
 n204639 , n37363 , n37364 , n204642 , n37366 , n37367 , n204645 , n204646 , n37370 , n37371 , 
 n204649 , n204650 , n37374 , n204652 , n204653 , n37377 , n204655 , n37379 , n37380 , n37381 , 
 n37382 , n37383 , n37384 , n204662 , n204663 , n204664 , n37388 , n204666 , n204667 , n204668 , 
 n204669 , n37393 , n204671 , n204672 , n37396 , n204674 , n204675 , n37399 , n37400 , n204678 , 
 n204679 , n37403 , n37404 , n37405 , n37406 , n37407 , n204685 , n204686 , n37410 , n204688 , 
 n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , 
 n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , 
 n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , 
 n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , 
 n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , 
 n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , 
 n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , 
 n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , 
 n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , 
 n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , 
 n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , 
 n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , 
 n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , 
 n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , 
 n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , 
 n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , 
 n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , 
 n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , 
 n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , 
 n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , 
 n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , 
 n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n204908 , 
 n37632 , n204910 , n204911 , n37635 , n204913 , n204914 , n37638 , n204916 , n204917 , n37641 , 
 n204919 , n37643 , n204921 , n204922 , n37646 , n37647 , n204925 , n204926 , n37650 , n37651 , 
 n204929 , n204930 , n37654 , n37655 , n204933 , n204934 , n37658 , n37659 , n204937 , n37661 , 
 n37662 , n37663 , n37664 , n37665 , n204943 , n37667 , n37668 , n37669 , n37670 , n37671 , 
 n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , 
 n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , 
 n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , 
 n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n204987 , n204988 , 
 n37712 , n204990 , n37714 , n37715 , n37716 , n204994 , n37718 , n204996 , n37720 , n204998 , 
 n37722 , n37723 , n205001 , n37725 , n205003 , n37727 , n37728 , n37729 , n37730 , n37731 , 
 n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n205017 , n205018 , 
 n37742 , n205020 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n205028 , 
 n205029 , n205030 , n37754 , n205032 , n205033 , n37757 , n37758 , n205036 , n37760 , n205038 , 
 n205039 , n205040 , n37764 , n37765 , n37766 , n37767 , n205045 , n37769 , n205047 , n205048 , 
 n37772 , n205050 , n205051 , n205052 , n205053 , n205054 , n37778 , n205056 , n205057 , n37781 , 
 n205059 , n205060 , n205061 , n37785 , n205063 , n205064 , n37788 , n205066 , n205067 , n37791 , 
 n205069 , n205070 , n37794 , n205072 , n37796 , n205074 , n205075 , n37799 , n205077 , n205078 , 
 n205079 , n205080 , n37804 , n205082 , n205083 , n37807 , n205085 , n205086 , n205087 , n37811 , 
 n205089 , n205090 , n37814 , n205092 , n205093 , n37817 , n205095 , n205096 , n205097 , n205098 , 
 n37822 , n205100 , n205101 , n37825 , n205103 , n37827 , n205105 , n205106 , n205107 , n205108 , 
 n37832 , n205110 , n205111 , n205112 , n37836 , n205114 , n205115 , n37839 , n205117 , n205118 , 
 n37842 , n205120 , n205121 , n37845 , n205123 , n205124 , n37848 , n205126 , n205127 , n37851 , 
 n205129 , n205130 , n37854 , n205132 , n205133 , n37857 , n205135 , n205136 , n37860 , n205138 , 
 n37862 , n205140 , n205141 , n37865 , n205143 , n205144 , n37868 , n205146 , n205147 , n37871 , 
 n205149 , n205150 , n205151 , n37875 , n205153 , n205154 , n37878 , n205156 , n205157 , n37881 , 
 n205159 , n205160 , n37884 , n37885 , n37886 , n37887 , n205165 , n205166 , n37890 , n37891 , 
 n37892 , n37893 , n205171 , n205172 , n37896 , n37897 , n205175 , n205176 , n37900 , n205178 , 
 n37902 , n37903 , n205181 , n205182 , n205183 , n37907 , n37908 , n205186 , n37910 , n205188 , 
 n205189 , n37913 , n37914 , n205192 , n205193 , n37917 , n205195 , n205196 , n37920 , n205198 , 
 n205199 , n37923 , n205201 , n37925 , n205203 , n37927 , n37928 , n205206 , n205207 , n205208 , 
 n37932 , n205210 , n205211 , n37935 , n205213 , n205214 , n37938 , n205216 , n205217 , n37941 , 
 n205219 , n205220 , n37944 , n205222 , n37946 , n37947 , n37948 , n37949 , n205227 , n37951 , 
 n37952 , n205230 , n205231 , n205232 , n37956 , n205234 , n37958 , n37959 , n205237 , n205238 , 
 n205239 , n37963 , n205241 , n205242 , n37966 , n205244 , n205245 , n37969 , n205247 , n205248 , 
 n37972 , n205250 , n37974 , n205252 , n37976 , n37977 , n205255 , n205256 , n205257 , n37981 , 
 n205259 , n205260 , n37984 , n205262 , n205263 , n37987 , n205265 , n205266 , n37990 , n205268 , 
 n205269 , n37993 , n205271 , n205272 , n37996 , n205274 , n205275 , n37999 , n38000 , n38001 , 
 n38002 , n38003 , n205281 , n205282 , n38006 , n205284 , n205285 , n38009 , n38010 , n38011 , 
 n38012 , n205290 , n205291 , n38015 , n205293 , n205294 , n38018 , n205296 , n205297 , n38021 , 
 n205299 , n205300 , n38024 , n205302 , n205303 , n38027 , n205305 , n205306 , n38030 , n205308 , 
 n205309 , n38033 , n38034 , n38035 , n38036 , n205314 , n205315 , n38039 , n205317 , n205318 , 
 n205319 , n38043 , n205321 , n38045 , n38046 , n205324 , n205325 , n38049 , n205327 , n205328 , 
 n38052 , n205330 , n38054 , n205332 , n205333 , n38057 , n205335 , n205336 , n38060 , n205338 , 
 n38062 , n205340 , n38064 , n38065 , n205343 , n205344 , n38068 , n205346 , n205347 , n38071 , 
 n205349 , n205350 , n38074 , n205352 , n205353 , n38077 , n38078 , n38079 , n38080 , n205358 , 
 n205359 , n38083 , n205361 , n38085 , n205363 , n38087 , n38088 , n205366 , n205367 , n205368 , 
 n38092 , n205370 , n205371 , n38095 , n205373 , n205374 , n38098 , n205376 , n205377 , n38101 , 
 n205379 , n205380 , n205381 , n38105 , n205383 , n38107 , n38108 , n205386 , n205387 , n205388 , 
 n38112 , n205390 , n205391 , n38115 , n205393 , n205394 , n38118 , n205396 , n205397 , n38121 , 
 n38122 , n38123 , n38124 , n38125 , n205403 , n205404 , n38128 , n205406 , n205407 , n38131 , 
 n205409 , n205410 , n38134 , n38135 , n38136 , n38137 , n38138 , n205416 , n205417 , n38141 , 
 n205419 , n205420 , n38144 , n38145 , n38146 , n38147 , n205425 , n205426 , n38150 , n205428 , 
 n205429 , n38153 , n205431 , n205432 , n38156 , n205434 , n205435 , n38159 , n205437 , n38161 , 
 n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n205447 , n205448 , 
 n38172 , n205450 , n38174 , n205452 , n38176 , n205454 , n38178 , n205456 , n205457 , n38181 , 
 n205459 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n205467 , n38191 , 
 n38192 , n205470 , n38194 , n205472 , n205473 , n205474 , n205475 , n38199 , n205477 , n205478 , 
 n38202 , n205480 , n205481 , n38205 , n205483 , n205484 , n38208 , n205486 , n205487 , n38211 , 
 n205489 , n205490 , n38214 , n38215 , n205493 , n38217 , n205495 , n38219 , n205497 , n38221 , 
 n205499 , n38223 , n205501 , n205502 , n38226 , n205504 , n205505 , n38229 , n38230 , n38231 , 
 n205509 , n38233 , n205511 , n205512 , n38236 , n38237 , n205515 , n205516 , n38240 , n205518 , 
 n205519 , n205520 , n38244 , n205522 , n205523 , n38247 , n205525 , n205526 , n38250 , n205528 , 
 n205529 , n38253 , n205531 , n205532 , n38256 , n205534 , n205535 , n38259 , n205537 , n205538 , 
 n38262 , n205540 , n205541 , n38265 , n38266 , n205544 , n205545 , n38269 , n205547 , n205548 , 
 n38272 , n205550 , n205551 , n38275 , n205553 , n38277 , n38278 , n38279 , n38280 , n205558 , 
 n205559 , n38283 , n38284 , n38285 , n38286 , n205564 , n205565 , n38289 , n38290 , n38291 , 
 n38292 , n205570 , n205571 , n38295 , n38296 , n38297 , n38298 , n205576 , n205577 , n38301 , 
 n38302 , n38303 , n38304 , n38305 , n205583 , n205584 , n38308 , n205586 , n205587 , n205588 , 
 n38312 , n205590 , n205591 , n38315 , n38316 , n205594 , n38318 , n205596 , n205597 , n38321 , 
 n38322 , n205600 , n205601 , n38325 , n205603 , n38327 , n38328 , n205606 , n205607 , n38331 , 
 n205609 , n205610 , n38334 , n205612 , n205613 , n38337 , n205615 , n205616 , n38340 , n205618 , 
 n38342 , n205620 , n38344 , n38345 , n205623 , n205624 , n38348 , n205626 , n205627 , n38351 , 
 n205629 , n38353 , n205631 , n205632 , n38356 , n205634 , n205635 , n205636 , n205637 , n38361 , 
 n205639 , n38363 , n205641 , n205642 , n38366 , n205644 , n38368 , n205646 , n205647 , n205648 , 
 n38372 , n205650 , n38374 , n205652 , n205653 , n205654 , n205655 , n38379 , n205657 , n205658 , 
 n38382 , n205660 , n205661 , n38385 , n38386 , n205664 , n205665 , n38389 , n205667 , n205668 , 
 n38392 , n205670 , n205671 , n38395 , n205673 , n205674 , n38398 , n205676 , n205677 , n38401 , 
 n205679 , n205680 , n38404 , n205682 , n205683 , n205684 , n205685 , n38409 , n205687 , n205688 , 
 n38412 , n205690 , n38414 , n38415 , n38416 , n205694 , n205695 , n38419 , n205697 , n205698 , 
 n205699 , n205700 , n38424 , n205702 , n205703 , n38427 , n205705 , n205706 , n38430 , n205708 , 
 n38432 , n205710 , n205711 , n38435 , n205713 , n38437 , n205715 , n205716 , n38440 , n205718 , 
 n205719 , n38443 , n205721 , n205722 , n38446 , n205724 , n205725 , n38449 , n205727 , n38451 , 
 n38452 , n38453 , n205731 , n38455 , n205733 , n38457 , n38458 , n205736 , n205737 , n38461 , 
 n205739 , n205740 , n205741 , n205742 , n38466 , n205744 , n205745 , n38469 , n205747 , n205748 , 
 n38472 , n205750 , n205751 , n38475 , n205753 , n38477 , n38478 , n38479 , n205757 , n205758 , 
 n38482 , n205760 , n38484 , n38485 , n205763 , n205764 , n205765 , n38489 , n205767 , n205768 , 
 n205769 , n38493 , n205771 , n205772 , n38496 , n205774 , n38498 , n38499 , n38500 , n38501 , 
 n205779 , n205780 , n205781 , n205782 , n38506 , n205784 , n205785 , n38509 , n205787 , n205788 , 
 n38512 , n205790 , n205791 , n205792 , n205793 , n38517 , n205795 , n205796 , n38520 , n205798 , 
 n38522 , n38523 , n205801 , n38525 , n205803 , n38527 , n38528 , n38529 , n38530 , n38531 , 
 n38532 , n38533 , n205811 , n38535 , n205813 , n205814 , n205815 , n205816 , n38540 , n205818 , 
 n205819 , n38543 , n205821 , n38545 , n205823 , n205824 , n205825 , n38549 , n205827 , n205828 , 
 n38552 , n38553 , n205831 , n205832 , n205833 , n205834 , n38558 , n205836 , n205837 , n205838 , 
 n205839 , n38563 , n205841 , n205842 , n205843 , n38567 , n205845 , n205846 , n38570 , n38571 , 
 n205849 , n205850 , n38574 , n205852 , n205853 , n205854 , n38578 , n205856 , n205857 , n38581 , 
 n38582 , n205860 , n205861 , n38585 , n38586 , n205864 , n205865 , n38589 , n205867 , n205868 , 
 n38592 , n205870 , n38594 , n205872 , n205873 , n38597 , n205875 , n205876 , n38600 , n205878 , 
 n205879 , n38603 , n205881 , n205882 , n205883 , n205884 , n205885 , n38609 , n205887 , n205888 , 
 n38612 , n38613 , n205891 , n205892 , n38616 , n205894 , n205895 , n38619 , n38620 , n205898 , 
 n205899 , n38623 , n205901 , n38625 , n205903 , n205904 , n38628 , n38629 , n38630 , n205908 , 
 n205909 , n38633 , n205911 , n205912 , n38636 , n205914 , n205915 , n205916 , n38640 , n205918 , 
 n205919 , n38643 , n205921 , n38645 , n205923 , n205924 , n38648 , n38649 , n205927 , n38651 , 
 n205929 , n205930 , n38654 , n205932 , n205933 , n205934 , n38658 , n205936 , n205937 , n38661 , 
 n205939 , n205940 , n38664 , n38665 , n205943 , n205944 , n38668 , n38669 , n38670 , n205948 , 
 n205949 , n38673 , n38674 , n205952 , n205953 , n38677 , n205955 , n205956 , n38680 , n205958 , 
 n205959 , n38683 , n205961 , n205962 , n38686 , n38687 , n205965 , n205966 , n205967 , n205968 , 
 n205969 , n38693 , n205971 , n205972 , n38696 , n205974 , n205975 , n38699 , n38700 , n205978 , 
 n205979 , n38703 , n205981 , n205982 , n38706 , n205984 , n205985 , n205986 , n38710 , n205988 , 
 n38712 , n38713 , n205991 , n38715 , n205993 , n38717 , n205995 , n205996 , n38720 , n205998 , 
 n205999 , n38723 , n206001 , n38725 , n206003 , n38727 , n38728 , n206006 , n38730 , n206008 , 
 n38732 , n206010 , n206011 , n38735 , n206013 , n206014 , n38738 , n38739 , n38740 , n206018 , 
 n206019 , n38743 , n38744 , n38745 , n206023 , n206024 , n38748 , n38749 , n38750 , n206028 , 
 n206029 , n38753 , n206031 , n206032 , n206033 , n206034 , n38758 , n206036 , n206037 , n206038 , 
 n206039 , n38763 , n206041 , n206042 , n38766 , n38767 , n206045 , n206046 , n38770 , n38771 , 
 n38772 , n38773 , n38774 , n206052 , n206053 , n38777 , n206055 , n206056 , n38780 , n38781 , 
 n38782 , n38783 , n206061 , n206062 , n38786 , n206064 , n206065 , n38789 , n206067 , n206068 , 
 n38792 , n206070 , n206071 , n38795 , n206073 , n206074 , n38798 , n206076 , n38800 , n206078 , 
 n38802 , n206080 , n206081 , n206082 , n206083 , n38807 , n206085 , n206086 , n38810 , n38811 , 
 n206089 , n206090 , n38814 , n38815 , n206093 , n206094 , n38818 , n206096 , n38820 , n206098 , 
 n206099 , n38823 , n38824 , n206102 , n206103 , n38827 , n38828 , n38829 , n38830 , n38831 , 
 n206109 , n206110 , n38834 , n38835 , n38836 , n206114 , n206115 , n38839 , n206117 , n206118 , 
 n38842 , n38843 , n38844 , n38845 , n206123 , n206124 , n38848 , n38849 , n206127 , n206128 , 
 n38852 , n38853 , n38854 , n38855 , n38856 , n206134 , n206135 , n38859 , n38860 , n38861 , 
 n206139 , n206140 , n38864 , n206142 , n206143 , n38867 , n38868 , n206146 , n206147 , n38871 , 
 n38872 , n38873 , n38874 , n206152 , n206153 , n38877 , n206155 , n206156 , n38880 , n206158 , 
 n206159 , n38883 , n206161 , n206162 , n38886 , n206164 , n206165 , n38889 , n206167 , n206168 , 
 n38892 , n206170 , n206171 , n38895 , n38896 , n38897 , n206175 , n206176 , n38900 , n38901 , 
 n38902 , n38903 , n206181 , n206182 , n38906 , n206184 , n206185 , n38909 , n206187 , n206188 , 
 n38912 , n206190 , n206191 , n38915 , n206193 , n206194 , n38918 , n206196 , n206197 , n38921 , 
 n206199 , n206200 , n38924 , n206202 , n206203 , n206204 , n38928 , n206206 , n38930 , n206208 , 
 n38932 , n206210 , n206211 , n38935 , n206213 , n206214 , n38938 , n206216 , n206217 , n38941 , 
 n206219 , n38943 , n38944 , n206222 , n38946 , n206224 , n38948 , n38949 , n38950 , n206228 , 
 n38952 , n206230 , n38954 , n206232 , n206233 , n38957 , n38958 , n206236 , n38960 , n206238 , 
 n38962 , n38963 , n206241 , n206242 , n38966 , n206244 , n206245 , n206246 , n38970 , n206248 , 
 n206249 , n38973 , n206251 , n206252 , n38976 , n206254 , n206255 , n38979 , n206257 , n206258 , 
 n38982 , n206260 , n38984 , n38985 , n206263 , n206264 , n38988 , n206266 , n206267 , n206268 , 
 n38992 , n206270 , n206271 , n38995 , n206273 , n206274 , n38998 , n206276 , n39000 , n206278 , 
 n39002 , n206280 , n206281 , n39005 , n206283 , n39007 , n39008 , n39009 , n39010 , n39011 , 
 n39012 , n39013 , n39014 , n206292 , n39016 , n206294 , n39018 , n206296 , n206297 , n39021 , 
 n206299 , n39023 , n206301 , n206302 , n39026 , n206304 , n39028 , n206306 , n206307 , n39031 , 
 n206309 , n206310 , n39034 , n206312 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , 
 n206319 , n39043 , n206321 , n206322 , n206323 , n39047 , n206325 , n206326 , n39050 , n206328 , 
 n39052 , n206330 , n206331 , n39055 , n206333 , n39057 , n206335 , n206336 , n206337 , n39061 , 
 n206339 , n206340 , n39064 , n206342 , n39066 , n39067 , n206345 , n39069 , n206347 , n39071 , 
 n39072 , n206350 , n39074 , n206352 , n206353 , n39077 , n206355 , n206356 , n39080 , n206358 , 
 n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n206367 , n206368 , 
 n206369 , n206370 , n39094 , n206372 , n206373 , n39097 , n206375 , n206376 , n39100 , n206378 , 
 n39102 , n206380 , n39104 , n206382 , n39106 , n206384 , n206385 , n206386 , n39110 , n206388 , 
 n39112 , n206390 , n206391 , n39115 , n206393 , n39117 , n39118 , n206396 , n39120 , n206398 , 
 n206399 , n39123 , n206401 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , 
 n39132 , n39133 , n39134 , n39135 , n39136 , n206414 , n206415 , n39139 , n206417 , n206418 , 
 n206419 , n39143 , n206421 , n206422 , n39146 , n206424 , n39148 , n206426 , n206427 , n206428 , 
 n39152 , n206430 , n206431 , n206432 , n39156 , n206434 , n39158 , n39159 , n206437 , n206438 , 
 n39162 , n206440 , n206441 , n39165 , n206443 , n39167 , n206445 , n206446 , n39170 , n206448 , 
 n206449 , n39173 , n206451 , n206452 , n39176 , n206454 , n206455 , n206456 , n39180 , n206458 , 
 n206459 , n39183 , n206461 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n206468 , 
 n206469 , n39193 , n206471 , n206472 , n206473 , n206474 , n39198 , n206476 , n206477 , n39201 , 
 n206479 , n206480 , n39204 , n206482 , n206483 , n206484 , n206485 , n39209 , n206487 , n206488 , 
 n39212 , n206490 , n39214 , n206492 , n206493 , n39217 , n206495 , n206496 , n39220 , n206498 , 
 n206499 , n39223 , n206501 , n206502 , n39226 , n206504 , n206505 , n39229 , n206507 , n206508 , 
 n39232 , n206510 , n206511 , n39235 , n206513 , n39237 , n39238 , n206516 , n39240 , n206518 , 
 n39242 , n39243 , n206521 , n39245 , n206523 , n206524 , n206525 , n39249 , n206527 , n206528 , 
 n39252 , n206530 , n206531 , n39255 , n206533 , n206534 , n39258 , n206536 , n206537 , n39261 , 
 n206539 , n39263 , n206541 , n39265 , n206543 , n206544 , n206545 , n206546 , n39270 , n206548 , 
 n206549 , n39273 , n206551 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , 
 n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n206566 , n206567 , n39291 , 
 n206569 , n39293 , n206571 , n206572 , n39296 , n206574 , n206575 , n39299 , n206577 , n206578 , 
 n206579 , n206580 , n39304 , n206582 , n206583 , n39307 , n206585 , n39309 , n39310 , n39311 , 
 n206589 , n206590 , n39314 , n206592 , n39316 , n39317 , n39318 , n206596 , n39320 , n206598 , 
 n39322 , n39323 , n206601 , n39325 , n206603 , n206604 , n39328 , n206606 , n206607 , n39331 , 
 n206609 , n39333 , n39334 , n39335 , n39336 , n206614 , n39338 , n206616 , n39340 , n206618 , 
 n39342 , n39343 , n206621 , n206622 , n39346 , n206624 , n39348 , n206626 , n206627 , n39351 , 
 n206629 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , 
 n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n206647 , n206648 , 
 n39372 , n39373 , n39374 , n39375 , n39376 , n206654 , n206655 , n206656 , n39380 , n206658 , 
 n206659 , n39383 , n206661 , n206662 , n39386 , n206664 , n206665 , n39389 , n206667 , n39391 , 
 n206669 , n206670 , n39394 , n39395 , n206673 , n206674 , n39398 , n39399 , n206677 , n206678 , 
 n39402 , n39403 , n206681 , n206682 , n39406 , n39407 , n206685 , n206686 , n39410 , n206688 , 
 n206689 , n39413 , n39414 , n206692 , n206693 , n39417 , n39418 , n206696 , n39420 , n39421 , 
 n206699 , n206700 , n206701 , n206702 , n206703 , n206704 , n39428 , n206706 , n206707 , n39431 , 
 n206709 , n206710 , n39434 , n206712 , n206713 , n39437 , n206715 , n206716 , n39440 , n206718 , 
 n206719 , n39443 , n206721 , n39445 , n39446 , n206724 , n39448 , n206726 , n39450 , n39451 , 
 n39452 , n206730 , n39454 , n206732 , n206733 , n39457 , n206735 , n39459 , n39460 , n39461 , 
 n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n206748 , 
 n39472 , n206750 , n206751 , n206752 , n39476 , n206754 , n206755 , n39479 , n206757 , n206758 , 
 n206759 , n39483 , n206761 , n39485 , n206763 , n206764 , n39488 , n206766 , n206767 , n39491 , 
 n206769 , n206770 , n39494 , n206772 , n39496 , n39497 , n206775 , n39499 , n206777 , n39501 , 
 n206779 , n206780 , n39504 , n39505 , n206783 , n206784 , n39508 , n206786 , n206787 , n39511 , 
 n206789 , n39513 , n206791 , n206792 , n39516 , n206794 , n206795 , n39519 , n206797 , n206798 , 
 n39522 , n206800 , n39524 , n206802 , n39526 , n206804 , n39528 , n206806 , n39530 , n39531 , 
 n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , 
 n206819 , n206820 , n206821 , n39545 , n206823 , n206824 , n39548 , n206826 , n206827 , n39551 , 
 n206829 , n39553 , n39554 , n206832 , n206833 , n206834 , n39558 , n206836 , n206837 , n39561 , 
 n206839 , n39563 , n206841 , n206842 , n39566 , n206844 , n39568 , n39569 , n206847 , n39571 , 
 n206849 , n39573 , n39574 , n206852 , n39576 , n206854 , n206855 , n39579 , n206857 , n206858 , 
 n39582 , n206860 , n206861 , n39585 , n206863 , n206864 , n39588 , n206866 , n206867 , n206868 , 
 n39592 , n206870 , n39594 , n39595 , n39596 , n39597 , n206875 , n39599 , n206877 , n39601 , 
 n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n206886 , n206887 , n206888 , 
 n39612 , n206890 , n39614 , n206892 , n206893 , n39617 , n206895 , n206896 , n39620 , n206898 , 
 n39622 , n39623 , n206901 , n206902 , n39626 , n206904 , n39628 , n206906 , n206907 , n39631 , 
 n206909 , n39633 , n39634 , n39635 , n39636 , n39637 , n206915 , n39639 , n206917 , n39641 , 
 n39642 , n206920 , n39644 , n206922 , n39646 , n206924 , n39648 , n39649 , n206927 , n39651 , 
 n206929 , n39653 , n39654 , n206932 , n206933 , n206934 , n39658 , n206936 , n206937 , n39661 , 
 n206939 , n206940 , n39664 , n39665 , n206943 , n39667 , n39668 , n206946 , n39670 , n39671 , 
 n206949 , n39673 , n206951 , n39675 , n39676 , n206954 , n39678 , n206956 , n39680 , n206958 , 
 n206959 , n39683 , n206961 , n39685 , n206963 , n206964 , n39688 , n206966 , n206967 , n206968 , 
 n39692 , n206970 , n206971 , n206972 , n39696 , n206974 , n39698 , n206976 , n206977 , n39701 , 
 n206979 , n206980 , n39704 , n206982 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , 
 n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n206995 , n206996 , n39720 , n39721 , 
 n206999 , n39723 , n39724 , n207002 , n207003 , n207004 , n39728 , n207006 , n207007 , n39731 , 
 n207009 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , 
 n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , 
 n39752 , n207030 , n39754 , n207032 , n207033 , n207034 , n39758 , n207036 , n207037 , n39761 , 
 n207039 , n207040 , n207041 , n207042 , n39766 , n207044 , n207045 , n39769 , n207047 , n207048 , 
 n207049 , n207050 , n39774 , n207052 , n207053 , n39777 , n207055 , n207056 , n39780 , n39781 , 
 n207059 , n39783 , n39784 , n207062 , n39786 , n39787 , n39788 , n207066 , n207067 , n39791 , 
 n207069 , n39793 , n39794 , n207072 , n207073 , n207074 , n39798 , n207076 , n207077 , n39801 , 
 n207079 , n207080 , n39804 , n39805 , n207083 , n39807 , n39808 , n207086 , n39810 , n39811 , 
 n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n207098 , 
 n207099 , n39823 , n207101 , n207102 , n39826 , n207104 , n207105 , n39829 , n207107 , n207108 , 
 n39832 , n207110 , n207111 , n39835 , n207113 , n39837 , n207115 , n207116 , n39840 , n207118 , 
 n207119 , n39843 , n207121 , n39845 , n39846 , n39847 , n207125 , n207126 , n207127 , n39851 , 
 n207129 , n207130 , n39854 , n207132 , n207133 , n207134 , n39858 , n207136 , n39860 , n39861 , 
 n207139 , n207140 , n39864 , n207142 , n39866 , n39867 , n39868 , n39869 , n39870 , n207148 , 
 n39872 , n207150 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , 
 n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n207165 , n39889 , n39890 , n207168 , 
 n39892 , n207170 , n207171 , n207172 , n207173 , n39897 , n207175 , n207176 , n207177 , n39901 , 
 n207179 , n207180 , n207181 , n207182 , n39906 , n207184 , n207185 , n39909 , n207187 , n39911 , 
 n207189 , n207190 , n39914 , n207192 , n207193 , n39917 , n207195 , n39919 , n207197 , n39921 , 
 n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , 
 n39932 , n39933 , n39934 , n39935 , n207213 , n207214 , n39938 , n207216 , n207217 , n39941 , 
 n207219 , n39943 , n39944 , n207222 , n39946 , n207224 , n207225 , n39949 , n207227 , n39951 , 
 n207229 , n39953 , n39954 , n207232 , n39956 , n207234 , n207235 , n39959 , n39960 , n207238 , 
 n207239 , n39963 , n207241 , n207242 , n39966 , n207244 , n207245 , n39969 , n207247 , n207248 , 
 n39972 , n207250 , n207251 , n39975 , n207253 , n39977 , n207255 , n39979 , n207257 , n207258 , 
 n39982 , n207260 , n207261 , n39985 , n207263 , n39987 , n39988 , n39989 , n39990 , n39991 , 
 n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n207277 , n40001 , 
 n207279 , n40003 , n40004 , n207282 , n40006 , n207284 , n40008 , n207286 , n207287 , n40011 , 
 n207289 , n40013 , n40014 , n40015 , n207293 , n40017 , n207295 , n40019 , n40020 , n207298 , 
 n40022 , n207300 , n40024 , n40025 , n207303 , n40027 , n207305 , n207306 , n40030 , n207308 , 
 n40032 , n207310 , n207311 , n40035 , n207313 , n40037 , n40038 , n40039 , n40040 , n40041 , 
 n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , 
 n40052 , n40053 , n40054 , n207332 , n207333 , n40057 , n207335 , n207336 , n207337 , n40061 , 
 n207339 , n207340 , n40064 , n207342 , n207343 , n40067 , n207345 , n207346 , n40070 , n207348 , 
 n40072 , n40073 , n207351 , n40075 , n207353 , n207354 , n40078 , n207356 , n40080 , n40081 , 
 n207359 , n40083 , n40084 , n207362 , n40086 , n40087 , n207365 , n40089 , n207367 , n207368 , 
 n40092 , n207370 , n207371 , n40095 , n207373 , n207374 , n40098 , n207376 , n207377 , n40101 , 
 n207379 , n207380 , n40104 , n207382 , n207383 , n207384 , n40108 , n207386 , n40110 , n40111 , 
 n207389 , n40113 , n207391 , n40115 , n40116 , n40117 , n40118 , n207396 , n40120 , n207398 , 
 n207399 , n207400 , n40124 , n207402 , n207403 , n207404 , n40128 , n207406 , n207407 , n40131 , 
 n207409 , n207410 , n40134 , n207412 , n40136 , n40137 , n40138 , n207416 , n40140 , n207418 , 
 n207419 , n40143 , n207421 , n40145 , n40146 , n207424 , n40148 , n207426 , n40150 , n207428 , 
 n207429 , n40153 , n40154 , n207432 , n40156 , n207434 , n207435 , n40159 , n207437 , n207438 , 
 n40162 , n207440 , n207441 , n40165 , n207443 , n207444 , n40168 , n207446 , n40170 , n40171 , 
 n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , 
 n40182 , n40183 , n40184 , n207462 , n207463 , n40187 , n207465 , n207466 , n40190 , n207468 , 
 n40192 , n40193 , n207471 , n40195 , n207473 , n40197 , n40198 , n207476 , n40200 , n207478 , 
 n207479 , n40203 , n207481 , n207482 , n40206 , n207484 , n40208 , n207486 , n207487 , n40211 , 
 n207489 , n40213 , n40214 , n207492 , n40216 , n207494 , n40218 , n207496 , n207497 , n40221 , 
 n207499 , n40223 , n40224 , n207502 , n40226 , n207504 , n207505 , n40229 , n207507 , n40231 , 
 n40232 , n40233 , n207511 , n40235 , n207513 , n207514 , n40238 , n207516 , n207517 , n40241 , 
 n207519 , n40243 , n207521 , n207522 , n40246 , n207524 , n207525 , n40249 , n207527 , n40251 , 
 n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n207537 , n40261 , 
 n207539 , n207540 , n40264 , n207542 , n40266 , n207544 , n207545 , n40269 , n207547 , n207548 , 
 n40272 , n40273 , n207551 , n40275 , n207553 , n207554 , n40278 , n207556 , n40280 , n40281 , 
 n207559 , n40283 , n207561 , n40285 , n40286 , n207564 , n40288 , n207566 , n207567 , n40291 , 
 n207569 , n207570 , n40294 , n207572 , n207573 , n40297 , n207575 , n207576 , n40300 , n207578 , 
 n207579 , n40303 , n207581 , n207582 , n207583 , n40307 , n207585 , n207586 , n40310 , n207588 , 
 n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n207595 , n207596 , n40320 , n207598 , 
 n207599 , n40323 , n207601 , n207602 , n40326 , n207604 , n40328 , n40329 , n207607 , n207608 , 
 n40332 , n207610 , n40334 , n207612 , n207613 , n40337 , n207615 , n207616 , n207617 , n40341 , 
 n207619 , n207620 , n40344 , n207622 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , 
 n207629 , n40353 , n207631 , n40355 , n207633 , n207634 , n40358 , n207636 , n40360 , n40361 , 
 n207639 , n40363 , n207641 , n40365 , n40366 , n207644 , n40368 , n207646 , n207647 , n40371 , 
 n207649 , n207650 , n40374 , n207652 , n207653 , n40377 , n207655 , n207656 , n207657 , n207658 , 
 n40382 , n207660 , n207661 , n40385 , n207663 , n207664 , n40388 , n40389 , n207667 , n40391 , 
 n40392 , n207670 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , 
 n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , 
 n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , 
 n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , 
 n207709 , n207710 , n40434 , n207712 , n207713 , n40437 , n207715 , n207716 , n207717 , n40441 , 
 n207719 , n207720 , n40444 , n207722 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , 
 n207729 , n40453 , n207731 , n40455 , n40456 , n207734 , n40458 , n207736 , n40460 , n207738 , 
 n40462 , n207740 , n207741 , n207742 , n40466 , n207744 , n207745 , n207746 , n40470 , n207748 , 
 n207749 , n40473 , n40474 , n207752 , n40476 , n207754 , n207755 , n40479 , n40480 , n207758 , 
 n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n207765 , n207766 , n207767 , n40491 , 
 n207769 , n207770 , n40494 , n207772 , n207773 , n207774 , n40498 , n207776 , n40500 , n40501 , 
 n40502 , n207780 , n40504 , n40505 , n207783 , n40507 , n207785 , n40509 , n207787 , n40511 , 
 n207789 , n40513 , n40514 , n207792 , n40516 , n207794 , n40518 , n40519 , n207797 , n40521 , 
 n207799 , n40523 , n40524 , n207802 , n40526 , n207804 , n207805 , n40529 , n207807 , n207808 , 
 n40532 , n207810 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , 
 n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , 
 n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , 
 n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n207847 , n40571 , 
 n207849 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n207857 , n40581 , 
 n207859 , n207860 , n40584 , n207862 , n207863 , n40587 , n207865 , n40589 , n207867 , n207868 , 
 n40592 , n40593 , n207871 , n40595 , n40596 , n207874 , n40598 , n40599 , n207877 , n207878 , 
 n40602 , n207880 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n207888 , 
 n40612 , n207890 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , 
 n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n207907 , n40631 , 
 n207909 , n40633 , n207911 , n207912 , n40636 , n207914 , n40638 , n207916 , n40640 , n207918 , 
 n207919 , n207920 , n207921 , n207922 , n207923 , n207924 , n207925 , n207926 , n40650 , n207928 , 
 n40652 , n207930 , n40654 , n207932 , n40656 , n207934 , n40658 , n207936 , n40660 , n207938 , 
 n40662 , n207940 , n40664 , n207942 , n40666 , n207944 , n40668 , n207946 , n40670 , n207948 , 
 n40672 , n207950 , n40674 , n207952 , n40676 , n207954 , n207955 , n207956 , n207957 , n207958 , 
 n40682 , n207960 , n207961 , n207962 , n207963 , n207964 , n40688 , n207966 , n207967 , n207968 , 
 n40692 , n207970 , n40694 , n207972 , n207973 , n207974 , n207975 , n207976 , n40700 , n207978 , 
 n207979 , n207980 , n40704 , n207982 , n40706 , n207984 , n40708 , n207986 , n40710 , n207988 , 
 n40712 , n207990 , n40714 , n207992 , n207993 , n207994 , n40718 , n207996 , n40720 , n207998 , 
 n40722 , n208000 , n40724 , n208002 , n40726 , n208004 , n40728 , n208006 , n40730 , n208008 , 
 n40732 , n208010 , n40734 , n208012 , n40736 , n208014 , n40738 , n208016 , n208017 , n208018 , 
 n208019 , n208020 , n40744 , n208022 , n40746 , n208024 , n40748 , n208026 , n40750 , n208028 , 
 n40752 , n208030 , n40754 , n208032 , n208033 , n208034 , n208035 , n208036 , n40760 , n208038 , 
 n40762 , n208040 , n40764 , n208042 , n40766 , n208044 , n40768 , n208046 , n40770 , n208048 , 
 n40772 , n208050 , n40774 , n208052 , n40776 , n208054 , n208055 , n208056 , n208057 , n208058 , 
 n40782 , n208060 , n208061 , n208062 , n208063 , n208064 , n40788 , n208066 , n40790 , n208068 , 
 n208069 , n208070 , n40794 , n208072 , n40796 , n208074 , n208075 , n208076 , n40800 , n208078 , 
 n40802 , n208080 , n40804 , n208082 , n40806 , n208084 , n40808 , n208086 , n40810 , n208088 , 
 n40812 , n208090 , n40814 , n208092 , n208093 , n208094 , n208095 , n208096 , n40820 , n208098 , 
 n40822 , n208100 , n208101 , n208102 , n40826 , n208104 , n208105 , n208106 , n40830 , n208108 , 
 n208109 , n208110 , n40834 , n208112 , n208113 , n208114 , n40838 , n208116 , n40840 , n208118 , 
 n40842 , n208120 , n208121 , n208122 , n208123 , n208124 , n40848 , n208126 , n40850 , n208128 , 
 n40852 , n208130 , n40854 , n208132 , n40856 , n208134 , n208135 , n208136 , n208137 , n208138 , 
 n208139 , n208140 , n40864 , n208142 , n208143 , n208144 , n40868 , n208146 , n208147 , n208148 , 
 n208149 , n208150 , n208151 , n208152 , n40876 , n208154 , n208155 , n208156 , n208157 , n208158 , 
 n40882 , n208160 , n40884 , n208162 , n40886 , n208164 , n40888 , n208166 , n40890 , n208168 , 
 n208169 , n208170 , n208171 , n208172 , n208173 , n208174 , n208175 , n208176 , n208177 , n208178 , 
 n208179 , n208180 , n208181 , n208182 , n208183 , n208184 , n208185 , n208186 , n208187 , n208188 , 
 n208189 , n208190 , n208191 , n208192 , n208193 , n208194 , n208195 , n208196 , n208197 , n208198 , 
 n208199 , n208200 , n208201 , n208202 , n208203 , n208204 , n208205 , n208206 , n208207 , n208208 , 
 n208209 , n208210 , n208211 , n208212 , n208213 , n208214 , n208215 , n208216 , n208217 , n208218 , 
 n208219 , n208220 , n208221 , n208222 , n208223 , n208224 , n208225 , n208226 , n208227 , n208228 , 
 n208229 , n208230 , n208231 , n208232 , n208233 , n208234 , n208235 , n208236 , n208237 , n208238 , 
 n208239 , n208240 , n208241 , n208242 , n208243 , n208244 , n208245 , n208246 , n208247 , n208248 , 
 n208249 , n208250 , n208251 , n208252 , n208253 , n208254 , n208255 , n208256 , n208257 , n208258 , 
 n208259 , n208260 , n208261 , n208262 , n208263 , n208264 , n208265 , n208266 , n208267 , n208268 , 
 n208269 , n208270 , n208271 , n208272 , n208273 , n208274 , n208275 , n208276 , n208277 , n208278 , 
 n208279 , n208280 , n208281 , n208282 , n208283 , n208284 , n208285 , n208286 , n208287 , n208288 , 
 n208289 , n208290 , n208291 , n208292 , n208293 , n41017 , n41018 , n208296 , n41020 , n208298 , 
 n41022 , n41023 , n208301 , n41025 , n208303 , n208304 , n41028 , n208306 , n41030 , n208308 , 
 n208309 , n41033 , n208311 , n208312 , n208313 , n41037 , n208315 , n208316 , n208317 , n41041 , 
 n208319 , n41043 , n41044 , n208322 , n208323 , n41047 , n208325 , n208326 , n41050 , n208328 , 
 n208329 , n208330 , n41054 , n208332 , n208333 , n41057 , n208335 , n41059 , n41060 , n208338 , 
 n41062 , n208340 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , 
 n41072 , n41073 , n41074 , n208352 , n208353 , n41077 , n208355 , n208356 , n41080 , n208358 , 
 n41082 , n41083 , n208361 , n41085 , n208363 , n41087 , n41088 , n208366 , n41090 , n208368 , 
 n208369 , n41093 , n208371 , n208372 , n41096 , n208374 , n208375 , n41099 , n208377 , n208378 , 
 n208379 , n41103 , n208381 , n208382 , n41106 , n208384 , n41108 , n208386 , n208387 , n41111 , 
 n41112 , n208390 , n41114 , n208392 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , 
 n41122 , n41123 , n208401 , n208402 , n41126 , n208404 , n41128 , n208406 , n41130 , n208408 , 
 n41132 , n41133 , n208411 , n41135 , n208413 , n41137 , n208415 , n41139 , n41140 , n41141 , 
 n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n208425 , n41149 , n41150 , n41151 , 
 n208429 , n41153 , n41154 , n208432 , n41156 , n208434 , n208435 , n41159 , n41160 , n208438 , 
 n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n208447 , n41171 , 
 n208449 , n208450 , n41174 , n208452 , n41176 , n41177 , n208455 , n41179 , n208457 , n41181 , 
 n208459 , n208460 , n41184 , n208462 , n41186 , n208464 , n208465 , n208466 , n41190 , n208468 , 
 n41192 , n208470 , n208471 , n208472 , n41196 , n208474 , n208475 , n41199 , n208477 , n208478 , 
 n41202 , n41203 , n208481 , n41205 , n41206 , n208484 , n41208 , n41209 , n208487 , n208488 , 
 n41212 , n208490 , n208491 , n41215 , n208493 , n41217 , n41218 , n41219 , n41220 , n41221 , 
 n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n208507 , n41231 , 
 n208509 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , 
 n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , 
 n208529 , n41253 , n208531 , n208532 , n41256 , n208534 , n208535 , n208536 , n208537 , n208538 , 
 n208539 , n208540 , n41264 , n208542 , n208543 , n208544 , n208545 , n208546 , n208547 , n41271 , 
 n208549 , n208550 , n41274 , n208552 , n208553 , n41277 , n208555 , n41279 , n208557 , n208558 , 
 n41282 , n208560 , n208561 , n41285 , n41286 , n208564 , n41288 , n41289 , n208567 , n208568 , 
 n208569 , n208570 , n208571 , n208572 , n208573 , n208574 , n41298 , n208576 , n41300 , n41301 , 
 n208579 , n208580 , n41304 , n208582 , n41306 , n41307 , n208585 , n41309 , n208587 , n208588 , 
 n41312 , n41313 , n208591 , n41315 , n41316 , n208594 , n41318 , n41319 , n208597 , n41321 , 
 n41322 , n208600 , n41324 , n208602 , n208603 , n208604 , n41328 , n208606 , n208607 , n41331 , 
 n208609 , n208610 , n208611 , n208612 , n208613 , n208614 , n208615 , n208616 , n208617 , n208618 , 
 n208619 , n208620 , n208621 , n208622 , n208623 , n208624 , n41348 , n208626 , n208627 , n41351 , 
 n208629 , n208630 , n41354 , n41355 , n208633 , n41357 , n41358 , n208636 , n208637 , n208638 , 
 n208639 , n208640 , n208641 , n208642 , n208643 , n208644 , n208645 , n208646 , n208647 , n208648 , 
 n208649 , n208650 , n208651 , n41375 , n208653 , n208654 , n41378 , n208656 , n208657 , n208658 , 
 n41382 , n208660 , n208661 , n41385 , n208663 , n208664 , n41388 , n208666 , n208667 , n41391 , 
 n208669 , n208670 , n41394 , n208672 , n41396 , n41397 , n208675 , n41399 , n41400 , n208678 , 
 n41402 , n41403 , n208681 , n41405 , n208683 , n208684 , n208685 , n208686 , n208687 , n208688 , 
 n41412 , n208690 , n208691 , n41415 , n208693 , n208694 , n41418 , n208696 , n208697 , n41421 , 
 n208699 , n208700 , n41424 , n208702 , n41426 , n208704 , n208705 , n41429 , n208707 , n208708 , 
 n41432 , n208710 , n208711 , n208712 , n41436 , n208714 , n41438 , n208716 , n208717 , n208718 , 
 n208719 , n208720 , n208721 , n208722 , n208723 , n208724 , n208725 , n208726 , n208727 , n208728 , 
 n208729 , n208730 , n208731 , n208732 , n208733 , n208734 , n208735 , n208736 , n208737 , n208738 , 
 n208739 , n208740 , n208741 , n208742 , n208743 , n208744 , n208745 , n208746 , n208747 , n208748 , 
 n208749 , n208750 , n208751 , n208752 , n208753 , n208754 , n208755 , n208756 , n208757 , n208758 , 
 n208759 , n208760 , n208761 , n208762 , n208763 , n208764 , n208765 , n208766 , n208767 , n208768 , 
 n208769 , n208770 , n208771 , n208772 , n208773 , n208774 , n208775 , n208776 , n208777 , n208778 , 
 n208779 , n208780 , n208781 , n208782 , n208783 , n208784 , n208785 , n208786 , n208787 , n208788 , 
 n208789 , n208790 , n208791 , n208792 , n208793 , n208794 , n208795 , n208796 , n208797 , n208798 , 
 n208799 , n208800 , n208801 , n208802 , n208803 , n208804 , n208805 , n208806 , n208807 , n208808 , 
 n208809 , n208810 , n208811 , n208812 , n208813 , n208814 , n208815 , n208816 , n208817 , n208818 , 
 n208819 , n208820 , n208821 , n208822 , n208823 , n208824 , n208825 , n208826 , n208827 , n208828 , 
 n208829 , n208830 , n208831 , n208832 , n208833 , n208834 , n208835 , n208836 , n208837 , n208838 , 
 n208839 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n208847 , n41571 , 
 n208849 , n41573 , n41574 , n208852 , n41576 , n208854 , n208855 , n208856 , n208857 , n41581 , 
 n208859 , n208860 , n208861 , n41585 , n208863 , n208864 , n41588 , n208866 , n208867 , n208868 , 
 n208869 , n41593 , n208871 , n208872 , n41596 , n208874 , n208875 , n41599 , n41600 , n208878 , 
 n41602 , n41603 , n208881 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , 
 n41612 , n41613 , n41614 , n41615 , n41616 , n208894 , n41618 , n41619 , n41620 , n208898 , 
 n41622 , n41623 , n41624 , n41625 , n41626 , n208904 , n41628 , n208906 , n41630 , n208908 , 
 n41632 , n208910 , n208911 , n41635 , n208913 , n208914 , n208915 , n208916 , n41640 , n208918 , 
 n208919 , n41643 , n208921 , n208922 , n41646 , n41647 , n208925 , n41649 , n41650 , n208928 , 
 n41652 , n41653 , n208931 , n208932 , n41656 , n208934 , n208935 , n41659 , n208937 , n208938 , 
 n41662 , n208940 , n41664 , n41665 , n208943 , n41667 , n208945 , n41669 , n41670 , n208948 , 
 n41672 , n208950 , n208951 , n41675 , n208953 , n208954 , n41678 , n208956 , n208957 , n208958 , 
 n41682 , n208960 , n208961 , n208962 , n41686 , n208964 , n208965 , n41689 , n41690 , n208968 , 
 n41692 , n208970 , n208971 , n41695 , n41696 , n208974 , n41698 , n41699 , n41700 , n41701 , 
 n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , 
 n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , 
 n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , 
 n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , 
 n41742 , n209020 , n209021 , n41745 , n209023 , n209024 , n41748 , n209026 , n209027 , n209028 , 
 n209029 , n41753 , n209031 , n209032 , n209033 , n209034 , n41758 , n209036 , n209037 , n209038 , 
 n41762 , n209040 , n41764 , n41765 , n209043 , n41767 , n209045 , n209046 , n41770 , n209048 , 
 n209049 , n41773 , n209051 , n209052 , n41776 , n209054 , n209055 , n41779 , n209057 , n41781 , 
 n209059 , n209060 , n41784 , n209062 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , 
 n209069 , n41793 , n209071 , n41795 , n41796 , n209074 , n41798 , n209076 , n209077 , n209078 , 
 n209079 , n209080 , n41804 , n209082 , n209083 , n209084 , n209085 , n209086 , n209087 , n209088 , 
 n209089 , n209090 , n209091 , n209092 , n209093 , n41817 , n209095 , n209096 , n41820 , n209098 , 
 n209099 , n41823 , n209101 , n209102 , n41826 , n209104 , n41828 , n209106 , n209107 , n41831 , 
 n41832 , n209110 , n41834 , n41835 , n209113 , n41837 , n41838 , n209116 , n209117 , n41841 , 
 n209119 , n209120 , n41844 , n209122 , n209123 , n209124 , n209125 , n209126 , n41850 , n209128 , 
 n209129 , n41853 , n209131 , n209132 , n209133 , n209134 , n41858 , n209136 , n209137 , n41861 , 
 n209139 , n209140 , n41864 , n41865 , n209143 , n41867 , n41868 , n209146 , n41870 , n41871 , 
 n209149 , n209150 , n41874 , n209152 , n209153 , n41877 , n209155 , n209156 , n209157 , n209158 , 
 n41882 , n209160 , n209161 , n41885 , n41886 , n209164 , n41888 , n41889 , n209167 , n41891 , 
 n41892 , n209170 , n41894 , n41895 , n209173 , n41897 , n41898 , n209176 , n41900 , n209178 , 
 n209179 , n41903 , n209181 , n209182 , n209183 , n209184 , n209185 , n41909 , n209187 , n209188 , 
 n209189 , n41913 , n209191 , n209192 , n209193 , n209194 , n209195 , n41919 , n209197 , n209198 , 
 n41922 , n209200 , n209201 , n41925 , n209203 , n209204 , n41928 , n209206 , n209207 , n41931 , 
 n209209 , n209210 , n41934 , n209212 , n41936 , n209214 , n209215 , n209216 , n209217 , n209218 , 
 n41942 , n209220 , n209221 , n209222 , n41946 , n209224 , n209225 , n209226 , n209227 , n209228 , 
 n41952 , n209230 , n209231 , n41955 , n209233 , n209234 , n41958 , n209236 , n209237 , n41961 , 
 n209239 , n209240 , n41964 , n209242 , n41966 , n41967 , n209245 , n41969 , n41970 , n209248 , 
 n41972 , n41973 , n209251 , n41975 , n41976 , n209254 , n41978 , n41979 , n209257 , n41981 , 
 n41982 , n209260 , n41984 , n209262 , n209263 , n209264 , n209265 , n209266 , n209267 , n209268 , 
 n209269 , n209270 , n209271 , n209272 , n209273 , n209274 , n209275 , n209276 , n209277 , n209278 , 
 n209279 , n209280 , n209281 , n209282 , n209283 , n209284 , n209285 , n209286 , n209287 , n209288 , 
 n209289 , n209290 , n209291 , n209292 , n209293 , n209294 , n209295 , n209296 , n209297 , n209298 , 
 n209299 , n209300 , n209301 , n209302 , n209303 , n209304 , n209305 , n209306 , n209307 , n209308 , 
 n209309 , n209310 , n209311 , n209312 , n209313 , n209314 , n209315 , n209316 , n209317 , n209318 , 
 n209319 , n209320 , n209321 , n209322 , n209323 , n209324 , n209325 , n209326 , n209327 , n209328 , 
 n209329 , n209330 , n209331 , n209332 , n209333 , n209334 , n209335 , n209336 , n209337 , n209338 , 
 n209339 , n209340 , n209341 , n209342 , n209343 , n209344 , n209345 , n209346 , n209347 , n209348 , 
 n209349 , n209350 , n209351 , n209352 , n209353 , n209354 , n209355 , n209356 , n209357 , n209358 , 
 n209359 , n209360 , n209361 , n209362 , n209363 , n209364 , n209365 , n209366 , n209367 , n209368 , 
 n209369 , n209370 , n209371 , n209372 , n209373 , n209374 , n209375 , n209376 , n209377 , n209378 , 
 n209379 , n209380 , n209381 , n209382 , n209383 , n209384 , n209385 , n209386 , n209387 , n209388 , 
 n209389 , n209390 , n209391 , n209392 , n209393 , n209394 , n209395 , n209396 , n209397 , n209398 , 
 n209399 , n209400 , n209401 , n209402 , n209403 , n209404 , n209405 , n209406 , n209407 , n209408 , 
 n209409 , n209410 , n209411 , n209412 , n209413 , n209414 , n209415 , n209416 , n209417 , n209418 , 
 n209419 , n209420 , n209421 , n209422 , n209423 , n209424 , n209425 , n209426 , n209427 , n209428 , 
 n209429 , n209430 , n209431 , n209432 , n209433 , n209434 , n209435 , n209436 , n209437 , n209438 , 
 n209439 , n209440 , n209441 , n209442 , n209443 , n209444 , n209445 , n209446 , n209447 , n209448 , 
 n209449 , n209450 , n209451 , n209452 , n209453 , n209454 , n209455 , n209456 , n209457 , n209458 , 
 n209459 , n209460 , n209461 , n209462 , n209463 , n209464 , n209465 , n209466 , n209467 , n209468 , 
 n209469 , n209470 , n209471 , n209472 , n209473 , n209474 , n209475 , n209476 , n209477 , n209478 , 
 n209479 , n209480 , n209481 , n209482 , n209483 , n209484 , n209485 , n209486 , n209487 , n209488 , 
 n209489 , n209490 , n209491 , n209492 , n209493 , n209494 , n209495 , n209496 , n209497 , n209498 , 
 n209499 , n209500 , n209501 , n209502 , n209503 , n209504 , n209505 , n209506 , n209507 , n209508 , 
 n209509 , n209510 , n209511 , n209512 , n209513 , n209514 , n209515 , n209516 , n209517 , n209518 , 
 n209519 , n209520 , n209521 , n209522 , n209523 , n209524 , n209525 , n209526 , n209527 , n209528 , 
 n209529 , n209530 , n209531 , n209532 , n209533 , n209534 , n209535 , n209536 , n209537 , n209538 , 
 n209539 , n209540 , n209541 , n209542 , n209543 , n209544 , n209545 , n209546 , n209547 , n209548 , 
 n209549 , n209550 , n209551 , n209552 , n209553 , n209554 , n209555 , n209556 , n209557 , n209558 , 
 n209559 , n209560 , n209561 , n209562 , n209563 , n209564 , n209565 , n209566 , n209567 , n209568 , 
 n209569 , n209570 , n209571 , n209572 , n209573 , n209574 , n209575 , n209576 , n209577 , n209578 , 
 n209579 , n209580 , n209581 , n209582 , n209583 , n209584 , n209585 , n209586 , n209587 , n209588 , 
 n209589 , n209590 , n209591 , n209592 , n209593 , n209594 , n209595 , n209596 , n209597 , n209598 , 
 n209599 , n209600 , n209601 , n209602 , n209603 , n209604 , n209605 , n209606 , n209607 , n209608 , 
 n209609 , n209610 , n209611 , n209612 , n209613 , n209614 , n209615 , n209616 , n209617 , n209618 , 
 n209619 , n209620 , n209621 , n209622 , n209623 , n209624 , n209625 , n209626 , n209627 , n209628 , 
 n209629 , n209630 , n209631 , n209632 , n209633 , n209634 , n209635 , n209636 , n209637 , n209638 , 
 n209639 , n209640 , n209641 , n209642 , n209643 , n209644 , n209645 , n209646 , n209647 , n209648 , 
 n209649 , n209650 , n209651 , n209652 , n209653 , n209654 , n209655 , n209656 , n209657 , n209658 , 
 n209659 , n209660 , n209661 , n209662 , n209663 , n209664 , n209665 , n209666 , n209667 , n209668 , 
 n209669 , n209670 , n209671 , n209672 , n209673 , n209674 , n209675 , n209676 , n209677 , n209678 , 
 n209679 , n209680 , n209681 , n209682 , n209683 , n209684 , n209685 , n209686 , n209687 , n209688 , 
 n209689 , n209690 , n209691 , n209692 , n209693 , n209694 , n209695 , n209696 , n209697 , n209698 , 
 n209699 , n209700 , n209701 , n209702 , n209703 , n209704 , n209705 , n209706 , n209707 , n209708 , 
 n209709 , n209710 , n209711 , n209712 , n209713 , n209714 , n209715 , n209716 , n209717 , n209718 , 
 n209719 , n209720 , n209721 , n209722 , n209723 , n209724 , n209725 , n209726 , n209727 , n209728 , 
 n209729 , n209730 , n209731 , n209732 , n209733 , n209734 , n209735 , n209736 , n209737 , n209738 , 
 n209739 , n209740 , n209741 , n209742 , n209743 , n209744 , n209745 , n209746 , n209747 , n209748 , 
 n209749 , n209750 , n209751 , n209752 , n209753 , n209754 , n209755 , n209756 , n209757 , n209758 , 
 n209759 , n209760 , n209761 , n209762 , n209763 , n209764 , n209765 , n209766 , n209767 , n209768 , 
 n209769 , n209770 , n209771 , n209772 , n209773 , n209774 , n209775 , n209776 , n209777 , n209778 , 
 n209779 , n209780 , n209781 , n209782 , n209783 , n209784 , n209785 , n209786 , n209787 , n209788 , 
 n209789 , n209790 , n209791 , n209792 , n209793 , n209794 , n209795 , n209796 , n209797 , n209798 , 
 n209799 , n209800 , n209801 , n209802 , n209803 , n209804 , n209805 , n209806 , n209807 , n209808 , 
 n209809 , n209810 , n209811 , n209812 , n209813 , n209814 , n209815 , n209816 , n209817 , n209818 , 
 n209819 , n209820 , n209821 , n209822 , n209823 , n209824 , n209825 , n209826 , n209827 , n209828 , 
 n209829 , n209830 , n209831 , n209832 , n209833 , n209834 , n209835 , n209836 , n209837 , n209838 , 
 n209839 , n209840 , n209841 , n209842 , n209843 , n209844 , n209845 , n209846 , n209847 , n209848 , 
 n209849 , n209850 , n209851 , n209852 , n209853 , n209854 , n209855 , n209856 , n209857 , n209858 , 
 n209859 , n209860 , n209861 , n209862 , n209863 , n209864 , n209865 , n209866 , n209867 , n209868 , 
 n209869 , n209870 , n209871 , n209872 , n209873 , n209874 , n209875 , n209876 , n209877 , n209878 , 
 n209879 , n209880 , n209881 , n209882 , n209883 , n209884 , n209885 , n209886 , n209887 , n209888 , 
 n209889 , n209890 , n209891 , n209892 , n209893 , n209894 , n209895 , n209896 , n209897 , n209898 , 
 n209899 , n209900 , n209901 , n209902 , n209903 , n209904 , n209905 , n209906 , n209907 , n209908 , 
 n209909 , n209910 , n209911 , n209912 , n209913 , n209914 , n209915 , n209916 , n209917 , n209918 , 
 n209919 , n209920 , n209921 , n209922 , n209923 , n209924 , n209925 , n209926 , n209927 , n209928 , 
 n209929 , n209930 , n209931 , n209932 , n209933 , n209934 , n209935 , n209936 , n209937 , n209938 , 
 n209939 , n209940 , n209941 , n209942 , n209943 , n209944 , n209945 , n209946 , n209947 , n209948 , 
 n209949 , n209950 , n209951 , n209952 , n209953 , n209954 , n209955 , n209956 , n209957 , n209958 , 
 n209959 , n209960 , n209961 , n209962 , n209963 , n209964 , n209965 , n209966 , n209967 , n209968 , 
 n209969 , n209970 , n209971 , n209972 , n209973 , n209974 , n209975 , n209976 , n209977 , n209978 , 
 n209979 , n209980 , n209981 , n209982 , n209983 , n209984 , n209985 , n209986 , n209987 , n209988 , 
 n209989 , n209990 , n209991 , n209992 , n209993 , n209994 , n209995 , n209996 , n209997 , n209998 , 
 n209999 , n210000 , n210001 , n210002 , n210003 , n210004 , n210005 , n210006 , n210007 , n210008 , 
 n210009 , n210010 , n210011 , n210012 , n210013 , n210014 , n210015 , n210016 , n210017 , n210018 , 
 n210019 , n210020 , n210021 , n210022 , n210023 , n210024 , n210025 , n210026 , n210027 , n210028 , 
 n210029 , n210030 , n210031 , n210032 , n210033 , n210034 , n210035 , n210036 , n210037 , n210038 , 
 n210039 , n210040 , n210041 , n210042 , n210043 , n210044 , n210045 , n210046 , n210047 , n210048 , 
 n210049 , n210050 , n210051 , n210052 , n210053 , n210054 , n210055 , n210056 , n210057 , n210058 , 
 n210059 , n210060 , n210061 , n210062 , n210063 , n210064 , n210065 , n210066 , n210067 , n210068 , 
 n210069 , n210070 , n210071 , n210072 , n210073 , n210074 , n210075 , n210076 , n210077 , n210078 , 
 n210079 , n210080 , n210081 , n210082 , n210083 , n210084 , n210085 , n210086 , n210087 , n210088 , 
 n210089 , n210090 , n210091 , n210092 , n210093 , n210094 , n210095 , n210096 , n210097 , n210098 , 
 n210099 , n210100 , n210101 , n210102 , n210103 , n210104 , n210105 , n210106 , n210107 , n210108 , 
 n210109 , n210110 , n210111 , n210112 , n210113 , n210114 , n210115 , n210116 , n210117 , n210118 , 
 n210119 , n210120 , n210121 , n210122 , n210123 , n210124 , n210125 , n210126 , n210127 , n210128 , 
 n210129 , n210130 , n210131 , n210132 , n210133 , n210134 , n210135 , n210136 , n210137 , n210138 , 
 n210139 , n210140 , n210141 , n210142 , n210143 , n210144 , n210145 , n210146 , n210147 , n210148 , 
 n210149 , n210150 , n210151 , n210152 , n210153 , n210154 , n210155 , n210156 , n210157 , n210158 , 
 n210159 , n210160 , n210161 , n210162 , n210163 , n210164 , n210165 , n210166 , n210167 , n210168 , 
 n210169 , n210170 , n210171 , n210172 , n210173 , n210174 , n210175 , n210176 , n210177 , n210178 , 
 n210179 , n210180 , n210181 , n210182 , n210183 , n210184 , n210185 , n210186 , n210187 , n210188 , 
 n210189 , n210190 , n210191 , n210192 , n210193 , n210194 , n210195 , n210196 , n210197 , n210198 , 
 n210199 , n210200 , n210201 , n210202 , n210203 , n210204 , n210205 , n210206 , n210207 , n210208 , 
 n210209 , n210210 , n210211 , n210212 , n210213 , n210214 , n210215 , n210216 , n210217 , n210218 , 
 n210219 , n210220 , n210221 , n210222 , n210223 , n210224 , n210225 , n210226 , n210227 , n210228 , 
 n210229 , n210230 , n210231 , n210232 , n210233 , n210234 , n210235 , n210236 , n210237 , n210238 , 
 n210239 , n210240 , n210241 , n210242 , n210243 , n210244 , n210245 , n210246 , n210247 , n210248 , 
 n210249 , n210250 , n210251 , n210252 , n210253 , n210254 , n210255 , n210256 , n210257 , n210258 , 
 n210259 , n210260 , n210261 , n210262 , n210263 , n210264 , n210265 , n210266 , n210267 , n210268 , 
 n210269 , n210270 , n210271 , n210272 , n210273 , n210274 , n210275 , n210276 , n210277 , n210278 , 
 n210279 , n210280 , n210281 , n210282 , n210283 , n210284 , n210285 , n210286 , n210287 , n210288 , 
 n210289 , n210290 , n210291 , n210292 , n210293 , n210294 , n210295 , n210296 , n210297 , n210298 , 
 n210299 , n210300 , n210301 , n210302 , n210303 , n210304 , n210305 , n210306 , n210307 , n210308 , 
 n210309 , n210310 , n210311 , n210312 , n210313 , n210314 , n210315 , n210316 , n210317 , n210318 , 
 n210319 , n210320 , n210321 , n210322 , n210323 , n210324 , n210325 , n210326 , n210327 , n210328 , 
 n210329 , n210330 , n210331 , n210332 , n210333 , n210334 , n210335 , n210336 , n210337 , n210338 , 
 n210339 , n210340 , n210341 , n210342 , n210343 , n210344 , n210345 , n210346 , n210347 , n210348 , 
 n210349 , n210350 , n210351 , n210352 , n210353 , n210354 , n210355 , n210356 , n210357 , n210358 , 
 n210359 , n210360 , n210361 , n210362 , n210363 , n210364 , n210365 , n210366 , n210367 , n210368 , 
 n210369 , n210370 , n210371 , n210372 , n210373 , n210374 , n210375 , n210376 , n210377 , n210378 , 
 n210379 , n210380 , n210381 , n210382 , n210383 , n210384 , n210385 , n210386 , n210387 , n210388 , 
 n210389 , n210390 , n210391 , n210392 , n210393 , n210394 , n210395 , n210396 , n210397 , n210398 , 
 n210399 , n210400 , n210401 , n210402 , n210403 , n210404 , n210405 , n210406 , n210407 , n210408 , 
 n210409 , n210410 , n210411 , n210412 , n210413 , n210414 , n210415 , n210416 , n210417 , n210418 , 
 n210419 , n210420 , n210421 , n210422 , n210423 , n210424 , n210425 , n210426 , n210427 , n210428 , 
 n210429 , n210430 , n210431 , n210432 , n210433 , n210434 , n210435 , n210436 , n210437 , n210438 , 
 n210439 , n210440 , n210441 , n210442 , n210443 , n210444 , n210445 , n210446 , n210447 , n210448 , 
 n210449 , n210450 , n210451 , n210452 , n210453 , n210454 , n210455 , n210456 , n210457 , n210458 , 
 n210459 , n210460 , n210461 , n210462 , n210463 , n210464 , n210465 , n210466 , n210467 , n210468 , 
 n210469 , n210470 , n210471 , n210472 , n210473 , n210474 , n210475 , n210476 , n210477 , n210478 , 
 n210479 , n210480 , n210481 , n210482 , n210483 , n210484 , n210485 , n210486 , n210487 , n210488 , 
 n210489 , n210490 , n210491 , n210492 , n210493 , n210494 , n210495 , n210496 , n210497 , n210498 , 
 n210499 , n210500 , n210501 , n210502 , n210503 , n210504 , n210505 , n210506 , n210507 , n210508 , 
 n210509 , n210510 , n210511 , n210512 , n210513 , n210514 , n210515 , n210516 , n210517 , n210518 , 
 n210519 , n210520 , n210521 , n210522 , n210523 , n210524 , n210525 , n210526 , n210527 , n210528 , 
 n210529 , n210530 , n210531 , n210532 , n210533 , n210534 , n210535 , n210536 , n210537 , n210538 , 
 n210539 , n210540 , n210541 , n210542 , n210543 , n210544 , n210545 , n210546 , n210547 , n210548 , 
 n210549 , n210550 , n210551 , n210552 , n210553 , n210554 , n210555 , n210556 , n210557 , n210558 , 
 n210559 , n210560 , n210561 , n210562 , n210563 , n210564 , n210565 , n210566 , n210567 , n210568 , 
 n210569 , n210570 , n210571 , n210572 , n210573 , n210574 , n210575 , n210576 , n210577 , n210578 , 
 n210579 , n210580 , n210581 , n210582 , n210583 , n210584 , n210585 , n210586 , n210587 , n210588 , 
 n210589 , n210590 , n210591 , n210592 , n210593 , n210594 , n210595 , n210596 , n210597 , n210598 , 
 n210599 , n210600 , n210601 , n210602 , n210603 , n210604 , n210605 , n210606 , n210607 , n210608 , 
 n210609 , n210610 , n210611 , n210612 , n210613 , n210614 , n210615 , n210616 , n210617 , n210618 , 
 n210619 , n210620 , n210621 , n210622 , n210623 , n210624 , n210625 , n210626 , n210627 , n210628 , 
 n210629 , n210630 , n210631 , n210632 , n210633 , n210634 , n210635 , n210636 , n210637 , n210638 , 
 n210639 , n210640 , n210641 , n210642 , n210643 , n210644 , n210645 , n210646 , n210647 , n210648 , 
 n210649 , n210650 , n210651 , n210652 , n210653 , n210654 , n210655 , n210656 , n210657 , n210658 , 
 n210659 , n210660 , n210661 , n210662 , n210663 , n210664 , n210665 , n210666 , n210667 , n210668 , 
 n210669 , n210670 , n210671 , n210672 , n210673 , n210674 , n210675 , n210676 , n210677 , n210678 , 
 n210679 , n210680 , n210681 , n210682 , n210683 , n210684 , n210685 , n210686 , n210687 , n210688 , 
 n210689 , n210690 , n210691 , n210692 , n210693 , n210694 , n210695 , n210696 , n210697 , n210698 , 
 n210699 , n210700 , n210701 , n210702 , n210703 , n210704 , n210705 , n210706 , n210707 , n210708 , 
 n210709 , n210710 , n210711 , n210712 , n210713 , n210714 , n210715 , n210716 , n210717 , n210718 , 
 n210719 , n210720 , n210721 , n210722 , n210723 , n210724 , n210725 , n210726 , n210727 , n210728 , 
 n210729 , n210730 , n210731 , n210732 , n210733 , n210734 , n210735 , n210736 , n210737 , n210738 , 
 n210739 , n210740 , n210741 , n210742 , n210743 , n210744 , n210745 , n210746 , n210747 , n210748 , 
 n210749 , n210750 , n210751 , n210752 , n210753 , n210754 , n210755 , n210756 , n210757 , n210758 , 
 n210759 , n210760 , n210761 , n210762 , n210763 , n210764 , n210765 , n210766 , n210767 , n210768 , 
 n210769 , n210770 , n210771 , n210772 , n210773 , n210774 , n210775 , n210776 , n210777 , n210778 , 
 n210779 , n210780 , n210781 , n210782 , n210783 , n210784 , n210785 , n210786 , n210787 , n210788 , 
 n210789 , n210790 , n210791 , n210792 , n210793 , n210794 , n210795 , n210796 , n210797 , n210798 , 
 n210799 , n210800 , n210801 , n210802 , n210803 , n210804 , n210805 , n210806 , n210807 , n210808 , 
 n210809 , n210810 , n210811 , n210812 , n210813 , n210814 , n210815 , n210816 , n210817 , n210818 , 
 n210819 , n210820 , n210821 , n210822 , n210823 , n210824 , n210825 , n210826 , n210827 , n210828 , 
 n210829 , n210830 , n210831 , n210832 , n210833 , n210834 , n210835 , n210836 , n210837 , n210838 , 
 n210839 , n210840 , n210841 , n210842 , n210843 , n210844 , n210845 , n210846 , n210847 , n210848 , 
 n210849 , n210850 , n210851 , n210852 , n210853 , n210854 , n210855 , n210856 , n210857 , n210858 , 
 n210859 , n210860 , n210861 , n210862 , n210863 , n210864 , n210865 , n210866 , n210867 , n210868 , 
 n210869 , n210870 , n210871 , n210872 , n210873 , n210874 , n210875 , n210876 , n210877 , n210878 , 
 n210879 , n210880 , n210881 , n210882 , n210883 , n210884 , n210885 , n210886 , n210887 , n210888 , 
 n210889 , n210890 , n210891 , n210892 , n210893 , n210894 , n210895 , n210896 , n210897 , n210898 , 
 n210899 , n210900 , n210901 , n210902 , n210903 , n210904 , n210905 , n210906 , n210907 , n210908 , 
 n210909 , n210910 , n210911 , n210912 , n210913 , n210914 , n210915 , n210916 , n210917 , n210918 , 
 n210919 , n210920 , n210921 , n210922 , n210923 , n210924 , n210925 , n210926 , n210927 , n210928 , 
 n210929 , n210930 , n210931 , n210932 , n210933 , n210934 , n210935 , n210936 , n210937 , n210938 , 
 n210939 , n210940 , n210941 , n210942 , n210943 , n210944 , n210945 , n210946 , n210947 , n210948 , 
 n210949 , n210950 , n210951 , n210952 , n210953 , n210954 , n210955 , n210956 , n210957 , n210958 , 
 n210959 , n210960 , n210961 , n210962 , n210963 , n210964 , n210965 , n210966 , n210967 , n210968 , 
 n210969 , n210970 , n210971 , n210972 , n210973 , n210974 , n210975 , n210976 , n210977 , n210978 , 
 n210979 , n210980 , n210981 , n210982 , n210983 , n210984 , n210985 , n210986 , n210987 , n210988 , 
 n210989 , n210990 , n210991 , n210992 , n210993 , n210994 , n210995 , n210996 , n210997 , n210998 , 
 n210999 , n211000 , n211001 , n211002 , n211003 , n211004 , n211005 , n211006 , n211007 , n211008 , 
 n211009 , n211010 , n211011 , n211012 , n211013 , n211014 , n211015 , n211016 , n211017 , n211018 , 
 n211019 , n211020 , n211021 , n211022 , n211023 , n211024 , n211025 , n211026 , n211027 , n211028 , 
 n211029 , n211030 , n211031 , n211032 , n211033 , n211034 , n211035 , n211036 , n211037 , n211038 , 
 n211039 , n211040 , n211041 , n211042 , n211043 , n211044 , n211045 , n211046 , n211047 , n211048 , 
 n211049 , n211050 , n211051 , n211052 , n211053 , n211054 , n211055 , n211056 , n211057 , n211058 , 
 n211059 , n211060 , n211061 , n211062 , n211063 , n211064 , n211065 , n211066 , n211067 , n211068 , 
 n211069 , n211070 , n211071 , n211072 , n211073 , n211074 , n211075 , n211076 , n211077 , n211078 , 
 n211079 , n211080 , n211081 , n211082 , n211083 , n211084 , n211085 , n211086 , n211087 , n211088 , 
 n211089 , n211090 , n211091 , n211092 , n211093 , n211094 , n211095 , n211096 , n211097 , n211098 , 
 n211099 , n211100 , n211101 , n211102 , n211103 , n211104 , n211105 , n211106 , n211107 , n211108 , 
 n211109 , n211110 , n211111 , n211112 , n211113 , n211114 , n211115 , n211116 , n211117 , n211118 , 
 n211119 , n211120 , n211121 , n211122 , n211123 , n211124 , n211125 , n211126 , n211127 , n211128 , 
 n211129 , n211130 , n211131 , n211132 , n211133 , n211134 , n211135 , n211136 , n211137 , n211138 , 
 n211139 , n211140 , n211141 , n211142 , n211143 , n211144 , n211145 , n211146 , n211147 , n211148 , 
 n211149 , n211150 , n211151 , n211152 , n211153 , n211154 , n211155 , n211156 , n211157 , n211158 , 
 n211159 , n211160 , n211161 , n211162 , n211163 , n211164 , n211165 , n211166 , n211167 , n211168 , 
 n211169 , n211170 , n211171 , n211172 , n211173 , n211174 , n211175 , n211176 , n211177 , n211178 , 
 n211179 , n211180 , n211181 , n211182 , n211183 , n211184 , n211185 , n211186 , n211187 , n211188 , 
 n211189 , n211190 , n211191 , n211192 , n211193 , n211194 , n211195 , n211196 , n211197 , n211198 , 
 n211199 , n211200 , n211201 , n211202 , n211203 , n211204 , n211205 , n211206 , n211207 , n211208 , 
 n211209 , n211210 , n211211 , n211212 , n211213 , n211214 , n211215 , n211216 , n211217 , n211218 , 
 n211219 , n211220 , n211221 , n211222 , n211223 , n211224 , n211225 , n211226 , n211227 , n211228 , 
 n211229 , n211230 , n211231 , n211232 , n211233 , n211234 , n211235 , n211236 , n211237 , n211238 , 
 n211239 , n211240 , n211241 , n211242 , n211243 , n211244 , n211245 , n211246 , n211247 , n211248 , 
 n211249 , n211250 , n211251 , n211252 , n211253 , n211254 , n211255 , n211256 , n211257 , n211258 , 
 n211259 , n211260 , n211261 , n211262 , n211263 , n211264 , n211265 , n211266 , n211267 , n211268 , 
 n211269 , n211270 , n211271 , n211272 , n211273 , n211274 , n211275 , n211276 , n211277 , n211278 , 
 n211279 , n211280 , n211281 , n211282 , n211283 , n211284 , n211285 , n211286 , n211287 , n211288 , 
 n211289 , n211290 , n211291 , n211292 , n211293 , n211294 , n211295 , n211296 , n211297 , n211298 , 
 n211299 , n211300 , n211301 , n211302 , n211303 , n211304 , n211305 , n211306 , n211307 , n211308 , 
 n211309 , n211310 , n211311 , n211312 , n211313 , n211314 , n211315 , n211316 , n211317 , n211318 , 
 n211319 , n211320 , n211321 , n211322 , n211323 , n211324 , n211325 , n211326 , n211327 , n211328 , 
 n211329 , n211330 , n211331 , n211332 , n211333 , n211334 , n211335 , n211336 , n211337 , n211338 , 
 n211339 , n211340 , n211341 , n211342 , n211343 , n211344 , n211345 , n211346 , n211347 , n211348 , 
 n211349 , n211350 , n211351 , n211352 , n211353 , n211354 , n211355 , n211356 , n211357 , n211358 , 
 n211359 , n211360 , n211361 , n211362 , n211363 , n211364 , n211365 , n211366 , n211367 , n211368 , 
 n211369 , n211370 , n211371 , n211372 , n211373 , n211374 , n211375 , n211376 , n211377 , n211378 , 
 n211379 , n211380 , n211381 , n211382 , n211383 , n211384 , n211385 , n211386 , n211387 , n211388 , 
 n211389 , n211390 , n211391 , n211392 , n211393 , n211394 , n211395 , n211396 , n211397 , n211398 , 
 n211399 , n211400 , n211401 , n211402 , n211403 , n211404 , n211405 , n211406 , n211407 , n211408 , 
 n211409 , n211410 , n211411 , n211412 , n211413 , n211414 , n211415 , n211416 , n211417 , n211418 , 
 n211419 , n211420 , n211421 , n211422 , n211423 , n211424 , n211425 , n211426 , n211427 , n211428 , 
 n211429 , n211430 , n211431 , n211432 , n211433 , n211434 , n211435 , n211436 , n211437 , n211438 , 
 n211439 , n211440 , n211441 , n211442 , n211443 , n211444 , n211445 , n211446 , n211447 , n211448 , 
 n211449 , n211450 , n211451 , n211452 , n211453 , n211454 , n211455 , n211456 , n211457 , n211458 , 
 n211459 , n211460 , n211461 , n211462 , n211463 , n211464 , n211465 , n211466 , n211467 , n211468 , 
 n211469 , n211470 , n211471 , n211472 , n211473 , n211474 , n211475 , n211476 , n211477 , n211478 , 
 n211479 , n211480 , n211481 , n211482 , n211483 , n211484 , n211485 , n211486 , n211487 , n211488 , 
 n211489 , n211490 , n211491 , n211492 , n211493 , n211494 , n211495 , n211496 , n211497 , n211498 , 
 n211499 , n211500 , n211501 , n211502 , n211503 , n211504 , n211505 , n211506 , n211507 , n211508 , 
 n211509 , n211510 , n211511 , n211512 , n211513 , n211514 , n211515 , n211516 , n211517 , n211518 , 
 n211519 , n211520 , n211521 , n211522 , n211523 , n211524 , n211525 , n211526 , n211527 , n211528 , 
 n211529 , n211530 , n211531 , n211532 , n211533 , n211534 , n211535 , n211536 , n211537 , n211538 , 
 n211539 , n211540 , n211541 , n211542 , n211543 , n211544 , n211545 , n211546 , n211547 , n211548 , 
 n211549 , n211550 , n211551 , n211552 , n211553 , n211554 , n211555 , n211556 , n211557 , n211558 , 
 n211559 , n211560 , n211561 , n211562 , n211563 , n211564 , n211565 , n211566 , n211567 , n211568 , 
 n211569 , n211570 , n211571 , n211572 , n211573 , n211574 , n211575 , n211576 , n211577 , n211578 , 
 n211579 , n211580 , n211581 , n211582 , n211583 , n211584 , n211585 , n211586 , n211587 , n211588 , 
 n211589 , n211590 , n211591 , n211592 , n211593 , n211594 , n211595 , n211596 , n211597 , n211598 , 
 n211599 , n211600 , n211601 , n211602 , n211603 , n211604 , n211605 , n211606 , n211607 , n211608 , 
 n211609 , n211610 , n211611 , n211612 , n211613 , n211614 , n211615 , n211616 , n211617 , n211618 , 
 n211619 , n211620 , n211621 , n211622 , n211623 , n211624 , n211625 , n211626 , n211627 , n211628 , 
 n211629 , n211630 , n211631 , n211632 , n211633 , n211634 , n211635 , n211636 , n211637 , n211638 , 
 n211639 , n211640 , n211641 , n211642 , n211643 , n211644 , n211645 , n211646 , n211647 , n211648 , 
 n211649 , n211650 , n211651 , n211652 , n211653 , n211654 , n211655 , n211656 , n211657 , n211658 , 
 n211659 , n211660 , n211661 , n211662 , n211663 , n211664 , n211665 , n211666 , n211667 , n211668 , 
 n211669 , n211670 , n211671 , n211672 , n211673 , n211674 , n211675 , n211676 , n211677 , n211678 , 
 n211679 , n211680 , n211681 , n211682 , n211683 , n211684 , n211685 , n211686 , n211687 , n211688 , 
 n211689 , n211690 , n211691 , n211692 , n211693 , n211694 , n211695 , n211696 , n211697 , n211698 , 
 n211699 , n211700 , n211701 , n211702 , n211703 , n211704 , n211705 , n211706 , n211707 , n211708 , 
 n211709 , n211710 , n211711 , n211712 , n211713 , n211714 , n211715 , n211716 , n211717 , n211718 , 
 n211719 , n211720 , n211721 , n211722 , n211723 , n211724 , n211725 , n211726 , n211727 , n211728 , 
 n211729 , n211730 , n211731 , n211732 , n211733 , n211734 , n211735 , n211736 , n211737 , n211738 , 
 n211739 , n211740 , n211741 , n211742 , n211743 , n211744 , n211745 , n211746 , n211747 , n211748 , 
 n211749 , n211750 , n211751 , n211752 , n211753 , n211754 , n211755 , n211756 , n211757 , n211758 , 
 n211759 , n211760 , n211761 , n211762 , n211763 , n211764 , n211765 , n211766 , n211767 , n211768 , 
 n211769 , n211770 , n211771 , n211772 , n211773 , n211774 , n211775 , n211776 , n211777 , n211778 , 
 n211779 , n211780 , n211781 , n211782 , n211783 , n211784 , n211785 , n211786 , n211787 , n211788 , 
 n211789 , n211790 , n211791 , n211792 , n211793 , n211794 , n211795 , n211796 , n211797 , n211798 , 
 n211799 , n211800 , n211801 , n211802 , n211803 , n211804 , n211805 , n211806 , n211807 , n211808 , 
 n211809 , n211810 , n211811 , n211812 , n211813 , n211814 , n211815 , n211816 , n211817 , n211818 , 
 n211819 , n211820 , n211821 , n211822 , n211823 , n211824 , n211825 , n211826 , n211827 , n211828 , 
 n211829 , n211830 , n211831 , n211832 , n211833 , n211834 , n211835 , n211836 , n211837 , n211838 , 
 n211839 , n211840 , n211841 , n211842 , n211843 , n211844 , n211845 , n211846 , n211847 , n211848 , 
 n211849 , n211850 , n211851 , n211852 , n211853 , n211854 , n211855 , n211856 , n211857 , n211858 , 
 n211859 , n211860 , n211861 , n211862 , n211863 , n211864 , n211865 , n211866 , n211867 , n211868 , 
 n211869 , n211870 , n211871 , n211872 , n211873 , n211874 , n211875 , n211876 , n211877 , n211878 , 
 n211879 , n211880 , n211881 , n211882 , n211883 , n211884 , n211885 , n211886 , n211887 , n211888 , 
 n211889 , n211890 , n211891 , n211892 , n211893 , n211894 , n211895 , n211896 , n211897 , n211898 , 
 n211899 , n211900 , n211901 , n211902 , n211903 , n211904 , n211905 , n211906 , n211907 , n211908 , 
 n211909 , n211910 , n211911 , n211912 , n211913 , n211914 , n211915 , n211916 , n211917 , n211918 , 
 n211919 , n211920 , n211921 , n211922 , n211923 , n211924 , n211925 , n211926 , n211927 , n211928 , 
 n211929 , n211930 , n211931 , n211932 , n211933 , n211934 , n211935 , n211936 , n211937 , n211938 , 
 n211939 , n211940 , n211941 , n211942 , n211943 , n211944 , n211945 , n211946 , n211947 , n211948 , 
 n211949 , n211950 , n211951 , n211952 , n211953 , n211954 , n211955 , n211956 , n211957 , n211958 , 
 n211959 , n211960 , n211961 , n211962 , n211963 , n211964 , n211965 , n211966 , n211967 , n211968 , 
 n211969 , n211970 , n211971 , n211972 , n211973 , n211974 , n211975 , n211976 , n211977 , n211978 , 
 n211979 , n211980 , n211981 , n211982 , n211983 , n211984 , n211985 , n211986 , n211987 , n211988 , 
 n211989 , n211990 , n211991 , n211992 , n211993 , n211994 , n211995 , n211996 , n211997 , n211998 , 
 n211999 , n212000 , n212001 , n212002 , n212003 , n212004 , n212005 , n212006 , n212007 , n212008 , 
 n212009 , n212010 , n212011 , n212012 , n212013 , n212014 , n212015 , n212016 , n212017 , n212018 , 
 n212019 , n212020 , n212021 , n212022 , n212023 , n212024 , n212025 , n212026 , n212027 , n212028 , 
 n212029 , n212030 , n212031 , n212032 , n212033 , n212034 , n212035 , n212036 , n212037 , n212038 , 
 n212039 , n212040 , n212041 , n212042 , n212043 , n212044 , n212045 , n212046 , n212047 , n212048 , 
 n212049 , n212050 , n212051 , n212052 , n212053 , n212054 , n212055 , n212056 , n212057 , n212058 , 
 n212059 , n212060 , n212061 , n212062 , n212063 , n212064 , n212065 , n212066 , n212067 , n212068 , 
 n212069 , n212070 , n212071 , n212072 , n212073 , n212074 , n212075 , n212076 , n212077 , n212078 , 
 n212079 , n212080 , n212081 , n212082 , n212083 , n212084 , n212085 , n212086 , n212087 , n212088 , 
 n212089 , n212090 , n212091 , n212092 , n212093 , n212094 , n212095 , n212096 , n212097 , n212098 , 
 n212099 , n212100 , n212101 , n212102 , n212103 , n212104 , n212105 , n212106 , n212107 , n212108 , 
 n212109 , n212110 , n212111 , n212112 , n212113 , n212114 , n212115 , n212116 , n212117 , n212118 , 
 n212119 , n212120 , n212121 , n212122 , n212123 , n212124 , n212125 , n212126 , n212127 , n212128 , 
 n212129 , n212130 , n212131 , n212132 , n212133 , n212134 , n212135 , n212136 , n212137 , n212138 , 
 n212139 , n212140 , n212141 , n212142 , n212143 , n212144 , n212145 , n212146 , n212147 , n212148 , 
 n212149 , n212150 , n212151 , n212152 , n212153 , n212154 , n212155 , n212156 , n212157 , n212158 , 
 n212159 , n212160 , n212161 , n212162 , n212163 , n212164 , n212165 , n212166 , n212167 , n212168 , 
 n212169 , n212170 , n212171 , n212172 , n212173 , n212174 , n212175 , n212176 , n212177 , n212178 , 
 n212179 , n212180 , n212181 , n212182 , n212183 , n212184 , n212185 , n212186 , n212187 , n212188 , 
 n212189 , n212190 , n212191 , n212192 , n212193 , n212194 , n212195 , n212196 , n212197 , n212198 , 
 n212199 , n212200 , n212201 , n212202 , n212203 , n212204 , n212205 , n212206 , n212207 , n212208 , 
 n212209 , n212210 , n212211 , n212212 , n212213 , n212214 , n212215 , n212216 , n212217 , n212218 , 
 n212219 , n212220 , n212221 , n212222 , n212223 , n212224 , n212225 , n212226 , n212227 , n212228 , 
 n212229 , n212230 , n212231 , n212232 , n212233 , n212234 , n212235 , n212236 , n212237 , n212238 , 
 n212239 , n212240 , n212241 , n212242 , n212243 , n212244 , n212245 , n212246 , n212247 , n212248 , 
 n212249 , n212250 , n212251 , n212252 , n212253 , n212254 , n212255 , n212256 , n212257 , n212258 , 
 n212259 , n212260 , n212261 , n212262 , n212263 , n212264 , n212265 , n212266 , n212267 , n212268 , 
 n212269 , n212270 , n212271 , n212272 , n212273 , n212274 , n212275 , n212276 , n212277 , n212278 , 
 n212279 , n212280 , n212281 , n212282 , n212283 , n212284 , n212285 , n212286 , n212287 , n212288 , 
 n212289 , n212290 , n212291 , n212292 , n212293 , n212294 , n212295 , n212296 , n212297 , n212298 , 
 n212299 , n212300 , n212301 , n212302 , n212303 , n212304 , n212305 , n212306 , n212307 , n212308 , 
 n212309 , n212310 , n212311 , n212312 , n212313 , n212314 , n212315 , n212316 , n212317 , n212318 , 
 n212319 , n212320 , n212321 , n212322 , n212323 , n212324 , n212325 , n212326 , n212327 , n212328 , 
 n212329 , n212330 , n212331 , n212332 , n212333 , n212334 , n212335 , n212336 , n212337 , n212338 , 
 n212339 , n212340 , n212341 , n212342 , n212343 , n212344 , n212345 , n212346 , n212347 , n212348 , 
 n212349 , n212350 , n212351 , n212352 , n212353 , n212354 , n212355 , n212356 , n212357 , n212358 , 
 n212359 , n212360 , n212361 , n212362 , n212363 , n212364 , n212365 , n212366 , n212367 , n212368 , 
 n212369 , n212370 , n212371 , n212372 , n212373 , n212374 , n212375 , n212376 , n212377 , n212378 , 
 n212379 , n212380 , n212381 , n212382 , n212383 , n212384 , n212385 , n212386 , n212387 , n212388 , 
 n212389 , n212390 , n212391 , n212392 , n212393 , n212394 , n212395 , n212396 , n212397 , n212398 , 
 n212399 , n212400 , n212401 , n212402 , n212403 , n212404 , n212405 , n212406 , n212407 , n212408 , 
 n212409 , n212410 , n212411 , n212412 , n212413 , n212414 , n212415 , n212416 , n212417 , n212418 , 
 n212419 , n212420 , n212421 , n212422 , n212423 , n212424 , n212425 , n212426 , n212427 , n212428 , 
 n212429 , n212430 , n212431 , n212432 , n212433 , n212434 , n212435 , n212436 , n212437 , n212438 , 
 n212439 , n212440 , n212441 , n212442 , n212443 , n212444 , n212445 , n212446 , n212447 , n212448 , 
 n212449 , n212450 , n212451 , n212452 , n212453 , n212454 , n212455 , n212456 , n212457 , n212458 , 
 n212459 , n212460 , n212461 , n212462 , n212463 , n212464 , n212465 , n212466 , n212467 , n212468 , 
 n212469 , n212470 , n212471 , n212472 , n212473 , n212474 , n212475 , n212476 , n212477 , n212478 , 
 n212479 , n212480 , n212481 , n212482 , n212483 , n212484 , n212485 , n212486 , n212487 , n212488 , 
 n212489 , n212490 , n212491 , n212492 , n212493 , n212494 , n212495 , n212496 , n212497 , n212498 , 
 n212499 , n212500 , n212501 , n212502 , n212503 , n212504 , n212505 , n212506 , n212507 , n212508 , 
 n212509 , n212510 , n212511 , n212512 , n212513 , n212514 , n212515 , n212516 , n212517 , n212518 , 
 n212519 , n212520 , n212521 , n212522 , n212523 , n212524 , n212525 , n212526 , n212527 , n212528 , 
 n212529 , n212530 , n212531 , n212532 , n212533 , n212534 , n212535 , n212536 , n212537 , n212538 , 
 n212539 , n212540 , n212541 , n212542 , n212543 , n212544 , n212545 , n212546 , n212547 , n212548 , 
 n212549 , n212550 , n212551 , n212552 , n212553 , n212554 , n212555 , n212556 , n212557 , n212558 , 
 n212559 , n212560 , n212561 , n212562 , n212563 , n212564 , n212565 , n212566 , n212567 , n212568 , 
 n212569 , n212570 , n212571 , n212572 , n212573 , n212574 , n212575 , n212576 , n212577 , n212578 , 
 n212579 , n212580 , n212581 , n212582 , n212583 , n212584 , n212585 , n212586 , n212587 , n212588 , 
 n212589 , n212590 , n212591 , n212592 , n212593 , n212594 , n212595 , n212596 , n212597 , n212598 , 
 n212599 , n212600 , n212601 , n212602 , n212603 , n212604 , n212605 , n212606 , n212607 , n212608 , 
 n212609 , n212610 , n212611 , n212612 , n212613 , n212614 , n212615 , n212616 , n212617 , n212618 , 
 n212619 , n212620 , n212621 , n212622 , n212623 , n212624 , n212625 , n212626 , n212627 , n212628 , 
 n212629 , n212630 , n212631 , n212632 , n212633 , n212634 , n212635 , n212636 , n212637 , n212638 , 
 n212639 , n212640 , n212641 , n212642 , n212643 , n212644 , n212645 , n212646 , n212647 , n212648 , 
 n212649 , n212650 , n212651 , n212652 , n212653 , n212654 , n212655 , n212656 , n212657 , n212658 , 
 n212659 , n212660 , n212661 , n212662 , n212663 , n212664 , n212665 , n212666 , n212667 , n212668 , 
 n212669 , n212670 , n212671 , n212672 , n212673 , n212674 , n212675 , n212676 , n212677 , n212678 , 
 n212679 , n212680 , n212681 , n212682 , n212683 , n212684 , n212685 , n212686 , n212687 , n212688 , 
 n212689 , n212690 , n212691 , n212692 , n212693 , n212694 , n212695 , n212696 , n212697 , n212698 , 
 n212699 , n212700 , n212701 , n212702 , n212703 , n212704 , n212705 , n212706 , n212707 , n212708 , 
 n212709 , n212710 , n212711 , n212712 , n212713 , n212714 , n212715 , n212716 , n212717 , n212718 , 
 n212719 , n212720 , n212721 , n212722 , n212723 , n212724 , n212725 , n212726 , n212727 , n212728 , 
 n212729 , n212730 , n212731 , n212732 , n212733 , n212734 , n212735 , n212736 , n212737 , n212738 , 
 n212739 , n212740 , n212741 , n212742 , n212743 , n212744 , n212745 , n212746 , n212747 , n212748 , 
 n212749 , n212750 , n212751 , n212752 , n212753 , n212754 , n212755 , n212756 , n212757 , n212758 , 
 n212759 , n212760 , n212761 , n212762 , n212763 , n212764 , n212765 , n212766 , n212767 , n212768 , 
 n212769 , n212770 , n212771 , n212772 , n212773 , n212774 , n212775 , n212776 , n212777 , n212778 , 
 n212779 , n212780 , n212781 , n212782 , n212783 , n212784 , n212785 , n212786 , n212787 , n212788 , 
 n212789 , n212790 , n212791 , n212792 , n212793 , n212794 , n212795 , n212796 , n212797 , n212798 , 
 n212799 , n212800 , n212801 , n212802 , n212803 , n212804 , n212805 , n212806 , n212807 , n212808 , 
 n212809 , n212810 , n212811 , n212812 , n212813 , n212814 , n212815 , n212816 , n212817 , n212818 , 
 n212819 , n212820 , n212821 , n212822 , n212823 , n212824 , n212825 , n212826 , n212827 , n212828 , 
 n212829 , n212830 , n212831 , n212832 , n212833 , n212834 , n212835 , n212836 , n212837 , n212838 , 
 n212839 , n212840 , n212841 , n212842 , n212843 , n212844 , n212845 , n212846 , n212847 , n212848 , 
 n212849 , n212850 , n212851 , n212852 , n212853 , n212854 , n212855 , n212856 , n212857 , n212858 , 
 n212859 , n212860 , n212861 , n212862 , n212863 , n212864 , n212865 , n212866 , n212867 , n212868 , 
 n212869 , n212870 , n212871 , n212872 , n212873 , n212874 , n212875 , n212876 , n212877 , n212878 , 
 n212879 , n212880 , n212881 , n212882 , n212883 , n212884 , n212885 , n212886 , n212887 , n212888 , 
 n212889 , n212890 , n212891 , n212892 , n212893 , n212894 , n212895 , n212896 , n212897 , n212898 , 
 n212899 , n212900 , n212901 , n212902 , n212903 , n212904 , n212905 , n212906 , n212907 , n212908 , 
 n212909 , n212910 , n212911 , n212912 , n212913 , n212914 , n212915 , n212916 , n212917 , n212918 , 
 n212919 , n212920 , n212921 , n212922 , n212923 , n212924 , n212925 , n212926 , n212927 , n212928 , 
 n212929 , n212930 , n212931 , n212932 , n212933 , n212934 , n212935 , n212936 , n212937 , n212938 , 
 n212939 , n212940 , n212941 , n212942 , n212943 , n212944 , n212945 , n212946 , n212947 , n212948 , 
 n212949 , n212950 , n212951 , n212952 , n212953 , n212954 , n212955 , n212956 , n212957 , n212958 , 
 n212959 , n212960 , n212961 , n212962 , n212963 , n212964 , n212965 , n212966 , n212967 , n212968 , 
 n212969 , n212970 , n212971 , n212972 , n212973 , n212974 , n212975 , n212976 , n212977 , n212978 , 
 n212979 , n212980 , n212981 , n212982 , n212983 , n212984 , n212985 , n212986 , n212987 , n212988 , 
 n212989 , n212990 , n212991 , n212992 , n212993 , n212994 , n212995 , n212996 , n212997 , n212998 , 
 n212999 , n213000 , n213001 , n213002 , n213003 , n213004 , n213005 , n213006 , n213007 , n213008 , 
 n213009 , n213010 , n213011 , n213012 , n213013 , n213014 , n213015 , n213016 , n213017 , n213018 , 
 n213019 , n213020 , n213021 , n213022 , n213023 , n213024 , n213025 , n213026 , n213027 , n213028 , 
 n213029 , n213030 , n213031 , n213032 , n213033 , n213034 , n213035 , n213036 , n213037 , n213038 , 
 n213039 , n213040 , n213041 , n213042 , n213043 , n213044 , n213045 , n213046 , n213047 , n213048 , 
 n213049 , n213050 , n213051 , n213052 , n213053 , n213054 , n213055 , n213056 , n213057 , n213058 , 
 n213059 , n213060 , n213061 , n213062 , n213063 , n213064 , n213065 , n213066 , n213067 , n213068 , 
 n213069 , n213070 , n213071 , n213072 , n213073 , n213074 , n213075 , n213076 , n213077 , n213078 , 
 n213079 , n213080 , n213081 , n213082 , n213083 , n213084 , n213085 , n213086 , n213087 , n213088 , 
 n213089 , n213090 , n213091 , n213092 , n213093 , n213094 , n213095 , n213096 , n213097 , n213098 , 
 n213099 , n213100 , n213101 , n213102 , n213103 , n213104 , n213105 , n213106 , n213107 , n213108 , 
 n213109 , n213110 , n213111 , n213112 , n213113 , n213114 , n213115 , n213116 , n213117 , n213118 , 
 n213119 , n213120 , n213121 , n213122 , n213123 , n213124 , n213125 , n213126 , n213127 , n213128 , 
 n213129 , n213130 , n213131 , n213132 , n213133 , n213134 , n213135 , n213136 , n213137 , n213138 , 
 n213139 , n213140 , n213141 , n213142 , n213143 , n213144 , n213145 , n213146 , n213147 , n213148 , 
 n213149 , n213150 , n213151 , n213152 , n213153 , n213154 , n213155 , n213156 , n213157 , n213158 , 
 n213159 , n213160 , n213161 , n213162 , n213163 , n213164 , n213165 , n213166 , n213167 , n213168 , 
 n213169 , n213170 , n213171 , n213172 , n213173 , n213174 , n213175 , n213176 , n213177 , n213178 , 
 n213179 , n213180 , n213181 , n213182 , n213183 , n213184 , n213185 , n213186 , n213187 , n213188 , 
 n213189 , n213190 , n213191 , n213192 , n213193 , n213194 , n213195 , n213196 , n213197 , n213198 , 
 n213199 , n213200 , n213201 , n213202 , n213203 , n213204 , n213205 , n213206 , n213207 , n213208 , 
 n213209 , n213210 , n213211 , n213212 , n213213 , n213214 , n213215 , n213216 , n213217 , n213218 , 
 n213219 , n213220 , n213221 , n213222 , n213223 , n213224 , n213225 , n213226 , n213227 , n213228 , 
 n213229 , n213230 , n213231 , n213232 , n213233 , n213234 , n213235 , n213236 , n213237 , n213238 , 
 n213239 , n213240 , n213241 , n213242 , n213243 , n213244 , n213245 , n213246 , n213247 , n213248 , 
 n213249 , n213250 , n213251 , n213252 , n213253 , n213254 , n213255 , n213256 , n213257 , n213258 , 
 n213259 , n213260 , n213261 , n213262 , n213263 , n213264 , n213265 , n213266 , n213267 , n213268 , 
 n213269 , n213270 , n213271 , n213272 , n213273 , n213274 , n213275 , n213276 , n213277 , n213278 , 
 n213279 , n213280 , n213281 , n213282 , n213283 , n213284 , n213285 , n213286 , n213287 , n213288 , 
 n213289 , n213290 , n213291 , n213292 , n213293 , n213294 , n213295 , n213296 , n213297 , n213298 , 
 n213299 , n213300 , n213301 , n213302 , n213303 , n213304 , n213305 , n213306 , n213307 , n213308 , 
 n213309 , n213310 , n213311 , n213312 , n213313 , n213314 , n213315 , n213316 , n213317 , n213318 , 
 n213319 , n213320 , n213321 , n213322 , n213323 , n213324 , n213325 , n213326 , n213327 , n213328 , 
 n213329 , n213330 , n213331 , n213332 , n213333 , n213334 , n213335 , n213336 , n213337 , n213338 , 
 n213339 , n213340 , n213341 , n213342 , n213343 , n213344 , n213345 , n213346 , n213347 , n213348 , 
 n213349 , n213350 , n213351 , n213352 , n213353 , n213354 , n213355 , n213356 , n213357 , n213358 , 
 n213359 , n213360 , n213361 , n213362 , n213363 , n213364 , n213365 , n213366 , n213367 , n213368 , 
 n213369 , n213370 , n213371 , n213372 , n213373 , n213374 , n213375 , n213376 , n213377 , n213378 , 
 n213379 , n213380 , n213381 , n213382 , n213383 , n213384 , n213385 , n213386 , n213387 , n213388 , 
 n213389 , n213390 , n213391 , n213392 , n213393 , n213394 , n213395 , n213396 , n213397 , n213398 , 
 n213399 , n213400 , n213401 , n213402 , n213403 , n213404 , n213405 , n213406 , n213407 , n213408 , 
 n213409 , n213410 , n213411 , n213412 , n213413 , n213414 , n213415 , n213416 , n213417 , n213418 , 
 n213419 , n213420 , n213421 , n213422 , n213423 , n213424 , n213425 , n213426 , n213427 , n213428 , 
 n213429 , n213430 , n213431 , n213432 , n213433 , n213434 , n213435 , n213436 , n213437 , n213438 , 
 n213439 , n213440 , n213441 , n213442 , n213443 , n213444 , n213445 , n213446 , n213447 , n213448 , 
 n213449 , n213450 , n213451 , n213452 , n213453 , n213454 , n213455 , n213456 , n213457 , n213458 , 
 n213459 , n213460 , n213461 , n213462 , n213463 , n213464 , n213465 , n213466 , n213467 , n213468 , 
 n213469 , n213470 , n213471 , n213472 , n213473 , n213474 , n213475 , n213476 , n213477 , n213478 , 
 n213479 , n213480 , n213481 , n213482 , n213483 , n213484 , n213485 , n213486 , n213487 , n213488 , 
 n213489 , n213490 , n213491 , n213492 , n213493 , n213494 , n213495 , n213496 , n213497 , n213498 , 
 n213499 , n213500 , n213501 , n213502 , n213503 , n213504 , n213505 , n213506 , n213507 , n213508 , 
 n213509 , n213510 , n213511 , n213512 , n213513 , n213514 , n213515 , n213516 , n213517 , n213518 , 
 n213519 , n213520 , n213521 , n213522 , n213523 , n213524 , n213525 , n213526 , n213527 , n213528 , 
 n213529 , n213530 , n213531 , n213532 , n213533 , n213534 , n213535 , n213536 , n213537 , n213538 , 
 n213539 , n213540 , n213541 , n213542 , n213543 , n213544 , n213545 , n213546 , n213547 , n213548 , 
 n213549 , n213550 , n213551 , n213552 , n213553 , n213554 , n213555 , n213556 , n213557 , n213558 , 
 n213559 , n213560 , n213561 , n213562 , n213563 , n213564 , n213565 , n213566 , n213567 , n213568 , 
 n213569 , n213570 , n213571 , n213572 , n213573 , n213574 , n213575 , n213576 , n213577 , n213578 , 
 n213579 , n213580 , n213581 , n213582 , n213583 , n213584 , n213585 , n213586 , n213587 , n213588 , 
 n213589 , n213590 , n213591 , n213592 , n213593 , n213594 , n213595 , n213596 , n213597 , n213598 , 
 n213599 , n213600 , n213601 , n213602 , n213603 , n213604 , n213605 , n213606 , n213607 , n213608 , 
 n213609 , n213610 , n213611 , n213612 , n213613 , n213614 , n213615 , n213616 , n213617 , n213618 , 
 n213619 , n213620 , n213621 , n213622 , n213623 , n213624 , n213625 , n213626 , n213627 , n213628 , 
 n213629 , n213630 , n213631 , n213632 , n213633 , n213634 , n213635 , n213636 , n213637 , n213638 , 
 n213639 , n213640 , n213641 , n213642 , n213643 , n213644 , n213645 , n213646 , n213647 , n213648 , 
 n213649 , n213650 , n213651 , n213652 , n213653 , n213654 , n213655 , n213656 , n213657 , n213658 , 
 n213659 , n213660 , n213661 , n213662 , n213663 , n213664 , n213665 , n213666 , n213667 , n213668 , 
 n213669 , n213670 , n213671 , n213672 , n213673 , n213674 , n213675 , n213676 , n213677 , n213678 , 
 n213679 , n213680 , n213681 , n213682 , n213683 , n213684 , n213685 , n213686 , n213687 , n213688 , 
 n213689 , n213690 , n213691 , n213692 , n213693 , n213694 , n213695 , n213696 , n213697 , n213698 , 
 n213699 , n213700 , n213701 , n213702 , n213703 , n213704 , n213705 , n213706 , n213707 , n213708 , 
 n213709 , n213710 , n213711 , n213712 , n213713 , n213714 , n213715 , n213716 , n213717 , n213718 , 
 n213719 , n213720 , n213721 , n213722 , n213723 , n213724 , n213725 , n213726 , n213727 , n213728 , 
 n213729 , n213730 , n213731 , n213732 , n213733 , n213734 , n213735 , n213736 , n213737 , n213738 , 
 n213739 , n213740 , n213741 , n213742 , n213743 , n213744 , n213745 , n213746 , n213747 , n213748 , 
 n213749 , n213750 , n213751 , n213752 , n213753 , n213754 , n213755 , n213756 , n213757 , n213758 , 
 n213759 , n213760 , n213761 , n213762 , n213763 , n213764 , n213765 , n213766 , n213767 , n213768 , 
 n213769 , n213770 , n213771 , n213772 , n213773 , n213774 , n213775 , n213776 , n213777 , n213778 , 
 n213779 , n213780 , n213781 , n213782 , n213783 , n213784 , n213785 , n213786 , n213787 , n213788 , 
 n213789 , n213790 , n213791 , n213792 , n213793 , n213794 , n213795 , n213796 , n213797 , n213798 , 
 n213799 , n213800 , n213801 , n213802 , n213803 , n213804 , n213805 , n213806 , n213807 , n213808 , 
 n213809 , n213810 , n213811 , n213812 , n213813 , n213814 , n213815 , n213816 , n213817 , n213818 , 
 n213819 , n213820 , n213821 , n213822 , n213823 , n213824 , n213825 , n213826 , n213827 , n213828 , 
 n213829 , n213830 , n213831 , n213832 , n213833 , n213834 , n213835 , n213836 , n213837 , n213838 , 
 n213839 , n213840 , n213841 , n213842 , n213843 , n213844 , n213845 , n213846 , n213847 , n213848 , 
 n213849 , n213850 , n213851 , n213852 , n213853 , n213854 , n213855 , n213856 , n213857 , n213858 , 
 n213859 , n213860 , n213861 , n213862 , n213863 , n213864 , n213865 , n213866 , n213867 , n213868 , 
 n213869 , n213870 , n213871 , n213872 , n213873 , n213874 , n213875 , n213876 , n213877 , n213878 , 
 n213879 , n213880 , n213881 , n213882 , n213883 , n213884 , n213885 , n213886 , n213887 , n213888 , 
 n213889 , n213890 , n213891 , n213892 , n213893 , n213894 , n213895 , n213896 , n213897 , n213898 , 
 n213899 , n213900 , n213901 , n213902 , n213903 , n213904 , n213905 , n213906 , n213907 , n213908 , 
 n213909 , n213910 , n213911 , n213912 , n213913 , n213914 , n213915 , n213916 , n213917 , n213918 , 
 n213919 , n213920 , n213921 , n213922 , n213923 , n213924 , n213925 , n213926 , n213927 , n213928 , 
 n213929 , n213930 , n213931 , n213932 , n213933 , n213934 , n213935 , n213936 , n213937 , n213938 , 
 n213939 , n213940 , n213941 , n213942 , n213943 , n213944 , n213945 , n213946 , n213947 , n213948 , 
 n213949 , n213950 , n213951 , n213952 , n213953 , n213954 , n213955 , n213956 , n213957 , n213958 , 
 n213959 , n213960 , n213961 , n213962 , n213963 , n213964 , n213965 , n213966 , n213967 , n213968 , 
 n213969 , n213970 , n213971 , n213972 , n213973 , n213974 , n213975 , n213976 , n213977 , n213978 , 
 n213979 , n213980 , n213981 , n213982 , n213983 , n213984 , n213985 , n213986 , n213987 , n213988 , 
 n213989 , n213990 , n213991 , n213992 , n213993 , n213994 , n213995 , n213996 , n213997 , n213998 , 
 n213999 , n214000 , n214001 , n214002 , n214003 , n214004 , n214005 , n214006 , n214007 , n214008 , 
 n214009 , n214010 , n214011 , n214012 , n214013 , n214014 , n214015 , n214016 , n214017 , n214018 , 
 n214019 , n214020 , n214021 , n214022 , n214023 , n214024 , n214025 , n214026 , n214027 , n214028 , 
 n214029 , n214030 , n214031 , n214032 , n214033 , n214034 , n214035 , n214036 , n214037 , n214038 , 
 n214039 , n214040 , n214041 , n214042 , n214043 , n214044 , n214045 , n214046 , n214047 , n214048 , 
 n214049 , n214050 , n214051 , n214052 , n214053 , n214054 , n214055 , n214056 , n214057 , n214058 , 
 n214059 , n214060 , n214061 , n214062 , n214063 , n214064 , n214065 , n214066 , n214067 , n214068 , 
 n214069 , n214070 , n214071 , n214072 , n214073 , n214074 , n214075 , n214076 , n214077 , n214078 , 
 n214079 , n214080 , n214081 , n214082 , n214083 , n214084 , n214085 , n214086 , n214087 , n214088 , 
 n214089 , n214090 , n214091 , n214092 , n214093 , n214094 , n214095 , n214096 , n214097 , n214098 , 
 n214099 , n214100 , n214101 , n214102 , n214103 , n214104 , n214105 , n214106 , n214107 , n214108 , 
 n214109 , n214110 , n214111 , n214112 , n214113 , n214114 , n214115 , n214116 , n214117 , n214118 , 
 n214119 , n214120 , n214121 , n214122 , n214123 , n214124 , n214125 , n214126 , n214127 , n214128 , 
 n214129 , n214130 , n214131 , n214132 , n214133 , n214134 , n214135 , n214136 , n214137 , n214138 , 
 n214139 , n214140 , n214141 , n214142 , n214143 , n214144 , n214145 , n214146 , n214147 , n214148 , 
 n214149 , n214150 , n214151 , n214152 , n214153 , n214154 , n214155 , n214156 , n214157 , n214158 , 
 n214159 , n214160 , n214161 , n214162 , n214163 , n214164 , n214165 , n214166 , n214167 , n214168 , 
 n214169 , n214170 , n214171 , n214172 , n214173 , n214174 , n214175 , n214176 , n214177 , n214178 , 
 n214179 , n214180 , n214181 , n214182 , n214183 , n214184 , n214185 , n214186 , n214187 , n214188 , 
 n214189 , n214190 , n214191 , n214192 , n214193 , n214194 , n214195 , n214196 , n214197 , n214198 , 
 n214199 , n214200 , n214201 , n214202 , n214203 , n214204 , n214205 , n214206 , n214207 , n214208 , 
 n214209 , n214210 , n214211 , n214212 , n214213 , n214214 , n214215 , n214216 , n214217 , n214218 , 
 n214219 , n214220 , n214221 , n214222 , n214223 , n214224 , n214225 , n214226 , n214227 , n214228 , 
 n214229 , n214230 , n214231 , n214232 , n214233 , n214234 , n214235 , n214236 , n214237 , n214238 , 
 n214239 , n214240 , n214241 , n214242 , n214243 , n214244 , n214245 , n214246 , n214247 , n214248 , 
 n214249 , n214250 , n214251 , n214252 , n214253 , n214254 , n214255 , n214256 , n214257 , n214258 , 
 n214259 , n214260 , n214261 , n214262 , n214263 , n214264 , n214265 , n214266 , n214267 , n214268 , 
 n214269 , n214270 , n214271 , n214272 , n214273 , n214274 , n214275 , n214276 , n214277 , n214278 , 
 n214279 , n214280 , n214281 , n214282 , n214283 , n214284 , n214285 , n214286 , n214287 , n214288 , 
 n214289 , n214290 , n214291 , n214292 , n214293 , n214294 , n214295 , n214296 , n214297 , n214298 , 
 n214299 , n214300 , n214301 , n214302 , n214303 , n214304 , n214305 , n214306 , n214307 , n214308 , 
 n214309 , n214310 , n214311 , n214312 , n214313 , n214314 , n214315 , n214316 , n214317 , n214318 , 
 n214319 , n214320 , n214321 , n214322 , n214323 , n214324 , n214325 , n214326 , n214327 , n214328 , 
 n214329 , n214330 , n214331 , n214332 , n214333 , n214334 , n214335 , n214336 , n214337 , n214338 , 
 n214339 , n214340 , n214341 , n214342 , n214343 , n214344 , n214345 , n214346 , n214347 , n214348 , 
 n214349 , n214350 , n214351 , n214352 , n214353 , n214354 , n214355 , n214356 , n214357 , n214358 , 
 n214359 , n214360 , n214361 , n214362 , n214363 , n214364 , n214365 , n214366 , n214367 , n214368 , 
 n214369 , n214370 , n214371 , n214372 , n214373 , n214374 , n214375 , n214376 , n214377 , n214378 , 
 n214379 , n214380 , n214381 , n214382 , n214383 , n214384 , n214385 , n214386 , n214387 , n214388 , 
 n214389 , n214390 , n214391 , n214392 , n214393 , n214394 , n214395 , n214396 , n214397 , n214398 , 
 n214399 , n214400 , n214401 , n214402 , n214403 , n214404 , n214405 , n214406 , n214407 , n214408 , 
 n214409 , n214410 , n214411 , n214412 , n214413 , n214414 , n214415 , n214416 , n214417 , n214418 , 
 n214419 , n214420 , n214421 , n214422 , n214423 , n214424 , n214425 , n214426 , n214427 , n214428 , 
 n214429 , n214430 , n214431 , n214432 , n214433 , n214434 , n214435 , n214436 , n214437 , n214438 , 
 n214439 , n214440 , n214441 , n214442 , n214443 , n214444 , n214445 , n214446 , n214447 , n214448 , 
 n214449 , n214450 , n214451 , n214452 , n214453 , n214454 , n214455 , n214456 , n214457 , n214458 , 
 n214459 , n214460 , n214461 , n214462 , n214463 , n214464 , n214465 , n214466 , n214467 , n214468 , 
 n214469 , n214470 , n214471 , n214472 , n214473 , n214474 , n214475 , n214476 , n214477 , n214478 , 
 n214479 , n214480 , n214481 , n214482 , n214483 , n214484 , n214485 , n214486 , n214487 , n214488 , 
 n214489 , n214490 , n214491 , n214492 , n214493 , n214494 , n214495 , n214496 , n214497 , n214498 , 
 n214499 , n214500 , n214501 , n214502 , n214503 , n214504 , n214505 , n214506 , n214507 , n214508 , 
 n214509 , n214510 , n214511 , n214512 , n214513 , n214514 , n214515 , n214516 , n214517 , n214518 , 
 n214519 , n214520 , n214521 , n214522 , n214523 , n214524 , n214525 , n214526 , n214527 , n214528 , 
 n214529 , n214530 , n214531 , n214532 , n214533 , n214534 , n214535 , n214536 , n214537 , n214538 , 
 n214539 , n214540 , n214541 , n214542 , n214543 , n214544 , n214545 , n214546 , n214547 , n214548 , 
 n214549 , n214550 , n214551 , n214552 , n214553 , n214554 , n214555 , n214556 , n214557 , n214558 , 
 n214559 , n214560 , n214561 , n214562 , n214563 , n214564 , n214565 , n214566 , n214567 , n214568 , 
 n214569 , n214570 , n214571 , n214572 , n214573 , n214574 , n214575 , n214576 , n214577 , n214578 , 
 n214579 , n214580 , n214581 , n214582 , n214583 , n214584 , n214585 , n214586 , n214587 , n214588 , 
 n214589 , n214590 , n214591 , n214592 , n214593 , n214594 , n214595 , n214596 , n214597 , n214598 , 
 n214599 , n214600 , n214601 , n214602 , n214603 , n214604 , n214605 , n214606 , n214607 , n214608 , 
 n214609 , n214610 , n214611 , n214612 , n214613 , n214614 , n214615 , n214616 , n214617 , n214618 , 
 n214619 , n214620 , n214621 , n214622 , n214623 , n214624 , n214625 , n214626 , n214627 , n214628 , 
 n214629 , n214630 , n214631 , n214632 , n214633 , n214634 , n214635 , n214636 , n214637 , n214638 , 
 n214639 , n214640 , n214641 , n214642 , n214643 , n214644 , n214645 , n214646 , n214647 , n214648 , 
 n214649 , n214650 , n214651 , n214652 , n214653 , n214654 , n214655 , n214656 , n214657 , n214658 , 
 n214659 , n214660 , n214661 , n214662 , n214663 , n214664 , n214665 , n214666 , n214667 , n214668 , 
 n214669 , n214670 , n214671 , n214672 , n214673 , n214674 , n214675 , n214676 , n214677 , n214678 , 
 n214679 , n214680 , n214681 , n214682 , n214683 , n214684 , n214685 , n214686 , n214687 , n214688 , 
 n214689 , n214690 , n214691 , n214692 , n214693 , n214694 , n214695 , n214696 , n214697 , n214698 , 
 n214699 , n214700 , n214701 , n214702 , n214703 , n214704 , n214705 , n214706 , n214707 , n214708 , 
 n214709 , n214710 , n214711 , n214712 , n214713 , n214714 , n214715 , n214716 , n214717 , n214718 , 
 n214719 , n214720 , n214721 , n214722 , n214723 , n214724 , n214725 , n214726 , n214727 , n214728 , 
 n214729 , n214730 , n214731 , n214732 , n214733 , n214734 , n214735 , n214736 , n214737 , n214738 , 
 n214739 , n214740 , n214741 , n214742 , n214743 , n214744 , n214745 , n214746 , n214747 , n214748 , 
 n214749 , n214750 , n214751 , n214752 , n214753 , n214754 , n214755 , n214756 , n214757 , n214758 , 
 n214759 , n214760 , n214761 , n214762 , n214763 , n214764 , n214765 , n214766 , n214767 , n214768 , 
 n214769 , n214770 , n214771 , n214772 , n214773 , n214774 , n214775 , n214776 , n214777 , n214778 , 
 n214779 , n214780 , n214781 , n214782 , n214783 , n214784 , n214785 , n214786 , n214787 , n214788 , 
 n214789 , n214790 , n214791 , n214792 , n214793 , n214794 , n214795 , n214796 , n214797 , n214798 , 
 n214799 , n214800 , n214801 , n214802 , n214803 , n214804 , n214805 , n214806 , n214807 , n214808 , 
 n214809 , n214810 , n214811 , n214812 , n214813 , n214814 , n214815 , n214816 , n214817 , n214818 , 
 n214819 , n214820 , n214821 , n214822 , n214823 , n214824 , n214825 , n214826 , n214827 , n214828 , 
 n214829 , n214830 , n214831 , n214832 , n214833 , n214834 , n214835 , n214836 , n214837 , n214838 , 
 n214839 , n214840 , n214841 , n214842 , n214843 , n214844 , n214845 , n214846 , n214847 , n214848 , 
 n214849 , n214850 , n214851 , n214852 , n214853 , n214854 , n214855 , n214856 , n214857 , n214858 , 
 n214859 , n214860 , n214861 , n214862 , n214863 , n214864 , n214865 , n214866 , n214867 , n214868 , 
 n214869 , n214870 , n214871 , n214872 , n214873 , n214874 , n214875 , n214876 , n214877 , n214878 , 
 n214879 , n214880 , n214881 , n214882 , n214883 , n214884 , n214885 , n214886 , n214887 , n214888 , 
 n214889 , n214890 , n214891 , n214892 , n214893 , n214894 , n214895 , n214896 , n214897 , n214898 , 
 n214899 , n214900 , n214901 , n214902 , n214903 , n214904 , n214905 , n214906 , n214907 , n214908 , 
 n214909 , n214910 , n214911 , n214912 , n214913 , n214914 , n214915 , n214916 , n214917 , n214918 , 
 n214919 , n214920 , n214921 , n214922 , n214923 , n214924 , n214925 , n214926 , n214927 , n214928 , 
 n214929 , n214930 , n214931 , n214932 , n214933 , n214934 , n214935 , n214936 , n214937 , n214938 , 
 n214939 , n214940 , n214941 , n214942 , n214943 , n214944 , n214945 , n214946 , n214947 , n214948 , 
 n214949 , n214950 , n214951 , n214952 , n214953 , n214954 , n214955 , n214956 , n214957 , n214958 , 
 n214959 , n214960 , n214961 , n214962 , n214963 , n214964 , n214965 , n214966 , n214967 , n214968 , 
 n214969 , n214970 , n214971 , n214972 , n214973 , n214974 , n214975 , n214976 , n214977 , n214978 , 
 n214979 , n214980 , n214981 , n214982 , n214983 , n214984 , n214985 , n214986 , n214987 , n214988 , 
 n214989 , n214990 , n214991 , n214992 , n214993 , n214994 , n214995 , n214996 , n214997 , n214998 , 
 n214999 , n215000 , n215001 , n215002 , n215003 , n215004 , n215005 , n215006 , n215007 , n215008 , 
 n215009 , n215010 , n215011 , n215012 , n215013 , n215014 , n215015 , n215016 , n215017 , n215018 , 
 n215019 , n215020 , n215021 , n215022 , n215023 , n215024 , n215025 , n215026 , n215027 , n215028 , 
 n215029 , n215030 , n215031 , n215032 , n215033 , n215034 , n215035 , n215036 , n215037 , n215038 , 
 n215039 , n215040 , n215041 , n215042 , n215043 , n215044 , n215045 , n215046 , n215047 , n215048 , 
 n215049 , n215050 , n215051 , n215052 , n215053 , n215054 , n215055 , n215056 , n215057 , n215058 , 
 n215059 , n215060 , n215061 , n215062 , n215063 , n215064 , n215065 , n215066 , n215067 , n215068 , 
 n215069 , n215070 , n215071 , n215072 , n215073 , n215074 , n215075 , n215076 , n215077 , n215078 , 
 n215079 , n215080 , n215081 , n215082 , n215083 , n215084 , n215085 , n215086 , n215087 , n215088 , 
 n215089 , n215090 , n215091 , n215092 , n215093 , n215094 , n215095 , n215096 , n215097 , n215098 , 
 n215099 , n215100 , n215101 , n215102 , n215103 , n215104 , n215105 , n215106 , n215107 , n215108 , 
 n215109 , n215110 , n215111 , n215112 , n215113 , n215114 , n215115 , n215116 , n215117 , n215118 , 
 n215119 , n215120 , n215121 , n215122 , n215123 , n215124 , n215125 , n215126 , n215127 , n215128 , 
 n215129 , n215130 , n215131 , n215132 , n215133 , n215134 , n215135 , n215136 , n215137 , n215138 , 
 n215139 , n215140 , n215141 , n215142 , n215143 , n215144 , n215145 , n215146 , n215147 , n215148 , 
 n215149 , n215150 , n215151 , n215152 , n215153 , n215154 , n215155 , n215156 , n215157 , n215158 , 
 n215159 , n215160 , n215161 , n215162 , n215163 , n215164 , n215165 , n215166 , n215167 , n215168 , 
 n215169 , n215170 , n215171 , n215172 , n215173 , n215174 , n215175 , n215176 , n215177 , n215178 , 
 n215179 , n215180 , n215181 , n215182 , n215183 , n215184 , n215185 , n215186 , n215187 , n215188 , 
 n215189 , n215190 , n215191 , n215192 , n215193 , n215194 , n215195 , n215196 , n215197 , n215198 , 
 n215199 , n215200 , n215201 , n215202 , n215203 , n215204 , n215205 , n215206 , n215207 , n215208 , 
 n215209 , n215210 , n215211 , n215212 , n215213 , n215214 , n215215 , n215216 , n215217 , n215218 , 
 n215219 , n215220 , n215221 , n215222 , n215223 , n215224 , n215225 , n215226 , n215227 , n215228 , 
 n215229 , n215230 , n215231 , n215232 , n215233 , n215234 , n215235 , n215236 , n215237 , n215238 , 
 n215239 , n215240 , n215241 , n215242 , n215243 , n215244 , n215245 , n215246 , n215247 , n215248 , 
 n215249 , n215250 , n215251 , n215252 , n215253 , n215254 , n215255 , n215256 , n215257 , n215258 , 
 n215259 , n215260 , n215261 , n215262 , n215263 , n215264 , n215265 , n215266 , n215267 , n215268 , 
 n215269 , n215270 , n215271 , n215272 , n215273 , n215274 , n215275 , n215276 , n215277 , n215278 , 
 n215279 , n215280 , n215281 , n215282 , n215283 , n215284 , n215285 , n215286 , n215287 , n215288 , 
 n215289 , n215290 , n215291 , n215292 , n215293 , n215294 , n215295 , n215296 , n215297 , n215298 , 
 n215299 , n215300 , n215301 , n215302 , n215303 , n215304 , n215305 , n215306 , n215307 , n215308 , 
 n215309 , n215310 , n215311 , n215312 , n215313 , n215314 , n215315 , n215316 , n215317 , n215318 , 
 n215319 , n215320 , n215321 , n215322 , n215323 , n215324 , n215325 , n215326 , n215327 , n215328 , 
 n215329 , n215330 , n215331 , n215332 , n215333 , n215334 , n215335 , n215336 , n215337 , n215338 , 
 n215339 , n215340 , n215341 , n215342 , n215343 , n215344 , n215345 , n215346 , n215347 , n215348 , 
 n215349 , n215350 , n215351 , n215352 , n215353 , n215354 , n215355 , n215356 , n215357 , n215358 , 
 n215359 , n215360 , n215361 , n215362 , n215363 , n215364 , n215365 , n215366 , n215367 , n215368 , 
 n215369 , n215370 , n215371 , n215372 , n215373 , n215374 , n215375 , n215376 , n215377 , n215378 , 
 n215379 , n215380 , n215381 , n215382 , n215383 , n215384 , n215385 , n215386 , n215387 , n215388 , 
 n215389 , n215390 , n215391 , n215392 , n215393 , n215394 , n215395 , n215396 , n215397 , n215398 , 
 n215399 , n215400 , n215401 , n215402 , n215403 , n215404 , n215405 , n215406 , n215407 , n215408 , 
 n215409 , n215410 , n215411 , n215412 , n215413 , n215414 , n215415 , n215416 , n215417 , n215418 , 
 n215419 , n215420 , n215421 , n215422 , n215423 , n215424 , n215425 , n215426 , n215427 , n215428 , 
 n215429 , n215430 , n215431 , n215432 , n215433 , n215434 , n215435 , n215436 , n215437 , n215438 , 
 n215439 , n215440 , n215441 , n215442 , n215443 , n215444 , n215445 , n215446 , n215447 , n215448 , 
 n215449 , n215450 , n215451 , n215452 , n215453 , n215454 , n215455 , n215456 , n215457 , n215458 , 
 n215459 , n215460 , n215461 , n215462 , n215463 , n215464 , n215465 , n215466 , n215467 , n215468 , 
 n215469 , n215470 , n215471 , n215472 , n215473 , n215474 , n215475 , n215476 , n215477 , n215478 , 
 n215479 , n215480 , n215481 , n215482 , n215483 , n215484 , n215485 , n215486 , n215487 , n215488 , 
 n215489 , n215490 , n215491 , n215492 , n215493 , n215494 , n215495 , n215496 , n215497 , n215498 , 
 n215499 , n215500 , n215501 , n215502 , n215503 , n215504 , n215505 , n215506 , n215507 , n215508 , 
 n215509 , n215510 , n215511 , n215512 , n215513 , n215514 , n215515 , n215516 , n215517 , n215518 , 
 n215519 , n215520 , n215521 , n215522 , n215523 , n215524 , n215525 , n215526 , n215527 , n215528 , 
 n215529 , n215530 , n215531 , n215532 , n215533 , n215534 , n215535 , n215536 , n215537 , n215538 , 
 n215539 , n215540 , n215541 , n215542 , n215543 , n215544 , n215545 , n215546 , n215547 , n215548 , 
 n215549 , n215550 , n215551 , n215552 , n215553 , n215554 , n215555 , n215556 , n215557 , n215558 , 
 n215559 , n215560 , n215561 , n215562 , n215563 , n215564 , n215565 , n215566 , n215567 , n215568 , 
 n215569 , n215570 , n215571 , n215572 , n215573 , n215574 , n215575 , n215576 , n215577 , n215578 , 
 n215579 , n215580 , n215581 , n215582 , n215583 , n215584 , n215585 , n215586 , n215587 , n215588 , 
 n215589 , n215590 , n215591 , n215592 , n215593 , n215594 , n215595 , n215596 , n215597 , n215598 , 
 n215599 , n215600 , n215601 , n215602 , n215603 , n215604 , n215605 , n215606 , n215607 , n215608 , 
 n215609 , n215610 , n215611 , n215612 , n215613 , n215614 , n215615 , n215616 , n215617 , n215618 , 
 n215619 , n215620 , n215621 , n215622 , n215623 , n215624 , n215625 , n215626 , n215627 , n215628 , 
 n215629 , n215630 , n215631 , n215632 , n215633 , n215634 , n215635 , n215636 , n215637 , n215638 , 
 n215639 , n215640 , n215641 , n215642 , n215643 , n215644 , n215645 , n215646 , n215647 , n215648 , 
 n215649 , n215650 , n215651 , n215652 , n215653 , n215654 , n215655 , n215656 , n215657 , n215658 , 
 n215659 , n215660 , n215661 , n215662 , n215663 , n215664 , n215665 , n215666 , n215667 , n215668 , 
 n215669 , n215670 , n215671 , n215672 , n215673 , n215674 , n215675 , n215676 , n215677 , n215678 , 
 n215679 , n215680 , n215681 , n215682 , n215683 , n215684 , n215685 , n215686 , n215687 , n215688 , 
 n215689 , n215690 , n215691 , n215692 , n215693 , n215694 , n215695 , n215696 , n215697 , n215698 , 
 n215699 , n215700 , n215701 , n215702 , n215703 , n215704 , n215705 , n215706 , n215707 , n215708 , 
 n215709 , n215710 , n215711 , n215712 , n215713 , n215714 , n215715 , n215716 , n215717 , n215718 , 
 n215719 , n215720 , n215721 , n215722 , n215723 , n215724 , n215725 , n215726 , n215727 , n215728 , 
 n215729 , n215730 , n215731 , n215732 , n215733 , n215734 , n215735 , n215736 , n215737 , n215738 , 
 n215739 , n215740 , n215741 , n215742 , n215743 , n215744 , n215745 , n215746 , n215747 , n215748 , 
 n215749 , n215750 , n215751 , n215752 , n215753 , n215754 , n215755 , n215756 , n215757 , n215758 , 
 n215759 , n215760 , n215761 , n215762 , n215763 , n215764 , n215765 , n215766 , n215767 , n215768 , 
 n215769 , n215770 , n215771 , n215772 , n215773 , n215774 , n215775 , n215776 , n215777 , n215778 , 
 n215779 , n215780 , n215781 , n215782 , n215783 , n215784 , n215785 , n215786 , n215787 , n215788 , 
 n215789 , n215790 , n215791 , n215792 , n215793 , n215794 , n215795 , n215796 , n215797 , n215798 , 
 n215799 , n215800 , n215801 , n215802 , n215803 , n215804 , n215805 , n215806 , n215807 , n215808 , 
 n215809 , n215810 , n215811 , n215812 , n215813 , n215814 , n215815 , n215816 , n215817 , n215818 , 
 n215819 , n215820 , n215821 , n215822 , n215823 , n215824 , n215825 , n215826 , n215827 , n215828 , 
 n215829 , n215830 , n215831 , n215832 , n215833 , n215834 , n215835 , n215836 , n215837 , n215838 , 
 n215839 , n215840 , n215841 , n215842 , n215843 , n215844 , n215845 , n215846 , n215847 , n215848 , 
 n215849 , n215850 , n215851 , n215852 , n215853 , n215854 , n215855 , n215856 , n215857 , n215858 , 
 n215859 , n215860 , n215861 , n215862 , n215863 , n215864 , n215865 , n215866 , n215867 , n215868 , 
 n215869 , n215870 , n215871 , n215872 , n215873 , n215874 , n215875 , n215876 , n215877 , n215878 , 
 n215879 , n215880 , n215881 , n215882 , n215883 , n215884 , n215885 , n215886 , n215887 , n215888 , 
 n215889 , n215890 , n215891 , n215892 , n215893 , n215894 , n215895 , n215896 , n215897 , n215898 , 
 n215899 , n215900 , n215901 , n215902 , n215903 , n215904 , n215905 , n215906 , n215907 , n215908 , 
 n215909 , n215910 , n215911 , n215912 , n215913 , n215914 , n215915 , n215916 , n215917 , n215918 , 
 n215919 , n215920 , n215921 , n215922 , n215923 , n215924 , n215925 , n215926 , n215927 , n215928 , 
 n215929 , n215930 , n215931 , n215932 , n215933 , n215934 , n215935 , n215936 , n215937 , n215938 , 
 n215939 , n215940 , n215941 , n215942 , n215943 , n215944 , n215945 , n215946 , n215947 , n215948 , 
 n215949 , n215950 , n215951 , n215952 , n215953 , n215954 , n215955 , n215956 , n215957 , n215958 , 
 n215959 , n215960 , n215961 , n215962 , n215963 , n215964 , n215965 , n215966 , n215967 , n215968 , 
 n215969 , n215970 , n215971 , n215972 , n215973 , n215974 , n215975 , n215976 , n215977 , n215978 , 
 n215979 , n215980 , n215981 , n215982 , n215983 , n215984 , n215985 , n215986 , n215987 , n215988 , 
 n215989 , n215990 , n215991 , n215992 , n215993 , n215994 , n215995 , n215996 , n215997 , n215998 , 
 n215999 , n216000 , n216001 , n216002 , n216003 , n216004 , n216005 , n216006 , n216007 , n216008 , 
 n216009 , n216010 , n216011 , n216012 , n216013 , n216014 , n216015 , n216016 , n216017 , n216018 , 
 n216019 , n216020 , n216021 , n216022 , n216023 , n216024 , n216025 , n216026 , n216027 , n216028 , 
 n216029 , n216030 , n216031 , n216032 , n216033 , n216034 , n216035 , n216036 , n216037 , n216038 , 
 n216039 , n216040 , n216041 , n216042 , n216043 , n216044 , n216045 , n216046 , n216047 , n216048 , 
 n216049 , n216050 , n216051 , n216052 , n216053 , n216054 , n216055 , n216056 , n216057 , n216058 , 
 n216059 , n216060 , n216061 , n216062 , n216063 , n216064 , n216065 , n216066 , n216067 , n216068 , 
 n216069 , n216070 , n216071 , n216072 , n216073 , n216074 , n216075 , n216076 , n216077 , n216078 , 
 n216079 , n216080 , n216081 , n216082 , n216083 , n216084 , n216085 , n216086 , n216087 , n216088 , 
 n216089 , n216090 , n216091 , n216092 , n216093 , n216094 , n216095 , n216096 , n216097 , n216098 , 
 n216099 , n216100 , n216101 , n216102 , n216103 , n216104 , n216105 , n216106 , n216107 , n216108 , 
 n216109 , n216110 , n216111 , n216112 , n216113 , n216114 , n216115 , n216116 , n216117 , n216118 , 
 n216119 , n216120 , n216121 , n216122 , n216123 , n216124 , n216125 , n216126 , n216127 , n216128 , 
 n216129 , n216130 , n216131 , n216132 , n216133 , n216134 , n216135 , n216136 , n216137 , n216138 , 
 n216139 , n216140 , n216141 , n216142 , n216143 , n216144 , n216145 , n216146 , n216147 , n216148 , 
 n216149 , n216150 , n216151 , n216152 , n216153 , n216154 , n216155 , n216156 , n216157 , n216158 , 
 n216159 , n216160 , n216161 , n216162 , n216163 , n216164 , n216165 , n216166 , n216167 , n216168 , 
 n216169 , n216170 , n216171 , n216172 , n216173 , n216174 , n216175 , n216176 , n216177 , n216178 , 
 n216179 , n216180 , n216181 , n216182 , n216183 , n216184 , n216185 , n216186 , n216187 , n216188 , 
 n216189 , n216190 , n216191 , n216192 , n216193 , n216194 , n216195 , n216196 , n216197 , n216198 , 
 n216199 , n216200 , n216201 , n216202 , n216203 , n216204 , n216205 , n216206 , n216207 , n216208 , 
 n216209 , n216210 , n216211 , n216212 , n216213 , n216214 , n216215 , n216216 , n216217 , n216218 , 
 n216219 , n216220 , n216221 , n216222 , n216223 , n216224 , n216225 , n216226 , n216227 , n216228 , 
 n216229 , n216230 , n216231 , n216232 , n216233 , n216234 , n216235 , n216236 , n216237 , n216238 , 
 n216239 , n216240 , n216241 , n216242 , n216243 , n216244 , n216245 , n216246 , n216247 , n216248 , 
 n216249 , n216250 , n216251 , n216252 , n216253 , n216254 , n216255 , n216256 , n216257 , n216258 , 
 n216259 , n216260 , n216261 , n216262 , n216263 , n216264 , n216265 , n216266 , n216267 , n216268 , 
 n216269 , n216270 , n216271 , n216272 , n216273 , n216274 , n216275 , n216276 , n216277 , n216278 , 
 n216279 , n216280 , n216281 , n216282 , n216283 , n216284 , n216285 , n216286 , n216287 , n216288 , 
 n216289 , n216290 , n216291 , n216292 , n216293 , n216294 , n216295 , n216296 , n216297 , n216298 , 
 n216299 , n216300 , n216301 , n216302 , n216303 , n216304 , n216305 , n216306 , n216307 , n216308 , 
 n216309 , n216310 , n216311 , n216312 , n216313 , n216314 , n216315 , n216316 , n216317 , n216318 , 
 n216319 , n216320 , n216321 , n216322 , n216323 , n216324 , n216325 , n216326 , n216327 , n216328 , 
 n216329 , n216330 , n216331 , n216332 , n216333 , n216334 , n216335 , n216336 , n216337 , n216338 , 
 n216339 , n216340 , n216341 , n216342 , n216343 , n216344 , n216345 , n216346 , n216347 , n216348 , 
 n216349 , n216350 , n216351 , n216352 , n216353 , n216354 , n216355 , n216356 , n216357 , n216358 , 
 n216359 , n216360 , n216361 , n216362 , n216363 , n216364 , n216365 , n216366 , n216367 , n216368 , 
 n216369 , n216370 , n216371 , n216372 , n216373 , n216374 , n216375 , n216376 , n216377 , n216378 , 
 n216379 , n216380 , n216381 , n216382 , n216383 , n216384 , n216385 , n216386 , n216387 , n216388 , 
 n216389 , n216390 , n216391 , n216392 , n216393 , n216394 , n216395 , n216396 , n216397 , n216398 , 
 n216399 , n216400 , n216401 , n216402 , n216403 , n216404 , n216405 , n216406 , n216407 , n216408 , 
 n216409 , n216410 , n216411 , n216412 , n216413 , n216414 , n216415 , n216416 , n216417 , n216418 , 
 n216419 , n216420 , n216421 , n216422 , n216423 , n216424 , n216425 , n216426 , n216427 , n216428 , 
 n216429 , n216430 , n216431 , n216432 , n216433 , n216434 , n216435 , n216436 , n216437 , n216438 , 
 n216439 , n216440 , n216441 , n216442 , n216443 , n216444 , n216445 , n216446 , n216447 , n216448 , 
 n216449 , n216450 , n216451 , n216452 , n216453 , n216454 , n216455 , n216456 , n216457 , n216458 , 
 n216459 , n216460 , n216461 , n216462 , n216463 , n216464 , n216465 , n216466 , n216467 , n216468 , 
 n216469 , n216470 , n216471 , n216472 , n216473 , n216474 , n216475 , n216476 , n216477 , n216478 , 
 n216479 , n216480 , n216481 , n216482 , n216483 , n216484 , n216485 , n216486 , n216487 , n216488 , 
 n216489 , n216490 , n216491 , n216492 , n216493 , n216494 , n216495 , n216496 , n216497 , n216498 , 
 n216499 , n216500 , n216501 , n216502 , n216503 , n216504 , n216505 , n216506 , n216507 , n216508 , 
 n216509 , n216510 , n216511 , n216512 , n216513 , n216514 , n216515 , n216516 , n216517 , n216518 , 
 n216519 , n216520 , n216521 , n216522 , n216523 , n216524 , n216525 , n216526 , n216527 , n216528 , 
 n216529 , n216530 , n216531 , n216532 , n216533 , n216534 , n216535 , n216536 , n216537 , n216538 , 
 n216539 , n216540 , n216541 , n216542 , n216543 , n216544 , n216545 , n216546 , n216547 , n216548 , 
 n216549 , n216550 , n216551 , n216552 , n216553 , n216554 , n216555 , n216556 , n216557 , n216558 , 
 n216559 , n216560 , n216561 , n216562 , n216563 , n216564 , n216565 , n216566 , n216567 , n216568 , 
 n216569 , n216570 , n216571 , n216572 , n216573 , n216574 , n216575 , n216576 , n216577 , n216578 , 
 n216579 , n216580 , n216581 , n216582 , n216583 , n216584 , n216585 , n216586 , n216587 , n216588 , 
 n216589 , n216590 , n216591 , n216592 , n216593 , n216594 , n216595 , n216596 , n216597 , n216598 , 
 n216599 , n216600 , n216601 , n216602 , n216603 , n216604 , n216605 , n216606 , n216607 , n216608 , 
 n216609 , n216610 , n216611 , n216612 , n216613 , n216614 , n216615 , n216616 , n216617 , n216618 , 
 n216619 , n216620 , n216621 , n216622 , n216623 , n216624 , n216625 , n216626 , n216627 , n216628 , 
 n216629 , n216630 , n216631 , n216632 , n216633 , n216634 , n216635 , n216636 , n216637 , n216638 , 
 n216639 , n216640 , n216641 , n216642 , n216643 , n216644 , n216645 , n216646 , n216647 , n216648 , 
 n216649 , n216650 , n216651 , n216652 , n216653 , n216654 , n216655 , n216656 , n216657 , n216658 , 
 n216659 , n216660 , n216661 , n216662 , n216663 , n216664 , n216665 , n216666 , n216667 , n216668 , 
 n216669 , n216670 , n216671 , n216672 , n216673 , n216674 , n216675 , n216676 , n216677 , n216678 , 
 n216679 , n216680 , n216681 , n216682 , n216683 , n216684 , n216685 , n216686 , n216687 , n216688 , 
 n216689 , n216690 , n216691 , n216692 , n216693 , n216694 , n216695 , n216696 , n216697 , n216698 , 
 n216699 , n216700 , n216701 , n216702 , n216703 , n216704 , n216705 , n216706 , n216707 , n216708 , 
 n216709 , n216710 , n216711 , n216712 , n216713 , n216714 , n216715 , n216716 , n216717 , n216718 , 
 n216719 , n216720 , n216721 , n216722 , n216723 , n216724 , n216725 , n216726 , n216727 , n216728 , 
 n216729 , n216730 , n216731 , n216732 , n216733 , n216734 , n216735 , n216736 , n216737 , n216738 , 
 n216739 , n216740 , n216741 , n216742 , n216743 , n216744 , n216745 , n216746 , n216747 , n216748 , 
 n216749 , n216750 , n216751 , n216752 , n216753 , n216754 , n216755 , n216756 , n216757 , n216758 , 
 n216759 , n216760 , n216761 , n216762 , n216763 , n216764 , n216765 , n216766 , n216767 , n216768 , 
 n216769 , n216770 , n216771 , n216772 , n216773 , n216774 , n216775 , n216776 , n216777 , n216778 , 
 n216779 , n216780 , n216781 , n216782 , n216783 , n216784 , n216785 , n216786 , n216787 , n216788 , 
 n216789 , n216790 , n216791 , n216792 , n216793 , n216794 , n216795 , n216796 , n216797 , n216798 , 
 n216799 , n216800 , n216801 , n216802 , n216803 , n216804 , n216805 , n216806 , n216807 , n216808 , 
 n216809 , n216810 , n216811 , n216812 , n216813 , n216814 , n216815 , n216816 , n216817 , n216818 , 
 n216819 , n216820 , n216821 , n216822 , n216823 , n216824 , n216825 , n216826 , n216827 , n216828 , 
 n216829 , n216830 , n216831 , n216832 , n216833 , n216834 , n216835 , n216836 , n216837 , n216838 , 
 n216839 , n216840 , n216841 , n216842 , n216843 , n216844 , n216845 , n216846 , n216847 , n216848 , 
 n216849 , n216850 , n216851 , n216852 , n216853 , n216854 , n216855 , n216856 , n216857 , n216858 , 
 n216859 , n216860 , n216861 , n216862 , n216863 , n216864 , n216865 , n216866 , n216867 , n216868 , 
 n216869 , n216870 , n216871 , n216872 , n216873 , n216874 , n216875 , n216876 , n216877 , n216878 , 
 n216879 , n216880 , n216881 , n216882 , n216883 , n216884 , n216885 , n216886 , n216887 , n216888 , 
 n216889 , n216890 , n216891 , n216892 , n216893 , n216894 , n216895 , n216896 , n216897 , n216898 , 
 n216899 , n216900 , n216901 , n216902 , n216903 , n216904 , n216905 , n216906 , n216907 , n216908 , 
 n216909 , n216910 , n216911 , n216912 , n216913 , n216914 , n216915 , n216916 , n216917 , n216918 , 
 n216919 , n216920 , n216921 , n216922 , n216923 , n216924 , n216925 , n216926 , n216927 , n216928 , 
 n216929 , n216930 , n216931 , n216932 , n216933 , n216934 , n216935 , n216936 , n216937 , n216938 , 
 n216939 , n216940 , n216941 , n216942 , n216943 , n216944 , n216945 , n216946 , n216947 , n216948 , 
 n216949 , n216950 , n216951 , n216952 , n216953 , n216954 , n216955 , n216956 , n216957 , n216958 , 
 n216959 , n216960 , n216961 , n216962 , n216963 , n216964 , n216965 , n216966 , n216967 , n216968 , 
 n216969 , n216970 , n216971 , n216972 , n216973 , n216974 , n216975 , n216976 , n216977 , n216978 , 
 n216979 , n216980 , n216981 , n216982 , n216983 , n216984 , n216985 , n216986 , n216987 , n216988 , 
 n216989 , n216990 , n216991 , n216992 , n216993 , n216994 , n216995 , n216996 , n216997 , n216998 , 
 n216999 , n217000 , n217001 , n217002 , n217003 , n217004 , n217005 , n217006 , n217007 , n217008 , 
 n217009 , n217010 , n217011 , n217012 , n217013 , n217014 , n217015 , n217016 , n217017 , n217018 , 
 n217019 , n217020 , n217021 , n217022 , n217023 , n217024 , n217025 , n217026 , n217027 , n217028 , 
 n217029 , n217030 , n217031 , n217032 , n217033 , n217034 , n217035 , n217036 , n217037 , n217038 , 
 n217039 , n217040 , n217041 , n217042 , n217043 , n217044 , n217045 , n217046 , n217047 , n217048 , 
 n217049 , n217050 , n217051 , n217052 , n217053 , n217054 , n217055 , n217056 , n217057 , n217058 , 
 n217059 , n217060 , n217061 , n217062 , n217063 , n217064 , n217065 , n217066 , n217067 , n217068 , 
 n217069 , n217070 , n217071 , n217072 , n217073 , n217074 , n217075 , n217076 , n217077 , n217078 , 
 n217079 , n217080 , n217081 , n217082 , n217083 , n217084 , n217085 , n217086 , n217087 , n217088 , 
 n217089 , n217090 , n217091 , n217092 , n217093 , n217094 , n217095 , n217096 , n217097 , n217098 , 
 n217099 , n217100 , n217101 , n217102 , n217103 , n217104 , n217105 , n217106 , n217107 , n217108 , 
 n217109 , n217110 , n217111 , n217112 , n217113 , n217114 , n217115 , n217116 , n217117 , n217118 , 
 n217119 , n217120 , n217121 , n217122 , n217123 , n217124 , n217125 , n217126 , n217127 , n217128 , 
 n217129 , n217130 , n217131 , n217132 , n217133 , n217134 , n217135 , n217136 , n217137 , n217138 , 
 n217139 , n217140 , n217141 , n217142 , n217143 , n217144 , n217145 , n217146 , n217147 , n217148 , 
 n217149 , n217150 , n217151 , n217152 , n217153 , n217154 , n217155 , n217156 , n217157 , n217158 , 
 n217159 , n217160 , n217161 , n217162 , n217163 , n217164 , n217165 , n217166 , n217167 , n217168 , 
 n217169 , n217170 , n217171 , n217172 , n217173 , n217174 , n217175 , n217176 , n217177 , n217178 , 
 n217179 , n217180 , n217181 , n217182 , n217183 , n217184 , n217185 , n217186 , n217187 , n217188 , 
 n217189 , n217190 , n217191 , n217192 , n217193 , n217194 , n217195 , n217196 , n217197 , n217198 , 
 n217199 , n217200 , n217201 , n217202 , n217203 , n217204 , n217205 , n217206 , n217207 , n217208 , 
 n217209 , n217210 , n217211 , n217212 , n217213 , n217214 , n217215 , n217216 , n217217 , n217218 , 
 n217219 , n217220 , n217221 , n217222 , n217223 , n217224 , n217225 , n217226 , n217227 , n217228 , 
 n217229 , n217230 , n217231 , n217232 , n217233 , n217234 , n217235 , n217236 , n217237 , n217238 , 
 n217239 , n217240 , n217241 , n217242 , n217243 , n217244 , n217245 , n217246 , n217247 , n217248 , 
 n217249 , n217250 , n217251 , n217252 , n217253 , n217254 , n217255 , n217256 , n217257 , n217258 , 
 n217259 , n217260 , n217261 , n217262 , n217263 , n217264 , n217265 , n217266 , n217267 , n217268 , 
 n217269 , n217270 , n217271 , n217272 , n217273 , n217274 , n217275 , n217276 , n217277 , n217278 , 
 n217279 , n217280 , n217281 , n217282 , n217283 , n217284 , n217285 , n217286 , n217287 , n217288 , 
 n217289 , n217290 , n217291 , n217292 , n217293 , n217294 , n217295 , n217296 , n217297 , n217298 , 
 n217299 , n217300 , n217301 , n217302 , n217303 , n217304 , n217305 , n217306 , n217307 , n217308 , 
 n217309 , n217310 , n217311 , n217312 , n217313 , n217314 , n217315 , n217316 , n217317 , n217318 , 
 n217319 , n217320 , n217321 , n217322 , n217323 , n217324 , n217325 , n217326 , n217327 , n217328 , 
 n217329 , n217330 , n217331 , n217332 , n217333 , n217334 , n217335 , n217336 , n217337 , n217338 , 
 n217339 , n217340 , n217341 , n217342 , n217343 , n217344 , n217345 , n217346 , n217347 , n217348 , 
 n217349 , n217350 , n217351 , n217352 , n217353 , n217354 , n217355 , n217356 , n217357 , n217358 , 
 n217359 , n217360 , n217361 , n217362 , n217363 , n217364 , n217365 , n217366 , n217367 , n217368 , 
 n217369 , n217370 , n217371 , n217372 , n217373 , n217374 , n217375 , n217376 , n217377 , n217378 , 
 n217379 , n217380 , n217381 , n217382 , n217383 , n217384 , n217385 , n217386 , n217387 , n217388 , 
 n217389 , n217390 , n217391 , n217392 , n217393 , n217394 , n217395 , n217396 , n217397 , n217398 , 
 n217399 , n217400 , n217401 , n217402 , n217403 , n217404 , n217405 , n217406 , n217407 , n217408 , 
 n217409 , n217410 , n217411 , n217412 , n217413 , n217414 , n217415 , n217416 , n217417 , n217418 , 
 n217419 , n217420 , n217421 , n217422 , n217423 , n217424 , n217425 , n217426 , n217427 , n217428 , 
 n217429 , n217430 , n217431 , n217432 , n217433 , n217434 , n217435 , n217436 , n217437 , n217438 , 
 n217439 , n217440 , n217441 , n217442 , n217443 , n217444 , n217445 , n217446 , n217447 , n217448 , 
 n217449 , n217450 , n217451 , n217452 , n217453 , n217454 , n217455 , n217456 , n217457 , n217458 , 
 n217459 , n217460 , n217461 , n217462 , n217463 , n217464 , n217465 , n217466 , n217467 , n217468 , 
 n217469 , n217470 , n217471 , n217472 , n217473 , n217474 , n217475 , n217476 , n217477 , n217478 , 
 n217479 , n217480 , n217481 , n217482 , n217483 , n217484 , n217485 , n217486 , n217487 , n217488 , 
 n217489 , n217490 , n217491 , n217492 , n217493 , n217494 , n217495 , n217496 , n217497 , n217498 , 
 n217499 , n217500 , n217501 , n217502 , n217503 , n217504 , n217505 , n217506 , n217507 , n217508 , 
 n217509 , n217510 , n217511 , n217512 , n217513 , n217514 , n217515 , n217516 , n217517 , n217518 , 
 n217519 , n217520 , n217521 , n217522 , n217523 , n217524 , n217525 , n217526 , n217527 , n217528 , 
 n217529 , n217530 , n217531 , n217532 , n217533 , n217534 , n217535 , n217536 , n217537 , n217538 , 
 n217539 , n217540 , n217541 , n217542 , n217543 , n217544 , n217545 , n217546 , n217547 , n217548 , 
 n217549 , n217550 , n217551 , n217552 , n217553 , n217554 , n217555 , n217556 , n217557 , n217558 , 
 n217559 , n217560 , n217561 , n217562 , n217563 , n217564 , n217565 , n217566 , n217567 , n217568 , 
 n217569 , n217570 , n217571 , n217572 , n217573 , n217574 , n217575 , n217576 , n217577 , n217578 , 
 n217579 , n217580 , n217581 , n217582 , n217583 , n217584 , n217585 , n217586 , n217587 , n217588 , 
 n217589 , n217590 , n217591 , n217592 , n217593 , n217594 , n217595 , n217596 , n217597 , n217598 , 
 n217599 , n217600 , n217601 , n217602 , n217603 , n217604 , n217605 , n217606 , n217607 , n217608 , 
 n217609 , n217610 , n217611 , n217612 , n217613 , n217614 , n217615 , n217616 , n217617 , n217618 , 
 n217619 , n217620 , n217621 , n217622 , n217623 , n217624 , n217625 , n217626 , n217627 , n217628 , 
 n217629 , n217630 , n217631 , n217632 , n217633 , n217634 , n217635 , n217636 , n217637 , n217638 , 
 n217639 , n217640 , n217641 , n217642 , n217643 , n217644 , n217645 , n217646 , n217647 , n217648 , 
 n217649 , n217650 , n217651 , n217652 , n217653 , n217654 , n217655 , n217656 , n217657 , n217658 , 
 n217659 , n217660 , n217661 , n217662 , n217663 , n217664 , n217665 , n217666 , n217667 , n217668 , 
 n217669 , n217670 , n217671 , n217672 , n217673 , n217674 , n217675 , n217676 , n217677 , n217678 , 
 n217679 , n217680 , n217681 , n217682 , n217683 , n217684 , n217685 , n217686 , n217687 , n217688 , 
 n217689 , n217690 , n217691 , n217692 , n217693 , n217694 , n217695 , n217696 , n217697 , n217698 , 
 n217699 , n217700 , n217701 , n217702 , n217703 , n217704 , n217705 , n217706 , n217707 , n217708 , 
 n217709 , n217710 , n217711 , n217712 , n217713 , n217714 , n217715 , n217716 , n217717 , n217718 , 
 n217719 , n217720 , n217721 , n217722 , n217723 , n217724 , n217725 , n217726 , n217727 , n217728 , 
 n217729 , n217730 , n217731 , n217732 , n217733 , n217734 , n217735 , n217736 , n217737 , n217738 , 
 n217739 , n217740 , n217741 , n217742 , n217743 , n217744 , n217745 , n217746 , n217747 , n217748 , 
 n217749 , n217750 , n217751 , n217752 , n217753 , n217754 , n217755 , n217756 , n217757 , n217758 , 
 n217759 , n217760 , n217761 , n217762 , n217763 , n217764 , n217765 , n217766 , n217767 , n217768 , 
 n217769 , n217770 , n217771 , n217772 , n217773 , n217774 , n217775 , n217776 , n217777 , n217778 , 
 n217779 , n217780 , n217781 , n217782 , n217783 , n217784 , n217785 , n217786 , n217787 , n217788 , 
 n217789 , n217790 , n217791 , n217792 , n217793 , n217794 , n217795 , n217796 , n217797 , n217798 , 
 n217799 , n217800 , n217801 , n217802 , n217803 , n217804 , n217805 , n217806 , n217807 , n217808 , 
 n217809 , n217810 , n217811 , n217812 , n217813 , n217814 , n217815 , n217816 , n217817 , n217818 , 
 n217819 , n217820 , n217821 , n217822 , n217823 , n217824 , n217825 , n217826 , n217827 , n217828 , 
 n217829 , n217830 , n217831 , n217832 , n217833 , n217834 , n217835 , n217836 , n217837 , n217838 , 
 n217839 , n217840 , n217841 , n217842 , n217843 , n217844 , n217845 , n217846 , n217847 , n217848 , 
 n217849 , n217850 , n217851 , n217852 , n217853 , n217854 , n217855 , n217856 , n217857 , n217858 , 
 n217859 , n217860 , n217861 , n217862 , n217863 , n217864 , n217865 , n217866 , n217867 , n217868 , 
 n217869 , n217870 , n217871 , n217872 , n217873 , n217874 , n217875 , n217876 , n217877 , n217878 , 
 n217879 , n217880 , n217881 , n217882 , n217883 , n217884 , n217885 , n217886 , n217887 , n217888 , 
 n217889 , n217890 , n217891 , n217892 , n217893 , n217894 , n217895 , n217896 , n217897 , n217898 , 
 n217899 , n217900 , n217901 , n217902 , n217903 , n217904 , n217905 , n217906 , n217907 , n217908 , 
 n217909 , n217910 , n217911 , n217912 , n217913 , n217914 , n217915 , n217916 , n217917 , n217918 , 
 n217919 , n217920 , n217921 , n217922 , n217923 , n217924 , n217925 , n217926 , n217927 , n217928 , 
 n217929 , n217930 , n217931 , n217932 , n217933 , n217934 , n217935 , n217936 , n217937 , n217938 , 
 n217939 , n217940 , n217941 , n217942 , n217943 , n217944 , n217945 , n217946 , n217947 , n217948 , 
 n217949 , n217950 , n217951 , n217952 , n217953 , n217954 , n217955 , n217956 , n217957 , n217958 , 
 n217959 , n217960 , n217961 , n217962 , n217963 , n217964 , n217965 , n217966 , n217967 , n217968 , 
 n217969 , n217970 , n217971 , n217972 , n217973 , n217974 , n217975 , n217976 , n217977 , n217978 , 
 n217979 , n217980 , n217981 , n217982 , n217983 , n217984 , n217985 , n217986 , n217987 , n217988 , 
 n217989 , n217990 , n217991 , n217992 , n217993 , n217994 , n217995 , n217996 , n217997 , n217998 , 
 n217999 , n218000 , n218001 , n218002 , n218003 , n218004 , n218005 , n218006 , n218007 , n218008 , 
 n218009 , n218010 , n218011 , n218012 , n218013 , n218014 , n218015 , n218016 , n218017 , n218018 , 
 n218019 , n218020 , n218021 , n218022 , n218023 , n218024 , n218025 , n218026 , n218027 , n218028 , 
 n218029 , n218030 , n218031 , n218032 , n218033 , n218034 , n218035 , n218036 , n218037 , n218038 , 
 n218039 , n218040 , n218041 , n218042 , n218043 , n218044 , n218045 , n218046 , n218047 , n218048 , 
 n218049 , n218050 , n218051 , n218052 , n218053 , n218054 , n218055 , n218056 , n218057 , n218058 , 
 n218059 , n218060 , n218061 , n218062 , n218063 , n218064 , n218065 , n218066 , n218067 , n218068 , 
 n218069 , n218070 , n218071 , n218072 , n218073 , n218074 , n218075 , n218076 , n218077 , n218078 , 
 n218079 , n218080 , n218081 , n218082 , n218083 , n218084 , n218085 , n218086 , n218087 , n218088 , 
 n218089 , n218090 , n218091 , n218092 , n218093 , n218094 , n218095 , n218096 , n218097 , n218098 , 
 n218099 , n218100 , n218101 , n218102 , n218103 , n218104 , n218105 , n218106 , n218107 , n218108 , 
 n218109 , n218110 , n218111 , n218112 , n218113 , n218114 , n218115 , n218116 , n218117 , n218118 , 
 n218119 , n218120 , n218121 , n218122 , n218123 , n218124 , n218125 , n218126 , n218127 , n218128 , 
 n218129 , n218130 , n218131 , n218132 , n218133 , n218134 , n218135 , n218136 , n218137 , n218138 , 
 n218139 , n218140 , n218141 , n218142 , n218143 , n218144 , n218145 , n218146 , n218147 , n218148 , 
 n218149 , n218150 , n218151 , n218152 , n218153 , n218154 , n218155 , n218156 , n218157 , n218158 , 
 n218159 , n218160 , n218161 , n218162 , n218163 , n218164 , n218165 , n218166 , n218167 , n218168 , 
 n218169 , n218170 , n218171 , n218172 , n218173 , n218174 , n218175 , n218176 , n218177 , n218178 , 
 n218179 , n218180 , n218181 , n218182 , n218183 , n218184 , n218185 , n218186 , n218187 , n218188 , 
 n218189 , n218190 , n218191 , n218192 , n218193 , n218194 , n218195 , n218196 , n218197 , n218198 , 
 n218199 , n218200 , n218201 , n218202 , n218203 , n218204 , n218205 , n218206 , n218207 , n218208 , 
 n218209 , n218210 , n218211 , n218212 , n218213 , n218214 , n218215 , n218216 , n218217 , n218218 , 
 n218219 , n218220 , n218221 , n218222 , n218223 , n218224 , n218225 , n218226 , n218227 , n218228 , 
 n218229 , n218230 , n218231 , n218232 , n218233 , n218234 , n218235 , n218236 , n218237 , n218238 , 
 n218239 , n218240 , n218241 , n218242 , n218243 , n218244 , n218245 , n218246 , n218247 , n218248 , 
 n218249 , n218250 , n218251 , n218252 , n218253 , n218254 , n218255 , n218256 , n218257 , n218258 , 
 n218259 , n218260 , n218261 , n218262 , n218263 , n218264 , n218265 , n218266 , n218267 , n218268 , 
 n218269 , n218270 , n218271 , n218272 , n218273 , n218274 , n218275 , n218276 , n218277 , n218278 , 
 n218279 , n218280 , n218281 , n218282 , n218283 , n218284 , n218285 , n218286 , n218287 , n218288 , 
 n218289 , n218290 , n218291 , n218292 , n218293 , n218294 , n218295 , n218296 , n218297 , n218298 , 
 n218299 , n218300 , n218301 , n218302 , n218303 , n218304 , n218305 , n218306 , n218307 , n218308 , 
 n218309 , n218310 , n218311 , n218312 , n218313 , n218314 , n218315 , n218316 , n218317 , n218318 , 
 n218319 , n218320 , n218321 , n218322 , n218323 , n218324 , n218325 , n218326 , n218327 , n218328 , 
 n218329 , n218330 , n218331 , n218332 , n218333 , n218334 , n218335 , n218336 , n218337 , n218338 , 
 n218339 , n218340 , n218341 , n218342 , n218343 , n218344 , n218345 , n218346 , n218347 , n218348 , 
 n218349 , n218350 , n218351 , n218352 , n218353 , n218354 , n218355 , n218356 , n218357 , n218358 , 
 n218359 , n218360 , n218361 , n218362 , n218363 , n218364 , n218365 , n218366 , n218367 , n218368 , 
 n218369 , n218370 , n218371 , n218372 , n218373 , n218374 , n218375 , n218376 , n218377 , n218378 , 
 n218379 , n218380 , n218381 , n218382 , n218383 , n218384 , n218385 , n218386 , n218387 , n218388 , 
 n218389 , n218390 , n218391 , n218392 , n218393 , n218394 , n218395 , n218396 , n218397 , n218398 , 
 n218399 , n218400 , n218401 , n218402 , n218403 , n218404 , n218405 , n218406 , n218407 , n218408 , 
 n218409 , n218410 , n218411 , n218412 , n218413 , n218414 , n218415 , n218416 , n218417 , n218418 , 
 n218419 , n218420 , n218421 , n218422 , n218423 , n218424 , n218425 , n218426 , n218427 , n218428 , 
 n218429 , n218430 , n218431 , n218432 , n218433 , n218434 , n218435 , n218436 , n218437 , n218438 , 
 n218439 , n218440 , n218441 , n218442 , n218443 , n218444 , n218445 , n218446 , n218447 , n218448 , 
 n218449 , n218450 , n218451 , n218452 , n218453 , n218454 , n218455 , n218456 , n218457 , n218458 , 
 n218459 , n218460 , n218461 , n218462 , n218463 , n218464 , n218465 , n218466 , n218467 , n218468 , 
 n218469 , n218470 , n218471 , n218472 , n218473 , n218474 , n218475 , n218476 , n218477 , n218478 , 
 n218479 , n218480 , n218481 , n218482 , n218483 , n218484 , n218485 , n218486 , n218487 , n218488 , 
 n218489 , n218490 , n218491 , n218492 , n218493 , n218494 , n218495 , n218496 , n218497 , n218498 , 
 n218499 , n218500 , n218501 , n218502 , n218503 , n218504 , n218505 , n218506 , n218507 , n218508 , 
 n218509 , n218510 , n218511 , n218512 , n218513 , n218514 , n218515 , n218516 , n218517 , n218518 , 
 n218519 , n218520 , n218521 , n218522 , n218523 , n218524 , n218525 , n218526 , n218527 , n218528 , 
 n218529 , n218530 , n218531 , n218532 , n218533 , n218534 , n218535 , n218536 , n218537 , n218538 , 
 n218539 , n218540 , n218541 , n218542 , n218543 , n218544 , n218545 , n218546 , n218547 , n218548 , 
 n218549 , n218550 , n218551 , n218552 , n218553 , n218554 , n218555 , n218556 , n218557 , n218558 , 
 n218559 , n218560 , n218561 , n218562 , n218563 , n218564 , n218565 , n218566 , n218567 , n218568 , 
 n218569 , n218570 , n218571 , n218572 , n218573 , n218574 , n218575 , n218576 , n218577 , n218578 , 
 n218579 , n218580 , n218581 , n218582 , n218583 , n218584 , n218585 , n218586 , n218587 , n218588 , 
 n218589 , n218590 , n218591 , n218592 , n218593 , n218594 , n218595 , n218596 , n218597 , n218598 , 
 n218599 , n218600 , n218601 , n218602 , n218603 , n218604 , n218605 , n218606 , n218607 , n218608 , 
 n218609 , n218610 , n218611 , n218612 , n218613 , n218614 , n218615 , n218616 , n218617 , n218618 , 
 n218619 , n218620 , n218621 , n218622 , n218623 , n218624 , n218625 , n218626 , n218627 , n218628 , 
 n218629 , n218630 , n218631 , n218632 , n218633 , n218634 , n218635 , n218636 , n218637 , n218638 , 
 n218639 , n218640 , n218641 , n218642 , n218643 , n218644 , n218645 , n218646 , n218647 , n218648 , 
 n218649 , n218650 , n218651 , n218652 , n218653 , n218654 , n218655 , n218656 , n218657 , n218658 , 
 n218659 , n218660 , n218661 , n218662 , n218663 , n218664 , n218665 , n218666 , n218667 , n218668 , 
 n218669 , n218670 , n218671 , n218672 , n218673 , n218674 , n218675 , n218676 , n218677 , n218678 , 
 n218679 , n218680 , n218681 , n218682 , n218683 , n218684 , n218685 , n218686 , n218687 , n218688 , 
 n218689 , n218690 , n218691 , n218692 , n218693 , n218694 , n218695 , n218696 , n218697 , n218698 , 
 n218699 , n218700 , n218701 , n218702 , n218703 , n218704 , n218705 , n218706 , n218707 , n218708 , 
 n218709 , n218710 , n218711 , n218712 , n218713 , n218714 , n218715 , n218716 , n218717 , n218718 , 
 n218719 , n218720 , n218721 , n218722 , n218723 , n218724 , n218725 , n218726 , n218727 , n218728 , 
 n218729 , n218730 , n218731 , n218732 , n218733 , n218734 , n218735 , n218736 , n218737 , n218738 , 
 n218739 , n218740 , n218741 , n218742 , n218743 , n218744 , n218745 , n218746 , n218747 , n218748 , 
 n218749 , n218750 , n218751 , n218752 , n218753 , n218754 , n218755 , n218756 , n218757 , n218758 , 
 n218759 , n218760 , n218761 , n218762 , n218763 , n218764 , n218765 , n218766 , n218767 , n218768 , 
 n218769 , n218770 , n218771 , n218772 , n218773 , n218774 , n218775 , n218776 , n218777 , n218778 , 
 n218779 , n218780 , n218781 , n218782 , n218783 , n218784 , n218785 , n218786 , n218787 , n218788 , 
 n218789 , n218790 , n218791 , n218792 , n218793 , n218794 , n218795 , n218796 , n218797 , n218798 , 
 n218799 , n218800 , n218801 , n218802 , n218803 , n218804 , n218805 , n218806 , n218807 , n218808 , 
 n218809 , n218810 , n218811 , n218812 , n218813 , n218814 , n218815 , n218816 , n218817 , n218818 , 
 n218819 , n218820 , n218821 , n218822 , n218823 , n218824 , n218825 , n218826 , n218827 , n218828 , 
 n218829 , n218830 , n218831 , n218832 , n218833 , n218834 , n218835 , n218836 , n218837 , n218838 , 
 n218839 , n218840 , n218841 , n218842 , n218843 , n218844 , n218845 , n218846 , n218847 , n218848 , 
 n218849 , n218850 , n218851 , n218852 , n218853 , n218854 , n218855 , n218856 , n218857 , n218858 , 
 n218859 , n218860 , n218861 , n218862 , n218863 , n218864 , n218865 , n218866 , n218867 , n218868 , 
 n218869 , n218870 , n218871 , n218872 , n218873 , n218874 , n218875 , n218876 , n218877 , n218878 , 
 n218879 , n218880 , n218881 , n218882 , n218883 , n218884 , n218885 , n218886 , n218887 , n218888 , 
 n218889 , n218890 , n218891 , n218892 , n218893 , n218894 , n218895 , n218896 , n218897 , n218898 , 
 n218899 , n218900 , n218901 , n218902 , n218903 , n218904 , n218905 , n218906 , n218907 , n218908 , 
 n218909 , n218910 , n218911 , n218912 , n218913 , n218914 , n218915 , n218916 , n218917 , n218918 , 
 n218919 , n218920 , n218921 , n218922 , n218923 , n218924 , n218925 , n218926 , n218927 , n218928 , 
 n218929 , n218930 , n218931 , n218932 , n218933 , n218934 , n218935 , n218936 , n218937 , n218938 , 
 n218939 , n218940 , n218941 , n218942 , n218943 , n218944 , n218945 , n218946 , n218947 , n218948 , 
 n218949 , n218950 , n218951 , n218952 , n218953 , n218954 , n218955 , n218956 , n218957 , n218958 , 
 n218959 , n218960 , n218961 , n218962 , n218963 , n218964 , n218965 , n218966 , n218967 , n218968 , 
 n218969 , n218970 , n218971 , n218972 , n218973 , n218974 , n218975 , n218976 , n218977 , n218978 , 
 n218979 , n218980 , n218981 , n218982 , n218983 , n218984 , n218985 , n218986 , n218987 , n218988 , 
 n218989 , n218990 , n218991 , n218992 , n218993 , n218994 , n218995 , n218996 , n218997 , n218998 , 
 n218999 , n219000 , n219001 , n219002 , n219003 , n219004 , n219005 , n219006 , n219007 , n219008 , 
 n219009 , n219010 , n219011 , n219012 , n219013 , n219014 , n219015 , n219016 , n219017 , n219018 , 
 n219019 , n219020 , n219021 , n219022 , n219023 , n219024 , n219025 , n219026 , n219027 , n219028 , 
 n219029 , n219030 , n219031 , n219032 , n219033 , n219034 , n219035 , n219036 , n219037 , n219038 , 
 n219039 , n219040 , n219041 , n219042 , n219043 , n219044 , n219045 , n219046 , n219047 , n219048 , 
 n219049 , n219050 , n219051 , n219052 , n219053 , n219054 , n219055 , n219056 , n219057 , n219058 , 
 n219059 , n219060 , n219061 , n219062 , n219063 , n219064 , n219065 , n219066 , n219067 , n219068 , 
 n219069 , n219070 , n219071 , n219072 , n219073 , n219074 , n219075 , n219076 , n219077 , n219078 , 
 n219079 , n219080 , n219081 , n219082 , n219083 , n219084 , n219085 , n219086 , n219087 , n219088 , 
 n219089 , n219090 , n219091 , n219092 , n219093 , n219094 , n219095 , n219096 , n219097 , n219098 , 
 n219099 , n219100 , n219101 , n219102 , n219103 , n219104 , n219105 , n219106 , n219107 , n219108 , 
 n219109 , n219110 , n219111 , n219112 , n219113 , n219114 , n219115 , n219116 , n219117 , n219118 , 
 n219119 , n219120 , n219121 , n219122 , n219123 , n219124 , n219125 , n219126 , n219127 , n219128 , 
 n219129 , n219130 , n219131 , n219132 , n219133 , n219134 , n219135 , n219136 , n219137 , n219138 , 
 n219139 , n219140 , n219141 , n219142 , n219143 , n219144 , n219145 , n219146 , n219147 , n219148 , 
 n219149 , n219150 , n219151 , n219152 , n219153 , n219154 , n219155 , n219156 , n219157 , n219158 , 
 n219159 , n219160 , n219161 , n219162 , n219163 , n219164 , n219165 , n219166 , n219167 , n219168 , 
 n219169 , n219170 , n219171 , n219172 , n219173 , n219174 , n219175 , n219176 , n219177 , n219178 , 
 n219179 , n219180 , n219181 , n219182 , n219183 , n219184 , n219185 , n219186 , n219187 , n219188 , 
 n219189 , n219190 , n219191 , n219192 , n219193 , n219194 , n219195 , n219196 , n219197 , n219198 , 
 n219199 , n219200 , n219201 , n219202 , n219203 , n219204 , n219205 , n219206 , n219207 , n219208 , 
 n219209 , n219210 , n219211 , n219212 , n219213 , n219214 , n219215 , n219216 , n219217 , n219218 , 
 n219219 , n219220 , n219221 , n219222 , n219223 , n219224 , n219225 , n219226 , n219227 , n219228 , 
 n219229 , n219230 , n219231 , n219232 , n219233 , n219234 , n219235 , n219236 , n219237 , n219238 , 
 n219239 , n219240 , n219241 , n219242 , n219243 , n219244 , n219245 , n219246 , n219247 , n219248 , 
 n219249 , n219250 , n219251 , n219252 , n219253 , n219254 , n219255 , n219256 , n219257 , n219258 , 
 n219259 , n219260 , n219261 , n219262 , n219263 , n219264 , n219265 , n219266 , n219267 , n219268 , 
 n219269 , n219270 , n219271 , n219272 , n219273 , n219274 , n219275 , n219276 , n219277 , n219278 , 
 n219279 , n219280 , n219281 , n219282 , n219283 , n219284 , n219285 , n219286 , n219287 , n219288 , 
 n219289 , n219290 , n219291 , n219292 , n219293 , n219294 , n219295 , n219296 , n219297 , n219298 , 
 n219299 , n219300 , n219301 , n219302 , n219303 , n219304 , n219305 , n219306 , n219307 , n219308 , 
 n219309 , n219310 , n219311 , n219312 , n219313 , n219314 , n219315 , n219316 , n219317 , n219318 , 
 n219319 , n219320 , n219321 , n219322 , n219323 , n219324 , n219325 , n219326 , n219327 , n219328 , 
 n219329 , n219330 , n219331 , n219332 , n219333 , n219334 , n219335 , n219336 , n219337 , n219338 , 
 n219339 , n219340 , n219341 , n219342 , n219343 , n219344 , n219345 , n219346 , n219347 , n219348 , 
 n219349 , n219350 , n219351 , n219352 , n219353 , n219354 , n219355 , n219356 , n219357 , n219358 , 
 n219359 , n219360 , n219361 , n219362 , n219363 , n219364 , n219365 , n219366 , n219367 , n219368 , 
 n219369 , n219370 , n219371 , n219372 , n219373 , n219374 , n219375 , n219376 , n219377 , n219378 , 
 n219379 , n219380 , n219381 , n219382 , n219383 , n219384 , n219385 , n219386 , n219387 , n219388 , 
 n219389 , n219390 , n219391 , n219392 , n219393 , n219394 , n219395 , n219396 , n219397 , n219398 , 
 n219399 , n219400 , n219401 , n219402 , n219403 , n219404 , n219405 , n219406 , n219407 , n219408 , 
 n219409 , n219410 , n219411 , n219412 , n219413 , n219414 , n219415 , n219416 , n219417 , n219418 , 
 n219419 , n219420 , n219421 , n219422 , n219423 , n219424 , n219425 , n219426 , n219427 , n219428 , 
 n219429 , n219430 , n219431 , n219432 , n219433 , n219434 , n219435 , n219436 , n219437 , n219438 , 
 n219439 , n219440 , n219441 , n219442 , n219443 , n219444 , n219445 , n219446 , n219447 , n219448 , 
 n219449 , n219450 , n219451 , n219452 , n219453 , n219454 , n219455 , n219456 , n219457 , n219458 , 
 n219459 , n219460 , n219461 , n219462 , n219463 , n219464 , n219465 , n219466 , n219467 , n219468 , 
 n219469 , n219470 , n219471 , n219472 , n219473 , n219474 , n219475 , n219476 , n219477 , n219478 , 
 n219479 , n219480 , n219481 , n219482 , n219483 , n219484 , n219485 , n219486 , n219487 , n219488 , 
 n219489 , n219490 , n219491 , n219492 , n219493 , n219494 , n219495 , n219496 , n219497 , n219498 , 
 n219499 , n219500 , n219501 , n219502 , n219503 , n219504 , n219505 , n219506 , n219507 , n219508 , 
 n219509 , n219510 , n219511 , n219512 , n219513 , n219514 , n219515 , n219516 , n219517 , n219518 , 
 n219519 , n219520 , n219521 , n219522 , n219523 , n219524 , n219525 , n219526 , n219527 , n219528 , 
 n219529 , n219530 , n219531 , n219532 , n219533 , n219534 , n219535 , n219536 , n219537 , n219538 , 
 n219539 , n219540 , n219541 , n219542 , n219543 , n219544 , n219545 , n219546 , n219547 , n219548 , 
 n219549 , n219550 , n219551 , n219552 , n219553 , n219554 , n219555 , n219556 , n219557 , n219558 , 
 n219559 , n219560 , n219561 , n219562 , n219563 , n219564 , n219565 , n219566 , n219567 , n219568 , 
 n219569 , n219570 , n219571 , n219572 , n219573 , n219574 , n219575 , n219576 , n219577 , n219578 , 
 n219579 , n219580 , n219581 , n219582 , n219583 , n219584 , n219585 , n219586 , n219587 , n219588 , 
 n219589 , n219590 , n219591 , n219592 , n219593 , n219594 , n219595 , n219596 , n219597 , n219598 , 
 n219599 , n219600 , n219601 , n219602 , n219603 , n219604 , n219605 , n219606 , n219607 , n219608 , 
 n219609 , n219610 , n219611 , n219612 , n219613 , n219614 , n219615 , n219616 , n219617 , n219618 , 
 n219619 , n219620 , n219621 , n219622 , n219623 , n219624 , n219625 , n219626 , n219627 , n219628 , 
 n219629 , n219630 , n219631 , n219632 , n219633 , n219634 , n219635 , n219636 , n219637 , n219638 , 
 n219639 , n219640 , n219641 , n219642 , n219643 , n219644 , n219645 , n219646 , n219647 , n219648 , 
 n219649 , n219650 , n219651 , n219652 , n219653 , n219654 , n219655 , n219656 , n219657 , n219658 , 
 n219659 , n219660 , n219661 , n219662 , n219663 , n219664 , n219665 , n219666 , n219667 , n219668 , 
 n219669 , n219670 , n219671 , n219672 , n219673 , n219674 , n219675 , n219676 , n219677 , n219678 , 
 n219679 , n219680 , n219681 , n219682 , n219683 , n219684 , n219685 , n219686 , n219687 , n219688 , 
 n219689 , n219690 , n219691 , n219692 , n219693 , n219694 , n219695 , n219696 , n219697 , n219698 , 
 n219699 , n219700 , n219701 , n219702 , n219703 , n219704 , n219705 , n219706 , n219707 , n219708 , 
 n219709 , n219710 , n219711 , n219712 , n219713 , n219714 , n219715 , n219716 , n219717 , n219718 , 
 n219719 , n219720 , n219721 , n219722 , n219723 , n219724 , n219725 , n219726 , n219727 , n219728 , 
 n219729 , n219730 , n219731 , n219732 , n219733 , n219734 , n219735 , n219736 , n219737 , n219738 , 
 n219739 , n219740 , n219741 , n219742 , n219743 , n219744 , n219745 , n219746 , n219747 , n219748 , 
 n219749 , n219750 , n219751 , n219752 , n219753 , n219754 , n219755 , n219756 , n219757 , n219758 , 
 n219759 , n219760 , n219761 , n219762 , n219763 , n219764 , n219765 , n219766 , n219767 , n219768 , 
 n219769 , n219770 , n219771 , n219772 , n219773 , n219774 , n219775 , n219776 , n219777 , n219778 , 
 n219779 , n219780 , n219781 , n219782 , n219783 , n219784 , n219785 , n219786 , n219787 , n219788 , 
 n219789 , n219790 , n219791 , n219792 , n219793 , n219794 , n219795 , n219796 , n219797 , n219798 , 
 n219799 , n219800 , n219801 , n219802 , n219803 , n219804 , n219805 , n219806 , n219807 , n219808 , 
 n219809 , n219810 , n219811 , n219812 , n219813 , n219814 , n219815 , n219816 , n219817 , n219818 , 
 n219819 , n219820 , n219821 , n219822 , n219823 , n219824 , n219825 , n219826 , n219827 , n219828 , 
 n219829 , n219830 , n219831 , n219832 , n219833 , n219834 , n219835 , n219836 , n219837 , n219838 , 
 n219839 , n219840 , n219841 , n219842 , n219843 , n219844 , n219845 , n219846 , n219847 , n219848 , 
 n219849 , n219850 , n219851 , n219852 , n219853 , n219854 , n219855 , n219856 , n219857 , n219858 , 
 n219859 , n219860 , n219861 , n219862 , n219863 , n219864 , n219865 , n219866 , n219867 , n219868 , 
 n219869 , n219870 , n219871 , n219872 , n219873 , n219874 , n219875 , n219876 , n219877 , n219878 , 
 n219879 , n219880 , n219881 , n219882 , n219883 , n219884 , n219885 , n219886 , n219887 , n219888 , 
 n219889 , n219890 , n219891 , n219892 , n219893 , n219894 , n219895 , n219896 , n219897 , n219898 , 
 n219899 , n219900 , n219901 , n219902 , n219903 , n219904 , n219905 , n219906 , n219907 , n219908 , 
 n219909 , n219910 , n219911 , n219912 , n219913 , n219914 , n219915 , n219916 , n219917 , n219918 , 
 n219919 , n219920 , n219921 , n219922 , n219923 , n219924 , n219925 , n219926 , n219927 , n219928 , 
 n219929 , n219930 , n219931 , n219932 , n219933 , n219934 , n219935 , n219936 , n219937 , n219938 , 
 n219939 , n219940 , n219941 , n219942 , n219943 , n219944 , n219945 , n219946 , n219947 , n219948 , 
 n219949 , n219950 , n219951 , n219952 , n219953 , n219954 , n219955 , n219956 , n219957 , n219958 , 
 n219959 , n219960 , n219961 , n219962 , n219963 , n219964 , n219965 , n219966 , n219967 , n219968 , 
 n219969 , n219970 , n219971 , n219972 , n219973 , n219974 , n219975 , n219976 , n219977 , n219978 , 
 n219979 , n219980 , n219981 , n219982 , n219983 , n219984 , n219985 , n219986 , n219987 , n219988 , 
 n219989 , n219990 , n219991 , n219992 , n219993 , n219994 , n219995 , n219996 , n219997 , n219998 , 
 n219999 , n220000 , n220001 , n220002 , n220003 , n220004 , n220005 , n220006 , n220007 , n220008 , 
 n220009 , n220010 , n220011 , n220012 , n220013 , n220014 , n220015 , n220016 , n220017 , n220018 , 
 n220019 , n220020 , n220021 , n220022 , n220023 , n220024 , n220025 , n220026 , n220027 , n220028 , 
 n220029 , n220030 , n220031 , n220032 , n220033 , n220034 , n220035 , n220036 , n220037 , n220038 , 
 n220039 , n220040 , n220041 , n220042 , n220043 , n220044 , n220045 , n220046 , n220047 , n220048 , 
 n220049 , n220050 , n220051 , n220052 , n220053 , n220054 , n220055 , n220056 , n220057 , n220058 , 
 n220059 , n220060 , n220061 , n220062 , n220063 , n220064 , n220065 , n220066 , n220067 , n220068 , 
 n220069 , n220070 , n220071 , n220072 , n220073 , n220074 , n220075 , n220076 , n220077 , n220078 , 
 n220079 , n220080 , n220081 , n220082 , n220083 , n220084 , n220085 , n220086 , n220087 , n220088 , 
 n220089 , n220090 , n220091 , n220092 , n220093 , n220094 , n220095 , n220096 , n220097 , n220098 , 
 n220099 , n220100 , n220101 , n220102 , n220103 , n220104 , n220105 , n220106 , n220107 , n220108 , 
 n220109 , n220110 , n220111 , n220112 , n220113 , n220114 , n220115 , n220116 , n220117 , n220118 , 
 n220119 , n220120 , n220121 , n220122 , n220123 , n220124 , n220125 , n220126 , n220127 , n220128 , 
 n220129 , n220130 , n220131 , n220132 , n220133 , n220134 , n220135 , n220136 , n220137 , n220138 , 
 n220139 , n220140 , n220141 , n220142 , n220143 , n220144 , n220145 , n220146 , n220147 , n220148 , 
 n220149 , n220150 , n220151 , n220152 , n220153 , n220154 , n220155 , n220156 , n220157 , n220158 , 
 n220159 , n220160 , n220161 , n220162 , n220163 , n220164 , n220165 , n220166 , n220167 , n220168 , 
 n220169 , n220170 , n220171 , n220172 , n220173 , n220174 , n220175 , n220176 , n220177 , n220178 , 
 n220179 , n220180 , n220181 , n220182 , n220183 , n220184 , n220185 , n220186 , n220187 , n220188 , 
 n220189 , n220190 , n220191 , n220192 , n220193 , n220194 , n220195 , n220196 , n220197 , n220198 , 
 n220199 , n220200 , n220201 , n220202 , n220203 , n220204 , n220205 , n220206 , n220207 , n220208 , 
 n220209 , n220210 , n220211 , n220212 , n220213 , n220214 , n220215 , n220216 , n220217 , n220218 , 
 n220219 , n220220 , n220221 , n220222 , n220223 , n220224 , n220225 , n220226 , n220227 , n220228 , 
 n220229 , n220230 , n220231 , n220232 , n220233 , n220234 , n220235 , n220236 , n220237 , n220238 , 
 n220239 , n220240 , n220241 , n220242 , n220243 , n220244 , n220245 , n220246 , n220247 , n220248 , 
 n220249 , n220250 , n220251 , n220252 , n220253 , n220254 , n220255 , n220256 , n220257 , n220258 , 
 n220259 , n220260 , n220261 , n220262 , n220263 , n220264 , n220265 , n220266 , n220267 , n220268 , 
 n220269 , n220270 , n220271 , n220272 , n220273 , n220274 , n220275 , n220276 , n220277 , n220278 , 
 n220279 , n220280 , n220281 , n220282 , n220283 , n220284 , n220285 , n220286 , n220287 , n220288 , 
 n220289 , n220290 , n220291 , n220292 , n220293 , n220294 , n220295 , n220296 , n220297 , n220298 , 
 n220299 , n220300 , n220301 , n220302 , n220303 , n220304 , n220305 , n220306 , n220307 , n220308 , 
 n220309 , n220310 , n220311 , n220312 , n220313 , n220314 , n220315 , n220316 , n220317 , n220318 , 
 n220319 , n220320 , n220321 , n220322 , n220323 , n220324 , n220325 , n220326 , n220327 , n220328 , 
 n220329 , n220330 , n220331 , n220332 , n220333 , n220334 , n220335 , n220336 , n220337 , n220338 , 
 n220339 , n220340 , n220341 , n220342 , n220343 , n220344 , n220345 , n220346 , n220347 , n220348 , 
 n220349 , n220350 , n220351 , n220352 , n220353 , n220354 , n220355 , n220356 , n220357 , n220358 , 
 n220359 , n220360 , n220361 , n220362 , n220363 , n220364 , n220365 , n220366 , n220367 , n220368 , 
 n220369 , n220370 , n220371 , n220372 , n220373 , n220374 , n220375 , n220376 , n220377 , n220378 , 
 n220379 , n220380 , n220381 , n220382 , n220383 , n220384 , n220385 , n220386 , n220387 , n220388 , 
 n220389 , n220390 , n220391 , n220392 , n220393 , n220394 , n220395 , n220396 , n220397 , n220398 , 
 n220399 , n220400 , n220401 , n220402 , n220403 , n220404 , n220405 , n220406 , n220407 , n220408 , 
 n220409 , n220410 , n220411 , n220412 , n220413 , n220414 , n220415 , n220416 , n220417 , n220418 , 
 n220419 , n220420 , n220421 , n220422 , n220423 , n220424 , n220425 , n220426 , n220427 , n220428 , 
 n220429 , n220430 , n220431 , n220432 , n220433 , n220434 , n220435 , n220436 , n220437 , n220438 , 
 n220439 , n220440 , n220441 , n220442 , n220443 , n220444 , n220445 , n220446 , n220447 , n220448 , 
 n220449 , n220450 , n220451 , n220452 , n220453 , n220454 , n220455 , n220456 , n220457 , n220458 , 
 n220459 , n220460 , n220461 , n220462 , n220463 , n220464 , n220465 , n220466 , n220467 , n220468 , 
 n220469 , n220470 , n220471 , n220472 , n220473 , n220474 , n220475 , n220476 , n220477 , n220478 , 
 n220479 , n220480 , n220481 , n220482 , n220483 , n220484 , n220485 , n220486 , n220487 , n220488 , 
 n220489 , n220490 , n220491 , n220492 , n220493 , n220494 , n220495 , n220496 , n220497 , n220498 , 
 n220499 , n220500 , n220501 , n220502 , n220503 , n220504 , n220505 , n220506 , n220507 , n220508 , 
 n220509 , n220510 , n220511 , n220512 , n220513 , n220514 , n220515 , n220516 , n220517 , n220518 , 
 n220519 , n220520 , n220521 , n220522 , n220523 , n220524 , n220525 , n220526 , n220527 , n220528 , 
 n220529 , n220530 , n220531 , n220532 , n220533 , n220534 , n220535 , n220536 , n220537 , n220538 , 
 n220539 , n220540 , n220541 , n220542 , n220543 , n220544 , n220545 , n220546 , n220547 , n220548 , 
 n220549 , n220550 , n220551 , n220552 , n220553 , n220554 , n220555 , n220556 , n220557 , n220558 , 
 n220559 , n220560 , n220561 , n220562 , n220563 , n220564 , n220565 , n220566 , n220567 , n220568 , 
 n220569 , n220570 , n220571 , n220572 , n220573 , n220574 , n220575 , n220576 , n220577 , n220578 , 
 n220579 , n220580 , n220581 , n220582 , n220583 , n220584 , n220585 , n220586 , n220587 , n220588 , 
 n220589 , n220590 , n220591 , n220592 , n220593 , n220594 , n220595 , n220596 , n220597 , n220598 , 
 n220599 , n220600 , n220601 , n220602 , n220603 , n220604 , n220605 , n220606 , n220607 , n220608 , 
 n220609 , n220610 , n220611 , n220612 , n220613 , n220614 , n220615 , n220616 , n220617 , n220618 , 
 n220619 , n220620 , n220621 , n220622 , n220623 , n220624 , n220625 , n220626 , n220627 , n220628 , 
 n220629 , n220630 , n220631 , n220632 , n220633 , n220634 , n220635 , n220636 , n220637 , n220638 , 
 n220639 , n220640 , n220641 , n220642 , n220643 , n220644 , n220645 , n220646 , n220647 , n220648 , 
 n220649 , n220650 , n220651 , n220652 , n220653 , n220654 , n220655 , n220656 , n220657 , n220658 , 
 n220659 , n220660 , n220661 , n220662 , n220663 , n220664 , n220665 , n220666 , n220667 , n220668 , 
 n220669 , n220670 , n220671 , n220672 , n220673 , n220674 , n220675 , n220676 , n220677 , n220678 , 
 n220679 , n220680 , n220681 , n220682 , n220683 , n220684 , n220685 , n220686 , n220687 , n220688 , 
 n220689 , n220690 , n220691 , n220692 , n220693 , n220694 , n220695 , n220696 , n220697 , n220698 , 
 n220699 , n220700 , n220701 , n220702 , n220703 , n220704 , n220705 , n220706 , n220707 , n220708 , 
 n220709 , n220710 , n220711 , n220712 , n220713 , n220714 , n220715 , n220716 , n220717 , n220718 , 
 n220719 , n220720 , n220721 , n220722 , n220723 , n220724 , n220725 , n220726 , n220727 , n220728 , 
 n220729 , n220730 , n220731 , n220732 , n220733 , n220734 , n220735 , n220736 , n220737 , n220738 , 
 n220739 , n220740 , n220741 , n220742 , n220743 , n220744 , n220745 , n220746 , n220747 , n220748 , 
 n220749 , n220750 , n220751 , n220752 , n220753 , n220754 , n220755 , n220756 , n220757 , n220758 , 
 n220759 , n220760 , n220761 , n220762 , n220763 , n220764 , n220765 , n220766 , n220767 , n220768 , 
 n220769 , n220770 , n220771 , n220772 , n220773 , n220774 , n220775 , n220776 , n220777 , n220778 , 
 n220779 , n220780 , n220781 , n220782 , n220783 , n220784 , n220785 , n220786 , n220787 , n220788 , 
 n220789 , n220790 , n220791 , n220792 , n220793 , n220794 , n220795 , n220796 , n220797 , n220798 , 
 n220799 , n220800 , n220801 , n220802 , n220803 , n220804 , n220805 , n220806 , n220807 , n220808 , 
 n220809 , n220810 , n220811 , n220812 , n220813 , n220814 , n220815 , n220816 , n220817 , n220818 , 
 n220819 , n220820 , n220821 , n220822 , n220823 , n220824 , n220825 , n220826 , n220827 , n220828 , 
 n220829 , n220830 , n220831 , n220832 , n220833 , n220834 , n220835 , n220836 , n220837 , n220838 , 
 n220839 , n220840 , n220841 , n220842 , n220843 , n220844 , n220845 , n220846 , n220847 , n220848 , 
 n220849 , n220850 , n220851 , n220852 , n220853 , n220854 , n220855 , n220856 , n220857 , n220858 , 
 n220859 , n220860 , n220861 , n220862 , n220863 , n220864 , n220865 , n220866 , n220867 , n220868 , 
 n220869 , n220870 , n220871 , n220872 , n220873 , n220874 , n220875 , n220876 , n220877 , n220878 , 
 n220879 , n220880 , n220881 , n220882 , n220883 , n220884 , n220885 , n220886 , n220887 , n220888 , 
 n220889 , n220890 , n220891 , n220892 , n220893 , n220894 , n220895 , n220896 , n220897 , n220898 , 
 n220899 , n220900 , n220901 , n220902 , n220903 , n220904 , n220905 , n220906 , n220907 , n220908 , 
 n220909 , n220910 , n220911 , n220912 , n220913 , n220914 , n220915 , n220916 , n220917 , n220918 , 
 n220919 , n220920 , n220921 , n220922 , n220923 , n220924 , n220925 , n220926 , n220927 , n220928 , 
 n220929 , n220930 , n220931 , n220932 , n220933 , n220934 , n220935 , n220936 , n220937 , n220938 , 
 n220939 , n220940 , n220941 , n220942 , n220943 , n220944 , n220945 , n220946 , n220947 , n220948 , 
 n220949 , n220950 , n220951 , n220952 , n220953 , n220954 , n220955 , n220956 , n220957 , n220958 , 
 n220959 , n220960 , n220961 , n220962 , n220963 , n220964 , n220965 , n220966 , n220967 , n220968 , 
 n220969 , n220970 , n220971 , n220972 , n220973 , n220974 , n220975 , n220976 , n220977 , n220978 , 
 n220979 , n220980 , n220981 , n220982 , n220983 , n220984 , n220985 , n220986 , n220987 , n220988 , 
 n220989 , n220990 , n220991 , n220992 , n220993 , n220994 , n220995 , n220996 , n220997 , n220998 , 
 n220999 , n221000 , n221001 , n221002 , n221003 , n221004 , n221005 , n221006 , n221007 , n221008 , 
 n221009 , n221010 , n221011 , n221012 , n221013 , n221014 , n221015 , n221016 , n221017 , n221018 , 
 n221019 , n221020 , n221021 , n221022 , n221023 , n221024 , n221025 , n221026 , n221027 , n221028 , 
 n221029 , n221030 , n221031 , n221032 , n221033 , n221034 , n221035 , n221036 , n221037 , n221038 , 
 n221039 , n221040 , n221041 , n221042 , n221043 , n221044 , n221045 , n221046 , n221047 , n221048 , 
 n221049 , n221050 , n221051 , n221052 , n221053 , n221054 , n221055 , n221056 , n221057 , n221058 , 
 n221059 , n221060 , n221061 , n221062 , n221063 , n221064 , n221065 , n221066 , n221067 , n221068 , 
 n221069 , n221070 , n221071 , n221072 , n221073 , n221074 , n221075 , n221076 , n221077 , n221078 , 
 n221079 , n221080 , n221081 , n221082 , n221083 , n221084 , n221085 , n221086 , n221087 , n221088 , 
 n221089 , n221090 , n221091 , n221092 , n221093 , n221094 , n221095 , n221096 , n221097 , n221098 , 
 n221099 , n221100 , n221101 , n221102 , n221103 , n221104 , n221105 , n221106 , n221107 , n221108 , 
 n221109 , n221110 , n221111 , n221112 , n221113 , n221114 , n221115 , n221116 , n221117 , n221118 , 
 n221119 , n221120 , n221121 , n221122 , n221123 , n221124 , n221125 , n221126 , n221127 , n221128 , 
 n221129 , n221130 , n221131 , n221132 , n221133 , n221134 , n221135 , n221136 , n221137 , n221138 , 
 n221139 , n221140 , n221141 , n221142 , n221143 , n221144 , n221145 , n221146 , n221147 , n221148 , 
 n221149 , n221150 , n221151 , n221152 , n221153 , n221154 , n221155 , n221156 , n221157 , n221158 , 
 n221159 , n221160 , n221161 , n221162 , n221163 , n221164 , n221165 , n221166 , n221167 , n221168 , 
 n221169 , n221170 , n221171 , n221172 , n221173 , n221174 , n221175 , n221176 , n221177 , n221178 , 
 n221179 , n221180 , n221181 , n221182 , n221183 , n221184 , n221185 , n221186 , n221187 , n221188 , 
 n221189 , n221190 , n221191 , n221192 , n221193 , n221194 , n221195 , n221196 , n221197 , n221198 , 
 n221199 , n221200 , n221201 , n221202 , n221203 , n221204 , n221205 , n221206 , n221207 , n221208 , 
 n221209 , n221210 , n221211 , n221212 , n221213 , n221214 , n221215 , n221216 , n221217 , n221218 , 
 n221219 , n221220 , n221221 , n221222 , n221223 , n221224 , n221225 , n221226 , n221227 , n221228 , 
 n221229 , n221230 , n221231 , n221232 , n221233 , n221234 , n221235 , n221236 , n221237 , n221238 , 
 n221239 , n221240 , n221241 , n221242 , n221243 , n221244 , n221245 , n221246 , n221247 , n221248 , 
 n221249 , n221250 , n221251 , n221252 , n221253 , n221254 , n221255 , n221256 , n221257 , n221258 , 
 n221259 , n221260 , n221261 , n221262 , n221263 , n221264 , n221265 , n221266 , n221267 , n221268 , 
 n221269 , n221270 , n221271 , n221272 , n221273 , n221274 , n221275 , n221276 , n221277 , n221278 , 
 n221279 , n221280 , n221281 , n221282 , n221283 , n221284 , n221285 , n221286 , n221287 , n221288 , 
 n221289 , n221290 , n221291 , n221292 , n221293 , n221294 , n221295 , n221296 , n221297 , n221298 , 
 n221299 , n221300 , n221301 , n221302 , n221303 , n221304 , n221305 , n221306 , n221307 , n221308 , 
 n221309 , n221310 , n221311 , n221312 , n221313 , n221314 , n221315 , n221316 , n221317 , n221318 , 
 n221319 , n221320 , n221321 , n221322 , n221323 , n221324 , n221325 , n221326 , n221327 , n221328 , 
 n221329 , n221330 , n221331 , n221332 , n221333 , n221334 , n221335 , n221336 , n221337 , n221338 , 
 n221339 , n221340 , n221341 , n221342 , n221343 , n221344 , n221345 , n221346 , n221347 , n221348 , 
 n221349 , n221350 , n221351 , n221352 , n221353 , n221354 , n221355 , n221356 , n221357 , n221358 , 
 n221359 , n221360 , n221361 , n221362 , n221363 , n221364 , n221365 , n221366 , n221367 , n221368 , 
 n221369 , n221370 , n221371 , n221372 , n221373 , n221374 , n221375 , n221376 , n221377 , n221378 , 
 n221379 , n221380 , n221381 , n221382 , n221383 , n221384 , n221385 , n221386 , n221387 , n221388 , 
 n221389 , n221390 , n221391 , n221392 , n221393 , n221394 , n221395 , n221396 , n221397 , n221398 , 
 n221399 , n221400 , n221401 , n221402 , n221403 , n221404 , n221405 , n221406 , n221407 , n221408 , 
 n221409 , n221410 , n221411 , n221412 , n221413 , n221414 , n221415 , n221416 , n221417 , n221418 , 
 n221419 , n221420 , n221421 , n221422 , n221423 , n221424 , n221425 , n221426 , n221427 , n221428 , 
 n221429 , n221430 , n221431 , n221432 , n221433 , n221434 , n221435 , n221436 , n221437 , n221438 , 
 n221439 , n221440 , n221441 , n221442 , n221443 , n221444 , n221445 , n221446 , n221447 , n221448 , 
 n221449 , n221450 , n221451 , n221452 , n221453 , n221454 , n221455 , n221456 , n221457 , n221458 , 
 n221459 , n221460 , n221461 , n221462 , n221463 , n221464 , n221465 , n221466 , n221467 , n221468 , 
 n221469 , n221470 , n221471 , n221472 , n221473 , n221474 , n221475 , n221476 , n221477 , n221478 , 
 n221479 , n221480 , n221481 , n221482 , n221483 , n221484 , n221485 , n221486 , n221487 , n221488 , 
 n221489 , n221490 , n221491 , n221492 , n221493 , n221494 , n221495 , n221496 , n221497 , n221498 , 
 n221499 , n221500 , n221501 , n221502 , n221503 , n221504 , n221505 , n221506 , n221507 , n221508 , 
 n221509 , n221510 , n221511 , n221512 , n221513 , n221514 , n221515 , n221516 , n221517 , n221518 , 
 n221519 , n221520 , n221521 , n221522 , n221523 , n221524 , n221525 , n221526 , n221527 , n221528 , 
 n221529 , n221530 , n221531 , n221532 , n221533 , n221534 , n221535 , n221536 , n221537 , n221538 , 
 n221539 , n221540 , n221541 , n221542 , n221543 , n221544 , n221545 , n221546 , n221547 , n221548 , 
 n221549 , n221550 , n221551 , n221552 , n221553 , n221554 , n221555 , n221556 , n221557 , n221558 , 
 n221559 , n221560 , n221561 , n221562 , n221563 , n221564 , n221565 , n221566 , n221567 , n221568 , 
 n221569 , n221570 , n221571 , n221572 , n221573 , n221574 , n221575 , n221576 , n221577 , n221578 , 
 n221579 , n221580 , n221581 , n221582 , n221583 , n221584 , n221585 , n221586 , n221587 , n221588 , 
 n221589 , n221590 , n221591 , n221592 , n221593 , n221594 , n221595 , n221596 , n221597 , n221598 , 
 n221599 , n221600 , n221601 , n221602 , n221603 , n221604 , n221605 , n221606 , n221607 , n221608 , 
 n221609 , n221610 , n221611 , n221612 , n221613 , n221614 , n221615 , n221616 , n221617 , n221618 , 
 n221619 , n221620 , n221621 , n221622 , n221623 , n221624 , n221625 , n221626 , n221627 , n221628 , 
 n221629 , n221630 , n221631 , n221632 , n221633 , n221634 , n221635 , n221636 , n221637 , n221638 , 
 n221639 , n221640 , n221641 , n221642 , n221643 , n221644 , n221645 , n221646 , n221647 , n221648 , 
 n221649 , n221650 , n221651 , n221652 , n221653 , n221654 , n221655 , n221656 , n221657 , n221658 , 
 n221659 , n221660 , n221661 , n221662 , n221663 , n221664 , n221665 , n221666 , n221667 , n221668 , 
 n221669 , n221670 , n221671 , n221672 , n221673 , n221674 , n221675 , n221676 , n221677 , n221678 , 
 n221679 , n221680 , n221681 , n221682 , n221683 , n221684 , n221685 , n221686 , n221687 , n221688 , 
 n221689 , n221690 , n221691 , n221692 , n221693 , n221694 , n221695 , n221696 , n221697 , n221698 , 
 n221699 , n221700 , n221701 , n221702 , n221703 , n221704 , n221705 , n221706 , n221707 , n221708 , 
 n221709 , n221710 , n221711 , n221712 , n221713 , n221714 , n221715 , n221716 , n221717 , n221718 , 
 n221719 , n221720 , n221721 , n221722 , n221723 , n221724 , n221725 , n221726 , n221727 , n221728 , 
 n221729 , n221730 , n221731 , n221732 , n221733 , n221734 , n221735 , n221736 , n221737 , n221738 , 
 n221739 , n221740 , n221741 , n221742 , n221743 , n221744 , n221745 , n221746 , n221747 , n221748 , 
 n221749 , n221750 , n221751 , n221752 , n221753 , n221754 , n221755 , n221756 , n221757 , n221758 , 
 n221759 , n221760 , n221761 , n221762 , n221763 , n221764 , n221765 , n221766 , n221767 , n221768 , 
 n221769 , n221770 , n221771 , n221772 , n221773 , n221774 , n221775 , n221776 , n221777 , n221778 , 
 n221779 , n221780 , n221781 , n221782 , n221783 , n221784 , n221785 , n221786 , n221787 , n221788 , 
 n221789 , n221790 , n221791 , n221792 , n221793 , n221794 , n221795 , n221796 , n221797 , n221798 , 
 n221799 , n221800 , n221801 , n221802 , n221803 , n221804 , n221805 , n221806 , n221807 , n221808 , 
 n221809 , n221810 , n221811 , n221812 , n221813 , n221814 , n221815 , n221816 , n221817 , n221818 , 
 n221819 , n221820 , n221821 , n221822 , n221823 , n221824 , n221825 , n221826 , n221827 , n221828 , 
 n221829 , n221830 , n221831 , n221832 , n221833 , n221834 , n221835 , n221836 , n221837 , n221838 , 
 n221839 , n221840 , n221841 , n221842 , n221843 , n221844 , n221845 , n221846 , n221847 , n221848 , 
 n221849 , n221850 , n221851 , n221852 , n221853 , n221854 , n221855 , n221856 , n221857 , n221858 , 
 n221859 , n221860 , n221861 , n221862 , n221863 , n221864 , n221865 , n221866 , n221867 , n221868 , 
 n221869 , n221870 , n221871 , n221872 , n221873 , n221874 , n221875 , n221876 , n221877 , n221878 , 
 n221879 , n221880 , n221881 , n221882 , n221883 , n221884 , n221885 , n221886 , n221887 , n221888 , 
 n221889 , n221890 , n221891 , n221892 , n221893 , n221894 , n221895 , n221896 , n221897 , n221898 , 
 n221899 , n221900 , n221901 , n221902 , n221903 , n221904 , n221905 , n221906 , n221907 , n221908 , 
 n221909 , n221910 , n221911 , n221912 , n221913 , n221914 , n221915 , n221916 , n221917 , n221918 , 
 n221919 , n221920 , n221921 , n221922 , n221923 , n221924 , n221925 , n221926 , n221927 , n221928 , 
 n221929 , n221930 , n221931 , n221932 , n221933 , n221934 , n221935 , n221936 , n221937 , n221938 , 
 n221939 , n221940 , n221941 , n221942 , n221943 , n221944 , n221945 , n221946 , n221947 , n221948 , 
 n221949 , n221950 , n221951 , n221952 , n221953 , n221954 , n221955 , n221956 , n221957 , n221958 , 
 n221959 , n221960 , n221961 , n221962 , n221963 , n221964 , n221965 , n221966 , n221967 , n221968 , 
 n221969 , n221970 , n221971 , n221972 , n221973 , n221974 , n221975 , n221976 , n221977 , n221978 , 
 n221979 , n221980 , n221981 , n221982 , n221983 , n221984 , n221985 , n221986 , n221987 , n221988 , 
 n221989 , n221990 , n221991 , n221992 , n221993 , n221994 , n221995 , n221996 , n221997 , n221998 , 
 n221999 , n222000 , n222001 , n222002 , n222003 , n222004 , n222005 , n222006 , n222007 , n222008 , 
 n222009 , n222010 , n222011 , n222012 , n222013 , n222014 , n222015 , n222016 , n222017 , n222018 , 
 n222019 , n222020 , n222021 , n222022 , n222023 , n222024 , n222025 , n222026 , n222027 , n222028 , 
 n222029 , n222030 , n222031 , n222032 , n222033 , n222034 , n222035 , n222036 , n222037 , n222038 , 
 n222039 , n222040 , n222041 , n222042 , n222043 , n222044 , n222045 , n222046 , n222047 , n222048 , 
 n222049 , n222050 , n222051 , n222052 , n222053 , n222054 , n222055 , n222056 , n222057 , n222058 , 
 n222059 , n222060 , n222061 , n222062 , n222063 , n222064 , n222065 , n222066 , n222067 , n222068 , 
 n222069 , n222070 , n222071 , n222072 , n222073 , n222074 , n222075 , n222076 , n222077 , n222078 , 
 n222079 , n222080 , n222081 , n222082 , n222083 , n222084 , n222085 , n222086 , n222087 , n222088 , 
 n222089 , n222090 , n222091 , n222092 , n222093 , n222094 , n222095 , n222096 , n222097 , n222098 , 
 n222099 , n222100 , n222101 , n222102 , n222103 , n222104 , n222105 , n222106 , n222107 , n222108 , 
 n222109 , n222110 , n222111 , n222112 , n222113 , n222114 , n222115 , n222116 , n222117 , n222118 , 
 n222119 , n222120 , n222121 , n222122 , n222123 , n222124 , n222125 , n222126 , n222127 , n222128 , 
 n222129 , n222130 , n222131 , n222132 , n222133 , n222134 , n222135 , n222136 , n222137 , n222138 , 
 n222139 , n222140 , n222141 , n222142 , n222143 , n222144 , n222145 , n222146 , n222147 , n222148 , 
 n222149 , n222150 , n222151 , n222152 , n222153 , n222154 , n222155 , n222156 , n222157 , n222158 , 
 n222159 , n222160 , n222161 , n222162 , n222163 , n222164 , n222165 , n222166 , n222167 , n222168 , 
 n222169 , n222170 , n222171 , n222172 , n222173 , n222174 , n222175 , n222176 , n222177 , n222178 , 
 n222179 , n222180 , n222181 , n222182 , n222183 , n222184 , n222185 , n222186 , n222187 , n222188 , 
 n222189 , n222190 , n222191 , n222192 , n222193 , n222194 , n222195 , n222196 , n222197 , n222198 , 
 n222199 , n222200 , n222201 , n222202 , n222203 , n222204 , n222205 , n222206 , n222207 , n222208 , 
 n222209 , n222210 , n222211 , n222212 , n222213 , n222214 , n222215 , n222216 , n222217 , n222218 , 
 n222219 , n222220 , n222221 , n222222 , n222223 , n222224 , n222225 , n222226 , n222227 , n222228 , 
 n222229 , n222230 , n222231 , n222232 , n222233 , n222234 , n222235 , n222236 , n222237 , n222238 , 
 n222239 , n222240 , n222241 , n222242 , n222243 , n222244 , n222245 , n222246 , n222247 , n222248 , 
 n222249 , n222250 , n222251 , n222252 , n222253 , n222254 , n222255 , n222256 , n222257 , n222258 , 
 n222259 , n222260 , n222261 , n222262 , n222263 , n222264 , n222265 , n222266 , n222267 , n222268 , 
 n222269 , n222270 , n222271 , n222272 , n222273 , n222274 , n222275 , n222276 , n222277 , n222278 , 
 n222279 , n222280 , n222281 , n222282 , n222283 , n222284 , n222285 , n222286 , n222287 , n222288 , 
 n222289 , n222290 , n222291 , n222292 , n222293 , n222294 , n222295 , n222296 , n222297 , n222298 , 
 n222299 , n222300 , n222301 , n222302 , n222303 , n222304 , n222305 , n222306 , n222307 , n222308 , 
 n222309 , n222310 , n222311 , n222312 , n222313 , n222314 , n222315 , n222316 , n222317 , n222318 , 
 n222319 , n222320 , n222321 , n222322 , n222323 , n222324 , n222325 , n222326 , n222327 , n222328 , 
 n222329 , n222330 , n222331 , n222332 , n222333 , n222334 , n222335 , n222336 , n222337 , n222338 , 
 n222339 , n222340 , n222341 , n222342 , n222343 , n222344 , n222345 , n222346 , n222347 , n222348 , 
 n222349 , n222350 , n222351 , n222352 , n222353 , n222354 , n222355 , n222356 , n222357 , n222358 , 
 n222359 , n222360 , n222361 , n222362 , n222363 , n222364 , n222365 , n222366 , n222367 , n222368 , 
 n222369 , n222370 , n222371 , n222372 , n222373 , n222374 , n222375 , n222376 , n222377 , n222378 , 
 n222379 , n222380 , n222381 , n222382 , n222383 , n222384 , n222385 , n222386 , n222387 , n222388 , 
 n222389 , n222390 , n222391 , n222392 , n222393 , n222394 , n222395 , n222396 , n222397 , n222398 , 
 n222399 , n222400 , n222401 , n222402 , n222403 , n222404 , n222405 , n222406 , n222407 , n222408 , 
 n222409 , n222410 , n222411 , n222412 , n222413 , n222414 , n222415 , n222416 , n222417 , n222418 , 
 n222419 , n222420 , n222421 , n222422 , n222423 , n222424 , n222425 , n222426 , n222427 , n222428 , 
 n222429 , n222430 , n222431 , n222432 , n222433 , n222434 , n222435 , n222436 , n222437 , n222438 , 
 n222439 , n222440 , n222441 , n222442 , n222443 , n222444 , n222445 , n222446 , n222447 , n222448 , 
 n222449 , n222450 , n222451 , n222452 , n222453 , n222454 , n222455 , n222456 , n222457 , n222458 , 
 n222459 , n222460 , n222461 , n222462 , n222463 , n222464 , n222465 , n222466 , n222467 , n222468 , 
 n222469 , n222470 , n222471 , n222472 , n222473 , n222474 , n222475 , n222476 , n222477 , n222478 , 
 n222479 , n222480 , n222481 , n222482 , n222483 , n222484 , n222485 , n222486 , n222487 , n222488 , 
 n222489 , n222490 , n222491 , n222492 , n222493 , n222494 , n222495 , n222496 , n222497 , n222498 , 
 n222499 , n222500 , n222501 , n222502 , n222503 , n222504 , n222505 , n222506 , n222507 , n222508 , 
 n222509 , n222510 , n222511 , n222512 , n222513 , n222514 , n222515 , n222516 , n222517 , n222518 , 
 n222519 , n222520 , n222521 , n222522 , n222523 , n222524 , n222525 , n222526 , n222527 , n222528 , 
 n222529 , n222530 , n222531 , n222532 , n222533 , n222534 , n222535 , n222536 , n222537 , n222538 , 
 n222539 , n222540 , n222541 , n222542 , n222543 , n222544 , n222545 , n222546 , n222547 , n222548 , 
 n222549 , n222550 , n222551 , n222552 , n222553 , n222554 , n222555 , n222556 , n222557 , n222558 , 
 n222559 , n222560 , n222561 , n222562 , n222563 , n222564 , n222565 , n222566 , n222567 , n222568 , 
 n222569 , n222570 , n222571 , n222572 , n222573 , n222574 , n222575 , n222576 , n222577 , n222578 , 
 n222579 , n222580 , n222581 , n222582 , n222583 , n222584 , n222585 , n222586 , n222587 , n222588 , 
 n222589 , n222590 , n222591 , n222592 , n222593 , n222594 , n222595 , n222596 , n222597 , n222598 , 
 n222599 , n222600 , n222601 , n222602 , n222603 , n222604 , n222605 , n222606 , n222607 , n222608 , 
 n222609 , n222610 , n222611 , n222612 , n222613 , n222614 , n222615 , n222616 , n222617 , n222618 , 
 n222619 , n222620 , n222621 , n222622 , n222623 , n222624 , n222625 , n222626 , n222627 , n222628 , 
 n222629 , n222630 , n222631 , n222632 , n222633 , n222634 , n222635 , n222636 , n222637 , n222638 , 
 n222639 , n222640 , n222641 , n222642 , n222643 , n222644 , n222645 , n222646 , n222647 , n222648 , 
 n222649 , n222650 , n222651 , n222652 , n222653 , n222654 , n222655 , n222656 , n222657 , n222658 , 
 n222659 , n222660 , n222661 , n222662 , n222663 , n222664 , n222665 , n222666 , n222667 , n222668 , 
 n222669 , n222670 , n222671 , n222672 , n222673 , n222674 , n222675 , n222676 , n222677 , n222678 , 
 n222679 , n222680 , n222681 , n222682 , n222683 , n222684 , n222685 , n222686 , n222687 , n222688 , 
 n222689 , n222690 , n222691 , n222692 , n222693 , n222694 , n222695 , n222696 , n222697 , n222698 , 
 n222699 , n222700 , n222701 , n222702 , n222703 , n222704 , n222705 , n222706 , n222707 , n222708 , 
 n222709 , n222710 , n222711 , n222712 , n222713 , n222714 , n222715 , n222716 , n222717 , n222718 , 
 n222719 , n222720 , n222721 , n222722 , n222723 , n222724 , n222725 , n222726 , n222727 , n222728 , 
 n222729 , n222730 , n222731 , n222732 , n222733 , n222734 , n222735 , n222736 , n222737 , n222738 , 
 n222739 , n222740 , n222741 , n222742 , n222743 , n222744 , n222745 , n222746 , n222747 , n222748 , 
 n222749 , n222750 , n222751 , n222752 , n222753 , n222754 , n222755 , n222756 , n222757 , n222758 , 
 n222759 , n222760 , n222761 , n222762 , n222763 , n222764 , n222765 , n222766 , n222767 , n222768 , 
 n222769 , n222770 , n222771 , n222772 , n222773 , n222774 , n222775 , n222776 , n222777 , n222778 , 
 n222779 , n222780 , n222781 , n222782 , n222783 , n222784 , n222785 , n222786 , n222787 , n222788 , 
 n222789 , n222790 , n222791 , n222792 , n222793 , n222794 , n222795 , n222796 , n222797 , n222798 , 
 n222799 , n222800 , n222801 , n222802 , n222803 , n222804 , n222805 , n222806 , n222807 , n222808 , 
 n222809 , n222810 , n222811 , n222812 , n222813 , n222814 , n222815 , n222816 , n222817 , n222818 , 
 n222819 , n222820 , n222821 , n222822 , n222823 , n222824 , n222825 , n222826 , n222827 , n222828 , 
 n222829 , n222830 , n222831 , n222832 , n222833 , n222834 , n222835 , n222836 , n222837 , n222838 , 
 n222839 , n222840 , n222841 , n222842 , n222843 , n222844 , n222845 , n222846 , n222847 , n222848 , 
 n222849 , n222850 , n222851 , n222852 , n222853 , n222854 , n222855 , n222856 , n222857 , n222858 , 
 n222859 , n222860 , n222861 , n222862 , n222863 , n222864 , n222865 , n222866 , n222867 , n222868 , 
 n222869 , n222870 , n222871 , n222872 , n222873 , n222874 , n222875 , n222876 , n222877 , n222878 , 
 n222879 , n222880 , n222881 , n222882 , n222883 , n222884 , n222885 , n222886 , n222887 , n222888 , 
 n222889 , n222890 , n222891 , n222892 , n222893 , n222894 , n222895 , n222896 , n222897 , n222898 , 
 n222899 , n222900 , n222901 , n222902 , n222903 , n222904 , n222905 , n222906 , n222907 , n222908 , 
 n222909 , n222910 , n222911 , n222912 , n222913 , n222914 , n222915 , n222916 , n222917 , n222918 , 
 n222919 , n222920 , n222921 , n222922 , n222923 , n222924 , n222925 , n222926 , n222927 , n222928 , 
 n222929 , n222930 , n222931 , n222932 , n222933 , n222934 , n222935 , n222936 , n222937 , n222938 , 
 n222939 , n222940 , n222941 , n222942 , n222943 , n222944 , n222945 , n222946 , n222947 , n222948 , 
 n222949 , n222950 , n222951 , n222952 , n222953 , n222954 , n222955 , n222956 , n222957 , n222958 , 
 n222959 , n222960 , n222961 , n222962 , n222963 , n222964 , n222965 , n222966 , n222967 , n222968 , 
 n222969 , n222970 , n222971 , n222972 , n222973 , n222974 , n222975 , n222976 , n222977 , n222978 , 
 n222979 , n222980 , n222981 , n222982 , n222983 , n222984 , n222985 , n222986 , n222987 , n222988 , 
 n222989 , n222990 , n222991 , n222992 , n222993 , n222994 , n222995 , n222996 , n222997 , n222998 , 
 n222999 , n223000 , n223001 , n223002 , n223003 , n223004 , n223005 , n223006 , n223007 , n223008 , 
 n223009 , n223010 , n223011 , n223012 , n223013 , n223014 , n223015 , n223016 , n223017 , n223018 , 
 n223019 , n223020 , n223021 , n223022 , n223023 , n223024 , n223025 , n223026 , n223027 , n223028 , 
 n223029 , n223030 , n223031 , n223032 , n223033 , n223034 , n223035 , n223036 , n223037 , n223038 , 
 n223039 , n223040 , n223041 , n223042 , n223043 , n223044 , n223045 , n223046 , n223047 , n223048 , 
 n223049 , n223050 , n223051 , n223052 , n223053 , n223054 , n223055 , n223056 , n223057 , n223058 , 
 n223059 , n223060 , n223061 , n223062 , n223063 , n223064 , n223065 , n223066 , n223067 , n223068 , 
 n223069 , n223070 , n223071 , n223072 , n223073 , n223074 , n223075 , n223076 , n223077 , n223078 , 
 n223079 , n223080 , n223081 , n223082 , n223083 , n223084 , n223085 , n223086 , n223087 , n223088 , 
 n223089 , n223090 , n223091 , n223092 , n223093 , n223094 , n223095 , n223096 , n223097 , n223098 , 
 n223099 , n223100 , n223101 , n223102 , n223103 , n223104 , n223105 , n223106 , n223107 , n223108 , 
 n223109 , n223110 , n223111 , n223112 , n223113 , n223114 , n223115 , n223116 , n223117 , n223118 , 
 n223119 , n223120 , n223121 , n223122 , n223123 , n223124 , n223125 , n223126 , n223127 , n223128 , 
 n223129 , n223130 , n223131 , n223132 , n223133 , n223134 , n223135 , n223136 , n223137 , n223138 , 
 n223139 , n223140 , n223141 , n223142 , n223143 , n223144 , n223145 , n223146 , n223147 , n223148 , 
 n223149 , n223150 , n223151 , n223152 , n223153 , n223154 , n223155 , n223156 , n223157 , n223158 , 
 n223159 , n223160 , n223161 , n223162 , n223163 , n223164 , n223165 , n223166 , n223167 , n223168 , 
 n223169 , n223170 , n223171 , n223172 , n223173 , n223174 , n223175 , n223176 , n223177 , n223178 , 
 n223179 , n223180 , n223181 , n223182 , n223183 , n223184 , n223185 , n223186 , n223187 , n223188 , 
 n223189 , n223190 , n223191 , n223192 , n223193 , n223194 , n223195 , n223196 , n223197 , n223198 , 
 n223199 , n223200 , n223201 , n223202 , n223203 , n223204 , n223205 , n223206 , n223207 , n223208 , 
 n223209 , n223210 , n223211 , n223212 , n223213 , n223214 , n223215 , n223216 , n223217 , n223218 , 
 n223219 , n223220 , n223221 , n223222 , n223223 , n223224 , n223225 , n223226 , n223227 , n223228 , 
 n223229 , n223230 , n223231 , n223232 , n223233 , n223234 , n223235 , n223236 , n223237 , n223238 , 
 n223239 , n223240 , n223241 , n223242 , n223243 , n223244 , n223245 , n223246 , n223247 , n223248 , 
 n223249 , n223250 , n223251 , n223252 , n223253 , n223254 , n223255 , n223256 , n223257 , n223258 , 
 n223259 , n223260 , n223261 , n223262 , n223263 , n223264 , n223265 , n223266 , n223267 , n223268 , 
 n223269 , n223270 , n223271 , n223272 , n223273 , n223274 , n223275 , n223276 , n223277 , n223278 , 
 n223279 , n223280 , n223281 , n223282 , n223283 , n223284 , n223285 , n223286 , n223287 , n223288 , 
 n223289 , n223290 , n223291 , n223292 , n223293 , n223294 , n223295 , n223296 , n223297 , n223298 , 
 n223299 , n223300 , n223301 , n223302 , n223303 , n223304 , n223305 , n223306 , n223307 , n223308 , 
 n223309 , n223310 , n223311 , n223312 , n223313 , n223314 , n223315 , n223316 , n223317 , n223318 , 
 n223319 , n223320 , n223321 , n223322 , n223323 , n223324 , n223325 , n223326 , n223327 , n223328 , 
 n223329 , n223330 , n223331 , n223332 , n223333 , n223334 , n223335 , n223336 , n223337 , n223338 , 
 n223339 , n223340 , n223341 , n223342 , n223343 , n223344 , n223345 , n223346 , n223347 , n223348 , 
 n223349 , n223350 , n223351 , n223352 , n223353 , n223354 , n223355 , n223356 , n223357 , n223358 , 
 n223359 , n223360 , n223361 , n223362 , n223363 , n223364 , n223365 , n223366 , n223367 , n223368 , 
 n223369 , n223370 , n223371 , n223372 , n223373 , n223374 , n223375 , n223376 , n223377 , n223378 , 
 n223379 , n223380 , n223381 , n223382 , n223383 , n223384 , n223385 , n223386 , n223387 , n223388 , 
 n223389 , n223390 , n223391 , n223392 , n223393 , n223394 , n223395 , n223396 , n223397 , n223398 , 
 n223399 , n223400 , n223401 , n223402 , n223403 , n223404 , n223405 , n223406 , n223407 , n223408 , 
 n223409 , n223410 , n223411 , n223412 , n223413 , n223414 , n223415 , n223416 , n223417 , n223418 , 
 n223419 , n223420 , n223421 , n223422 , n223423 , n223424 , n223425 , n223426 , n223427 , n223428 , 
 n223429 , n223430 , n223431 , n223432 , n223433 , n223434 , n223435 , n223436 , n223437 , n223438 , 
 n223439 , n223440 , n223441 , n223442 , n223443 , n223444 , n223445 , n223446 , n223447 , n223448 , 
 n223449 , n223450 , n223451 , n223452 , n223453 , n223454 , n223455 , n223456 , n223457 , n223458 , 
 n223459 , n223460 , n223461 , n223462 , n223463 , n223464 , n223465 , n223466 , n223467 , n223468 , 
 n223469 , n223470 , n223471 , n223472 , n223473 , n223474 , n223475 , n223476 , n223477 , n223478 , 
 n223479 , n223480 , n223481 , n223482 , n223483 , n223484 , n223485 , n223486 , n223487 , n223488 , 
 n223489 , n223490 , n223491 , n223492 , n223493 , n223494 , n223495 , n223496 , n223497 , n223498 , 
 n223499 , n223500 , n223501 , n223502 , n223503 , n223504 , n223505 , n223506 , n223507 , n223508 , 
 n223509 , n223510 , n223511 , n223512 , n223513 , n223514 , n223515 , n223516 , n223517 , n223518 , 
 n223519 , n223520 , n223521 , n223522 , n223523 , n223524 , n223525 , n223526 , n223527 , n223528 , 
 n223529 , n223530 , n223531 , n223532 , n223533 , n223534 , n223535 , n223536 , n223537 , n223538 , 
 n223539 , n223540 , n223541 , n223542 , n223543 , n223544 , n223545 , n223546 , n223547 , n223548 , 
 n223549 , n223550 , n223551 , n223552 , n223553 , n223554 , n223555 , n223556 , n223557 , n223558 , 
 n223559 , n223560 , n223561 , n223562 , n223563 , n223564 , n223565 , n223566 , n223567 , n223568 , 
 n223569 , n223570 , n223571 , n223572 , n223573 , n223574 , n223575 , n223576 , n223577 , n223578 , 
 n223579 , n223580 , n223581 , n223582 , n223583 , n223584 , n223585 , n223586 , n223587 , n223588 , 
 n223589 , n223590 , n223591 , n223592 , n223593 , n223594 , n223595 , n223596 , n223597 , n223598 , 
 n223599 , n223600 , n223601 , n223602 , n223603 , n223604 , n223605 , n223606 , n223607 , n223608 , 
 n223609 , n223610 , n223611 , n223612 , n223613 , n223614 , n223615 , n223616 , n223617 , n223618 , 
 n223619 , n223620 , n223621 , n223622 , n223623 , n223624 , n223625 , n223626 , n223627 , n223628 , 
 n223629 , n223630 , n223631 , n223632 , n223633 , n223634 , n223635 , n223636 , n223637 , n223638 , 
 n223639 , n223640 , n223641 , n223642 , n223643 , n223644 , n223645 , n223646 , n223647 , n223648 , 
 n223649 , n223650 , n223651 , n223652 , n223653 , n223654 , n223655 , n223656 , n223657 , n223658 , 
 n223659 , n223660 , n223661 , n223662 , n223663 , n223664 , n223665 , n223666 , n223667 , n223668 , 
 n223669 , n223670 , n223671 , n223672 , n223673 , n223674 , n223675 , n223676 , n223677 , n223678 , 
 n223679 , n223680 , n223681 , n223682 , n223683 , n223684 , n223685 , n223686 , n223687 , n223688 , 
 n223689 , n223690 , n223691 , n223692 , n223693 , n223694 , n223695 , n223696 , n223697 , n223698 , 
 n223699 , n223700 , n223701 , n223702 , n223703 , n223704 , n223705 , n223706 , n223707 , n223708 , 
 n223709 , n223710 , n223711 , n223712 , n223713 , n223714 , n223715 , n223716 , n223717 , n223718 , 
 n223719 , n223720 , n223721 , n223722 , n223723 , n223724 , n223725 , n223726 , n223727 , n223728 , 
 n223729 , n223730 , n223731 , n223732 , n223733 , n223734 , n223735 , n223736 , n223737 , n223738 , 
 n223739 , n223740 , n223741 , n223742 , n223743 , n223744 , n223745 , n223746 , n223747 , n223748 , 
 n223749 , n223750 , n223751 , n223752 , n223753 , n223754 , n223755 , n223756 , n223757 , n223758 , 
 n223759 , n223760 , n223761 , n223762 , n223763 , n223764 , n223765 , n223766 , n223767 , n223768 , 
 n223769 , n223770 , n223771 , n223772 , n223773 , n223774 , n223775 , n223776 , n223777 , n223778 , 
 n223779 , n223780 , n223781 , n223782 , n223783 , n223784 , n223785 , n223786 , n223787 , n223788 , 
 n223789 , n223790 , n223791 , n223792 , n223793 , n223794 , n223795 , n223796 , n223797 , n223798 , 
 n223799 , n223800 , n223801 , n223802 , n223803 , n223804 , n223805 , n223806 , n223807 , n223808 , 
 n223809 , n223810 , n223811 , n223812 , n223813 , n223814 , n223815 , n223816 , n223817 , n223818 , 
 n223819 , n223820 , n223821 , n223822 , n223823 , n223824 , n223825 , n223826 , n223827 , n223828 , 
 n223829 , n223830 , n223831 , n223832 , n223833 , n223834 , n223835 , n223836 , n223837 , n223838 , 
 n223839 , n223840 , n223841 , n223842 , n223843 , n223844 , n223845 , n223846 , n223847 , n223848 , 
 n223849 , n223850 , n223851 , n223852 , n223853 , n223854 , n223855 , n223856 , n223857 , n223858 , 
 n223859 , n223860 , n223861 , n223862 , n223863 , n223864 , n223865 , n223866 , n223867 , n223868 , 
 n223869 , n223870 , n223871 , n223872 , n223873 , n223874 , n223875 , n223876 , n223877 , n223878 , 
 n223879 , n223880 , n223881 , n223882 , n223883 , n223884 , n223885 , n223886 , n223887 , n223888 , 
 n223889 , n223890 , n223891 , n223892 , n223893 , n223894 , n223895 , n223896 , n223897 , n223898 , 
 n223899 , n223900 , n223901 , n223902 , n223903 , n223904 , n223905 , n223906 , n223907 , n223908 , 
 n223909 , n223910 , n223911 , n223912 , n223913 , n223914 , n223915 , n223916 , n223917 , n223918 , 
 n223919 , n223920 , n223921 , n223922 , n223923 , n223924 , n223925 , n223926 , n223927 , n223928 , 
 n223929 , n223930 , n223931 , n223932 , n223933 , n223934 , n223935 , n223936 , n223937 , n223938 , 
 n223939 , n223940 , n223941 , n223942 , n223943 , n223944 , n223945 , n223946 , n223947 , n223948 , 
 n223949 , n223950 , n223951 , n223952 , n223953 , n223954 , n223955 , n223956 , n223957 , n223958 , 
 n223959 , n223960 , n223961 , n223962 , n223963 , n223964 , n223965 , n223966 , n223967 , n223968 , 
 n223969 , n223970 , n223971 , n223972 , n223973 , n223974 , n223975 , n223976 , n223977 , n223978 , 
 n223979 , n223980 , n223981 , n223982 , n223983 , n223984 , n223985 , n223986 , n223987 , n223988 , 
 n223989 , n223990 , n223991 , n223992 , n223993 , n223994 , n223995 , n223996 , n223997 , n223998 , 
 n223999 , n224000 , n224001 , n224002 , n224003 , n224004 , n224005 , n224006 , n224007 , n224008 , 
 n224009 , n224010 , n224011 , n224012 , n224013 , n224014 , n224015 , n224016 , n224017 , n224018 , 
 n224019 , n224020 , n224021 , n224022 , n224023 , n224024 , n224025 , n224026 , n224027 , n224028 , 
 n224029 , n224030 , n224031 , n224032 , n224033 , n224034 , n224035 , n224036 , n224037 , n224038 , 
 n224039 , n224040 , n224041 , n224042 , n224043 , n224044 , n224045 , n224046 , n224047 , n224048 , 
 n224049 , n224050 , n224051 , n224052 , n224053 , n224054 , n224055 , n224056 , n224057 , n224058 , 
 n224059 , n224060 , n224061 , n224062 , n224063 , n224064 , n224065 , n224066 , n224067 , n224068 , 
 n224069 , n224070 , n224071 , n224072 , n224073 , n224074 , n224075 , n224076 , n224077 , n224078 , 
 n224079 , n224080 , n224081 , n224082 , n224083 , n224084 , n224085 , n224086 , n224087 , n224088 , 
 n224089 , n224090 , n224091 , n224092 , n224093 , n224094 , n224095 , n224096 , n224097 , n224098 , 
 n224099 , n224100 , n224101 , n224102 , n224103 , n224104 , n224105 , n224106 , n224107 , n224108 , 
 n224109 , n224110 , n224111 , n224112 , n224113 , n224114 , n224115 , n224116 , n224117 , n224118 , 
 n224119 , n224120 , n224121 , n224122 , n224123 , n224124 , n224125 , n224126 , n224127 , n224128 , 
 n224129 , n224130 , n224131 , n224132 , n224133 , n224134 , n224135 , n224136 , n224137 , n224138 , 
 n224139 , n224140 , n224141 , n224142 , n224143 , n224144 , n224145 , n224146 , n224147 , n224148 , 
 n224149 , n224150 , n224151 , n224152 , n224153 , n224154 , n224155 , n224156 , n224157 , n224158 , 
 n224159 , n224160 , n224161 , n224162 , n224163 , n224164 , n224165 , n224166 , n224167 , n224168 , 
 n224169 , n224170 , n224171 , n224172 , n224173 , n224174 , n224175 , n224176 , n224177 , n224178 , 
 n224179 , n224180 , n224181 , n224182 , n224183 , n224184 , n224185 , n224186 , n224187 , n224188 , 
 n224189 , n224190 , n224191 , n224192 , n224193 , n224194 , n224195 , n224196 , n224197 , n224198 , 
 n224199 , n224200 , n224201 , n224202 , n224203 , n224204 , n224205 , n224206 , n224207 , n224208 , 
 n224209 , n224210 , n224211 , n224212 , n224213 , n224214 , n224215 , n224216 , n224217 , n224218 , 
 n224219 , n224220 , n224221 , n224222 , n224223 , n224224 , n224225 , n224226 , n224227 , n224228 , 
 n224229 , n224230 , n224231 , n224232 , n224233 , n224234 , n224235 , n224236 , n224237 , n224238 , 
 n224239 , n224240 , n224241 , n224242 , n224243 , n224244 , n224245 , n224246 , n224247 , n224248 , 
 n224249 , n224250 , n224251 , n224252 , n224253 , n224254 , n224255 , n224256 , n224257 , n224258 , 
 n224259 , n224260 , n224261 , n224262 , n224263 , n224264 , n224265 , n224266 , n224267 , n224268 , 
 n224269 , n224270 , n224271 , n224272 , n224273 , n224274 , n224275 , n224276 , n224277 , n224278 , 
 n224279 , n224280 , n224281 , n224282 , n224283 , n224284 , n224285 , n224286 , n224287 , n224288 , 
 n224289 , n224290 , n224291 , n224292 , n224293 , n224294 , n224295 , n224296 , n224297 , n224298 , 
 n224299 , n224300 , n224301 , n224302 , n224303 , n224304 , n224305 , n224306 , n224307 , n224308 , 
 n224309 , n224310 , n224311 , n224312 , n224313 , n224314 , n224315 , n224316 , n224317 , n224318 , 
 n224319 , n224320 , n224321 , n224322 , n224323 , n224324 , n224325 , n224326 , n224327 , n224328 , 
 n224329 , n224330 , n224331 , n224332 , n224333 , n224334 , n224335 , n224336 , n224337 , n224338 , 
 n224339 , n224340 , n224341 , n224342 , n224343 , n224344 , n224345 , n224346 , n224347 , n224348 , 
 n224349 , n224350 , n224351 , n224352 , n224353 , n224354 , n224355 , n224356 , n224357 , n224358 , 
 n224359 , n224360 , n224361 , n224362 , n224363 , n224364 , n224365 , n224366 , n224367 , n224368 , 
 n224369 , n224370 , n224371 , n224372 , n224373 , n224374 , n224375 , n224376 , n224377 , n224378 , 
 n224379 , n224380 , n224381 , n224382 , n224383 , n224384 , n224385 , n224386 , n224387 , n224388 , 
 n224389 , n224390 , n224391 , n224392 , n224393 , n224394 , n224395 , n224396 , n224397 , n224398 , 
 n224399 , n224400 , n224401 , n224402 , n224403 , n224404 , n224405 , n224406 , n224407 , n224408 , 
 n224409 , n224410 , n224411 , n224412 , n224413 , n224414 , n224415 , n224416 , n224417 , n224418 , 
 n224419 , n224420 , n224421 , n224422 , n224423 , n224424 , n224425 , n224426 , n224427 , n224428 , 
 n224429 , n224430 , n224431 , n224432 , n224433 , n224434 , n224435 , n224436 , n224437 , n224438 , 
 n224439 , n224440 , n224441 , n224442 , n224443 , n224444 , n224445 , n224446 , n224447 , n224448 , 
 n224449 , n224450 , n224451 , n224452 , n224453 , n224454 , n224455 , n224456 , n224457 , n224458 , 
 n224459 , n224460 , n224461 , n224462 , n224463 , n224464 , n224465 , n224466 , n224467 , n224468 , 
 n224469 , n224470 , n224471 , n224472 , n224473 , n224474 , n224475 , n224476 , n224477 , n224478 , 
 n224479 , n224480 , n224481 , n224482 , n224483 , n224484 , n224485 , n224486 , n224487 , n224488 , 
 n224489 , n224490 , n224491 , n224492 , n224493 , n224494 , n224495 , n224496 , n224497 , n224498 , 
 n224499 , n224500 , n224501 , n224502 , n224503 , n224504 , n224505 , n224506 , n224507 , n224508 , 
 n224509 , n224510 , n224511 , n224512 , n224513 , n224514 , n224515 , n224516 , n224517 , n224518 , 
 n224519 , n224520 , n224521 , n224522 , n224523 , n224524 , n224525 , n224526 , n224527 , n224528 , 
 n224529 , n224530 , n224531 , n224532 , n224533 , n224534 , n224535 , n224536 , n224537 , n224538 , 
 n224539 , n224540 , n224541 , n224542 , n224543 , n224544 , n224545 , n224546 , n224547 , n224548 , 
 n224549 , n224550 , n224551 , n224552 , n224553 , n224554 , n224555 , n224556 , n224557 , n224558 , 
 n224559 , n224560 , n224561 , n224562 , n224563 , n224564 , n224565 , n224566 , n224567 , n224568 , 
 n224569 , n224570 , n224571 , n224572 , n224573 , n224574 , n224575 , n224576 , n224577 , n224578 , 
 n224579 , n224580 , n224581 , n224582 , n224583 , n224584 , n224585 , n224586 , n224587 , n224588 , 
 n224589 , n224590 , n224591 , n224592 , n224593 , n224594 , n224595 , n224596 , n224597 , n224598 , 
 n224599 , n224600 , n224601 , n224602 , n224603 , n224604 , n224605 , n224606 , n224607 , n224608 , 
 n224609 , n224610 , n224611 , n224612 , n224613 , n224614 , n224615 , n224616 , n224617 , n224618 , 
 n224619 , n224620 , n224621 , n224622 , n224623 , n224624 , n224625 , n224626 , n224627 , n224628 , 
 n224629 , n224630 , n224631 , n224632 , n224633 , n224634 , n224635 , n224636 , n224637 , n224638 , 
 n224639 , n224640 , n224641 , n224642 , n224643 , n224644 , n224645 , n224646 , n224647 , n224648 , 
 n224649 , n224650 , n224651 , n224652 , n224653 , n224654 , n224655 , n224656 , n224657 , n224658 , 
 n224659 , n224660 , n224661 , n224662 , n224663 , n224664 , n224665 , n224666 , n224667 , n224668 , 
 n224669 , n224670 , n224671 , n224672 , n224673 , n224674 , n224675 , n224676 , n224677 , n224678 , 
 n224679 , n224680 , n224681 , n224682 , n224683 , n224684 , n224685 , n224686 , n224687 , n224688 , 
 n224689 , n224690 , n224691 , n224692 , n224693 , n224694 , n224695 , n224696 , n224697 , n224698 , 
 n224699 , n224700 , n224701 , n224702 , n224703 , n224704 , n224705 , n224706 , n224707 , n224708 , 
 n224709 , n224710 , n224711 , n224712 , n224713 , n224714 , n224715 , n224716 , n224717 , n224718 , 
 n224719 , n224720 , n224721 , n224722 , n224723 , n224724 , n224725 , n224726 , n224727 , n224728 , 
 n224729 , n224730 , n224731 , n224732 , n224733 , n224734 , n224735 , n224736 , n224737 , n224738 , 
 n224739 , n224740 , n224741 , n224742 , n224743 , n224744 , n224745 , n224746 , n224747 , n224748 , 
 n224749 , n224750 , n224751 , n224752 , n224753 , n224754 , n224755 , n224756 , n224757 , n224758 , 
 n224759 , n224760 , n224761 , n224762 , n224763 , n224764 , n224765 , n224766 , n224767 , n224768 , 
 n224769 , n224770 , n224771 , n224772 , n224773 , n224774 , n224775 , n224776 , n224777 , n224778 , 
 n224779 , n224780 , n224781 , n224782 , n224783 , n224784 , n224785 , n224786 , n224787 , n224788 , 
 n224789 , n224790 , n224791 , n224792 , n224793 , n224794 , n224795 , n224796 , n224797 , n224798 , 
 n224799 , n224800 , n224801 , n224802 , n224803 , n224804 , n224805 , n224806 , n224807 , n224808 , 
 n224809 , n224810 , n224811 , n224812 , n224813 , n224814 , n224815 , n224816 , n224817 , n224818 , 
 n224819 , n224820 , n224821 , n224822 , n224823 , n224824 , n224825 , n224826 , n224827 , n224828 , 
 n224829 , n224830 , n224831 , n224832 , n224833 , n224834 , n224835 , n224836 , n224837 , n224838 , 
 n224839 , n224840 , n224841 , n224842 , n224843 , n224844 , n224845 , n224846 , n224847 , n224848 , 
 n224849 , n224850 , n224851 , n224852 , n224853 , n224854 , n224855 , n224856 , n224857 , n224858 , 
 n224859 , n224860 , n224861 , n224862 , n224863 , n224864 , n224865 , n224866 , n224867 , n224868 , 
 n224869 , n224870 , n224871 , n224872 , n224873 , n224874 , n224875 , n224876 , n224877 , n224878 , 
 n224879 , n224880 , n224881 , n224882 , n224883 , n224884 , n224885 , n224886 , n224887 , n224888 , 
 n224889 , n224890 , n224891 , n224892 , n224893 , n224894 , n224895 , n224896 , n224897 , n224898 , 
 n224899 , n224900 , n224901 , n224902 , n224903 , n224904 , n224905 , n224906 , n224907 , n224908 , 
 n224909 , n224910 , n224911 , n224912 , n224913 , n224914 , n224915 , n224916 , n224917 , n224918 , 
 n224919 , n224920 , n224921 , n224922 , n224923 , n224924 , n224925 , n224926 , n224927 , n224928 , 
 n224929 , n224930 , n224931 , n224932 , n224933 , n224934 , n224935 , n224936 , n224937 , n224938 , 
 n224939 , n224940 , n224941 , n224942 , n224943 , n224944 , n224945 , n224946 , n224947 , n224948 , 
 n224949 , n224950 , n224951 , n224952 , n224953 , n224954 , n224955 , n224956 , n224957 , n224958 , 
 n224959 , n224960 , n224961 , n224962 , n224963 , n224964 , n224965 , n224966 , n224967 , n224968 , 
 n224969 , n224970 , n224971 , n224972 , n224973 , n224974 , n224975 , n224976 , n224977 , n224978 , 
 n224979 , n224980 , n224981 , n224982 , n224983 , n224984 , n224985 , n224986 , n224987 , n224988 , 
 n224989 , n224990 , n224991 , n224992 , n224993 , n224994 , n224995 , n224996 , n224997 , n224998 , 
 n224999 , n225000 , n225001 , n225002 , n225003 , n225004 , n225005 , n225006 , n225007 , n225008 , 
 n225009 , n225010 , n225011 , n225012 , n225013 , n225014 , n225015 , n225016 , n225017 , n225018 , 
 n225019 , n225020 , n225021 , n225022 , n225023 , n225024 , n225025 , n225026 , n225027 , n225028 , 
 n225029 , n225030 , n225031 , n225032 , n225033 , n225034 , n225035 , n225036 , n225037 , n225038 , 
 n225039 , n225040 , n225041 , n225042 , n225043 , n225044 , n225045 , n225046 , n225047 , n225048 , 
 n225049 , n225050 , n225051 , n225052 , n225053 , n225054 , n225055 , n225056 , n225057 , n225058 , 
 n225059 , n225060 , n225061 , n225062 , n225063 , n225064 , n225065 , n225066 , n225067 , n225068 , 
 n225069 , n225070 , n225071 , n225072 , n225073 , n225074 , n225075 , n225076 , n225077 , n225078 , 
 n225079 , n225080 , n225081 , n225082 , n225083 , n225084 , n225085 , n225086 , n225087 , n225088 , 
 n225089 , n225090 , n225091 , n225092 , n225093 , n225094 , n225095 , n225096 , n225097 , n225098 , 
 n225099 , n225100 , n225101 , n225102 , n225103 , n225104 , n225105 , n225106 , n225107 , n225108 , 
 n225109 , n225110 , n225111 , n225112 , n225113 , n225114 , n225115 , n225116 , n225117 , n225118 , 
 n225119 , n225120 , n225121 , n225122 , n225123 , n225124 , n225125 , n225126 , n225127 , n225128 , 
 n225129 , n225130 , n225131 , n225132 , n225133 , n225134 , n225135 , n225136 , n225137 , n225138 , 
 n225139 , n225140 , n225141 , n225142 , n225143 , n225144 , n225145 , n225146 , n225147 , n225148 , 
 n225149 , n225150 , n225151 , n225152 , n225153 , n225154 , n225155 , n225156 , n225157 , n225158 , 
 n225159 , n225160 , n225161 , n225162 , n225163 , n225164 , n225165 , n225166 , n225167 , n225168 , 
 n225169 , n225170 , n225171 , n225172 , n225173 , n225174 , n225175 , n225176 , n225177 , n225178 , 
 n225179 , n225180 , n225181 , n225182 , n225183 , n225184 , n225185 , n225186 , n225187 , n225188 , 
 n225189 , n225190 , n225191 , n225192 , n225193 , n225194 , n225195 , n225196 , n225197 , n225198 , 
 n225199 , n225200 , n225201 , n225202 , n225203 , n225204 , n225205 , n225206 , n225207 , n225208 , 
 n225209 , n225210 , n225211 , n225212 , n225213 , n225214 , n225215 , n225216 , n225217 , n225218 , 
 n225219 , n225220 , n225221 , n225222 , n225223 , n225224 , n225225 , n225226 , n225227 , n225228 , 
 n225229 , n225230 , n225231 , n225232 , n225233 , n225234 , n225235 , n225236 , n225237 , n225238 , 
 n225239 , n225240 , n225241 , n225242 , n225243 , n225244 , n225245 , n225246 , n225247 , n225248 , 
 n225249 , n225250 , n225251 , n225252 , n225253 , n225254 , n225255 , n225256 , n225257 , n225258 , 
 n225259 , n225260 , n225261 , n225262 , n225263 , n225264 , n225265 , n225266 , n225267 , n225268 , 
 n225269 , n225270 , n225271 , n225272 , n225273 , n225274 , n225275 , n225276 , n225277 , n225278 , 
 n225279 , n225280 , n225281 , n225282 , n225283 , n225284 , n225285 , n225286 , n225287 , n225288 , 
 n225289 , n225290 , n225291 , n225292 , n225293 , n225294 , n225295 , n225296 , n225297 , n225298 , 
 n225299 , n225300 , n225301 , n225302 , n225303 , n225304 , n225305 , n225306 , n225307 , n225308 , 
 n225309 , n225310 , n225311 , n225312 , n225313 , n225314 , n225315 , n225316 , n225317 , n225318 , 
 n225319 , n225320 , n225321 , n225322 , n225323 , n225324 , n225325 , n225326 , n225327 , n225328 , 
 n225329 , n225330 , n225331 , n225332 , n225333 , n225334 , n225335 , n225336 , n225337 , n225338 , 
 n225339 , n225340 , n225341 , n225342 , n225343 , n225344 , n225345 , n225346 , n225347 , n225348 , 
 n225349 , n225350 , n225351 , n225352 , n225353 , n225354 , n225355 , n225356 , n225357 , n225358 , 
 n225359 , n225360 , n225361 , n225362 , n225363 , n225364 , n225365 , n225366 , n225367 , n225368 , 
 n225369 , n225370 , n225371 , n225372 , n225373 , n225374 , n225375 , n225376 , n225377 , n225378 , 
 n225379 , n225380 , n225381 , n225382 , n225383 , n225384 , n225385 , n225386 , n225387 , n225388 , 
 n225389 , n225390 , n225391 , n225392 , n225393 , n225394 , n225395 , n225396 , n225397 , n225398 , 
 n225399 , n225400 , n225401 , n225402 , n225403 , n225404 , n225405 , n225406 , n225407 , n225408 , 
 n225409 , n225410 , n225411 , n225412 , n225413 , n225414 , n225415 , n225416 , n225417 , n225418 , 
 n225419 , n225420 , n225421 , n225422 , n225423 , n225424 , n225425 , n225426 , n225427 , n225428 , 
 n225429 , n225430 , n225431 , n225432 , n225433 , n225434 , n225435 , n225436 , n225437 , n225438 , 
 n225439 , n225440 , n225441 , n225442 , n225443 , n225444 , n225445 , n225446 , n225447 , n225448 , 
 n225449 , n225450 , n225451 , n225452 , n225453 , n225454 , n225455 , n225456 , n225457 , n225458 , 
 n225459 , n225460 , n225461 , n225462 , n225463 , n225464 , n225465 , n225466 , n225467 , n225468 , 
 n225469 , n225470 , n225471 , n225472 , n225473 , n225474 , n225475 , n225476 , n225477 , n225478 , 
 n225479 , n225480 , n225481 , n225482 , n225483 , n225484 , n225485 , n225486 , n225487 , n225488 , 
 n225489 , n225490 , n225491 , n225492 , n225493 , n225494 , n225495 , n225496 , n225497 , n225498 , 
 n225499 , n225500 , n225501 , n225502 , n225503 , n225504 , n225505 , n225506 , n225507 , n225508 , 
 n225509 , n225510 , n225511 , n225512 , n225513 , n225514 , n225515 , n225516 , n225517 , n225518 , 
 n225519 , n225520 , n225521 , n225522 , n225523 , n225524 , n225525 , n225526 , n225527 , n225528 , 
 n225529 , n225530 , n225531 , n225532 , n225533 , n225534 , n225535 , n225536 , n225537 , n225538 , 
 n225539 , n225540 , n225541 , n225542 , n225543 , n225544 , n225545 , n225546 , n225547 , n225548 , 
 n225549 , n225550 , n225551 , n225552 , n225553 , n225554 , n225555 , n225556 , n225557 , n225558 , 
 n225559 , n225560 , n225561 , n225562 , n225563 , n225564 , n225565 , n225566 , n225567 , n225568 , 
 n225569 , n225570 , n225571 , n225572 , n225573 , n225574 , n225575 , n225576 , n225577 , n225578 , 
 n225579 , n225580 , n225581 , n225582 , n225583 , n225584 , n225585 , n225586 , n225587 , n225588 , 
 n225589 , n225590 , n225591 , n225592 , n225593 , n225594 , n225595 , n225596 , n225597 , n225598 , 
 n225599 , n225600 , n225601 , n225602 , n225603 , n225604 , n225605 , n225606 , n225607 , n225608 , 
 n225609 , n225610 , n225611 , n225612 , n225613 , n225614 , n225615 , n225616 , n225617 , n225618 , 
 n225619 , n225620 , n225621 , n225622 , n225623 , n225624 , n225625 , n225626 , n225627 , n225628 , 
 n225629 , n225630 , n225631 , n225632 , n225633 , n225634 , n225635 , n225636 , n225637 , n225638 , 
 n225639 , n225640 , n225641 , n225642 , n225643 , n225644 , n225645 , n225646 , n225647 , n225648 , 
 n225649 , n225650 , n225651 , n225652 , n225653 , n225654 , n225655 , n225656 , n225657 , n225658 , 
 n225659 , n225660 , n225661 , n225662 , n225663 , n225664 , n225665 , n225666 , n225667 , n225668 , 
 n225669 , n225670 , n225671 , n225672 , n225673 , n225674 , n225675 , n225676 , n225677 , n225678 , 
 n225679 , n225680 , n225681 , n225682 , n225683 , n225684 , n225685 , n225686 , n225687 , n225688 , 
 n225689 , n225690 , n225691 , n225692 , n225693 , n225694 , n225695 , n225696 , n225697 , n225698 , 
 n225699 , n225700 , n225701 , n225702 , n225703 , n225704 , n225705 , n225706 , n225707 , n225708 , 
 n225709 , n225710 , n225711 , n225712 , n225713 , n225714 , n225715 , n225716 , n225717 , n225718 , 
 n225719 , n225720 , n225721 , n225722 , n225723 , n225724 , n225725 , n225726 , n225727 , n225728 , 
 n225729 , n225730 , n225731 , n225732 , n225733 , n225734 , n225735 , n225736 , n225737 , n225738 , 
 n225739 , n225740 , n225741 , n225742 , n225743 , n225744 , n225745 , n225746 , n225747 , n225748 , 
 n225749 , n225750 , n225751 , n225752 , n225753 , n225754 , n225755 , n225756 , n225757 , n225758 , 
 n225759 , n225760 , n225761 , n225762 , n225763 , n225764 , n225765 , n225766 , n225767 , n225768 , 
 n225769 , n225770 , n225771 , n225772 , n225773 , n225774 , n225775 , n225776 , n225777 , n225778 , 
 n225779 , n225780 , n225781 , n225782 , n225783 , n225784 , n225785 , n225786 , n225787 , n225788 , 
 n225789 , n225790 , n225791 , n225792 , n225793 , n225794 , n225795 , n225796 , n225797 , n225798 , 
 n225799 , n225800 , n225801 , n225802 , n225803 , n225804 , n225805 , n225806 , n225807 , n225808 , 
 n225809 , n225810 , n225811 , n225812 , n225813 , n225814 , n225815 , n225816 , n225817 , n225818 , 
 n225819 , n225820 , n225821 , n225822 , n225823 , n225824 , n225825 , n225826 , n225827 , n225828 , 
 n225829 , n225830 , n225831 , n225832 , n225833 , n225834 , n225835 , n225836 , n225837 , n225838 , 
 n225839 , n225840 , n225841 , n225842 , n225843 , n225844 , n225845 , n225846 , n225847 , n225848 , 
 n225849 , n225850 , n225851 , n225852 , n225853 , n225854 , n225855 , n225856 , n225857 , n225858 , 
 n225859 , n225860 , n225861 , n225862 , n225863 , n225864 , n225865 , n225866 , n225867 , n225868 , 
 n225869 , n225870 , n225871 , n225872 , n225873 , n225874 , n225875 , n225876 , n225877 , n225878 , 
 n225879 , n225880 , n225881 , n225882 , n225883 , n225884 , n225885 , n225886 , n225887 , n225888 , 
 n225889 , n225890 , n225891 , n225892 , n225893 , n225894 , n225895 , n225896 , n225897 , n225898 , 
 n225899 , n225900 , n225901 , n225902 , n225903 , n225904 , n225905 , n225906 , n225907 , n225908 , 
 n225909 , n225910 , n225911 , n225912 , n225913 , n225914 , n225915 , n225916 , n225917 , n225918 , 
 n225919 , n225920 , n225921 , n225922 , n225923 , n225924 , n225925 , n225926 , n225927 , n225928 , 
 n225929 , n225930 , n225931 , n225932 , n225933 , n225934 , n225935 , n225936 , n225937 , n225938 , 
 n225939 , n225940 , n225941 , n225942 , n225943 , n225944 , n225945 , n225946 , n225947 , n225948 , 
 n225949 , n225950 , n225951 , n225952 , n225953 , n225954 , n225955 , n225956 , n225957 , n225958 , 
 n225959 , n225960 , n225961 , n225962 , n225963 , n225964 , n225965 , n225966 , n225967 , n225968 , 
 n225969 , n225970 , n225971 , n225972 , n225973 , n225974 , n225975 , n225976 , n225977 , n225978 , 
 n225979 , n225980 , n225981 , n225982 , n225983 , n225984 , n225985 , n225986 , n225987 , n225988 , 
 n225989 , n225990 , n225991 , n225992 , n225993 , n225994 , n225995 , n225996 , n225997 , n225998 , 
 n225999 , n226000 , n226001 , n226002 , n226003 , n226004 , n226005 , n226006 , n226007 , n226008 , 
 n226009 , n226010 , n226011 , n226012 , n226013 , n226014 , n226015 , n226016 , n226017 , n226018 , 
 n226019 , n226020 , n226021 , n226022 , n226023 , n226024 , n226025 , n226026 , n226027 , n226028 , 
 n226029 , n226030 , n226031 , n226032 , n226033 , n226034 , n226035 , n226036 , n226037 , n226038 , 
 n226039 , n226040 , n226041 , n226042 , n226043 , n226044 , n226045 , n226046 , n226047 , n226048 , 
 n226049 , n226050 , n226051 , n226052 , n226053 , n226054 , n226055 , n226056 , n226057 , n226058 , 
 n226059 , n226060 , n226061 , n226062 , n226063 , n226064 , n226065 , n226066 , n226067 , n226068 , 
 n226069 , n226070 , n226071 , n226072 , n226073 , n226074 , n226075 , n226076 , n226077 , n226078 , 
 n226079 , n226080 , n226081 , n226082 , n226083 , n226084 , n226085 , n226086 , n226087 , n226088 , 
 n226089 , n226090 , n226091 , n226092 , n226093 , n226094 , n226095 , n226096 , n226097 , n226098 , 
 n226099 , n226100 , n226101 , n226102 , n226103 , n226104 , n226105 , n226106 , n226107 , n226108 , 
 n226109 , n226110 , n226111 , n226112 , n226113 , n226114 , n226115 , n226116 , n226117 , n226118 , 
 n226119 , n226120 , n226121 , n226122 , n226123 , n226124 , n226125 , n226126 , n226127 , n226128 , 
 n226129 , n226130 , n226131 , n226132 , n226133 , n226134 , n226135 , n226136 , n226137 , n226138 , 
 n226139 , n226140 , n226141 , n226142 , n226143 , n226144 , n226145 , n226146 , n226147 , n226148 , 
 n226149 , n226150 , n226151 , n226152 , n226153 , n226154 , n226155 , n226156 , n226157 , n226158 , 
 n226159 , n226160 , n226161 , n226162 , n226163 , n226164 , n226165 , n226166 , n226167 , n226168 , 
 n226169 , n226170 , n226171 , n226172 , n226173 , n226174 , n226175 , n226176 , n226177 , n226178 , 
 n226179 , n226180 , n226181 , n226182 , n226183 , n226184 , n226185 , n226186 , n226187 , n226188 , 
 n226189 , n226190 , n226191 , n226192 , n226193 , n226194 , n226195 , n226196 , n226197 , n226198 , 
 n226199 , n226200 , n226201 , n226202 , n226203 , n226204 , n226205 , n226206 , n226207 , n226208 , 
 n226209 , n226210 , n226211 , n226212 , n226213 , n226214 , n226215 , n226216 , n226217 , n226218 , 
 n226219 , n226220 , n226221 , n226222 , n226223 , n226224 , n226225 , n226226 , n226227 , n226228 , 
 n226229 , n226230 , n226231 , n226232 , n226233 , n226234 , n226235 , n226236 , n226237 , n226238 , 
 n226239 , n226240 , n226241 , n226242 , n226243 , n226244 , n226245 , n226246 , n226247 , n226248 , 
 n226249 , n226250 , n226251 , n226252 , n226253 , n226254 , n226255 , n226256 , n226257 , n226258 , 
 n226259 , n226260 , n226261 , n226262 , n226263 , n226264 , n226265 , n226266 , n226267 , n226268 , 
 n226269 , n226270 , n226271 , n226272 , n226273 , n226274 , n226275 , n226276 , n226277 , n226278 , 
 n226279 , n226280 , n226281 , n226282 , n226283 , n226284 , n226285 , n226286 , n226287 , n226288 , 
 n226289 , n226290 , n226291 , n226292 , n226293 , n226294 , n226295 , n226296 , n226297 , n226298 , 
 n226299 , n226300 , n226301 , n226302 , n226303 , n226304 , n226305 , n226306 , n226307 , n226308 , 
 n226309 , n226310 , n226311 , n226312 , n226313 , n226314 , n226315 , n226316 , n226317 , n226318 , 
 n226319 , n226320 , n226321 , n226322 , n226323 , n226324 , n226325 , n226326 , n226327 , n226328 , 
 n226329 , n226330 , n226331 , n226332 , n226333 , n226334 , n226335 , n226336 , n226337 , n226338 , 
 n226339 , n226340 , n226341 , n226342 , n226343 , n226344 , n226345 , n226346 , n226347 , n226348 , 
 n226349 , n226350 , n226351 , n226352 , n226353 , n226354 , n226355 , n226356 , n226357 , n226358 , 
 n226359 , n226360 , n226361 , n226362 , n226363 , n226364 , n226365 , n226366 , n226367 , n226368 , 
 n226369 , n226370 , n226371 , n226372 , n226373 , n226374 , n226375 , n226376 , n226377 , n226378 , 
 n226379 , n226380 , n226381 , n226382 , n226383 , n226384 , n226385 , n226386 , n226387 , n226388 , 
 n226389 , n226390 , n226391 , n226392 , n226393 , n226394 , n226395 , n226396 , n226397 , n226398 , 
 n226399 , n226400 , n226401 , n226402 , n226403 , n226404 , n226405 , n226406 , n226407 , n226408 , 
 n226409 , n226410 , n226411 , n226412 , n226413 , n226414 , n226415 , n226416 , n226417 , n226418 , 
 n226419 , n226420 , n226421 , n226422 , n226423 , n226424 , n226425 , n226426 , n226427 , n226428 , 
 n226429 , n226430 , n226431 , n226432 , n226433 , n226434 , n226435 , n226436 , n226437 , n226438 , 
 n226439 , n226440 , n226441 , n226442 , n226443 , n226444 , n226445 , n226446 , n226447 , n226448 , 
 n226449 , n226450 , n226451 , n226452 , n226453 , n226454 , n226455 , n226456 , n226457 , n226458 , 
 n226459 , n226460 , n226461 , n226462 , n226463 , n226464 , n226465 , n226466 , n226467 , n226468 , 
 n226469 , n226470 , n226471 , n226472 , n226473 , n226474 , n226475 , n226476 , n226477 , n226478 , 
 n226479 , n226480 , n226481 , n226482 , n226483 , n226484 , n226485 , n226486 , n226487 , n226488 , 
 n226489 , n226490 , n226491 , n226492 , n226493 , n226494 , n226495 , n226496 , n226497 , n226498 , 
 n226499 , n226500 , n226501 , n226502 , n226503 , n226504 , n226505 , n226506 , n226507 , n226508 , 
 n226509 , n226510 , n226511 , n226512 , n226513 , n226514 , n226515 , n226516 , n226517 , n226518 , 
 n226519 , n226520 , n226521 , n226522 , n226523 , n226524 , n226525 , n226526 , n226527 , n226528 , 
 n226529 , n226530 , n226531 , n226532 , n226533 , n226534 , n226535 , n226536 , n226537 , n226538 , 
 n226539 , n226540 , n226541 , n226542 , n226543 , n226544 , n226545 , n226546 , n226547 , n226548 , 
 n226549 , n226550 , n226551 , n226552 , n226553 , n226554 , n226555 , n226556 , n226557 , n226558 , 
 n226559 , n226560 , n226561 , n226562 , n226563 , n226564 , n226565 , n226566 , n226567 , n226568 , 
 n226569 , n226570 , n226571 , n226572 , n226573 , n226574 , n226575 , n226576 , n226577 , n226578 , 
 n226579 , n226580 , n226581 , n226582 , n226583 , n226584 , n226585 , n226586 , n226587 , n226588 , 
 n226589 , n226590 , n226591 , n226592 , n226593 , n226594 , n226595 , n226596 , n226597 , n226598 , 
 n226599 , n226600 , n226601 , n226602 , n226603 , n226604 , n226605 , n226606 , n226607 , n226608 , 
 n226609 , n226610 , n226611 , n226612 , n226613 , n226614 , n226615 , n226616 , n226617 , n226618 , 
 n226619 , n226620 , n226621 , n226622 , n226623 , n226624 , n226625 , n226626 , n226627 , n226628 , 
 n226629 , n226630 , n226631 , n226632 , n226633 , n226634 , n226635 , n226636 , n226637 , n226638 , 
 n226639 , n226640 , n226641 , n226642 , n226643 , n226644 , n226645 , n226646 , n226647 , n226648 , 
 n226649 , n226650 , n226651 , n226652 , n226653 , n226654 , n226655 , n226656 , n226657 , n226658 , 
 n226659 , n226660 , n226661 , n226662 , n226663 , n226664 , n226665 , n226666 , n226667 , n226668 , 
 n226669 , n226670 , n226671 , n226672 , n226673 , n226674 , n226675 , n226676 , n226677 , n226678 , 
 n226679 , n226680 , n226681 , n226682 , n226683 , n226684 , n226685 , n226686 , n226687 , n226688 , 
 n226689 , n226690 , n226691 , n226692 , n226693 , n226694 , n226695 , n226696 , n226697 , n226698 , 
 n226699 , n226700 , n226701 , n226702 , n226703 , n226704 , n226705 , n226706 , n226707 , n226708 , 
 n226709 , n226710 , n226711 , n226712 , n226713 , n226714 , n226715 , n226716 , n226717 , n226718 , 
 n226719 , n226720 , n226721 , n226722 , n226723 , n226724 , n226725 , n226726 , n226727 , n226728 , 
 n226729 , n226730 , n226731 , n226732 , n226733 , n226734 , n226735 , n226736 , n226737 , n226738 , 
 n226739 , n226740 , n226741 , n226742 , n226743 , n226744 , n226745 , n226746 , n226747 , n226748 , 
 n226749 , n226750 , n226751 , n226752 , n226753 , n226754 , n226755 , n226756 , n226757 , n226758 , 
 n226759 , n226760 , n226761 , n226762 , n226763 , n226764 , n226765 , n226766 , n226767 , n226768 , 
 n226769 , n226770 , n226771 , n226772 , n226773 , n226774 , n226775 , n226776 , n226777 , n226778 , 
 n226779 , n226780 , n226781 , n226782 , n226783 , n226784 , n226785 , n226786 , n226787 , n226788 , 
 n226789 , n226790 , n226791 , n226792 , n226793 , n226794 , n226795 , n226796 , n226797 , n226798 , 
 n226799 , n226800 , n226801 , n226802 , n226803 , n226804 , n226805 , n226806 , n226807 , n226808 , 
 n226809 , n226810 , n226811 , n226812 , n226813 , n226814 , n226815 , n226816 , n226817 , n226818 , 
 n226819 , n226820 , n226821 , n226822 , n226823 , n226824 , n226825 , n226826 , n226827 , n226828 , 
 n226829 , n226830 , n226831 , n226832 , n226833 , n226834 , n226835 , n226836 , n226837 , n226838 , 
 n226839 , n226840 , n226841 , n226842 , n226843 , n226844 , n226845 , n226846 , n226847 , n226848 , 
 n226849 , n226850 , n226851 , n226852 , n226853 , n226854 , n226855 , n226856 , n226857 , n226858 , 
 n226859 , n226860 , n226861 , n226862 , n226863 , n226864 , n226865 , n226866 , n226867 , n226868 , 
 n226869 , n226870 , n226871 , n226872 , n226873 , n226874 , n226875 , n226876 , n226877 , n226878 , 
 n226879 , n226880 , n226881 , n226882 , n226883 , n226884 , n226885 , n226886 , n226887 , n226888 , 
 n226889 , n226890 , n226891 , n226892 , n226893 , n226894 , n226895 , n226896 , n226897 , n226898 , 
 n226899 , n226900 , n226901 , n226902 , n226903 , n226904 , n226905 , n226906 , n226907 , n226908 , 
 n226909 , n226910 , n226911 , n226912 , n226913 , n226914 , n226915 , n226916 , n226917 , n226918 , 
 n226919 , n226920 , n226921 , n226922 , n226923 , n226924 , n226925 , n226926 , n226927 , n226928 , 
 n226929 , n226930 , n226931 , n226932 , n226933 , n226934 , n226935 , n226936 , n226937 , n226938 , 
 n226939 , n226940 , n226941 , n226942 , n226943 , n226944 , n226945 , n226946 , n226947 , n226948 , 
 n226949 , n226950 , n226951 , n226952 , n226953 , n226954 , n226955 , n226956 , n226957 , n226958 , 
 n226959 , n226960 , n226961 , n226962 , n226963 , n226964 , n226965 , n226966 , n226967 , n226968 , 
 n226969 , n226970 , n226971 , n226972 , n226973 , n226974 , n226975 , n226976 , n226977 , n226978 , 
 n226979 , n226980 , n226981 , n226982 , n226983 , n226984 , n226985 , n226986 , n226987 , n226988 , 
 n226989 , n226990 , n226991 , n226992 , n226993 , n226994 , n226995 , n226996 , n226997 , n226998 , 
 n226999 , n227000 , n227001 , n227002 , n227003 , n227004 , n227005 , n227006 , n227007 , n227008 , 
 n227009 , n227010 , n227011 , n227012 , n227013 , n227014 , n227015 , n227016 , n227017 , n227018 , 
 n227019 , n227020 , n227021 , n227022 , n227023 , n227024 , n227025 , n227026 , n227027 , n227028 , 
 n227029 , n227030 , n227031 , n227032 , n227033 , n227034 , n227035 , n227036 , n227037 , n227038 , 
 n227039 , n227040 , n227041 , n227042 , n227043 , n227044 , n227045 , n227046 , n227047 , n227048 , 
 n227049 , n227050 , n227051 , n227052 , n227053 , n227054 , n227055 , n227056 , n227057 , n227058 , 
 n227059 , n227060 , n227061 , n227062 , n227063 , n227064 , n227065 , n227066 , n227067 , n227068 , 
 n227069 , n227070 , n227071 , n227072 , n227073 , n227074 , n227075 , n227076 , n227077 , n227078 , 
 n227079 , n227080 , n227081 , n227082 , n227083 , n227084 , n227085 , n227086 , n227087 , n227088 , 
 n227089 , n227090 , n227091 , n227092 , n227093 , n227094 , n227095 , n227096 , n227097 , n227098 , 
 n227099 , n227100 , n227101 , n227102 , n227103 , n227104 , n227105 , n227106 , n227107 , n227108 , 
 n227109 , n227110 , n227111 , n227112 , n227113 , n227114 , n227115 , n227116 , n227117 , n227118 , 
 n227119 , n227120 , n227121 , n227122 , n227123 , n227124 , n227125 , n227126 , n227127 , n227128 , 
 n227129 , n227130 , n227131 , n227132 , n227133 , n227134 , n227135 , n227136 , n227137 , n227138 , 
 n227139 , n227140 , n227141 , n227142 , n227143 , n227144 , n227145 , n227146 , n227147 , n227148 , 
 n227149 , n227150 , n227151 , n227152 , n227153 , n227154 , n227155 , n227156 , n227157 , n227158 , 
 n227159 , n227160 , n227161 , n227162 , n227163 , n227164 , n227165 , n227166 , n227167 , n227168 , 
 n227169 , n227170 , n227171 , n227172 , n227173 , n227174 , n227175 , n227176 , n227177 , n227178 , 
 n227179 , n227180 , n227181 , n227182 , n227183 , n227184 , n227185 , n227186 , n227187 , n227188 , 
 n227189 , n227190 , n227191 , n227192 , n227193 , n227194 , n227195 , n227196 , n227197 , n227198 , 
 n227199 , n227200 , n227201 , n227202 , n227203 , n227204 , n227205 , n227206 , n227207 , n227208 , 
 n227209 , n227210 , n227211 , n227212 , n227213 , n227214 , n227215 , n227216 , n227217 , n227218 , 
 n227219 , n227220 , n227221 , n227222 , n227223 , n227224 , n227225 , n227226 , n227227 , n227228 , 
 n227229 , n227230 , n227231 , n227232 , n227233 , n227234 , n227235 , n227236 , n227237 , n227238 , 
 n227239 , n227240 , n227241 , n227242 , n227243 , n227244 , n227245 , n227246 , n227247 , n227248 , 
 n227249 , n227250 , n227251 , n227252 , n227253 , n227254 , n227255 , n227256 , n227257 , n227258 , 
 n227259 , n227260 , n227261 , n227262 , n227263 , n227264 , n227265 , n227266 , n227267 , n227268 , 
 n227269 , n227270 , n227271 , n227272 , n227273 , n227274 , n227275 , n227276 , n227277 , n227278 , 
 n227279 , n227280 , n227281 , n227282 , n227283 , n227284 , n227285 , n227286 , n227287 , n227288 , 
 n227289 , n227290 , n227291 , n227292 , n227293 , n227294 , n227295 , n227296 , n227297 , n227298 , 
 n227299 , n227300 , n227301 , n227302 , n227303 , n227304 , n227305 , n227306 , n227307 , n227308 , 
 n227309 , n227310 , n227311 , n227312 , n227313 , n227314 , n227315 , n227316 , n227317 , n227318 , 
 n227319 , n227320 , n227321 , n227322 , n227323 , n227324 , n227325 , n227326 , n227327 , n227328 , 
 n227329 , n227330 , n227331 , n227332 , n227333 , n227334 , n227335 , n227336 , n227337 , n227338 , 
 n227339 , n227340 , n227341 , n227342 , n227343 , n227344 , n227345 , n227346 , n227347 , n227348 , 
 n227349 , n227350 , n227351 , n227352 , n227353 , n227354 , n227355 , n227356 , n227357 , n227358 , 
 n227359 , n227360 , n227361 , n227362 , n227363 , n227364 , n227365 , n227366 , n227367 , n227368 , 
 n227369 , n227370 , n227371 , n227372 , n227373 , n227374 , n227375 , n227376 , n227377 , n227378 , 
 n227379 , n227380 , n227381 , n227382 , n227383 , n227384 , n227385 , n227386 , n227387 , n227388 , 
 n227389 , n227390 , n227391 , n227392 , n227393 , n227394 , n227395 , n227396 , n227397 , n227398 , 
 n227399 , n227400 , n227401 , n227402 , n227403 , n227404 , n227405 , n227406 , n227407 , n227408 , 
 n227409 , n227410 , n227411 , n227412 , n227413 , n227414 , n227415 , n227416 , n227417 , n227418 , 
 n227419 , n227420 , n227421 , n227422 , n227423 , n227424 , n227425 , n227426 , n227427 , n227428 , 
 n227429 , n227430 , n227431 , n227432 , n227433 , n227434 , n227435 , n227436 , n227437 , n227438 , 
 n227439 , n227440 , n227441 , n227442 , n227443 , n227444 , n227445 , n227446 , n227447 , n227448 , 
 n227449 , n227450 , n227451 , n227452 , n227453 , n227454 , n227455 , n227456 , n227457 , n227458 , 
 n227459 , n227460 , n227461 , n227462 , n227463 , n227464 , n227465 , n227466 , n227467 , n227468 , 
 n227469 , n227470 , n227471 , n227472 , n227473 , n227474 , n227475 , n227476 , n227477 , n227478 , 
 n227479 , n227480 , n227481 , n227482 , n227483 , n227484 , n227485 , n227486 , n227487 , n227488 , 
 n227489 , n227490 , n227491 , n227492 , n227493 , n227494 , n227495 , n227496 , n227497 , n227498 , 
 n227499 , n227500 , n227501 , n227502 , n227503 , n227504 , n227505 , n227506 , n227507 , n227508 , 
 n227509 , n227510 , n227511 , n227512 , n227513 , n227514 , n227515 , n227516 , n227517 , n227518 , 
 n227519 , n227520 , n227521 , n227522 , n227523 , n227524 , n227525 , n227526 , n227527 , n227528 , 
 n227529 , n227530 , n227531 , n227532 , n227533 , n227534 , n227535 , n227536 , n227537 , n227538 , 
 n227539 , n227540 , n227541 , n227542 , n227543 , n227544 , n227545 , n227546 , n227547 , n227548 , 
 n227549 , n227550 , n227551 , n227552 , n227553 , n227554 , n227555 , n227556 , n227557 , n227558 , 
 n227559 , n227560 , n227561 , n227562 , n227563 , n227564 , n227565 , n227566 , n227567 , n227568 , 
 n227569 , n227570 , n227571 , n227572 , n227573 , n227574 , n227575 , n227576 , n227577 , n227578 , 
 n227579 , n227580 , n227581 , n227582 , n227583 , n227584 , n227585 , n227586 , n227587 , n227588 , 
 n227589 , n227590 , n227591 , n227592 , n227593 , n227594 , n227595 , n227596 , n227597 , n227598 , 
 n227599 , n227600 , n227601 , n227602 , n227603 , n227604 , n227605 , n227606 , n227607 , n227608 , 
 n227609 , n227610 , n227611 , n227612 , n227613 , n227614 , n227615 , n227616 , n227617 , n227618 , 
 n227619 , n227620 , n227621 , n227622 , n227623 , n227624 , n227625 , n227626 , n227627 , n227628 , 
 n227629 , n227630 , n227631 , n227632 , n227633 , n227634 , n227635 , n227636 , n227637 , n227638 , 
 n227639 , n227640 , n227641 , n227642 , n227643 , n227644 , n227645 , n227646 , n227647 , n227648 , 
 n227649 , n227650 , n227651 , n227652 , n227653 , n227654 , n227655 , n227656 , n227657 , n227658 , 
 n227659 , n227660 , n227661 , n227662 , n227663 , n227664 , n227665 , n227666 , n227667 , n227668 , 
 n227669 , n227670 , n227671 , n227672 , n227673 , n227674 , n227675 , n227676 , n227677 , n227678 , 
 n227679 , n227680 , n227681 , n227682 , n227683 , n227684 , n227685 , n227686 , n227687 , n227688 , 
 n227689 , n227690 , n227691 , n227692 , n227693 , n227694 , n227695 , n227696 , n227697 , n227698 , 
 n227699 , n227700 , n227701 , n227702 , n227703 , n227704 , n227705 , n227706 , n227707 , n227708 , 
 n227709 , n227710 , n227711 , n227712 , n227713 , n227714 , n227715 , n227716 , n227717 , n227718 , 
 n227719 , n227720 , n227721 , n227722 , n227723 , n227724 , n227725 , n227726 , n227727 , n227728 , 
 n227729 , n227730 , n227731 , n227732 , n227733 , n227734 , n227735 , n227736 , n227737 , n227738 , 
 n227739 , n227740 , n227741 , n227742 , n227743 , n227744 , n227745 , n227746 , n227747 , n227748 , 
 n227749 , n227750 , n227751 , n227752 , n227753 , n227754 , n227755 , n227756 , n227757 , n227758 , 
 n227759 , n227760 , n227761 , n227762 , n227763 , n227764 , n227765 , n227766 , n227767 , n227768 , 
 n227769 , n227770 , n227771 , n227772 , n227773 , n227774 , n227775 , n227776 , n227777 , n227778 , 
 n227779 , n227780 , n227781 , n227782 , n227783 , n227784 , n227785 , n227786 , n227787 , n227788 , 
 n227789 , n227790 , n227791 , n227792 , n227793 , n227794 , n227795 , n227796 , n227797 , n227798 , 
 n227799 , n227800 , n227801 , n227802 , n227803 , n227804 , n227805 , n227806 , n227807 , n227808 , 
 n227809 , n227810 , n227811 , n227812 , n227813 , n227814 , n227815 , n227816 , n227817 , n227818 , 
 n227819 , n227820 , n227821 , n227822 , n227823 , n227824 , n227825 , n227826 , n227827 , n227828 , 
 n227829 , n227830 , n227831 , n227832 , n227833 , n227834 , n227835 , n227836 , n227837 , n227838 , 
 n227839 , n227840 , n227841 , n227842 , n227843 , n227844 , n227845 , n227846 , n227847 , n227848 , 
 n227849 , n227850 , n227851 , n227852 , n227853 , n227854 , n227855 , n227856 , n227857 , n227858 , 
 n227859 , n227860 , n227861 , n227862 , n227863 , n227864 , n227865 , n227866 , n227867 , n227868 , 
 n227869 , n227870 , n227871 , n227872 , n227873 , n227874 , n227875 , n227876 , n227877 , n227878 , 
 n227879 , n227880 , n227881 , n227882 , n227883 , n227884 , n227885 , n227886 , n227887 , n227888 , 
 n227889 , n227890 , n227891 , n227892 , n227893 , n227894 , n227895 , n227896 , n227897 , n227898 , 
 n227899 , n227900 , n227901 , n227902 , n227903 , n227904 , n227905 , n227906 , n227907 , n227908 , 
 n227909 , n227910 , n227911 , n227912 , n227913 , n227914 , n227915 , n227916 , n227917 , n227918 , 
 n227919 , n227920 , n227921 , n227922 , n227923 , n227924 , n227925 , n227926 , n227927 , n227928 , 
 n227929 , n227930 , n227931 , n227932 , n227933 , n227934 , n227935 , n227936 , n227937 , n227938 , 
 n227939 , n227940 , n227941 , n227942 , n227943 , n227944 , n227945 , n227946 , n227947 , n227948 , 
 n227949 , n227950 , n227951 , n227952 , n227953 , n227954 , n227955 , n227956 , n227957 , n227958 , 
 n227959 , n227960 , n227961 , n227962 , n227963 , n227964 , n227965 , n227966 , n227967 , n227968 , 
 n227969 , n227970 , n227971 , n227972 , n227973 , n227974 , n227975 , n227976 , n227977 , n227978 , 
 n227979 , n227980 , n227981 , n227982 , n227983 , n227984 , n227985 , n227986 , n227987 , n227988 , 
 n227989 , n227990 , n227991 , n227992 , n227993 , n227994 , n227995 , n227996 , n227997 , n227998 , 
 n227999 , n228000 , n228001 , n228002 , n228003 , n228004 , n228005 , n228006 , n228007 , n228008 , 
 n228009 , n228010 , n228011 , n228012 , n228013 , n228014 , n228015 , n228016 , n228017 , n228018 , 
 n228019 , n228020 , n228021 , n228022 , n228023 , n228024 , n228025 , n228026 , n228027 , n228028 , 
 n228029 , n228030 , n228031 , n228032 , n228033 , n228034 , n228035 , n228036 , n228037 , n228038 , 
 n228039 , n228040 , n228041 , n228042 , n228043 , n228044 , n228045 , n228046 , n228047 , n228048 , 
 n228049 , n228050 , n228051 , n228052 , n228053 , n228054 , n228055 , n228056 , n228057 , n228058 , 
 n228059 , n228060 , n228061 , n228062 , n228063 , n228064 , n228065 , n228066 , n228067 , n228068 , 
 n228069 , n228070 , n228071 , n228072 , n228073 , n228074 , n228075 , n228076 , n228077 , n228078 , 
 n228079 , n228080 , n228081 , n228082 , n228083 , n228084 , n228085 , n228086 , n228087 , n228088 , 
 n228089 , n228090 , n228091 , n228092 , n228093 , n228094 , n228095 , n228096 , n228097 , n228098 , 
 n228099 , n228100 , n228101 , n228102 , n228103 , n228104 , n228105 , n228106 , n228107 , n228108 , 
 n228109 , n228110 , n228111 , n228112 , n228113 , n228114 , n228115 , n228116 , n228117 , n228118 , 
 n228119 , n228120 , n228121 , n228122 , n228123 , n228124 , n228125 , n228126 , n228127 , n228128 , 
 n228129 , n228130 , n228131 , n228132 , n228133 , n228134 , n228135 , n228136 , n228137 , n228138 , 
 n228139 , n228140 , n228141 , n228142 , n228143 , n228144 , n228145 , n228146 , n228147 , n228148 , 
 n228149 , n228150 , n228151 , n228152 , n228153 , n228154 , n228155 , n228156 , n228157 , n228158 , 
 n228159 , n228160 , n228161 , n228162 , n228163 , n228164 , n228165 , n228166 , n228167 , n228168 , 
 n228169 , n228170 , n228171 , n228172 , n228173 , n228174 , n228175 , n228176 , n228177 , n228178 , 
 n228179 , n228180 , n228181 , n228182 , n228183 , n228184 , n228185 , n228186 , n228187 , n228188 , 
 n228189 , n228190 , n228191 , n228192 , n228193 , n228194 , n228195 , n228196 , n228197 , n228198 , 
 n228199 , n228200 , n228201 , n228202 , n228203 , n228204 , n228205 , n228206 , n228207 , n228208 , 
 n228209 , n228210 , n228211 , n228212 , n228213 , n228214 , n228215 , n228216 , n228217 , n228218 , 
 n228219 , n228220 , n228221 , n228222 , n228223 , n228224 , n228225 , n228226 , n228227 , n228228 , 
 n228229 , n228230 , n228231 , n228232 , n228233 , n228234 , n228235 , n228236 , n228237 , n228238 , 
 n228239 , n228240 , n228241 , n228242 , n228243 , n228244 , n228245 , n228246 , n228247 , n228248 , 
 n228249 , n228250 , n228251 , n228252 , n228253 , n228254 , n228255 , n228256 , n228257 , n228258 , 
 n228259 , n228260 , n228261 , n228262 , n228263 , n228264 , n228265 , n228266 , n228267 , n228268 , 
 n228269 , n228270 , n228271 , n228272 , n228273 , n228274 , n228275 , n228276 , n228277 , n228278 , 
 n228279 , n228280 , n228281 , n228282 , n228283 , n228284 , n228285 , n228286 , n228287 , n228288 , 
 n228289 , n228290 , n228291 , n228292 , n228293 , n228294 , n228295 , n228296 , n228297 , n228298 , 
 n228299 , n228300 , n228301 , n228302 , n228303 , n228304 , n228305 , n228306 , n228307 , n228308 , 
 n228309 , n228310 , n228311 , n228312 , n228313 , n228314 , n228315 , n228316 , n228317 , n228318 , 
 n228319 , n228320 , n228321 , n228322 , n228323 , n228324 , n228325 , n228326 , n228327 , n228328 , 
 n228329 , n228330 , n228331 , n228332 , n228333 , n228334 , n228335 , n228336 , n228337 , n228338 , 
 n228339 , n228340 , n228341 , n228342 , n228343 , n228344 , n228345 , n228346 , n228347 , n228348 , 
 n228349 , n228350 , n228351 , n228352 , n228353 , n228354 , n228355 , n228356 , n228357 , n228358 , 
 n228359 , n228360 , n228361 , n228362 , n228363 , n228364 , n228365 , n228366 , n228367 , n228368 , 
 n228369 , n228370 , n228371 , n228372 , n228373 , n228374 , n228375 , n228376 , n228377 , n228378 , 
 n228379 , n228380 , n228381 , n228382 , n228383 , n228384 , n228385 , n228386 , n228387 , n228388 , 
 n228389 , n228390 , n228391 , n228392 , n228393 , n228394 , n228395 , n228396 , n228397 , n228398 , 
 n228399 , n228400 , n228401 , n228402 , n228403 , n228404 , n228405 , n228406 , n228407 , n228408 , 
 n228409 , n228410 , n228411 , n228412 , n228413 , n228414 , n228415 , n228416 , n228417 , n228418 , 
 n228419 , n228420 , n228421 , n228422 , n228423 , n228424 , n228425 , n228426 , n228427 , n228428 , 
 n228429 , n228430 , n228431 , n228432 , n228433 , n228434 , n228435 , n228436 , n228437 , n228438 , 
 n228439 , n228440 , n228441 , n228442 , n228443 , n228444 , n228445 , n228446 , n228447 , n228448 , 
 n228449 , n228450 , n228451 , n228452 , n228453 , n228454 , n228455 , n228456 , n228457 , n228458 , 
 n228459 , n228460 , n228461 , n228462 , n228463 , n228464 , n228465 , n228466 , n228467 , n228468 , 
 n228469 , n228470 , n228471 , n228472 , n228473 , n228474 , n228475 , n228476 , n228477 , n228478 , 
 n228479 , n228480 , n228481 , n228482 , n228483 , n228484 , n228485 , n228486 , n228487 , n228488 , 
 n228489 , n228490 , n228491 , n228492 , n228493 , n228494 , n228495 , n228496 , n228497 , n228498 , 
 n228499 , n228500 , n228501 , n228502 , n228503 , n228504 , n228505 , n228506 , n228507 , n228508 , 
 n228509 , n228510 , n228511 , n228512 , n228513 , n228514 , n228515 , n228516 , n228517 , n228518 , 
 n228519 , n228520 , n228521 , n228522 , n228523 , n228524 , n228525 , n228526 , n228527 , n228528 , 
 n228529 , n228530 , n228531 , n228532 , n228533 , n228534 , n228535 , n228536 , n228537 , n228538 , 
 n228539 , n228540 , n228541 , n228542 , n228543 , n228544 , n228545 , n228546 , n228547 , n228548 , 
 n228549 , n228550 , n228551 , n228552 , n228553 , n228554 , n228555 , n228556 , n228557 , n228558 , 
 n228559 , n228560 , n228561 , n228562 , n228563 , n228564 , n228565 , n228566 , n228567 , n228568 , 
 n228569 , n228570 , n228571 , n228572 , n228573 , n228574 , n228575 , n228576 , n228577 , n228578 , 
 n228579 , n228580 , n228581 , n228582 , n228583 , n228584 , n228585 , n228586 , n228587 , n228588 , 
 n228589 , n228590 , n228591 , n228592 , n228593 , n228594 , n228595 , n228596 , n228597 , n228598 , 
 n228599 , n228600 , n228601 , n228602 , n228603 , n228604 , n228605 , n228606 , n228607 , n228608 , 
 n228609 , n228610 , n228611 , n228612 , n228613 , n228614 , n228615 , n228616 , n228617 , n228618 , 
 n228619 , n228620 , n228621 , n228622 , n228623 , n228624 , n228625 , n228626 , n228627 , n228628 , 
 n228629 , n228630 , n228631 , n228632 , n228633 , n228634 , n228635 , n228636 , n228637 , n228638 , 
 n228639 , n228640 , n228641 , n228642 , n228643 , n228644 , n228645 , n228646 , n228647 , n228648 , 
 n228649 , n228650 , n228651 , n228652 , n228653 , n228654 , n228655 , n228656 , n228657 , n228658 , 
 n228659 , n228660 , n228661 , n228662 , n228663 , n228664 , n228665 , n228666 , n228667 , n228668 , 
 n228669 , n228670 , n228671 , n228672 , n228673 , n228674 , n228675 , n228676 , n228677 , n228678 , 
 n228679 , n228680 , n228681 , n228682 , n228683 , n228684 , n228685 , n228686 , n228687 , n228688 , 
 n228689 , n228690 , n228691 , n228692 , n228693 , n228694 , n228695 , n228696 , n228697 , n228698 , 
 n228699 , n228700 , n228701 , n228702 , n228703 , n228704 , n228705 , n228706 , n228707 , n228708 , 
 n228709 , n228710 , n228711 , n228712 , n228713 , n228714 , n228715 , n228716 , n228717 , n228718 , 
 n228719 , n228720 , n228721 , n228722 , n228723 , n228724 , n228725 , n228726 , n228727 , n228728 , 
 n228729 , n228730 , n228731 , n228732 , n228733 , n228734 , n228735 , n228736 , n228737 , n228738 , 
 n228739 , n228740 , n228741 , n228742 , n228743 , n228744 , n228745 , n228746 , n228747 , n228748 , 
 n228749 , n228750 , n228751 , n228752 , n228753 , n228754 , n228755 , n228756 , n228757 , n228758 , 
 n228759 , n228760 , n228761 , n228762 , n228763 , n228764 , n228765 , n228766 , n228767 , n228768 , 
 n228769 , n228770 , n228771 , n228772 , n228773 , n228774 , n228775 , n228776 , n228777 , n228778 , 
 n228779 , n228780 , n228781 , n228782 , n228783 , n228784 , n228785 , n228786 , n228787 , n228788 , 
 n228789 , n228790 , n228791 , n228792 , n228793 , n228794 , n228795 , n228796 , n228797 , n228798 , 
 n228799 , n228800 , n228801 , n228802 , n228803 , n228804 , n228805 , n228806 , n228807 , n228808 , 
 n228809 , n228810 , n228811 , n228812 , n228813 , n228814 , n228815 , n228816 , n228817 , n228818 , 
 n228819 , n228820 , n228821 , n228822 , n228823 , n228824 , n228825 , n228826 , n228827 , n228828 , 
 n228829 , n228830 , n228831 , n228832 , n228833 , n228834 , n228835 , n228836 , n228837 , n228838 , 
 n228839 , n228840 , n228841 , n228842 , n228843 , n228844 , n228845 , n228846 , n228847 , n228848 , 
 n228849 , n228850 , n228851 , n228852 , n228853 , n228854 , n228855 , n228856 , n228857 , n228858 , 
 n228859 , n228860 , n228861 , n228862 , n228863 , n228864 , n228865 , n228866 , n228867 , n228868 , 
 n228869 , n228870 , n228871 , n228872 , n228873 , n228874 , n228875 , n228876 , n228877 , n228878 , 
 n228879 , n228880 , n228881 , n228882 , n228883 , n228884 , n228885 , n228886 , n228887 , n228888 , 
 n228889 , n228890 , n228891 , n228892 , n228893 , n228894 , n228895 , n228896 , n228897 , n228898 , 
 n228899 , n228900 , n228901 , n228902 , n228903 , n228904 , n228905 , n228906 , n228907 , n228908 , 
 n228909 , n228910 , n228911 , n228912 , n228913 , n228914 , n228915 , n228916 , n228917 , n228918 , 
 n228919 , n228920 , n228921 , n228922 , n228923 , n228924 , n228925 , n228926 , n228927 , n228928 , 
 n228929 , n228930 , n228931 , n228932 , n228933 , n228934 , n228935 , n228936 , n228937 , n228938 , 
 n228939 , n228940 , n228941 , n228942 , n228943 , n228944 , n228945 , n228946 , n228947 , n228948 , 
 n228949 , n228950 , n228951 , n228952 , n228953 , n228954 , n228955 , n228956 , n228957 , n228958 , 
 n228959 , n228960 , n228961 , n228962 , n228963 , n228964 , n228965 , n228966 , n228967 , n228968 , 
 n228969 , n228970 , n228971 , n228972 , n228973 , n228974 , n228975 , n228976 , n228977 , n228978 , 
 n228979 , n228980 , n228981 , n228982 , n228983 , n228984 , n228985 , n228986 , n228987 , n228988 , 
 n228989 , n228990 , n228991 , n228992 , n228993 , n228994 , n228995 , n228996 , n228997 , n228998 , 
 n228999 , n229000 , n229001 , n229002 , n229003 , n229004 , n229005 , n229006 , n229007 , n229008 , 
 n229009 , n229010 , n229011 , n229012 , n229013 , n229014 , n229015 , n229016 , n229017 , n229018 , 
 n229019 , n229020 , n229021 , n229022 , n229023 , n229024 , n229025 , n229026 , n229027 , n229028 , 
 n229029 , n229030 , n229031 , n229032 , n229033 , n229034 , n229035 , n229036 , n229037 , n229038 , 
 n229039 , n229040 , n229041 , n229042 , n229043 , n229044 , n229045 , n229046 , n229047 , n229048 , 
 n229049 , n229050 , n229051 , n229052 , n229053 , n229054 , n229055 , n229056 , n229057 , n229058 , 
 n229059 , n229060 , n229061 , n229062 , n229063 , n229064 , n229065 , n229066 , n229067 , n229068 , 
 n229069 , n229070 , n229071 , n229072 , n229073 , n229074 , n229075 , n229076 , n229077 , n229078 , 
 n229079 , n229080 , n229081 , n229082 , n229083 , n229084 , n229085 , n229086 , n229087 , n229088 , 
 n229089 , n229090 , n229091 , n229092 , n229093 , n229094 , n229095 , n229096 , n229097 , n229098 , 
 n229099 , n229100 , n229101 , n229102 , n229103 , n229104 , n229105 , n229106 , n229107 , n229108 , 
 n229109 , n229110 , n229111 , n229112 , n229113 , n229114 , n229115 , n229116 , n229117 , n229118 , 
 n229119 , n229120 , n229121 , n229122 , n229123 , n229124 , n229125 , n229126 , n229127 , n229128 , 
 n229129 , n229130 , n229131 , n229132 , n229133 , n229134 , n229135 , n229136 , n229137 , n229138 , 
 n229139 , n229140 , n229141 , n229142 , n229143 , n229144 , n229145 , n229146 , n229147 , n229148 , 
 n229149 , n229150 , n229151 , n229152 , n229153 , n229154 , n229155 , n229156 , n229157 , n229158 , 
 n229159 , n229160 , n229161 , n229162 , n229163 , n229164 , n229165 , n229166 , n229167 , n229168 , 
 n229169 , n229170 , n229171 , n229172 , n229173 , n229174 , n229175 , n229176 , n229177 , n229178 , 
 n229179 , n229180 , n229181 , n229182 , n229183 , n229184 , n229185 , n229186 , n229187 , n229188 , 
 n229189 , n229190 , n229191 , n229192 , n229193 , n229194 , n229195 , n229196 , n229197 , n229198 , 
 n229199 , n229200 , n229201 , n229202 , n229203 , n229204 , n229205 , n229206 , n229207 , n229208 , 
 n229209 , n229210 , n229211 , n229212 , n229213 , n229214 , n229215 , n229216 , n229217 , n229218 , 
 n229219 , n229220 , n229221 , n229222 , n229223 , n229224 , n229225 , n229226 , n229227 , n229228 , 
 n229229 , n229230 , n229231 , n229232 , n229233 , n229234 , n229235 , n229236 , n229237 , n229238 , 
 n229239 , n229240 , n229241 , n229242 , n229243 , n229244 , n229245 , n229246 , n229247 , n229248 , 
 n229249 , n229250 , n229251 , n229252 , n229253 , n229254 , n229255 , n229256 , n229257 , n229258 , 
 n229259 , n229260 , n229261 , n229262 , n229263 , n229264 , n229265 , n229266 , n229267 , n229268 , 
 n229269 , n229270 , n229271 , n229272 , n229273 , n229274 , n229275 , n229276 , n229277 , n229278 , 
 n229279 , n229280 , n229281 , n229282 , n229283 , n229284 , n229285 , n229286 , n229287 , n229288 , 
 n229289 , n229290 , n229291 , n229292 , n229293 , n229294 , n229295 , n229296 , n229297 , n229298 , 
 n229299 , n229300 , n229301 , n229302 , n229303 , n229304 , n229305 , n229306 , n229307 , n229308 , 
 n229309 , n229310 , n229311 , n229312 , n229313 , n229314 , n229315 , n229316 , n229317 , n229318 , 
 n229319 , n229320 , n229321 , n229322 , n229323 , n229324 , n229325 , n229326 , n229327 , n229328 , 
 n229329 , n229330 , n229331 , n229332 , n229333 , n229334 , n229335 , n229336 , n229337 , n229338 , 
 n229339 , n229340 , n229341 , n229342 , n229343 , n229344 , n229345 , n229346 , n229347 , n229348 , 
 n229349 , n229350 , n229351 , n229352 , n229353 , n229354 , n229355 , n229356 , n229357 , n229358 , 
 n229359 , n229360 , n229361 , n229362 , n229363 , n229364 , n229365 , n229366 , n229367 , n229368 , 
 n229369 , n229370 , n229371 , n229372 , n229373 , n229374 , n229375 , n229376 , n229377 , n229378 , 
 n229379 , n229380 , n229381 , n229382 , n229383 , n229384 , n229385 , n229386 , n229387 , n229388 , 
 n229389 , n229390 , n229391 , n229392 , n229393 , n229394 , n229395 , n229396 , n229397 , n229398 , 
 n229399 , n229400 , n229401 , n229402 , n229403 , n229404 , n229405 , n229406 , n229407 , n229408 , 
 n229409 , n229410 , n229411 , n229412 , n229413 , n229414 , n229415 , n229416 , n229417 , n229418 , 
 n229419 , n229420 , n229421 , n229422 , n229423 , n229424 , n229425 , n229426 , n229427 , n229428 , 
 n229429 , n229430 , n229431 , n229432 , n229433 , n229434 , n229435 , n229436 , n229437 , n229438 , 
 n229439 , n229440 , n229441 , n229442 , n229443 , n229444 , n229445 , n229446 , n229447 , n229448 , 
 n229449 , n229450 , n229451 , n229452 , n229453 , n229454 , n229455 , n229456 , n229457 , n229458 , 
 n229459 , n229460 , n229461 , n229462 , n229463 , n229464 , n229465 , n229466 , n229467 , n229468 , 
 n229469 , n229470 , n229471 , n229472 , n229473 , n229474 , n229475 , n229476 , n229477 , n229478 , 
 n229479 , n229480 , n229481 , n229482 , n229483 , n229484 , n229485 , n229486 , n229487 , n229488 , 
 n229489 , n229490 , n229491 , n229492 , n229493 , n229494 , n229495 , n229496 , n229497 , n229498 , 
 n229499 , n229500 , n229501 , n229502 , n229503 , n229504 , n229505 , n229506 , n229507 , n229508 , 
 n229509 , n229510 , n229511 , n229512 , n229513 , n229514 , n229515 , n229516 , n229517 , n229518 , 
 n229519 , n229520 , n229521 , n229522 , n229523 , n229524 , n229525 , n229526 , n229527 , n229528 , 
 n229529 , n229530 , n229531 , n229532 , n229533 , n229534 , n229535 , n229536 , n229537 , n229538 , 
 n229539 , n229540 , n229541 , n229542 , n229543 , n229544 , n229545 , n229546 , n229547 , n229548 , 
 n229549 , n229550 , n229551 , n229552 , n229553 , n229554 , n229555 , n229556 , n229557 , n229558 , 
 n229559 , n229560 , n229561 , n229562 , n229563 , n229564 , n229565 , n229566 , n229567 , n229568 , 
 n229569 , n229570 , n229571 , n229572 , n229573 , n229574 , n229575 , n229576 , n229577 , n229578 , 
 n229579 , n229580 , n229581 , n229582 , n229583 , n229584 , n229585 , n229586 , n229587 , n229588 , 
 n229589 , n229590 , n229591 , n229592 , n229593 , n229594 , n229595 , n229596 , n229597 , n229598 , 
 n229599 , n229600 , n229601 , n229602 , n229603 , n229604 , n229605 , n229606 , n229607 , n229608 , 
 n229609 , n229610 , n229611 , n229612 , n229613 , n229614 , n229615 , n229616 , n229617 , n229618 , 
 n229619 , n229620 , n229621 , n229622 , n229623 , n229624 , n229625 , n229626 , n229627 , n229628 , 
 n229629 , n229630 , n229631 , n229632 , n229633 , n229634 , n229635 , n229636 , n229637 , n229638 , 
 n229639 , n229640 , n229641 , n229642 , n229643 , n229644 , n229645 , n229646 , n229647 , n229648 , 
 n229649 , n229650 , n229651 , n229652 , n229653 , n229654 , n229655 , n229656 , n229657 , n229658 , 
 n229659 , n229660 , n229661 , n229662 , n229663 , n229664 , n229665 , n229666 , n229667 , n229668 , 
 n229669 , n229670 , n229671 , n229672 , n229673 , n229674 , n229675 , n229676 , n229677 , n229678 , 
 n229679 , n229680 , n229681 , n229682 , n229683 , n229684 , n229685 , n229686 , n229687 , n229688 , 
 n229689 , n229690 , n229691 , n229692 , n229693 , n229694 , n229695 , n229696 , n229697 , n229698 , 
 n229699 , n229700 , n229701 , n229702 , n229703 , n229704 , n229705 , n229706 , n229707 , n229708 , 
 n229709 , n229710 , n229711 , n229712 , n229713 , n229714 , n229715 , n229716 , n229717 , n229718 , 
 n229719 , n229720 , n229721 , n229722 , n229723 , n229724 , n229725 , n229726 , n229727 , n229728 , 
 n229729 , n229730 , n229731 , n229732 , n229733 , n229734 , n229735 , n229736 , n229737 , n229738 , 
 n229739 , n229740 , n229741 , n229742 , n229743 , n229744 , n229745 , n229746 , n229747 , n229748 , 
 n229749 , n229750 , n229751 , n229752 , n229753 , n229754 , n229755 , n229756 , n229757 , n229758 , 
 n229759 , n229760 , n229761 , n229762 , n229763 , n229764 , n229765 , n229766 , n229767 , n229768 , 
 n229769 , n229770 , n229771 , n229772 , n229773 , n229774 , n229775 , n229776 , n229777 , n229778 , 
 n229779 , n229780 , n229781 , n229782 , n229783 , n229784 , n229785 , n229786 , n229787 , n229788 , 
 n229789 , n229790 , n229791 , n229792 , n229793 , n229794 , n229795 , n229796 , n229797 , n229798 , 
 n229799 , n229800 , n229801 , n229802 , n229803 , n229804 , n229805 , n229806 , n229807 , n229808 , 
 n229809 , n229810 , n229811 , n229812 , n229813 , n229814 , n229815 , n229816 , n229817 , n229818 , 
 n229819 , n229820 , n229821 , n229822 , n229823 , n229824 , n229825 , n229826 , n229827 , n229828 , 
 n229829 , n229830 , n229831 , n229832 , n229833 , n229834 , n229835 , n229836 , n229837 , n229838 , 
 n229839 , n229840 , n229841 , n229842 , n229843 , n229844 , n229845 , n229846 , n229847 , n229848 , 
 n229849 , n229850 , n229851 , n229852 , n229853 , n229854 , n229855 , n229856 , n229857 , n229858 , 
 n229859 , n229860 , n229861 , n229862 , n229863 , n229864 , n229865 , n229866 , n229867 , n229868 , 
 n229869 , n229870 , n229871 , n229872 , n229873 , n229874 , n229875 , n229876 , n229877 , n229878 , 
 n229879 , n229880 , n229881 , n229882 , n229883 , n229884 , n229885 , n229886 , n229887 , n229888 , 
 n229889 , n229890 , n229891 , n229892 , n229893 , n229894 , n229895 , n229896 , n229897 , n229898 , 
 n229899 , n229900 , n229901 , n229902 , n229903 , n229904 , n229905 , n229906 , n229907 , n229908 , 
 n229909 , n229910 , n229911 , n229912 , n229913 , n229914 , n229915 , n229916 , n229917 , n229918 , 
 n229919 , n229920 , n229921 , n229922 , n229923 , n229924 , n229925 , n229926 , n229927 , n229928 , 
 n229929 , n229930 , n229931 , n229932 , n229933 , n229934 , n229935 , n229936 , n229937 , n229938 , 
 n229939 , n229940 , n229941 , n229942 , n229943 , n229944 , n229945 , n229946 , n229947 , n229948 , 
 n229949 , n229950 , n229951 , n229952 , n229953 , n229954 , n229955 , n229956 , n229957 , n229958 , 
 n229959 , n229960 , n229961 , n229962 , n229963 , n229964 , n229965 , n229966 , n229967 , n229968 , 
 n229969 , n229970 , n229971 , n229972 , n229973 , n229974 , n229975 , n229976 , n229977 , n229978 , 
 n229979 , n229980 , n229981 , n229982 , n229983 , n229984 , n229985 , n229986 , n229987 , n229988 , 
 n229989 , n229990 , n229991 , n229992 , n229993 , n229994 , n229995 , n229996 , n229997 , n229998 , 
 n229999 , n230000 , n230001 , n230002 , n230003 , n230004 , n230005 , n230006 , n230007 , n230008 , 
 n230009 , n230010 , n230011 , n230012 , n230013 , n230014 , n230015 , n230016 , n230017 , n230018 , 
 n230019 , n230020 , n230021 , n230022 , n230023 , n230024 , n230025 , n230026 , n230027 , n230028 , 
 n230029 , n230030 , n230031 , n230032 , n230033 , n230034 , n230035 , n230036 , n230037 , n230038 , 
 n230039 , n230040 , n230041 , n230042 , n230043 , n230044 , n230045 , n230046 , n230047 , n230048 , 
 n230049 , n230050 , n230051 , n230052 , n230053 , n230054 , n230055 , n230056 , n230057 , n230058 , 
 n230059 , n230060 , n230061 , n230062 , n230063 , n230064 , n230065 , n230066 , n230067 , n230068 , 
 n230069 , n230070 , n230071 , n230072 , n230073 , n230074 , n230075 , n230076 , n230077 , n230078 , 
 n230079 , n230080 , n230081 , n230082 , n230083 , n230084 , n230085 , n230086 , n230087 , n230088 , 
 n230089 , n230090 , n230091 , n230092 , n230093 , n230094 , n230095 , n230096 , n230097 , n230098 , 
 n230099 , n230100 , n230101 , n230102 , n230103 , n230104 , n230105 , n230106 , n230107 , n230108 , 
 n230109 , n230110 , n230111 , n230112 , n230113 , n230114 , n230115 , n230116 , n230117 , n230118 , 
 n230119 , n230120 , n230121 , n230122 , n230123 , n230124 , n230125 , n230126 , n230127 , n230128 , 
 n230129 , n230130 , n230131 , n230132 , n230133 , n230134 , n230135 , n230136 , n230137 , n230138 , 
 n230139 , n230140 , n230141 , n230142 , n230143 , n230144 , n230145 , n230146 , n230147 , n230148 , 
 n230149 , n230150 , n230151 , n230152 , n230153 , n230154 , n230155 , n230156 , n230157 , n230158 , 
 n230159 , n230160 , n230161 , n230162 , n230163 , n230164 , n230165 , n230166 , n230167 , n230168 , 
 n230169 , n230170 , n230171 , n230172 , n230173 , n230174 , n230175 , n230176 , n230177 , n230178 , 
 n230179 , n230180 , n230181 , n230182 , n230183 , n230184 , n230185 , n230186 , n230187 , n230188 , 
 n230189 , n230190 , n230191 , n230192 , n230193 , n230194 , n230195 , n230196 , n230197 , n230198 , 
 n230199 , n230200 , n230201 , n230202 , n230203 , n230204 , n230205 , n230206 , n230207 , n230208 , 
 n230209 , n230210 , n230211 , n230212 , n230213 , n230214 , n230215 , n230216 , n230217 , n230218 , 
 n230219 , n230220 , n230221 , n230222 , n230223 , n230224 , n230225 , n230226 , n230227 , n230228 , 
 n230229 , n230230 , n230231 , n230232 , n230233 , n230234 , n230235 , n230236 , n230237 , n230238 , 
 n230239 , n230240 , n230241 , n230242 , n230243 , n230244 , n230245 , n230246 , n230247 , n230248 , 
 n230249 , n230250 , n230251 , n230252 , n230253 , n230254 , n230255 , n230256 , n230257 , n230258 , 
 n230259 , n230260 , n230261 , n230262 , n230263 , n230264 , n230265 , n230266 , n230267 , n230268 , 
 n230269 , n230270 , n230271 , n230272 , n230273 , n230274 , n230275 , n230276 , n230277 , n230278 , 
 n230279 , n230280 , n230281 , n230282 , n230283 , n230284 , n230285 , n230286 , n230287 , n230288 , 
 n230289 , n230290 , n230291 , n230292 , n230293 , n230294 , n230295 , n230296 , n230297 , n230298 , 
 n230299 , n230300 , n230301 , n230302 , n230303 , n230304 , n230305 , n230306 , n230307 , n230308 , 
 n230309 , n230310 , n230311 , n230312 , n230313 , n230314 , n230315 , n230316 , n230317 , n230318 , 
 n230319 , n230320 , n230321 , n230322 , n230323 , n230324 , n230325 , n230326 , n230327 , n230328 , 
 n230329 , n230330 , n230331 , n230332 , n230333 , n230334 , n230335 , n230336 , n230337 , n230338 , 
 n230339 , n230340 , n230341 , n230342 , n230343 , n230344 , n230345 , n230346 , n230347 , n230348 , 
 n230349 , n230350 , n230351 , n230352 , n230353 , n230354 , n230355 , n230356 , n230357 , n230358 , 
 n230359 , n230360 , n230361 , n230362 , n230363 , n230364 , n230365 , n230366 , n230367 , n230368 , 
 n230369 , n230370 , n230371 , n230372 , n230373 , n230374 , n230375 , n230376 , n230377 , n230378 , 
 n230379 , n230380 , n230381 , n230382 , n230383 , n230384 , n230385 , n230386 , n230387 , n230388 , 
 n230389 , n230390 , n230391 , n230392 , n230393 , n230394 , n230395 , n230396 , n230397 , n230398 , 
 n230399 , n230400 , n230401 , n230402 , n230403 , n230404 , n230405 , n230406 , n230407 , n230408 , 
 n230409 , n230410 , n230411 , n230412 , n230413 , n230414 , n230415 , n230416 , n230417 , n230418 , 
 n230419 , n230420 , n230421 , n230422 , n230423 , n230424 , n230425 , n230426 , n230427 , n230428 , 
 n230429 , n230430 , n230431 , n230432 , n230433 , n230434 , n230435 , n230436 , n230437 , n230438 , 
 n230439 , n230440 , n230441 , n230442 , n230443 , n230444 , n230445 , n230446 , n230447 , n230448 , 
 n230449 , n230450 , n230451 , n230452 , n230453 , n230454 , n230455 , n230456 , n230457 , n230458 , 
 n230459 , n230460 , n230461 , n230462 , n230463 , n230464 , n230465 , n230466 , n230467 , n230468 , 
 n230469 , n230470 , n230471 , n230472 , n230473 , n230474 , n230475 , n230476 , n230477 , n230478 , 
 n230479 , n230480 , n230481 , n230482 , n230483 , n230484 , n230485 , n230486 , n230487 , n230488 , 
 n230489 , n230490 , n230491 , n230492 , n230493 , n230494 , n230495 , n230496 , n230497 , n230498 , 
 n230499 , n230500 , n230501 , n230502 , n230503 , n230504 , n230505 , n230506 , n230507 , n230508 , 
 n230509 , n230510 , n230511 , n230512 , n230513 , n230514 , n230515 , n230516 , n230517 , n230518 , 
 n230519 , n230520 , n230521 , n230522 , n230523 , n230524 , n230525 , n230526 , n230527 , n230528 , 
 n230529 , n230530 , n230531 , n230532 , n230533 , n230534 , n230535 , n230536 , n230537 , n230538 , 
 n230539 , n230540 , n230541 , n230542 , n230543 , n230544 , n230545 , n230546 , n230547 , n230548 , 
 n230549 , n230550 , n230551 , n230552 , n230553 , n230554 , n230555 , n230556 , n230557 , n230558 , 
 n230559 , n230560 , n230561 , n230562 , n230563 , n230564 , n230565 , n230566 , n230567 , n230568 , 
 n230569 , n230570 , n230571 , n230572 , n230573 , n230574 , n230575 , n230576 , n230577 , n230578 , 
 n230579 , n230580 , n230581 , n230582 , n230583 , n230584 , n230585 , n230586 , n230587 , n230588 , 
 n230589 , n230590 , n230591 , n230592 , n230593 , n230594 , n230595 , n230596 , n230597 , n230598 , 
 n230599 , n230600 , n230601 , n230602 , n230603 , n230604 , n230605 , n230606 , n230607 , n230608 , 
 n230609 , n230610 , n230611 , n230612 , n230613 , n230614 , n230615 , n230616 , n230617 , n230618 , 
 n230619 , n230620 , n230621 , n230622 , n230623 , n230624 , n230625 , n230626 , n230627 , n230628 , 
 n230629 , n230630 , n230631 , n230632 , n230633 , n230634 , n230635 , n230636 , n230637 , n230638 , 
 n230639 , n230640 , n230641 , n230642 , n230643 , n230644 , n230645 , n230646 , n230647 , n230648 , 
 n230649 , n230650 , n230651 , n230652 , n230653 , n230654 , n230655 , n230656 , n230657 , n230658 , 
 n230659 , n230660 , n230661 , n230662 , n230663 , n230664 , n230665 , n230666 , n230667 , n230668 , 
 n230669 , n230670 , n230671 , n230672 , n230673 , n230674 , n230675 , n230676 , n230677 , n230678 , 
 n230679 , n230680 , n230681 , n230682 , n230683 , n230684 , n230685 , n230686 , n230687 , n230688 , 
 n230689 , n230690 , n230691 , n230692 , n230693 , n230694 , n230695 , n230696 , n230697 , n230698 , 
 n230699 , n230700 , n230701 , n230702 , n230703 , n230704 , n230705 , n230706 , n230707 , n230708 , 
 n230709 , n230710 , n230711 , n230712 , n230713 , n230714 , n230715 , n230716 , n230717 , n230718 , 
 n230719 , n230720 , n230721 , n230722 , n230723 , n230724 , n230725 , n230726 , n230727 , n230728 , 
 n230729 , n230730 , n230731 , n230732 , n230733 , n230734 , n230735 , n230736 , n230737 , n230738 , 
 n230739 , n230740 , n230741 , n230742 , n230743 , n230744 , n230745 , n230746 , n230747 , n230748 , 
 n230749 , n230750 , n230751 , n230752 , n230753 , n230754 , n230755 , n230756 , n230757 , n230758 , 
 n230759 , n230760 , n230761 , n230762 , n230763 , n230764 , n230765 , n230766 , n230767 , n230768 , 
 n230769 , n230770 , n230771 , n230772 , n230773 , n230774 , n230775 , n230776 , n230777 , n230778 , 
 n230779 , n230780 , n230781 , n230782 , n230783 , n230784 , n230785 , n230786 , n230787 , n230788 , 
 n230789 , n230790 , n230791 , n230792 , n230793 , n230794 , n230795 , n230796 , n230797 , n230798 , 
 n230799 , n230800 , n230801 , n230802 , n230803 , n230804 , n230805 , n230806 , n230807 , n230808 , 
 n230809 , n230810 , n230811 , n230812 , n230813 , n230814 , n230815 , n230816 , n230817 , n230818 , 
 n230819 , n230820 , n230821 , n230822 , n230823 , n230824 , n230825 , n230826 , n230827 , n230828 , 
 n230829 , n230830 , n230831 , n230832 , n230833 , n230834 , n230835 , n230836 , n230837 , n230838 , 
 n230839 , n230840 , n230841 , n230842 , n230843 , n230844 , n230845 , n230846 , n230847 , n230848 , 
 n230849 , n230850 , n230851 , n230852 , n230853 , n230854 , n230855 , n230856 , n230857 , n230858 , 
 n230859 , n230860 , n230861 , n230862 , n230863 , n230864 , n230865 , n230866 , n230867 , n230868 , 
 n230869 , n230870 , n230871 , n230872 , n230873 , n230874 , n230875 , n230876 , n230877 , n230878 , 
 n230879 , n230880 , n230881 , n230882 , n230883 , n230884 , n230885 , n230886 , n230887 , n230888 , 
 n230889 , n230890 , n230891 , n230892 , n230893 , n230894 , n230895 , n230896 , n230897 , n230898 , 
 n230899 , n230900 , n230901 , n230902 , n230903 , n230904 , n230905 , n230906 , n230907 , n230908 , 
 n230909 , n230910 , n230911 , n230912 , n230913 , n230914 , n230915 , n230916 , n230917 , n230918 , 
 n230919 , n230920 , n230921 , n230922 , n230923 , n230924 , n230925 , n230926 , n230927 , n230928 , 
 n230929 , n230930 , n230931 , n230932 , n230933 , n230934 , n230935 , n230936 , n230937 , n230938 , 
 n230939 , n230940 , n230941 , n230942 , n230943 , n230944 , n230945 , n230946 , n230947 , n230948 , 
 n230949 , n230950 , n230951 , n230952 , n230953 , n230954 , n230955 , n230956 , n230957 , n230958 , 
 n230959 , n230960 , n230961 , n230962 , n230963 , n230964 , n230965 , n230966 , n230967 , n230968 , 
 n230969 , n230970 , n230971 , n230972 , n230973 , n230974 , n230975 , n230976 , n230977 , n230978 , 
 n230979 , n230980 , n230981 , n230982 , n230983 , n230984 , n230985 , n230986 , n230987 , n230988 , 
 n230989 , n230990 , n230991 , n230992 , n230993 , n230994 , n230995 , n230996 , n230997 , n230998 , 
 n230999 , n231000 , n231001 , n231002 , n231003 , n231004 , n231005 , n231006 , n231007 , n231008 , 
 n231009 , n231010 , n231011 , n231012 , n231013 , n231014 , n231015 , n231016 , n231017 , n231018 , 
 n231019 , n231020 , n231021 , n231022 , n231023 , n231024 , n231025 , n231026 , n231027 , n231028 , 
 n231029 , n231030 , n231031 , n231032 , n231033 , n231034 , n231035 , n231036 , n231037 , n231038 , 
 n231039 , n231040 , n231041 , n231042 , n231043 , n231044 , n231045 , n231046 , n231047 , n231048 , 
 n231049 , n231050 , n231051 , n231052 , n231053 , n231054 , n231055 , n231056 , n231057 , n231058 , 
 n231059 , n231060 , n231061 , n231062 , n231063 , n231064 , n231065 , n231066 , n231067 , n231068 , 
 n231069 , n231070 , n231071 , n231072 , n231073 , n231074 , n231075 , n231076 , n231077 , n231078 , 
 n231079 , n231080 , n231081 , n231082 , n231083 , n231084 , n231085 , n231086 , n231087 , n231088 , 
 n231089 , n231090 , n231091 , n231092 , n231093 , n231094 , n231095 , n231096 , n231097 , n231098 , 
 n231099 , n231100 , n231101 , n231102 , n231103 , n231104 , n231105 , n231106 , n231107 , n231108 , 
 n231109 , n231110 , n231111 , n231112 , n231113 , n231114 , n231115 , n231116 , n231117 , n231118 , 
 n231119 , n231120 , n231121 , n231122 , n231123 , n231124 , n231125 , n231126 , n231127 , n231128 , 
 n231129 , n231130 , n231131 , n231132 , n231133 , n231134 , n231135 , n231136 , n231137 , n231138 , 
 n231139 , n231140 , n231141 , n231142 , n231143 , n231144 , n231145 , n231146 , n231147 , n231148 , 
 n231149 , n231150 , n231151 , n231152 , n231153 , n231154 , n231155 , n231156 , n231157 , n231158 , 
 n231159 , n231160 , n231161 , n231162 , n231163 , n231164 , n231165 , n231166 , n231167 , n231168 , 
 n231169 , n231170 , n231171 , n231172 , n231173 , n231174 , n231175 , n231176 , n231177 , n231178 , 
 n231179 , n231180 , n231181 , n231182 , n231183 , n231184 , n231185 , n231186 , n231187 , n231188 , 
 n231189 , n231190 , n231191 , n231192 , n231193 , n231194 , n231195 , n231196 , n231197 , n231198 , 
 n231199 , n231200 , n231201 , n231202 , n231203 , n231204 , n231205 , n231206 , n231207 , n231208 , 
 n231209 , n231210 , n231211 , n231212 , n231213 , n231214 , n231215 , n231216 , n231217 , n231218 , 
 n231219 , n231220 , n231221 , n231222 , n231223 , n231224 , n231225 , n231226 , n231227 , n231228 , 
 n231229 , n231230 , n231231 , n231232 , n231233 , n231234 , n231235 , n231236 , n231237 , n231238 , 
 n231239 , n231240 , n231241 , n231242 , n231243 , n231244 , n231245 , n231246 , n231247 , n231248 , 
 n231249 , n231250 , n231251 , n231252 , n231253 , n231254 , n231255 , n231256 , n231257 , n231258 , 
 n231259 , n231260 , n231261 , n231262 , n231263 , n231264 , n231265 , n231266 , n231267 , n231268 , 
 n231269 , n231270 , n231271 , n231272 , n231273 , n231274 , n231275 , n231276 , n231277 , n231278 , 
 n231279 , n231280 , n231281 , n231282 , n231283 , n231284 , n231285 , n231286 , n231287 , n231288 , 
 n231289 , n231290 , n231291 , n231292 , n231293 , n231294 , n231295 , n231296 , n231297 , n231298 , 
 n231299 , n231300 , n231301 , n231302 , n231303 , n231304 , n231305 , n231306 , n231307 , n231308 , 
 n231309 , n231310 , n231311 , n231312 , n231313 , n231314 , n231315 , n231316 , n231317 , n231318 , 
 n231319 , n231320 , n231321 , n231322 , n231323 , n231324 , n231325 , n231326 , n231327 , n231328 , 
 n231329 , n231330 , n231331 , n231332 , n231333 , n231334 , n231335 , n231336 , n231337 , n231338 , 
 n231339 , n231340 , n231341 , n231342 , n231343 , n231344 , n231345 , n231346 , n231347 , n231348 , 
 n231349 , n231350 , n231351 , n231352 , n231353 , n231354 , n231355 , n231356 , n231357 , n231358 , 
 n231359 , n231360 , n231361 , n231362 , n231363 , n231364 , n231365 , n231366 , n231367 , n231368 , 
 n231369 , n231370 , n231371 , n231372 , n231373 , n231374 , n231375 , n231376 , n231377 , n231378 , 
 n231379 , n231380 , n231381 , n231382 , n231383 , n231384 , n231385 , n231386 , n231387 , n231388 , 
 n231389 , n231390 , n231391 , n231392 , n231393 , n231394 , n231395 , n231396 , n231397 , n231398 , 
 n231399 , n231400 , n231401 , n231402 , n231403 , n231404 , n231405 , n231406 , n231407 , n231408 , 
 n231409 , n231410 , n231411 , n231412 , n231413 , n231414 , n231415 , n231416 , n231417 , n231418 , 
 n231419 , n231420 , n231421 , n231422 , n231423 , n231424 , n231425 , n231426 , n231427 , n231428 , 
 n231429 , n231430 , n231431 , n231432 , n231433 , n231434 , n231435 , n231436 , n231437 , n231438 , 
 n231439 , n231440 , n231441 , n231442 , n231443 , n231444 , n231445 , n231446 , n231447 , n231448 , 
 n231449 , n231450 , n231451 , n231452 , n231453 , n231454 , n231455 , n231456 , n231457 , n231458 , 
 n231459 , n231460 , n231461 , n231462 , n231463 , n231464 , n231465 , n231466 , n231467 , n231468 , 
 n231469 , n231470 , n231471 , n231472 , n231473 , n231474 , n231475 , n231476 , n231477 , n231478 , 
 n231479 , n231480 , n231481 , n231482 , n231483 , n231484 , n231485 , n231486 , n231487 , n231488 , 
 n231489 , n231490 , n231491 , n231492 , n231493 , n231494 , n231495 , n231496 , n231497 , n231498 , 
 n231499 , n231500 , n231501 , n231502 , n231503 , n231504 , n231505 , n231506 , n231507 , n231508 , 
 n231509 , n231510 , n231511 , n231512 , n231513 , n231514 , n231515 , n231516 , n231517 , n231518 , 
 n231519 , n231520 , n231521 , n231522 , n231523 , n231524 , n231525 , n231526 , n231527 , n231528 , 
 n231529 , n231530 , n231531 , n231532 , n231533 , n231534 , n231535 , n231536 , n231537 , n231538 , 
 n231539 , n231540 , n231541 , n231542 , n231543 , n231544 , n231545 , n231546 , n231547 , n231548 , 
 n231549 , n231550 , n231551 , n231552 , n231553 , n231554 , n231555 , n231556 , n231557 , n231558 , 
 n231559 , n231560 , n231561 , n231562 , n231563 , n231564 , n231565 , n231566 , n231567 , n231568 , 
 n231569 , n231570 , n231571 , n231572 , n231573 , n231574 , n231575 , n231576 , n231577 , n231578 , 
 n231579 , n231580 , n231581 , n231582 , n231583 , n231584 , n231585 , n231586 , n231587 , n231588 , 
 n231589 , n231590 , n231591 , n231592 , n231593 , n231594 , n231595 , n231596 , n231597 , n231598 , 
 n231599 , n231600 , n231601 , n231602 , n231603 , n231604 , n231605 , n231606 , n231607 , n231608 , 
 n231609 , n231610 , n231611 , n231612 , n231613 , n231614 , n231615 , n231616 , n231617 , n231618 , 
 n231619 , n231620 , n231621 , n231622 , n231623 , n231624 , n231625 , n231626 , n231627 , n231628 , 
 n231629 , n231630 , n231631 , n231632 , n231633 , n231634 , n231635 , n231636 , n231637 , n231638 , 
 n231639 , n231640 , n231641 , n231642 , n231643 , n231644 , n231645 , n231646 , n231647 , n231648 , 
 n231649 , n231650 , n231651 , n231652 , n231653 , n231654 , n231655 , n231656 , n231657 , n231658 , 
 n231659 , n231660 , n231661 , n231662 , n231663 , n231664 , n231665 , n231666 , n231667 , n231668 , 
 n231669 , n231670 , n231671 , n231672 , n231673 , n231674 , n231675 , n231676 , n231677 , n231678 , 
 n231679 , n231680 , n231681 , n231682 , n231683 , n231684 , n231685 , n231686 , n231687 , n231688 , 
 n231689 , n231690 , n231691 , n231692 , n231693 , n231694 , n231695 , n231696 , n231697 , n231698 , 
 n231699 , n231700 , n231701 , n231702 , n231703 , n231704 , n231705 , n231706 , n231707 , n231708 , 
 n231709 , n231710 , n231711 , n231712 , n231713 , n231714 , n231715 , n231716 , n231717 , n231718 , 
 n231719 , n231720 , n231721 , n231722 , n231723 , n231724 , n231725 , n231726 , n231727 , n231728 , 
 n231729 , n231730 , n231731 , n231732 , n231733 , n231734 , n231735 , n231736 , n231737 , n231738 , 
 n231739 , n231740 , n231741 , n231742 , n231743 , n231744 , n231745 , n231746 , n231747 , n231748 , 
 n231749 , n231750 , n231751 , n231752 , n231753 , n231754 , n231755 , n231756 , n231757 , n231758 , 
 n231759 , n231760 , n231761 , n231762 , n231763 , n231764 , n231765 , n231766 , n231767 , n231768 , 
 n231769 , n231770 , n231771 , n231772 , n231773 , n231774 , n231775 , n231776 , n231777 , n231778 , 
 n231779 , n231780 , n231781 , n231782 , n231783 , n231784 , n231785 , n231786 , n231787 , n231788 , 
 n231789 , n231790 , n231791 , n231792 , n231793 , n231794 , n231795 , n231796 , n231797 , n231798 , 
 n231799 , n231800 , n231801 , n231802 , n231803 , n231804 , n231805 , n231806 , n231807 , n231808 , 
 n231809 , n231810 , n231811 , n231812 , n231813 , n231814 , n231815 , n231816 , n231817 , n231818 , 
 n231819 , n231820 , n231821 , n231822 , n231823 , n231824 , n231825 , n231826 , n231827 , n231828 , 
 n231829 , n231830 , n231831 , n231832 , n231833 , n231834 , n231835 , n231836 , n231837 , n231838 , 
 n231839 , n231840 , n231841 , n231842 , n231843 , n231844 , n231845 , n231846 , n231847 , n231848 , 
 n231849 , n231850 , n231851 , n231852 , n231853 , n231854 , n231855 , n231856 , n231857 , n231858 , 
 n231859 , n231860 , n231861 , n231862 , n231863 , n231864 , n231865 , n231866 , n231867 , n231868 , 
 n231869 , n231870 , n231871 , n231872 , n231873 , n231874 , n231875 , n231876 , n231877 , n231878 , 
 n231879 , n231880 , n231881 , n231882 , n231883 , n231884 , n231885 , n231886 , n231887 , n231888 , 
 n231889 , n231890 , n231891 , n231892 , n231893 , n231894 , n231895 , n231896 , n231897 , n231898 , 
 n231899 , n231900 , n231901 , n231902 , n231903 , n231904 , n231905 , n231906 , n231907 , n231908 , 
 n231909 , n231910 , n231911 , n231912 , n231913 , n231914 , n231915 , n231916 , n231917 , n231918 , 
 n231919 , n231920 , n231921 , n231922 , n231923 , n231924 , n231925 , n231926 , n231927 , n231928 , 
 n231929 , n231930 , n231931 , n231932 , n231933 , n231934 , n231935 , n231936 , n231937 , n231938 , 
 n231939 , n231940 , n231941 , n231942 , n231943 , n231944 , n231945 , n231946 , n231947 , n231948 , 
 n231949 , n231950 , n231951 , n231952 , n231953 , n231954 , n231955 , n231956 , n231957 , n231958 , 
 n231959 , n231960 , n231961 , n231962 , n231963 , n231964 , n231965 , n231966 , n231967 , n231968 , 
 n231969 , n231970 , n231971 , n231972 , n231973 , n231974 , n231975 , n231976 , n231977 , n231978 , 
 n231979 , n231980 , n231981 , n231982 , n231983 , n231984 , n231985 , n231986 , n231987 , n231988 , 
 n231989 , n231990 , n231991 , n231992 , n231993 , n231994 , n231995 , n231996 , n231997 , n231998 , 
 n231999 , n232000 , n232001 , n232002 , n232003 , n232004 , n232005 , n232006 , n232007 , n232008 , 
 n232009 , n232010 , n232011 , n232012 , n232013 , n232014 , n232015 , n232016 , n232017 , n232018 , 
 n232019 , n232020 , n232021 , n232022 , n232023 , n232024 , n232025 , n232026 , n232027 , n232028 , 
 n232029 , n232030 , n232031 , n232032 , n232033 , n232034 , n232035 , n232036 , n232037 , n232038 , 
 n232039 , n232040 , n232041 , n232042 , n232043 , n232044 , n232045 , n232046 , n232047 , n232048 , 
 n232049 , n232050 , n232051 , n232052 , n232053 , n232054 , n232055 , n232056 , n232057 , n232058 , 
 n232059 , n232060 , n232061 , n232062 , n232063 , n232064 , n232065 , n232066 , n232067 , n232068 , 
 n232069 , n232070 , n232071 , n232072 , n232073 , n232074 , n232075 , n232076 , n232077 , n232078 , 
 n232079 , n232080 , n232081 , n232082 , n232083 , n232084 , n232085 , n232086 , n232087 , n232088 , 
 n232089 , n232090 , n232091 , n232092 , n232093 , n232094 , n232095 , n232096 , n232097 , n232098 , 
 n232099 , n232100 , n232101 , n232102 , n232103 , n232104 , n232105 , n232106 , n232107 , n232108 , 
 n232109 , n232110 , n232111 , n232112 , n232113 , n232114 , n232115 , n232116 , n232117 , n232118 , 
 n232119 , n232120 , n232121 , n232122 , n232123 , n232124 , n232125 , n232126 , n232127 , n232128 , 
 n232129 , n232130 , n232131 , n232132 , n232133 , n232134 , n232135 , n232136 , n232137 , n232138 , 
 n232139 , n232140 , n232141 , n232142 , n232143 , n232144 , n232145 , n232146 , n232147 , n232148 , 
 n232149 , n232150 , n232151 , n232152 , n232153 , n232154 , n232155 , n232156 , n232157 , n232158 , 
 n232159 , n232160 , n232161 , n232162 , n232163 , n232164 , n232165 , n232166 , n232167 , n232168 , 
 n232169 , n232170 , n232171 , n232172 , n232173 , n232174 , n232175 , n232176 , n232177 , n232178 , 
 n232179 , n232180 , n232181 , n232182 , n232183 , n232184 , n232185 , n232186 , n232187 , n232188 , 
 n232189 , n232190 , n232191 , n232192 , n232193 , n232194 , n232195 , n232196 , n232197 , n232198 , 
 n232199 , n232200 , n232201 , n232202 , n232203 , n232204 , n232205 , n232206 , n232207 , n232208 , 
 n232209 , n232210 , n232211 , n232212 , n232213 , n232214 , n232215 , n232216 , n232217 , n232218 , 
 n232219 , n232220 , n232221 , n232222 , n232223 , n232224 , n232225 , n232226 , n232227 , n232228 , 
 n232229 , n232230 , n232231 , n232232 , n232233 , n232234 , n232235 , n232236 , n232237 , n232238 , 
 n232239 , n232240 , n232241 , n232242 , n232243 , n232244 , n232245 , n232246 , n232247 , n232248 , 
 n232249 , n232250 , n232251 , n232252 , n232253 , n232254 , n232255 , n232256 , n232257 , n232258 , 
 n232259 , n232260 , n232261 , n232262 , n232263 , n232264 , n232265 , n232266 , n232267 , n232268 , 
 n232269 , n232270 , n232271 , n232272 , n232273 , n232274 , n232275 , n232276 , n232277 , n232278 , 
 n232279 , n232280 , n232281 , n232282 , n232283 , n232284 , n232285 , n232286 , n232287 , n232288 , 
 n232289 , n232290 , n232291 , n232292 , n232293 , n232294 , n232295 , n232296 , n232297 , n232298 , 
 n232299 , n232300 , n232301 , n232302 , n232303 , n232304 , n232305 , n232306 , n232307 , n232308 , 
 n232309 , n232310 , n232311 , n232312 , n232313 , n232314 , n232315 , n232316 , n232317 , n232318 , 
 n232319 , n232320 , n232321 , n232322 , n232323 , n232324 , n232325 , n232326 , n232327 , n232328 , 
 n232329 , n232330 , n232331 , n232332 , n232333 , n232334 , n232335 , n232336 , n232337 , n232338 , 
 n232339 , n232340 , n232341 , n232342 , n232343 , n232344 , n232345 , n232346 , n232347 , n232348 , 
 n232349 , n232350 , n232351 , n232352 , n232353 , n232354 , n232355 , n232356 , n232357 , n232358 , 
 n232359 , n232360 , n232361 , n232362 , n232363 , n232364 , n232365 , n232366 , n232367 , n232368 , 
 n232369 , n232370 , n232371 , n232372 , n232373 , n232374 , n232375 , n232376 , n232377 , n232378 , 
 n232379 , n232380 , n232381 , n232382 , n232383 , n232384 , n232385 , n232386 , n232387 , n232388 , 
 n232389 , n232390 , n232391 , n232392 , n232393 , n232394 , n232395 , n232396 , n232397 , n232398 , 
 n232399 , n232400 , n232401 , n232402 , n232403 , n232404 , n232405 , n232406 , n232407 , n232408 , 
 n232409 , n232410 , n232411 , n232412 , n232413 , n232414 , n232415 , n232416 , n232417 , n232418 , 
 n232419 , n232420 , n232421 , n232422 , n232423 , n232424 , n232425 , n232426 , n232427 , n232428 , 
 n232429 , n232430 , n232431 , n232432 , n232433 , n232434 , n232435 , n232436 , n232437 , n232438 , 
 n232439 , n232440 , n232441 , n232442 , n232443 , n232444 , n232445 , n232446 , n232447 , n232448 , 
 n232449 , n232450 , n232451 , n232452 , n232453 , n232454 , n232455 , n232456 , n232457 , n232458 , 
 n232459 , n232460 , n232461 , n232462 , n232463 , n232464 , n232465 , n232466 , n232467 , n232468 , 
 n232469 , n232470 , n232471 , n232472 , n232473 , n232474 , n232475 , n232476 , n232477 , n232478 , 
 n232479 , n232480 , n232481 , n232482 , n232483 , n232484 , n232485 , n232486 , n232487 , n232488 , 
 n232489 , n232490 , n232491 , n232492 , n232493 , n232494 , n232495 , n232496 , n232497 , n232498 , 
 n232499 , n232500 , n232501 , n232502 , n232503 , n232504 , n232505 , n232506 , n232507 , n232508 , 
 n232509 , n232510 , n232511 , n232512 , n232513 , n232514 , n232515 , n232516 , n232517 , n232518 , 
 n232519 , n232520 , n232521 , n232522 , n232523 , n232524 , n232525 , n232526 , n232527 , n232528 , 
 n232529 , n232530 , n232531 , n232532 , n232533 , n232534 , n232535 , n232536 , n232537 , n232538 , 
 n232539 , n232540 , n232541 , n232542 , n232543 , n232544 , n232545 , n232546 , n232547 , n232548 , 
 n232549 , n232550 , n232551 , n232552 , n232553 , n232554 , n232555 , n232556 , n232557 , n232558 , 
 n232559 , n232560 , n232561 , n232562 , n232563 , n232564 , n232565 , n232566 , n232567 , n232568 , 
 n232569 , n232570 , n232571 , n232572 , n232573 , n232574 , n232575 , n232576 , n232577 , n232578 , 
 n232579 , n232580 , n232581 , n232582 , n232583 , n232584 , n232585 , n232586 , n232587 , n232588 , 
 n232589 , n232590 , n232591 , n232592 , n232593 , n232594 , n232595 , n232596 , n232597 , n232598 , 
 n232599 , n232600 , n232601 , n232602 , n232603 , n232604 , n232605 , n232606 , n232607 , n232608 , 
 n232609 , n232610 , n232611 , n232612 , n232613 , n232614 , n232615 , n232616 , n232617 , n232618 , 
 n232619 , n232620 , n232621 , n232622 , n232623 , n232624 , n232625 , n232626 , n232627 , n232628 , 
 n232629 , n232630 , n232631 , n232632 , n232633 , n232634 , n232635 , n232636 , n232637 , n232638 , 
 n232639 , n232640 , n232641 , n232642 , n232643 , n232644 , n232645 , n232646 , n232647 , n232648 , 
 n232649 , n232650 , n232651 , n232652 , n232653 , n232654 , n232655 , n232656 , n232657 , n232658 , 
 n232659 , n232660 , n232661 , n232662 , n232663 , n232664 , n232665 , n232666 , n232667 , n232668 , 
 n232669 , n232670 , n232671 , n232672 , n232673 , n232674 , n232675 , n232676 , n232677 , n232678 , 
 n232679 , n232680 , n232681 , n232682 , n232683 , n232684 , n232685 , n232686 , n232687 , n232688 , 
 n232689 , n232690 , n232691 , n232692 , n232693 , n232694 , n232695 , n232696 , n232697 , n232698 , 
 n232699 , n232700 , n232701 , n232702 , n232703 , n232704 , n232705 , n232706 , n232707 , n232708 , 
 n232709 , n232710 , n232711 , n232712 , n232713 , n232714 , n232715 , n232716 , n232717 , n232718 , 
 n232719 , n232720 , n232721 , n232722 , n232723 , n232724 , n232725 , n232726 , n232727 , n232728 , 
 n232729 , n232730 , n232731 , n232732 , n232733 , n232734 , n232735 , n232736 , n232737 , n232738 , 
 n232739 , n232740 , n232741 , n232742 , n232743 , n232744 , n232745 , n232746 , n232747 , n232748 , 
 n232749 , n232750 , n232751 , n232752 , n232753 , n232754 , n232755 , n232756 , n232757 , n232758 , 
 n232759 , n232760 , n232761 , n232762 , n232763 , n232764 , n232765 , n232766 , n232767 , n232768 , 
 n232769 , n232770 , n232771 , n232772 , n232773 , n232774 , n232775 , n232776 , n232777 , n232778 , 
 n232779 , n232780 , n232781 , n232782 , n232783 , n232784 , n232785 , n232786 , n232787 , n232788 , 
 n232789 , n232790 , n232791 , n232792 , n232793 , n232794 , n232795 , n232796 , n232797 , n232798 , 
 n232799 , n232800 , n232801 , n232802 , n232803 , n232804 , n232805 , n232806 , n232807 , n232808 , 
 n232809 , n232810 , n232811 , n232812 , n232813 , n232814 , n232815 , n232816 , n232817 , n232818 , 
 n232819 , n232820 , n232821 , n232822 , n232823 , n232824 , n232825 , n232826 , n232827 , n232828 , 
 n232829 , n232830 , n232831 , n232832 , n232833 , n232834 , n232835 , n232836 , n232837 , n232838 , 
 n232839 , n232840 , n232841 , n232842 , n232843 , n232844 , n232845 , n232846 , n232847 , n232848 , 
 n232849 , n232850 , n232851 , n232852 , n232853 , n232854 , n232855 , n232856 , n232857 , n232858 , 
 n232859 , n232860 , n232861 , n232862 , n232863 , n232864 , n232865 , n232866 , n232867 , n232868 , 
 n232869 , n232870 , n232871 , n232872 , n232873 , n232874 , n232875 , n232876 , n232877 , n232878 , 
 n232879 , n232880 , n232881 , n232882 , n232883 , n232884 , n232885 , n232886 , n232887 , n232888 , 
 n232889 , n232890 , n232891 , n232892 , n232893 , n232894 , n232895 , n232896 , n232897 , n232898 , 
 n232899 , n232900 , n232901 , n232902 , n232903 , n232904 , n232905 , n232906 , n232907 , n232908 , 
 n232909 , n232910 , n232911 , n232912 , n232913 , n232914 , n232915 , n232916 , n232917 , n232918 , 
 n232919 , n232920 , n232921 , n232922 , n232923 , n232924 , n232925 , n232926 , n232927 , n232928 , 
 n232929 , n232930 , n232931 , n232932 , n232933 , n232934 , n232935 , n232936 , n232937 , n232938 , 
 n232939 , n232940 , n232941 , n232942 , n232943 , n232944 , n232945 , n232946 , n232947 , n232948 , 
 n232949 , n232950 , n232951 , n232952 , n232953 , n232954 , n232955 , n232956 , n232957 , n232958 , 
 n232959 , n232960 , n232961 , n232962 , n232963 , n232964 , n232965 , n232966 , n232967 , n232968 , 
 n232969 , n232970 , n232971 , n232972 , n232973 , n232974 , n232975 , n232976 , n232977 , n232978 , 
 n232979 , n232980 , n232981 , n232982 , n232983 , n232984 , n232985 , n232986 , n232987 , n232988 , 
 n232989 , n232990 , n232991 , n232992 , n232993 , n232994 , n232995 , n232996 , n232997 , n232998 , 
 n232999 , n233000 , n233001 , n233002 , n233003 , n233004 , n233005 , n233006 , n233007 , n233008 , 
 n233009 , n233010 , n233011 , n233012 , n233013 , n233014 , n233015 , n233016 , n233017 , n233018 , 
 n233019 , n233020 , n233021 , n233022 , n233023 , n233024 , n233025 , n233026 , n233027 , n233028 , 
 n233029 , n233030 , n233031 , n233032 , n233033 , n233034 , n233035 , n233036 , n233037 , n233038 , 
 n233039 , n233040 , n233041 , n233042 , n233043 , n233044 , n233045 , n233046 , n233047 , n233048 , 
 n233049 , n233050 , n233051 , n233052 , n233053 , n233054 , n233055 , n233056 , n233057 , n233058 , 
 n233059 , n233060 , n233061 , n233062 , n233063 , n233064 , n233065 , n233066 , n233067 , n233068 , 
 n233069 , n233070 , n233071 , n233072 , n233073 , n233074 , n233075 , n233076 , n233077 , n233078 , 
 n233079 , n233080 , n233081 , n233082 , n233083 , n233084 , n233085 , n233086 , n233087 , n233088 , 
 n233089 , n233090 , n233091 , n233092 , n233093 , n233094 , n233095 , n233096 , n233097 , n233098 , 
 n233099 , n233100 , n233101 , n233102 , n233103 , n233104 , n233105 , n233106 , n233107 , n233108 , 
 n233109 , n233110 , n233111 , n233112 , n233113 , n233114 , n233115 , n233116 , n233117 , n233118 , 
 n233119 , n233120 , n233121 , n233122 , n233123 , n233124 , n233125 , n233126 , n233127 , n233128 , 
 n233129 , n233130 , n233131 , n233132 , n233133 , n233134 , n233135 , n233136 , n233137 , n233138 , 
 n233139 , n233140 , n233141 , n233142 , n233143 , n233144 , n233145 , n233146 , n233147 , n233148 , 
 n233149 , n233150 , n233151 , n233152 , n233153 , n233154 , n233155 , n233156 , n233157 , n233158 , 
 n233159 , n233160 , n233161 , n233162 , n233163 , n233164 , n233165 , n233166 , n233167 , n233168 , 
 n233169 , n233170 , n233171 , n233172 , n233173 , n233174 , n233175 , n233176 , n233177 , n233178 , 
 n233179 , n233180 , n233181 , n233182 , n233183 , n233184 , n233185 , n233186 , n233187 , n233188 , 
 n233189 , n233190 , n233191 , n233192 , n233193 , n233194 , n233195 , n233196 , n233197 , n233198 , 
 n233199 , n233200 , n233201 , n233202 , n233203 , n233204 , n233205 , n233206 , n233207 , n233208 , 
 n233209 , n233210 , n233211 , n233212 , n233213 , n233214 , n233215 , n233216 , n233217 , n233218 , 
 n233219 , n233220 , n233221 , n233222 , n233223 , n233224 , n233225 , n233226 , n233227 , n233228 , 
 n233229 , n233230 , n233231 , n233232 , n233233 , n233234 , n233235 , n233236 , n233237 , n233238 , 
 n233239 , n233240 , n233241 , n233242 , n233243 , n233244 , n233245 , n233246 , n233247 , n233248 , 
 n233249 , n233250 , n233251 , n233252 , n233253 , n233254 , n233255 , n233256 , n233257 , n233258 , 
 n233259 , n233260 , n233261 , n233262 , n233263 , n233264 , n233265 , n233266 , n233267 , n233268 , 
 n233269 , n233270 , n233271 , n233272 , n233273 , n233274 , n233275 , n233276 , n233277 , n233278 , 
 n233279 , n233280 , n233281 , n233282 , n233283 , n233284 , n233285 , n233286 , n233287 , n233288 , 
 n233289 , n233290 , n233291 , n233292 , n233293 , n233294 , n233295 , n233296 , n233297 , n233298 , 
 n233299 , n233300 , n233301 , n233302 , n233303 , n233304 , n233305 , n233306 , n233307 , n233308 , 
 n233309 , n233310 , n233311 , n233312 , n233313 , n233314 , n233315 , n233316 , n233317 , n233318 , 
 n233319 , n233320 , n233321 , n233322 , n233323 , n233324 , n233325 , n233326 , n233327 , n233328 , 
 n233329 , n233330 , n233331 , n233332 , n233333 , n233334 , n233335 , n233336 , n233337 , n233338 , 
 n233339 , n233340 , n233341 , n233342 , n233343 , n233344 , n233345 , n233346 , n233347 , n233348 , 
 n233349 , n233350 , n233351 , n233352 , n233353 , n233354 , n233355 , n233356 , n233357 , n233358 , 
 n233359 , n233360 , n233361 , n233362 , n233363 , n233364 , n233365 , n233366 , n233367 , n233368 , 
 n233369 , n233370 , n233371 , n233372 , n233373 , n233374 , n233375 , n233376 , n233377 , n233378 , 
 n233379 , n233380 , n233381 , n233382 , n233383 , n233384 , n233385 , n233386 , n233387 , n233388 , 
 n233389 , n233390 , n233391 , n233392 , n233393 , n233394 , n233395 , n233396 , n233397 , n233398 , 
 n233399 , n233400 , n233401 , n233402 , n233403 , n233404 , n233405 , n233406 , n233407 , n233408 , 
 n233409 , n233410 , n233411 , n233412 , n233413 , n233414 , n233415 , n233416 , n233417 , n233418 , 
 n233419 , n233420 , n233421 , n233422 , n233423 , n233424 , n233425 , n233426 , n233427 , n233428 , 
 n233429 , n233430 , n233431 , n233432 , n233433 , n233434 , n233435 , n233436 , n233437 , n233438 , 
 n233439 , n233440 , n233441 , n233442 , n233443 , n233444 , n233445 , n233446 , n233447 , n233448 , 
 n233449 , n233450 , n233451 , n233452 , n233453 , n233454 , n233455 , n233456 , n233457 , n233458 , 
 n233459 , n233460 , n233461 , n233462 , n233463 , n233464 , n233465 , n233466 , n233467 , n233468 , 
 n233469 , n233470 , n233471 , n233472 , n233473 , n233474 , n233475 , n233476 , n233477 , n233478 , 
 n233479 , n233480 , n233481 , n233482 , n233483 , n233484 , n233485 , n233486 , n233487 , n233488 , 
 n233489 , n233490 , n233491 , n233492 , n233493 , n233494 , n233495 , n233496 , n233497 , n233498 , 
 n233499 , n233500 , n233501 , n233502 , n233503 , n233504 , n233505 , n233506 , n233507 , n233508 , 
 n233509 , n233510 , n233511 , n233512 , n233513 , n233514 , n233515 , n233516 , n233517 , n233518 , 
 n233519 , n233520 , n233521 , n233522 , n233523 , n233524 , n233525 , n233526 , n233527 , n233528 , 
 n233529 , n233530 , n233531 , n233532 , n233533 , n233534 , n233535 , n233536 , n233537 , n233538 , 
 n233539 , n233540 , n233541 , n233542 , n233543 , n233544 , n233545 , n233546 , n233547 , n233548 , 
 n233549 , n233550 , n233551 , n233552 , n233553 , n233554 , n233555 , n233556 , n233557 , n233558 , 
 n233559 , n233560 , n233561 , n233562 , n233563 , n233564 , n233565 , n233566 , n233567 , n233568 , 
 n233569 , n233570 , n233571 , n233572 , n233573 , n233574 , n233575 , n233576 , n233577 , n233578 , 
 n233579 , n233580 , n233581 , n233582 , n233583 , n233584 , n233585 , n233586 , n233587 , n233588 , 
 n233589 , n233590 , n233591 , n233592 , n233593 , n233594 , n233595 , n233596 , n233597 , n233598 , 
 n233599 , n233600 , n233601 , n233602 , n233603 , n233604 , n233605 , n233606 , n233607 , n233608 , 
 n233609 , n233610 , n233611 , n233612 , n233613 , n233614 , n233615 , n233616 , n233617 , n233618 , 
 n233619 , n233620 , n233621 , n233622 , n233623 , n233624 , n233625 , n233626 , n233627 , n233628 , 
 n233629 , n233630 , n233631 , n233632 , n233633 , n233634 , n233635 , n233636 , n233637 , n233638 , 
 n233639 , n233640 , n233641 , n233642 , n233643 , n233644 , n233645 , n233646 , n233647 , n233648 , 
 n233649 , n233650 , n233651 , n233652 , n233653 , n233654 , n233655 , n233656 , n233657 , n233658 , 
 n233659 , n233660 , n233661 , n233662 , n233663 , n233664 , n233665 , n233666 , n233667 , n233668 , 
 n233669 , n233670 , n233671 , n233672 , n233673 , n233674 , n233675 , n233676 , n233677 , n233678 , 
 n233679 , n233680 , n233681 , n233682 , n233683 , n233684 , n233685 , n233686 , n233687 , n233688 , 
 n233689 , n233690 , n233691 , n233692 , n233693 , n233694 , n233695 , n233696 , n233697 , n233698 , 
 n233699 , n233700 , n233701 , n233702 , n233703 , n233704 , n233705 , n233706 , n233707 , n233708 , 
 n233709 , n233710 , n233711 , n233712 , n233713 , n233714 , n233715 , n233716 , n233717 , n233718 , 
 n233719 , n233720 , n233721 , n233722 , n233723 , n233724 , n233725 , n233726 , n233727 , n233728 , 
 n233729 , n233730 , n233731 , n233732 , n233733 , n233734 , n233735 , n233736 , n233737 , n233738 , 
 n233739 , n233740 , n233741 , n233742 , n233743 , n233744 , n233745 , n233746 , n233747 , n233748 , 
 n233749 , n233750 , n233751 , n233752 , n233753 , n233754 , n233755 , n233756 , n233757 , n233758 , 
 n233759 , n233760 , n233761 , n233762 , n233763 , n233764 , n233765 , n233766 , n233767 , n233768 , 
 n233769 , n233770 , n233771 , n233772 , n233773 , n233774 , n233775 , n233776 , n233777 , n233778 , 
 n233779 , n233780 , n233781 , n233782 , n233783 , n233784 , n233785 , n233786 , n233787 , n233788 , 
 n233789 , n233790 , n233791 , n233792 , n233793 , n233794 , n233795 , n233796 , n233797 , n233798 , 
 n233799 , n233800 , n233801 , n233802 , n233803 , n233804 , n233805 , n233806 , n233807 , n233808 , 
 n233809 , n233810 , n233811 , n233812 , n233813 , n233814 , n233815 , n233816 , n233817 , n233818 , 
 n233819 , n233820 , n233821 , n233822 , n233823 , n233824 , n233825 , n233826 , n233827 , n233828 , 
 n233829 , n233830 , n233831 , n233832 , n233833 , n233834 , n233835 , n233836 , n233837 , n233838 , 
 n233839 , n233840 , n233841 , n233842 , n233843 , n233844 , n233845 , n233846 , n233847 , n233848 , 
 n233849 , n233850 , n233851 , n233852 , n233853 , n233854 , n233855 , n233856 , n233857 , n233858 , 
 n233859 , n233860 , n233861 , n233862 , n233863 , n233864 , n233865 , n233866 , n233867 , n233868 , 
 n233869 , n233870 , n233871 , n233872 , n233873 , n233874 , n233875 , n233876 , n233877 , n233878 , 
 n233879 , n233880 , n233881 , n233882 , n233883 , n233884 , n233885 , n233886 , n233887 , n233888 , 
 n233889 , n233890 , n233891 , n233892 , n233893 , n233894 , n233895 , n233896 , n233897 , n233898 , 
 n233899 , n233900 , n233901 , n233902 , n233903 , n233904 , n233905 , n233906 , n233907 , n233908 , 
 n233909 , n233910 , n233911 , n233912 , n233913 , n233914 , n233915 , n233916 , n233917 , n233918 , 
 n233919 , n233920 , n233921 , n233922 , n233923 , n233924 , n233925 , n233926 , n233927 , n233928 , 
 n233929 , n233930 , n233931 , n233932 , n233933 , n233934 , n233935 , n233936 , n233937 , n233938 , 
 n233939 , n233940 , n233941 , n233942 , n233943 , n233944 , n233945 , n233946 , n233947 , n233948 , 
 n233949 , n233950 , n233951 , n233952 , n233953 , n233954 , n233955 , n233956 , n233957 , n233958 , 
 n233959 , n233960 , n233961 , n233962 , n233963 , n233964 , n233965 , n233966 , n233967 , n233968 , 
 n233969 , n233970 , n233971 , n233972 , n233973 , n233974 , n233975 , n233976 , n233977 , n233978 , 
 n233979 , n233980 , n233981 , n233982 , n233983 , n233984 , n233985 , n233986 , n233987 , n233988 , 
 n233989 , n233990 , n233991 , n233992 , n233993 , n233994 , n233995 , n233996 , n233997 , n233998 , 
 n233999 , n234000 , n234001 , n234002 , n234003 , n234004 , n234005 , n234006 , n234007 , n234008 , 
 n234009 , n234010 , n234011 , n234012 , n234013 , n234014 , n234015 , n234016 , n234017 , n234018 , 
 n234019 , n234020 , n234021 , n234022 , n234023 , n234024 , n234025 , n234026 , n234027 , n234028 , 
 n234029 , n234030 , n234031 , n234032 , n234033 , n234034 , n234035 , n234036 , n234037 , n234038 , 
 n234039 , n234040 , n234041 , n234042 , n234043 , n234044 , n234045 , n234046 , n234047 , n234048 , 
 n234049 , n234050 , n234051 , n234052 , n234053 , n234054 , n234055 , n234056 , n234057 , n234058 , 
 n234059 , n234060 , n234061 , n234062 , n234063 , n234064 , n234065 , n234066 , n234067 , n234068 , 
 n234069 , n234070 , n234071 , n234072 , n234073 , n234074 , n234075 , n234076 , n234077 , n234078 , 
 n234079 , n234080 , n234081 , n234082 , n234083 , n234084 , n234085 , n234086 , n234087 , n234088 , 
 n234089 , n234090 , n234091 , n234092 , n234093 , n234094 , n234095 , n234096 , n234097 , n234098 , 
 n234099 , n234100 , n234101 , n234102 , n234103 , n234104 , n234105 , n234106 , n234107 , n234108 , 
 n234109 , n234110 , n234111 , n234112 , n234113 , n234114 , n234115 , n234116 , n234117 , n234118 , 
 n234119 , n234120 , n234121 , n234122 , n234123 , n234124 , n234125 , n234126 , n234127 , n234128 , 
 n234129 , n234130 , n234131 , n234132 , n234133 , n234134 , n234135 , n234136 , n234137 , n234138 , 
 n234139 , n234140 , n234141 , n234142 , n234143 , n234144 , n234145 , n234146 , n234147 , n234148 , 
 n234149 , n234150 , n234151 , n234152 , n234153 , n234154 , n234155 , n234156 , n234157 , n234158 , 
 n234159 , n234160 , n234161 , n234162 , n234163 , n234164 , n234165 , n234166 , n234167 , n234168 , 
 n234169 , n234170 , n234171 , n234172 , n234173 , n234174 , n234175 , n234176 , n234177 , n234178 , 
 n234179 , n234180 , n234181 , n234182 , n234183 , n234184 , n234185 , n234186 , n234187 , n234188 , 
 n234189 , n234190 , n234191 , n234192 , n234193 , n234194 , n234195 , n234196 , n234197 , n234198 , 
 n234199 , n234200 , n234201 , n234202 , n234203 , n234204 , n234205 , n234206 , n234207 , n234208 , 
 n234209 , n234210 , n234211 , n234212 , n234213 , n234214 , n234215 , n234216 , n234217 , n234218 , 
 n234219 , n234220 , n234221 , n234222 , n234223 , n234224 , n234225 , n234226 , n234227 , n234228 , 
 n234229 , n234230 , n234231 , n234232 , n234233 , n234234 , n234235 , n234236 , n234237 , n234238 , 
 n234239 , n234240 , n234241 , n234242 , n234243 , n234244 , n234245 , n234246 , n234247 , n234248 , 
 n234249 , n234250 , n234251 , n234252 , n234253 , n234254 , n234255 , n234256 , n234257 , n234258 , 
 n234259 , n234260 , n234261 , n234262 , n234263 , n234264 , n234265 , n234266 , n234267 , n234268 , 
 n234269 , n234270 , n234271 , n234272 , n234273 , n234274 , n234275 , n234276 , n234277 , n234278 , 
 n234279 , n234280 , n234281 , n234282 , n234283 , n234284 , n234285 , n234286 , n234287 , n234288 , 
 n234289 , n234290 , n234291 , n234292 , n234293 , n234294 , n234295 , n234296 , n234297 , n234298 , 
 n234299 , n234300 , n234301 , n234302 , n234303 , n234304 , n234305 , n234306 , n234307 , n234308 , 
 n234309 , n234310 , n234311 , n234312 , n234313 , n234314 , n234315 , n234316 , n234317 , n234318 , 
 n234319 , n234320 , n234321 , n234322 , n234323 , n234324 , n234325 , n234326 , n234327 , n234328 , 
 n234329 , n234330 , n234331 , n234332 , n234333 , n234334 , n234335 , n234336 , n234337 , n234338 , 
 n234339 , n234340 , n234341 , n234342 , n234343 , n234344 , n234345 , n234346 , n234347 , n234348 , 
 n234349 , n234350 , n234351 , n234352 , n234353 , n234354 , n234355 , n234356 , n234357 , n234358 , 
 n234359 , n234360 , n234361 , n234362 , n234363 , n234364 , n234365 , n234366 , n234367 , n234368 , 
 n234369 , n234370 , n234371 , n234372 , n234373 , n234374 , n234375 , n234376 , n234377 , n234378 , 
 n234379 , n234380 , n234381 , n234382 , n234383 , n234384 , n234385 , n234386 , n234387 , n234388 , 
 n234389 , n234390 , n234391 , n234392 , n234393 , n234394 , n234395 , n234396 , n234397 , n234398 , 
 n234399 , n234400 , n234401 , n234402 , n234403 , n234404 , n234405 , n234406 , n234407 , n234408 , 
 n234409 , n234410 , n234411 , n234412 , n234413 , n234414 , n234415 , n234416 , n234417 , n234418 , 
 n234419 , n234420 , n234421 , n234422 , n234423 , n234424 , n234425 , n234426 , n234427 , n234428 , 
 n234429 , n234430 , n234431 , n234432 , n234433 , n234434 , n234435 , n234436 , n234437 , n234438 , 
 n234439 , n234440 , n234441 , n234442 , n234443 , n234444 , n234445 , n234446 , n234447 , n234448 , 
 n234449 , n234450 , n234451 , n234452 , n234453 , n234454 , n234455 , n234456 , n234457 , n234458 , 
 n234459 , n234460 , n234461 , n234462 , n234463 , n234464 , n234465 , n234466 , n234467 , n234468 , 
 n234469 , n234470 , n234471 , n234472 , n234473 , n234474 , n234475 , n234476 , n234477 , n234478 , 
 n234479 , n234480 , n234481 , n234482 , n234483 , n234484 , n234485 , n234486 , n234487 , n234488 , 
 n234489 , n234490 , n234491 , n234492 , n234493 , n234494 , n234495 , n234496 , n234497 , n234498 , 
 n234499 , n234500 , n234501 , n234502 , n234503 , n234504 , n234505 , n234506 , n234507 , n234508 , 
 n234509 , n234510 , n234511 , n234512 , n234513 , n234514 , n234515 , n234516 , n234517 , n234518 , 
 n234519 , n234520 , n234521 , n234522 , n234523 , n234524 , n234525 , n234526 , n234527 , n234528 , 
 n234529 , n234530 , n234531 , n234532 , n234533 , n234534 , n234535 , n234536 , n234537 , n234538 , 
 n234539 , n234540 , n234541 , n234542 , n234543 , n234544 , n234545 , n234546 , n234547 , n234548 , 
 n234549 , n234550 , n234551 , n234552 , n234553 , n234554 , n234555 , n234556 , n234557 , n234558 , 
 n234559 , n234560 , n234561 , n234562 , n234563 , n234564 , n234565 , n234566 , n234567 , n234568 , 
 n234569 , n234570 , n234571 , n234572 , n234573 , n234574 , n234575 , n234576 , n234577 , n234578 , 
 n234579 , n234580 , n234581 , n234582 , n234583 , n234584 , n234585 , n234586 , n234587 , n234588 , 
 n234589 , n234590 , n234591 , n234592 , n234593 , n234594 , n234595 , n234596 , n234597 , n234598 , 
 n234599 , n234600 , n234601 , n234602 , n234603 , n234604 , n234605 , n234606 , n234607 , n234608 , 
 n234609 , n234610 , n234611 , n234612 , n234613 , n234614 , n234615 , n234616 , n234617 , n234618 , 
 n234619 , n234620 , n234621 , n234622 , n234623 , n234624 , n234625 , n234626 , n234627 , n234628 , 
 n234629 , n234630 , n234631 , n234632 , n234633 , n234634 , n234635 , n234636 , n234637 , n234638 , 
 n234639 , n234640 , n234641 , n234642 , n234643 , n234644 , n234645 , n234646 , n234647 , n234648 , 
 n234649 , n234650 , n234651 , n234652 , n234653 , n234654 , n234655 , n234656 , n234657 , n234658 , 
 n234659 , n234660 , n234661 , n234662 , n234663 , n234664 , n234665 , n234666 , n234667 , n234668 , 
 n234669 , n234670 , n234671 , n234672 , n234673 , n234674 , n234675 , n234676 , n234677 , n234678 , 
 n234679 , n234680 , n234681 , n234682 , n234683 , n234684 , n234685 , n234686 , n234687 , n234688 , 
 n234689 , n234690 , n234691 , n234692 , n234693 , n234694 , n234695 , n234696 , n234697 , n234698 , 
 n234699 , n234700 , n234701 , n234702 , n234703 , n234704 , n234705 , n234706 , n234707 , n234708 , 
 n234709 , n234710 , n234711 , n234712 , n234713 , n234714 , n234715 , n234716 , n234717 , n234718 , 
 n234719 , n234720 , n234721 , n234722 , n234723 , n234724 , n234725 , n234726 , n234727 , n234728 , 
 n234729 , n234730 , n234731 , n234732 , n234733 , n234734 , n234735 , n234736 , n234737 , n234738 , 
 n234739 , n234740 , n234741 , n234742 , n234743 , n234744 , n234745 , n234746 , n234747 , n234748 , 
 n234749 , n234750 , n234751 , n234752 , n234753 , n234754 , n234755 , n234756 , n234757 , n234758 , 
 n234759 , n234760 , n234761 , n234762 , n234763 , n234764 , n234765 , n234766 , n234767 , n234768 , 
 n234769 , n234770 , n234771 , n234772 , n234773 , n234774 , n234775 , n234776 , n234777 , n234778 , 
 n234779 , n234780 , n234781 , n234782 , n234783 , n234784 , n234785 , n234786 , n234787 , n234788 , 
 n234789 , n234790 , n234791 , n234792 , n234793 , n234794 , n234795 , n234796 , n234797 , n234798 , 
 n234799 , n234800 , n234801 , n234802 , n234803 , n234804 , n234805 , n234806 , n234807 , n234808 , 
 n234809 , n234810 , n234811 , n234812 , n234813 , n234814 , n234815 , n234816 , n234817 , n234818 , 
 n234819 , n234820 , n234821 , n234822 , n234823 , n234824 , n234825 , n234826 , n234827 , n234828 , 
 n234829 , n234830 , n234831 , n234832 , n234833 , n234834 , n234835 , n234836 , n234837 , n234838 , 
 n234839 , n234840 , n234841 , n234842 , n234843 , n234844 , n234845 , n234846 , n234847 , n234848 , 
 n234849 , n234850 , n234851 , n234852 , n234853 , n234854 , n234855 , n234856 , n234857 , n234858 , 
 n234859 , n234860 , n234861 , n234862 , n234863 , n234864 , n234865 , n234866 , n234867 , n234868 , 
 n234869 , n234870 , n234871 , n234872 , n234873 , n234874 , n234875 , n234876 , n234877 , n234878 , 
 n234879 , n234880 , n234881 , n234882 , n234883 , n234884 , n234885 , n234886 , n234887 , n234888 , 
 n234889 , n234890 , n234891 , n234892 , n234893 , n234894 , n234895 , n234896 , n234897 , n234898 , 
 n234899 , n234900 , n234901 , n234902 , n234903 , n234904 , n234905 , n234906 , n234907 , n234908 , 
 n234909 , n234910 , n234911 , n234912 , n234913 , n234914 , n234915 , n234916 , n234917 , n234918 , 
 n234919 , n234920 , n234921 , n234922 , n234923 , n234924 , n234925 , n234926 , n234927 , n234928 , 
 n234929 , n234930 , n234931 , n234932 , n234933 , n234934 , n234935 , n234936 , n234937 , n234938 , 
 n234939 , n234940 , n234941 , n234942 , n234943 , n234944 , n234945 , n234946 , n234947 , n234948 , 
 n234949 , n234950 , n234951 , n234952 , n234953 , n234954 , n234955 , n234956 , n234957 , n234958 , 
 n234959 , n234960 , n234961 , n234962 , n234963 , n234964 , n234965 , n234966 , n234967 , n234968 , 
 n234969 , n234970 , n234971 , n234972 , n234973 , n234974 , n234975 , n234976 , n234977 , n234978 , 
 n234979 , n234980 , n234981 , n234982 , n234983 , n234984 , n234985 , n234986 , n234987 , n234988 , 
 n234989 , n234990 , n234991 , n234992 , n234993 , n234994 , n234995 , n234996 , n234997 , n234998 , 
 n234999 , n235000 , n235001 , n235002 , n235003 , n235004 , n235005 , n235006 , n235007 , n235008 , 
 n235009 , n235010 , n235011 , n235012 , n235013 , n235014 , n235015 , n235016 , n235017 , n235018 , 
 n235019 , n235020 , n235021 , n235022 , n235023 , n235024 , n235025 , n235026 , n235027 , n235028 , 
 n235029 , n235030 , n235031 , n235032 , n235033 , n235034 , n235035 , n235036 , n235037 , n235038 , 
 n235039 , n235040 , n235041 , n235042 , n235043 , n235044 , n235045 , n235046 , n235047 , n235048 , 
 n235049 , n235050 , n235051 , n235052 , n235053 , n235054 , n235055 , n235056 , n235057 , n235058 , 
 n235059 , n235060 , n235061 , n235062 , n235063 , n235064 , n235065 , n235066 , n235067 , n235068 , 
 n235069 , n235070 , n235071 , n235072 , n235073 , n235074 , n235075 , n235076 , n235077 , n235078 , 
 n235079 , n235080 , n235081 , n235082 , n235083 , n235084 , n235085 , n235086 , n235087 , n235088 , 
 n235089 , n235090 , n235091 , n235092 , n235093 , n235094 , n235095 , n235096 , n235097 , n235098 , 
 n235099 , n235100 , n235101 , n235102 , n235103 , n235104 , n235105 , n235106 , n235107 , n235108 , 
 n235109 , n235110 , n235111 , n235112 , n235113 , n235114 , n235115 , n235116 , n235117 , n235118 , 
 n235119 , n235120 , n235121 , n235122 , n235123 , n235124 , n235125 , n235126 , n235127 , n235128 , 
 n235129 , n235130 , n235131 , n235132 , n235133 , n235134 , n235135 , n235136 , n235137 , n235138 , 
 n235139 , n235140 , n235141 , n235142 , n235143 , n235144 , n235145 , n235146 , n235147 , n235148 , 
 n235149 , n235150 , n235151 , n235152 , n235153 , n235154 , n235155 , n235156 , n235157 , n235158 , 
 n235159 , n235160 , n235161 , n235162 , n235163 , n235164 , n235165 , n235166 , n235167 , n235168 , 
 n235169 , n235170 , n235171 , n235172 , n235173 , n235174 , n235175 , n235176 , n235177 , n235178 , 
 n235179 , n235180 , n235181 , n235182 , n235183 , n235184 , n235185 , n235186 , n235187 , n235188 , 
 n235189 , n235190 , n235191 , n235192 , n235193 , n235194 , n235195 , n235196 , n235197 , n235198 , 
 n235199 , n235200 , n235201 , n235202 , n235203 , n235204 , n235205 , n235206 , n235207 , n235208 , 
 n235209 , n235210 , n235211 , n235212 , n235213 , n235214 , n235215 , n235216 , n235217 , n235218 , 
 n235219 , n235220 , n235221 , n235222 , n235223 , n235224 , n235225 , n235226 , n235227 , n235228 , 
 n235229 , n235230 , n235231 , n235232 , n235233 , n235234 , n235235 , n235236 , n235237 , n235238 , 
 n235239 , n235240 , n235241 , n235242 , n235243 , n235244 , n235245 , n235246 , n235247 , n235248 , 
 n235249 , n235250 , n235251 , n235252 , n235253 , n235254 , n235255 , n235256 , n235257 , n235258 , 
 n235259 , n235260 , n235261 , n235262 , n235263 , n235264 , n235265 , n235266 , n235267 , n235268 , 
 n235269 , n235270 , n235271 , n235272 , n235273 , n235274 , n235275 , n235276 , n235277 , n235278 , 
 n235279 , n235280 , n235281 , n235282 , n235283 , n235284 , n235285 , n235286 , n235287 , n235288 , 
 n235289 , n235290 , n235291 , n235292 , n235293 , n235294 , n235295 , n235296 , n235297 , n235298 , 
 n235299 , n235300 , n235301 , n235302 , n235303 , n235304 , n235305 , n235306 , n235307 , n235308 , 
 n235309 , n235310 , n235311 , n235312 , n235313 , n235314 , n235315 , n235316 , n235317 , n235318 , 
 n235319 , n235320 , n235321 , n235322 , n235323 , n235324 , n235325 , n235326 , n235327 , n235328 , 
 n235329 , n235330 , n235331 , n235332 , n235333 , n235334 , n235335 , n235336 , n235337 , n235338 , 
 n235339 , n235340 , n235341 , n235342 , n235343 , n235344 , n235345 , n235346 , n235347 , n235348 , 
 n235349 , n235350 , n235351 , n235352 , n235353 , n235354 , n235355 , n235356 , n235357 , n235358 , 
 n235359 , n235360 , n235361 , n235362 , n235363 , n235364 , n235365 , n235366 , n235367 , n235368 , 
 n235369 , n235370 , n235371 , n235372 , n235373 , n235374 , n235375 , n235376 , n235377 , n235378 , 
 n235379 , n235380 , n235381 , n235382 , n235383 , n235384 , n235385 , n235386 , n235387 , n235388 , 
 n235389 , n235390 , n235391 , n235392 , n235393 , n235394 , n235395 , n235396 , n235397 , n235398 , 
 n235399 , n235400 , n235401 , n235402 , n235403 , n235404 , n235405 , n235406 , n235407 , n235408 , 
 n235409 , n235410 , n235411 , n235412 , n235413 , n235414 , n235415 , n235416 , n235417 , n235418 , 
 n235419 , n235420 , n235421 , n235422 , n235423 , n235424 , n235425 , n235426 , n235427 , n235428 , 
 n235429 , n235430 , n235431 , n235432 , n235433 , n235434 , n235435 , n235436 , n235437 , n235438 , 
 n235439 , n235440 , n235441 , n235442 , n235443 , n235444 , n235445 , n235446 , n235447 , n235448 , 
 n235449 , n235450 , n235451 , n235452 , n235453 , n235454 , n235455 , n235456 , n235457 , n235458 , 
 n235459 , n235460 , n235461 , n235462 , n235463 , n235464 , n235465 , n235466 , n235467 , n235468 , 
 n235469 , n235470 , n235471 , n235472 , n235473 , n235474 , n235475 , n235476 , n235477 , n235478 , 
 n235479 , n235480 , n235481 , n235482 , n235483 , n235484 , n235485 , n235486 , n235487 , n235488 , 
 n235489 , n235490 , n235491 , n235492 , n235493 , n235494 , n235495 , n235496 , n235497 , n235498 , 
 n235499 , n235500 , n235501 , n235502 , n235503 , n235504 , n235505 , n235506 , n235507 , n235508 , 
 n235509 , n235510 , n235511 , n235512 , n235513 , n235514 , n235515 , n235516 , n235517 , n235518 , 
 n235519 , n235520 , n235521 , n235522 , n235523 , n235524 , n235525 , n235526 , n235527 , n235528 , 
 n235529 , n235530 , n235531 , n235532 , n235533 , n235534 , n235535 , n235536 , n235537 , n235538 , 
 n235539 , n235540 , n235541 , n235542 , n235543 , n235544 , n235545 , n235546 , n235547 , n235548 , 
 n235549 , n235550 , n235551 , n235552 , n235553 , n235554 , n235555 , n235556 , n235557 , n235558 , 
 n235559 , n235560 , n235561 , n235562 , n235563 , n235564 , n235565 , n235566 , n235567 , n235568 , 
 n235569 , n235570 , n235571 , n235572 , n235573 , n235574 , n235575 , n235576 , n235577 , n235578 , 
 n235579 , n235580 , n235581 , n235582 , n235583 , n235584 , n235585 , n235586 , n235587 , n235588 , 
 n235589 , n235590 , n235591 , n235592 , n235593 , n235594 , n235595 , n235596 , n235597 , n235598 , 
 n235599 , n235600 , n235601 , n235602 , n235603 , n235604 , n235605 , n235606 , n235607 , n235608 , 
 n235609 , n235610 , n235611 , n235612 , n235613 , n235614 , n235615 , n235616 , n235617 , n235618 , 
 n235619 , n235620 , n235621 , n235622 , n235623 , n235624 , n235625 , n235626 , n235627 , n235628 , 
 n235629 , n235630 , n235631 , n235632 , n235633 , n235634 , n235635 , n235636 , n235637 , n235638 , 
 n235639 , n235640 , n235641 , n235642 , n235643 , n235644 , n235645 , n235646 , n235647 , n235648 , 
 n235649 , n235650 , n235651 , n235652 , n235653 , n235654 , n235655 , n235656 , n235657 , n235658 , 
 n235659 , n235660 , n235661 , n235662 , n235663 , n235664 , n235665 , n235666 , n235667 , n235668 , 
 n235669 , n235670 , n235671 , n235672 , n235673 , n235674 , n235675 , n235676 , n235677 , n235678 , 
 n235679 , n235680 , n235681 , n235682 , n235683 , n235684 , n235685 , n235686 , n235687 , n235688 , 
 n235689 , n235690 , n235691 , n235692 , n235693 , n235694 , n235695 , n235696 , n235697 , n235698 , 
 n235699 , n235700 , n235701 , n235702 , n235703 , n235704 , n235705 , n235706 , n235707 , n235708 , 
 n235709 , n235710 , n235711 , n235712 , n235713 , n235714 , n235715 , n235716 , n235717 , n235718 , 
 n235719 , n235720 , n235721 , n235722 , n235723 , n235724 , n235725 , n235726 , n235727 , n235728 , 
 n235729 , n235730 , n235731 , n235732 , n235733 , n235734 , n235735 , n235736 , n235737 , n235738 , 
 n235739 , n235740 , n235741 , n235742 , n235743 , n235744 , n235745 , n235746 , n235747 , n235748 , 
 n235749 , n235750 , n235751 , n235752 , n235753 , n235754 , n235755 , n235756 , n235757 , n235758 , 
 n235759 , n235760 , n235761 , n235762 , n235763 , n235764 , n235765 , n235766 , n235767 , n235768 , 
 n235769 , n235770 , n235771 , n235772 , n235773 , n235774 , n235775 , n235776 , n235777 , n235778 , 
 n235779 , n235780 , n235781 , n235782 , n235783 , n235784 , n235785 , n235786 , n235787 , n235788 , 
 n235789 , n235790 , n235791 , n235792 , n235793 , n235794 , n235795 , n235796 , n235797 , n235798 , 
 n235799 , n235800 , n235801 , n235802 , n235803 , n235804 , n235805 , n235806 , n235807 , n235808 , 
 n235809 , n235810 , n235811 , n235812 , n235813 , n235814 , n235815 , n235816 , n235817 , n235818 , 
 n235819 , n235820 , n235821 , n235822 , n235823 , n235824 , n235825 , n235826 , n235827 , n235828 , 
 n235829 , n235830 , n235831 , n235832 , n235833 , n235834 , n235835 , n235836 , n235837 , n235838 , 
 n235839 , n235840 , n235841 , n235842 , n235843 , n235844 , n235845 , n235846 , n235847 , n235848 , 
 n235849 , n235850 , n235851 , n235852 , n235853 , n235854 , n235855 , n235856 , n235857 , n235858 , 
 n235859 , n235860 , n235861 , n235862 , n235863 , n235864 , n235865 , n235866 , n235867 , n235868 , 
 n235869 , n235870 , n235871 , n235872 , n235873 , n235874 , n235875 , n235876 , n235877 , n235878 , 
 n235879 , n235880 , n235881 , n235882 , n235883 , n235884 , n235885 , n235886 , n235887 , n235888 , 
 n235889 , n235890 , n235891 , n235892 , n235893 , n235894 , n235895 , n235896 , n235897 , n235898 , 
 n235899 , n235900 , n235901 , n235902 , n235903 , n235904 , n235905 , n235906 , n235907 , n235908 , 
 n235909 , n235910 , n235911 , n235912 , n235913 , n235914 , n235915 , n235916 , n235917 , n235918 , 
 n235919 , n235920 , n235921 , n235922 , n235923 , n235924 , n235925 , n235926 , n235927 , n235928 , 
 n235929 , n235930 , n235931 , n235932 , n235933 , n235934 , n235935 , n235936 , n235937 , n235938 , 
 n235939 , n235940 , n235941 , n235942 , n235943 , n235944 , n235945 , n235946 , n235947 , n235948 , 
 n235949 , n235950 , n235951 , n235952 , n235953 , n235954 , n235955 , n235956 , n235957 , n235958 , 
 n235959 , n235960 , n235961 , n235962 , n235963 , n235964 , n235965 , n235966 , n235967 , n235968 , 
 n235969 , n235970 , n235971 , n235972 , n235973 , n235974 , n235975 , n235976 , n235977 , n235978 , 
 n235979 , n235980 , n235981 , n235982 , n235983 , n235984 , n235985 , n235986 , n235987 , n235988 , 
 n235989 , n235990 , n235991 , n235992 , n235993 , n235994 , n235995 , n235996 , n235997 , n235998 , 
 n235999 , n236000 , n236001 , n236002 , n236003 , n236004 , n236005 , n236006 , n236007 , n236008 , 
 n236009 , n236010 , n236011 , n236012 , n236013 , n236014 , n236015 , n236016 , n236017 , n236018 , 
 n236019 , n236020 , n236021 , n236022 , n236023 , n236024 , n236025 , n236026 , n236027 , n236028 , 
 n236029 , n236030 , n236031 , n236032 , n236033 , n236034 , n236035 , n236036 , n236037 , n236038 , 
 n236039 , n236040 , n236041 , n236042 , n236043 , n236044 , n236045 , n236046 , n236047 , n236048 , 
 n236049 , n236050 , n236051 , n236052 , n236053 , n236054 , n236055 , n236056 , n236057 , n236058 , 
 n236059 , n236060 , n236061 , n236062 , n236063 , n236064 , n236065 , n236066 , n236067 , n236068 , 
 n236069 , n236070 , n236071 , n236072 , n236073 , n236074 , n236075 , n236076 , n236077 , n236078 , 
 n236079 , n236080 , n236081 , n236082 , n236083 , n236084 , n236085 , n236086 , n236087 , n236088 , 
 n236089 , n236090 , n236091 , n236092 , n236093 , n236094 , n236095 , n236096 , n236097 , n236098 , 
 n236099 , n236100 , n236101 , n236102 , n236103 , n236104 , n236105 , n236106 , n236107 , n236108 , 
 n236109 , n236110 , n236111 , n236112 , n236113 , n236114 , n236115 , n236116 , n236117 , n236118 , 
 n236119 , n236120 , n236121 , n236122 , n236123 , n236124 , n236125 , n236126 , n236127 , n236128 , 
 n236129 , n236130 , n236131 , n236132 , n236133 , n236134 , n236135 , n236136 , n236137 , n236138 , 
 n236139 , n236140 , n236141 , n236142 , n236143 , n236144 , n236145 , n236146 , n236147 , n236148 , 
 n236149 , n236150 , n236151 , n236152 , n236153 , n236154 , n236155 , n236156 , n236157 , n236158 , 
 n236159 , n236160 , n236161 , n236162 , n236163 , n236164 , n236165 , n236166 , n236167 , n236168 , 
 n236169 , n236170 , n236171 , n236172 , n236173 , n236174 , n236175 , n236176 , n236177 , n236178 , 
 n236179 , n236180 , n236181 , n236182 , n236183 , n236184 , n236185 , n236186 , n236187 , n236188 , 
 n236189 , n236190 , n236191 , n236192 , n236193 , n236194 , n236195 , n236196 , n236197 , n236198 , 
 n236199 , n236200 , n236201 , n236202 , n236203 , n236204 , n236205 , n236206 , n236207 , n236208 , 
 n236209 , n236210 , n236211 , n236212 , n236213 , n236214 , n236215 , n236216 , n236217 , n236218 , 
 n236219 , n236220 , n236221 , n236222 , n236223 , n236224 , n236225 , n236226 , n236227 , n236228 , 
 n236229 , n236230 , n236231 , n236232 , n236233 , n236234 , n236235 , n236236 , n236237 , n236238 , 
 n236239 , n236240 , n236241 , n236242 , n236243 , n236244 , n236245 , n236246 , n236247 , n236248 , 
 n236249 , n236250 , n236251 , n236252 , n236253 , n236254 , n236255 , n236256 , n236257 , n236258 , 
 n236259 , n236260 , n236261 , n236262 , n236263 , n236264 , n236265 , n236266 , n236267 , n236268 , 
 n236269 , n236270 , n236271 , n236272 , n236273 , n236274 , n236275 , n236276 , n236277 , n236278 , 
 n236279 , n236280 , n236281 , n236282 , n236283 , n236284 , n236285 , n236286 , n236287 , n236288 , 
 n236289 , n236290 , n236291 , n236292 , n236293 , n236294 , n236295 , n236296 , n236297 , n236298 , 
 n236299 , n236300 , n236301 , n236302 , n236303 , n236304 , n236305 , n236306 , n236307 , n236308 , 
 n236309 , n236310 , n236311 , n236312 , n236313 , n236314 , n236315 , n236316 , n236317 , n236318 , 
 n236319 , n236320 , n236321 , n236322 , n236323 , n236324 , n236325 , n236326 , n236327 , n236328 , 
 n236329 , n236330 , n236331 , n236332 , n236333 , n236334 , n236335 , n236336 , n236337 , n236338 , 
 n236339 , n236340 , n236341 , n236342 , n236343 , n236344 , n236345 , n236346 , n236347 , n236348 , 
 n236349 , n236350 , n236351 , n236352 , n236353 , n236354 , n236355 , n236356 , n236357 , n236358 , 
 n236359 , n236360 , n236361 , n236362 , n236363 , n236364 , n236365 , n236366 , n236367 , n236368 , 
 n236369 , n236370 , n236371 , n236372 , n236373 , n236374 , n236375 , n236376 , n236377 , n236378 , 
 n236379 , n236380 , n236381 , n236382 , n236383 , n236384 , n236385 , n236386 , n236387 , n236388 , 
 n236389 , n236390 , n236391 , n236392 , n236393 , n236394 , n236395 , n236396 , n236397 , n236398 , 
 n236399 , n236400 , n236401 , n236402 , n236403 , n236404 , n236405 , n236406 , n236407 , n236408 , 
 n236409 , n236410 , n236411 , n236412 , n236413 , n236414 , n236415 , n236416 , n236417 , n236418 , 
 n236419 , n236420 , n236421 , n236422 , n236423 , n236424 , n236425 , n236426 , n236427 , n236428 , 
 n236429 , n236430 , n236431 , n236432 , n236433 , n236434 , n236435 , n236436 , n236437 , n236438 , 
 n236439 , n236440 , n236441 , n236442 , n236443 , n236444 , n236445 , n236446 , n236447 , n236448 , 
 n236449 , n236450 , n236451 , n236452 , n236453 , n236454 , n236455 , n236456 , n236457 , n236458 , 
 n236459 , n236460 , n236461 , n236462 , n236463 , n236464 , n236465 , n236466 , n236467 , n236468 , 
 n236469 , n236470 , n236471 , n236472 , n236473 , n236474 , n236475 , n236476 , n236477 , n236478 , 
 n236479 , n236480 , n236481 , n236482 , n236483 , n236484 , n236485 , n236486 , n236487 , n236488 , 
 n236489 , n236490 , n236491 , n236492 , n236493 , n236494 , n236495 , n236496 , n236497 , n236498 , 
 n236499 , n236500 , n236501 , n236502 , n236503 , n236504 , n236505 , n236506 , n236507 , n236508 , 
 n236509 , n236510 , n236511 , n236512 , n236513 , n236514 , n236515 , n236516 , n236517 , n236518 , 
 n236519 , n236520 , n236521 , n236522 , n236523 , n236524 , n236525 , n236526 , n236527 , n236528 , 
 n236529 , n236530 , n236531 , n236532 , n236533 , n236534 , n236535 , n236536 , n236537 , n236538 , 
 n236539 , n236540 , n236541 , n236542 , n236543 , n236544 , n236545 , n236546 , n236547 , n236548 , 
 n236549 , n236550 , n236551 , n236552 , n236553 , n236554 , n236555 , n236556 , n236557 , n236558 , 
 n236559 , n236560 , n236561 , n236562 , n236563 , n236564 , n236565 , n236566 , n236567 , n236568 , 
 n236569 , n236570 , n236571 , n236572 , n236573 , n236574 , n236575 , n236576 , n236577 , n236578 , 
 n236579 , n236580 , n236581 , n236582 , n236583 , n236584 , n236585 , n236586 , n236587 , n236588 , 
 n236589 , n236590 , n236591 , n236592 , n236593 , n236594 , n236595 , n236596 , n236597 , n236598 , 
 n236599 , n236600 , n236601 , n236602 , n236603 , n236604 , n236605 , n236606 , n236607 , n236608 , 
 n236609 , n236610 , n236611 , n236612 , n236613 , n236614 , n236615 , n236616 , n236617 , n236618 , 
 n236619 , n236620 , n236621 , n236622 , n236623 , n236624 , n236625 , n236626 , n236627 , n236628 , 
 n236629 , n236630 , n236631 , n236632 , n236633 , n236634 , n236635 , n236636 , n236637 , n236638 , 
 n236639 , n236640 , n236641 , n236642 , n236643 , n236644 , n236645 , n236646 , n236647 , n236648 , 
 n236649 , n236650 , n236651 , n236652 , n236653 , n236654 , n236655 , n236656 , n236657 , n236658 , 
 n236659 , n236660 , n236661 , n236662 , n236663 , n236664 , n236665 , n236666 , n236667 , n236668 , 
 n236669 , n236670 , n236671 , n236672 , n236673 , n236674 , n236675 , n236676 , n236677 , n236678 , 
 n236679 , n236680 , n236681 , n236682 , n236683 , n236684 , n236685 , n236686 , n236687 , n236688 , 
 n236689 , n236690 , n236691 , n236692 , n236693 , n236694 , n236695 , n236696 , n236697 , n236698 , 
 n236699 , n236700 , n236701 , n236702 , n236703 , n236704 , n236705 , n236706 , n236707 , n236708 , 
 n236709 , n236710 , n236711 , n236712 , n236713 , n236714 , n236715 , n236716 , n236717 , n236718 , 
 n236719 , n236720 , n236721 , n236722 , n236723 , n236724 , n236725 , n236726 , n236727 , n236728 , 
 n236729 , n236730 , n236731 , n236732 , n236733 , n236734 , n236735 , n236736 , n236737 , n236738 , 
 n236739 , n236740 , n236741 , n236742 , n236743 , n236744 , n236745 , n236746 , n236747 , n236748 , 
 n236749 , n236750 , n236751 , n236752 , n236753 , n236754 , n236755 , n236756 , n236757 , n236758 , 
 n236759 , n236760 , n236761 , n236762 , n236763 , n236764 , n236765 , n236766 , n236767 , n236768 , 
 n236769 , n236770 , n236771 , n236772 , n236773 , n236774 , n236775 , n236776 , n236777 , n236778 , 
 n236779 , n236780 , n236781 , n236782 , n236783 , n236784 , n236785 , n236786 , n236787 , n236788 , 
 n236789 , n236790 , n236791 , n236792 , n236793 , n236794 , n236795 , n236796 , n236797 , n236798 , 
 n236799 , n236800 , n236801 , n236802 , n236803 , n236804 , n236805 , n236806 , n236807 , n236808 , 
 n236809 , n236810 , n236811 , n236812 , n236813 , n236814 , n236815 , n236816 , n236817 , n236818 , 
 n236819 , n236820 , n236821 , n236822 , n236823 , n236824 , n236825 , n236826 , n236827 , n236828 , 
 n236829 , n236830 , n236831 , n236832 , n236833 , n236834 , n236835 , n236836 , n236837 , n236838 , 
 n236839 , n236840 , n236841 , n236842 , n236843 , n236844 , n236845 , n236846 , n236847 , n236848 , 
 n236849 , n236850 , n236851 , n236852 , n236853 , n236854 , n236855 , n236856 , n236857 , n236858 , 
 n236859 , n236860 , n236861 , n236862 , n236863 , n236864 , n236865 , n236866 , n236867 , n236868 , 
 n236869 , n236870 , n236871 , n236872 , n236873 , n236874 , n236875 , n236876 , n236877 , n236878 , 
 n236879 , n236880 , n236881 , n236882 , n236883 , n236884 , n236885 , n236886 , n236887 , n236888 , 
 n236889 , n236890 , n236891 , n236892 , n236893 , n236894 , n236895 , n236896 , n236897 , n236898 , 
 n236899 , n236900 , n236901 , n236902 , n236903 , n236904 , n236905 , n236906 , n236907 , n236908 , 
 n236909 , n236910 , n236911 , n236912 , n236913 , n236914 , n236915 , n236916 , n236917 , n236918 , 
 n236919 , n236920 , n236921 , n236922 , n236923 , n236924 , n236925 , n236926 , n236927 , n236928 , 
 n236929 , n236930 , n236931 , n236932 , n236933 , n236934 , n236935 , n236936 , n236937 , n236938 , 
 n236939 , n236940 , n236941 , n236942 , n236943 , n236944 , n236945 , n236946 , n236947 , n236948 , 
 n236949 , n236950 , n236951 , n236952 , n236953 , n236954 , n236955 , n236956 , n236957 , n236958 , 
 n236959 , n236960 , n236961 , n236962 , n236963 , n236964 , n236965 , n236966 , n236967 , n236968 , 
 n236969 , n236970 , n236971 , n236972 , n236973 , n236974 , n236975 , n236976 , n236977 , n236978 , 
 n236979 , n236980 , n236981 , n236982 , n236983 , n236984 , n236985 , n236986 , n236987 , n236988 , 
 n236989 , n236990 , n236991 , n236992 , n236993 , n236994 , n236995 , n236996 , n236997 , n236998 , 
 n236999 , n237000 , n237001 , n237002 , n237003 , n237004 , n237005 , n237006 , n237007 , n237008 , 
 n237009 , n237010 , n237011 , n237012 , n237013 , n237014 , n237015 , n237016 , n237017 , n237018 , 
 n237019 , n237020 , n237021 , n237022 , n237023 , n237024 , n237025 , n237026 , n237027 , n237028 , 
 n237029 , n237030 , n237031 , n237032 , n237033 , n237034 , n237035 , n237036 , n237037 , n237038 , 
 n237039 , n237040 , n237041 , n237042 , n237043 , n237044 , n237045 , n237046 , n237047 , n237048 , 
 n237049 , n237050 , n237051 , n237052 , n237053 , n237054 , n237055 , n237056 , n237057 , n237058 , 
 n237059 , n237060 , n237061 , n237062 , n237063 , n237064 , n237065 , n237066 , n237067 , n237068 , 
 n237069 , n237070 , n237071 , n237072 , n237073 , n237074 , n237075 , n237076 , n237077 , n237078 , 
 n237079 , n237080 , n237081 , n237082 , n237083 , n237084 , n237085 , n237086 , n237087 , n237088 , 
 n237089 , n237090 , n237091 , n237092 , n237093 , n237094 , n237095 , n237096 , n237097 , n237098 , 
 n237099 , n237100 , n237101 , n237102 , n237103 , n237104 , n237105 , n237106 , n237107 , n237108 , 
 n237109 , n237110 , n237111 , n237112 , n237113 , n237114 , n237115 , n237116 , n237117 , n237118 , 
 n237119 , n237120 , n237121 , n237122 , n237123 , n237124 , n237125 , n237126 , n237127 , n237128 , 
 n237129 , n237130 , n237131 , n237132 , n237133 , n237134 , n237135 , n237136 , n237137 , n237138 , 
 n237139 , n237140 , n237141 , n237142 , n237143 , n237144 , n237145 , n237146 , n237147 , n237148 , 
 n237149 , n237150 , n237151 , n237152 , n237153 , n237154 , n237155 , n237156 , n237157 , n237158 , 
 n237159 , n237160 , n237161 , n237162 , n237163 , n237164 , n237165 , n237166 , n237167 , n237168 , 
 n237169 , n237170 , n237171 , n237172 , n237173 , n237174 , n237175 , n237176 , n237177 , n237178 , 
 n237179 , n237180 , n237181 , n237182 , n237183 , n237184 , n237185 , n237186 , n237187 , n237188 , 
 n237189 , n237190 , n237191 , n237192 , n237193 , n237194 , n237195 , n237196 , n237197 , n237198 , 
 n237199 , n237200 , n237201 , n237202 , n237203 , n237204 , n237205 , n237206 , n237207 , n237208 , 
 n237209 , n237210 , n237211 , n237212 , n237213 , n237214 , n237215 , n237216 , n237217 , n237218 , 
 n237219 , n237220 , n237221 , n237222 , n237223 , n237224 , n237225 , n237226 , n237227 , n237228 , 
 n237229 , n237230 , n237231 , n237232 , n237233 , n237234 , n237235 , n237236 , n237237 , n237238 , 
 n237239 , n237240 , n237241 , n237242 , n237243 , n237244 , n237245 , n237246 , n237247 , n237248 , 
 n237249 , n237250 , n237251 , n237252 , n237253 , n237254 , n237255 , n237256 , n237257 , n237258 , 
 n237259 , n237260 , n237261 , n237262 , n237263 , n237264 , n237265 , n237266 , n237267 , n237268 , 
 n237269 , n237270 , n237271 , n237272 , n237273 , n237274 , n237275 , n237276 , n237277 , n237278 , 
 n237279 , n237280 , n237281 , n237282 , n237283 , n237284 , n237285 , n237286 , n237287 , n237288 , 
 n237289 , n237290 , n237291 , n237292 , n237293 , n237294 , n237295 , n237296 , n237297 , n237298 , 
 n237299 , n237300 , n237301 , n237302 , n237303 , n237304 , n237305 , n237306 , n237307 , n237308 , 
 n237309 , n237310 , n237311 , n237312 , n237313 , n237314 , n237315 , n237316 , n237317 , n237318 , 
 n237319 , n237320 , n237321 , n237322 , n237323 , n237324 , n237325 , n237326 , n237327 , n237328 , 
 n237329 , n237330 , n237331 , n237332 , n237333 , n237334 , n237335 , n237336 , n237337 , n237338 , 
 n237339 , n237340 , n237341 , n237342 , n237343 , n237344 , n237345 , n237346 , n237347 , n237348 , 
 n237349 , n237350 , n237351 , n237352 , n237353 , n237354 , n237355 , n237356 , n237357 , n237358 , 
 n237359 , n237360 , n237361 , n237362 , n237363 , n237364 , n237365 , n237366 , n237367 , n237368 , 
 n237369 , n237370 , n237371 , n237372 , n237373 , n237374 , n237375 , n237376 , n237377 , n237378 , 
 n237379 , n237380 , n237381 , n237382 , n237383 , n237384 , n237385 , n237386 , n237387 , n237388 , 
 n237389 , n237390 , n237391 , n237392 , n237393 , n237394 , n237395 , n237396 , n237397 , n237398 , 
 n237399 , n237400 , n237401 , n237402 , n237403 , n237404 , n237405 , n237406 , n237407 , n237408 , 
 n237409 , n237410 , n237411 , n237412 , n237413 , n237414 , n237415 , n237416 , n237417 , n237418 , 
 n237419 , n237420 , n237421 , n237422 , n237423 , n237424 , n237425 , n237426 , n237427 , n237428 , 
 n237429 , n237430 , n237431 , n237432 , n237433 , n237434 , n237435 , n237436 , n237437 , n237438 , 
 n237439 , n237440 , n237441 , n237442 , n237443 , n237444 , n237445 , n237446 , n237447 , n237448 , 
 n237449 , n237450 , n237451 , n237452 , n237453 , n237454 , n237455 , n237456 , n237457 , n237458 , 
 n237459 , n237460 , n237461 , n237462 , n237463 , n237464 , n237465 , n237466 , n237467 , n237468 , 
 n237469 , n237470 , n237471 , n237472 , n237473 , n237474 , n237475 , n237476 , n237477 , n237478 , 
 n237479 , n237480 , n237481 , n237482 , n237483 , n237484 , n237485 , n237486 , n237487 , n237488 , 
 n237489 , n237490 , n237491 , n237492 , n237493 , n237494 , n237495 , n237496 , n237497 , n237498 , 
 n237499 , n237500 , n237501 , n237502 , n237503 , n237504 , n237505 , n237506 , n237507 , n237508 , 
 n237509 , n237510 , n237511 , n237512 , n237513 , n237514 , n237515 , n237516 , n237517 , n237518 , 
 n237519 , n237520 , n237521 , n237522 , n237523 , n237524 , n237525 , n237526 , n237527 , n237528 , 
 n237529 , n237530 , n237531 , n237532 , n237533 , n237534 , n237535 , n237536 , n237537 , n237538 , 
 n237539 , n237540 , n237541 , n237542 , n237543 , n237544 , n237545 , n237546 , n237547 , n237548 , 
 n237549 , n237550 , n237551 , n237552 , n237553 , n237554 , n237555 , n237556 , n237557 , n237558 , 
 n237559 , n237560 , n237561 , n237562 , n237563 , n237564 , n237565 , n237566 , n237567 , n237568 , 
 n237569 , n237570 , n237571 , n237572 , n237573 , n237574 , n237575 , n237576 , n237577 , n237578 , 
 n237579 , n237580 , n237581 , n237582 , n237583 , n237584 , n237585 , n237586 , n237587 , n237588 , 
 n237589 , n237590 , n237591 , n237592 , n237593 , n237594 , n237595 , n237596 , n237597 , n237598 , 
 n237599 , n237600 , n237601 , n237602 , n237603 , n237604 , n237605 , n237606 , n237607 , n237608 , 
 n237609 , n237610 , n237611 , n237612 , n237613 , n237614 , n237615 , n237616 , n237617 , n237618 , 
 n237619 , n237620 , n237621 , n237622 , n237623 , n237624 , n237625 , n237626 , n237627 , n237628 , 
 n237629 , n237630 , n237631 , n237632 , n237633 , n237634 , n237635 , n237636 , n237637 , n237638 , 
 n237639 , n237640 , n237641 , n237642 , n237643 , n237644 , n237645 , n237646 , n237647 , n237648 , 
 n237649 , n237650 , n237651 , n237652 , n237653 , n237654 , n237655 , n237656 , n237657 , n237658 , 
 n237659 , n237660 , n237661 , n237662 , n237663 , n237664 , n237665 , n237666 , n237667 , n237668 , 
 n237669 , n237670 , n237671 , n237672 , n237673 , n237674 , n237675 , n237676 , n237677 , n237678 , 
 n237679 , n237680 , n237681 , n237682 , n237683 , n237684 , n237685 , n237686 , n237687 , n237688 , 
 n237689 , n237690 , n237691 , n237692 , n237693 , n237694 , n237695 , n237696 , n237697 , n237698 , 
 n237699 , n237700 , n237701 , n237702 , n237703 , n237704 , n237705 , n237706 , n237707 , n237708 , 
 n237709 , n237710 , n237711 , n237712 , n237713 , n237714 , n237715 , n237716 , n237717 , n237718 , 
 n237719 , n237720 , n237721 , n237722 , n237723 , n237724 , n237725 , n237726 , n237727 , n237728 , 
 n237729 , n237730 , n237731 , n237732 , n237733 , n237734 , n237735 , n237736 , n237737 , n237738 , 
 n237739 , n237740 , n237741 , n237742 , n237743 , n237744 , n237745 , n237746 , n237747 , n237748 , 
 n237749 , n237750 , n237751 , n237752 , n237753 , n237754 , n237755 , n237756 , n237757 , n237758 , 
 n237759 , n237760 , n237761 , n237762 , n237763 , n237764 , n237765 , n237766 , n237767 , n237768 , 
 n237769 , n237770 , n237771 , n237772 , n237773 , n237774 , n237775 , n237776 , n237777 , n237778 , 
 n237779 , n237780 , n237781 , n237782 , n237783 , n237784 , n237785 , n237786 , n237787 , n237788 , 
 n237789 , n237790 , n237791 , n237792 , n237793 , n237794 , n237795 , n237796 , n237797 , n237798 , 
 n237799 , n237800 , n237801 , n237802 , n237803 , n237804 , n237805 , n237806 , n237807 , n237808 , 
 n237809 , n237810 , n237811 , n237812 , n237813 , n237814 , n237815 , n237816 , n237817 , n237818 , 
 n237819 , n237820 , n237821 , n237822 , n237823 , n237824 , n237825 , n237826 , n237827 , n237828 , 
 n237829 , n237830 , n237831 , n237832 , n237833 , n237834 , n237835 , n237836 , n237837 , n237838 , 
 n237839 , n237840 , n237841 , n237842 , n237843 , n237844 , n237845 , n237846 , n237847 , n237848 , 
 n237849 , n237850 , n237851 , n237852 , n237853 , n237854 , n237855 , n237856 , n237857 , n237858 , 
 n237859 , n237860 , n237861 , n237862 , n237863 , n237864 , n237865 , n237866 , n237867 , n237868 , 
 n237869 , n237870 , n237871 , n237872 , n237873 , n237874 , n237875 , n237876 , n237877 , n237878 , 
 n237879 , n237880 , n237881 , n237882 , n237883 , n237884 , n237885 , n237886 , n237887 , n237888 , 
 n237889 , n237890 , n237891 , n237892 , n237893 , n237894 , n237895 , n237896 , n237897 , n237898 , 
 n237899 , n237900 , n237901 , n237902 , n237903 , n237904 , n237905 , n237906 , n237907 , n237908 , 
 n237909 , n237910 , n237911 , n237912 , n237913 , n237914 , n237915 , n237916 , n237917 , n237918 , 
 n237919 , n237920 , n237921 , n237922 , n237923 , n237924 , n237925 , n237926 , n237927 , n237928 , 
 n237929 , n237930 , n237931 , n237932 , n237933 , n237934 , n237935 , n237936 , n237937 , n237938 , 
 n237939 , n237940 , n237941 , n237942 , n237943 , n237944 , n237945 , n237946 , n237947 , n237948 , 
 n237949 , n237950 , n237951 , n237952 , n237953 , n237954 , n237955 , n237956 , n237957 , n237958 , 
 n237959 , n237960 , n237961 , n237962 , n237963 , n237964 , n237965 , n237966 , n237967 , n237968 , 
 n237969 , n237970 , n237971 , n237972 , n237973 , n237974 , n237975 , n237976 , n237977 , n237978 , 
 n237979 , n237980 , n237981 , n237982 , n237983 , n237984 , n237985 , n237986 , n237987 , n237988 , 
 n237989 , n237990 , n237991 , n237992 , n237993 , n237994 , n237995 , n237996 , n237997 , n237998 , 
 n237999 , n238000 , n238001 , n238002 , n238003 , n238004 , n238005 , n238006 , n238007 , n238008 , 
 n238009 , n238010 , n238011 , n238012 , n238013 , n238014 , n238015 , n238016 , n238017 , n238018 , 
 n238019 , n238020 , n238021 , n238022 , n238023 , n238024 , n238025 , n238026 , n238027 , n238028 , 
 n238029 , n238030 , n238031 , n238032 , n238033 , n238034 , n238035 , n238036 , n238037 , n238038 , 
 n238039 , n238040 , n238041 , n238042 , n238043 , n238044 , n238045 , n238046 , n238047 , n238048 , 
 n238049 , n238050 , n238051 , n238052 , n238053 , n238054 , n238055 , n238056 , n238057 , n238058 , 
 n238059 , n238060 , n238061 , n238062 , n238063 , n238064 , n238065 , n238066 , n238067 , n238068 , 
 n238069 , n238070 , n238071 , n238072 , n238073 , n238074 , n238075 , n238076 , n238077 , n238078 , 
 n238079 , n238080 , n238081 , n238082 , n238083 , n238084 , n238085 , n238086 , n238087 , n238088 , 
 n238089 , n238090 , n238091 , n238092 , n238093 , n238094 , n238095 , n238096 , n238097 , n238098 , 
 n238099 , n238100 , n238101 , n238102 , n238103 , n238104 , n238105 , n238106 , n238107 , n238108 , 
 n238109 , n238110 , n238111 , n238112 , n238113 , n238114 , n238115 , n238116 , n238117 , n238118 , 
 n238119 , n238120 , n238121 , n238122 , n238123 , n238124 , n238125 , n238126 , n238127 , n238128 , 
 n238129 , n238130 , n238131 , n238132 , n238133 , n238134 , n238135 , n238136 , n238137 , n238138 , 
 n238139 , n238140 , n238141 , n238142 , n238143 , n238144 , n238145 , n238146 , n238147 , n238148 , 
 n238149 , n238150 , n238151 , n238152 , n238153 , n238154 , n238155 , n238156 , n238157 , n238158 , 
 n238159 , n238160 , n238161 , n238162 , n238163 , n238164 , n238165 , n238166 , n238167 , n238168 , 
 n238169 , n238170 , n238171 , n238172 , n238173 , n238174 , n238175 , n238176 , n238177 , n238178 , 
 n238179 , n238180 , n238181 , n238182 , n238183 , n238184 , n238185 , n238186 , n238187 , n238188 , 
 n238189 , n238190 , n238191 , n238192 , n238193 , n238194 , n238195 , n238196 , n238197 , n238198 , 
 n238199 , n238200 , n238201 , n238202 , n238203 , n238204 , n238205 , n238206 , n238207 , n238208 , 
 n238209 , n238210 , n238211 , n238212 , n238213 , n238214 , n238215 , n238216 , n238217 , n238218 , 
 n238219 , n238220 , n238221 , n238222 , n238223 , n238224 , n238225 , n238226 , n238227 , n238228 , 
 n238229 , n238230 , n238231 , n238232 , n238233 , n238234 , n238235 , n238236 , n238237 , n238238 , 
 n238239 , n238240 , n238241 , n238242 , n238243 , n238244 , n238245 , n238246 , n238247 , n238248 , 
 n238249 , n238250 , n238251 , n238252 , n238253 , n238254 , n238255 , n238256 , n238257 , n238258 , 
 n238259 , n238260 , n238261 , n238262 , n238263 , n238264 , n238265 , n238266 , n238267 , n238268 , 
 n238269 , n238270 , n238271 , n238272 , n238273 , n238274 , n238275 , n238276 , n238277 , n238278 , 
 n238279 , n238280 , n238281 , n238282 , n238283 , n238284 , n238285 , n238286 , n238287 , n238288 , 
 n238289 , n238290 , n238291 , n238292 , n238293 , n238294 , n238295 , n238296 , n238297 , n238298 , 
 n238299 , n238300 , n238301 , n238302 , n238303 , n238304 , n238305 , n238306 , n238307 , n238308 , 
 n238309 , n238310 , n238311 , n238312 , n238313 , n238314 , n238315 , n238316 , n238317 , n238318 , 
 n238319 , n238320 , n238321 , n238322 , n238323 , n238324 , n238325 , n238326 , n238327 , n238328 , 
 n238329 , n238330 , n238331 , n238332 , n238333 , n238334 , n238335 , n238336 , n238337 , n238338 , 
 n238339 , n238340 , n238341 , n238342 , n238343 , n238344 , n238345 , n238346 , n238347 , n238348 , 
 n238349 , n238350 , n238351 , n238352 , n238353 , n238354 , n238355 , n238356 , n238357 , n238358 , 
 n238359 , n238360 , n238361 , n238362 , n238363 , n238364 , n238365 , n238366 , n238367 , n238368 , 
 n238369 , n238370 , n238371 , n238372 , n238373 , n238374 , n238375 , n238376 , n238377 , n238378 , 
 n238379 , n238380 , n238381 , n238382 , n238383 , n238384 , n238385 , n238386 , n238387 , n238388 , 
 n238389 , n238390 , n238391 , n238392 , n238393 , n238394 , n238395 , n238396 , n238397 , n238398 , 
 n238399 , n238400 , n238401 , n238402 , n238403 , n238404 , n238405 , n238406 , n238407 , n238408 , 
 n238409 , n238410 , n238411 , n238412 , n238413 , n238414 , n238415 , n238416 , n238417 , n238418 , 
 n238419 , n238420 , n238421 , n238422 , n238423 , n238424 , n238425 , n238426 , n238427 , n238428 , 
 n238429 , n238430 , n238431 , n238432 , n238433 , n238434 , n238435 , n238436 , n238437 , n238438 , 
 n238439 , n238440 , n238441 , n238442 , n238443 , n238444 , n238445 , n238446 , n238447 , n238448 , 
 n238449 , n238450 , n238451 , n238452 , n238453 , n238454 , n238455 , n238456 , n238457 , n238458 , 
 n238459 , n238460 , n238461 , n238462 , n238463 , n238464 , n238465 , n238466 , n238467 , n238468 , 
 n238469 , n238470 , n238471 , n238472 , n238473 , n238474 , n238475 , n238476 , n238477 , n238478 , 
 n238479 , n238480 , n238481 , n238482 , n238483 , n238484 , n238485 , n238486 , n238487 , n238488 , 
 n238489 , n238490 , n238491 , n238492 , n238493 , n238494 , n238495 , n238496 , n238497 , n238498 , 
 n238499 , n238500 , n238501 , n238502 , n238503 , n238504 , n238505 , n238506 , n238507 , n238508 , 
 n238509 , n238510 , n238511 , n238512 , n238513 , n238514 , n238515 , n238516 , n238517 , n238518 , 
 n238519 , n238520 , n238521 , n238522 , n238523 , n238524 , n238525 , n238526 , n238527 , n238528 , 
 n238529 , n238530 , n238531 , n238532 , n238533 , n238534 , n238535 , n238536 , n238537 , n238538 , 
 n238539 , n238540 , n238541 , n238542 , n238543 , n238544 , n238545 , n238546 , n238547 , n238548 , 
 n238549 , n238550 , n238551 , n238552 , n238553 , n238554 , n238555 , n238556 , n238557 , n238558 , 
 n238559 , n238560 , n238561 , n238562 , n238563 , n238564 , n238565 , n238566 , n238567 , n238568 , 
 n238569 , n238570 , n238571 , n238572 , n238573 , n238574 , n238575 , n238576 , n238577 , n238578 , 
 n238579 , n238580 , n238581 , n238582 , n238583 , n238584 , n238585 , n238586 , n238587 , n238588 , 
 n238589 , n238590 , n238591 , n238592 , n238593 , n238594 , n238595 , n238596 , n238597 , n238598 , 
 n238599 , n238600 , n238601 , n238602 , n238603 , n238604 , n238605 , n238606 , n238607 , n238608 , 
 n238609 , n238610 , n238611 , n238612 , n238613 , n238614 , n238615 , n238616 , n238617 , n238618 , 
 n238619 , n238620 , n238621 , n238622 , n238623 , n238624 , n238625 , n238626 , n238627 , n238628 , 
 n238629 , n238630 , n238631 , n238632 , n238633 , n238634 , n238635 , n238636 , n238637 , n238638 , 
 n238639 , n238640 , n238641 , n238642 , n238643 , n238644 , n238645 , n238646 , n238647 , n238648 , 
 n238649 , n238650 , n238651 , n238652 , n238653 , n238654 , n238655 , n238656 , n238657 , n238658 , 
 n238659 , n238660 , n238661 , n238662 , n238663 , n238664 , n238665 , n238666 , n238667 , n238668 , 
 n238669 , n238670 , n238671 , n238672 , n238673 , n238674 , n238675 , n238676 , n238677 , n238678 , 
 n238679 , n238680 , n238681 , n238682 , n238683 , n238684 , n238685 , n238686 , n238687 , n238688 , 
 n238689 , n238690 , n238691 , n238692 , n238693 , n238694 , n238695 , n238696 , n238697 , n238698 , 
 n238699 , n238700 , n238701 , n238702 , n238703 , n238704 , n238705 , n238706 , n238707 , n238708 , 
 n238709 , n238710 , n238711 , n238712 , n238713 , n238714 , n238715 , n238716 , n238717 , n238718 , 
 n238719 , n238720 , n238721 , n238722 , n238723 , n238724 , n238725 , n238726 , n238727 , n238728 , 
 n238729 , n238730 , n238731 , n238732 , n238733 , n238734 , n238735 , n238736 , n238737 , n238738 , 
 n238739 , n238740 , n238741 , n238742 , n238743 , n238744 , n238745 , n238746 , n238747 , n238748 , 
 n238749 , n238750 , n238751 , n238752 , n238753 , n238754 , n238755 , n238756 , n238757 , n238758 , 
 n238759 , n238760 , n238761 , n238762 , n238763 , n238764 , n238765 , n238766 , n238767 , n238768 , 
 n238769 , n238770 , n238771 , n238772 , n238773 , n238774 , n238775 , n238776 , n238777 , n238778 , 
 n238779 , n238780 , n238781 , n238782 , n238783 , n238784 , n238785 , n238786 , n238787 , n238788 , 
 n238789 , n238790 , n238791 , n238792 , n238793 , n238794 , n238795 , n238796 , n238797 , n238798 , 
 n238799 , n238800 , n238801 , n238802 , n238803 , n238804 , n238805 , n238806 , n238807 , n238808 , 
 n238809 , n238810 , n238811 , n238812 , n238813 , n238814 , n238815 , n238816 , n238817 , n238818 , 
 n238819 , n238820 , n238821 , n238822 , n238823 , n238824 , n238825 , n238826 , n238827 , n238828 , 
 n238829 , n238830 , n238831 , n238832 , n238833 , n238834 , n238835 , n238836 , n238837 , n238838 , 
 n238839 , n238840 , n238841 , n238842 , n238843 , n238844 , n238845 , n238846 , n238847 , n238848 , 
 n238849 , n238850 , n238851 , n238852 , n238853 , n238854 , n238855 , n238856 , n238857 , n238858 , 
 n238859 , n238860 , n238861 , n238862 , n238863 , n238864 , n238865 , n238866 , n238867 , n238868 , 
 n238869 , n238870 , n238871 , n238872 , n238873 , n238874 , n238875 , n238876 , n238877 , n238878 , 
 n238879 , n238880 , n238881 , n238882 , n238883 , n238884 , n238885 , n238886 , n238887 , n238888 , 
 n238889 , n238890 , n238891 , n238892 , n238893 , n238894 , n238895 , n238896 , n238897 , n238898 , 
 n238899 , n238900 , n238901 , n238902 , n238903 , n238904 , n238905 , n238906 , n238907 , n238908 , 
 n238909 , n238910 , n238911 , n238912 , n238913 , n238914 , n238915 , n238916 , n238917 , n238918 , 
 n238919 , n238920 , n238921 , n238922 , n238923 , n238924 , n238925 , n238926 , n238927 , n238928 , 
 n238929 , n238930 , n238931 , n238932 , n238933 , n238934 , n238935 , n238936 , n238937 , n238938 , 
 n238939 , n238940 , n238941 , n238942 , n238943 , n238944 , n238945 , n238946 , n238947 , n238948 , 
 n238949 , n238950 , n238951 , n238952 , n238953 , n238954 , n238955 , n238956 , n238957 , n238958 , 
 n238959 , n238960 , n238961 , n238962 , n238963 , n238964 , n238965 , n238966 , n238967 , n238968 , 
 n238969 , n238970 , n238971 , n238972 , n238973 , n238974 , n238975 , n238976 , n238977 , n238978 , 
 n238979 , n238980 , n238981 , n238982 , n238983 , n238984 , n238985 , n238986 , n238987 , n238988 , 
 n238989 , n238990 , n238991 , n238992 , n238993 , n238994 , n238995 , n238996 , n238997 , n238998 , 
 n238999 , n239000 , n239001 , n239002 , n239003 , n239004 , n239005 , n239006 , n239007 , n239008 , 
 n239009 , n239010 , n239011 , n239012 , n239013 , n239014 , n239015 , n239016 , n239017 , n239018 , 
 n239019 , n239020 , n239021 , n239022 , n239023 , n239024 , n239025 , n239026 , n239027 , n239028 , 
 n239029 , n239030 , n239031 , n239032 , n239033 , n239034 , n239035 , n239036 , n239037 , n239038 , 
 n239039 , n239040 , n239041 , n239042 , n239043 , n239044 , n239045 , n239046 , n239047 , n239048 , 
 n239049 , n239050 , n239051 , n239052 , n239053 , n239054 , n239055 , n239056 , n239057 , n239058 , 
 n239059 , n239060 , n239061 , n239062 , n239063 , n239064 , n239065 , n239066 , n239067 , n239068 , 
 n239069 , n239070 , n239071 , n239072 , n239073 , n239074 , n239075 , n239076 , n239077 , n239078 , 
 n239079 , n239080 , n239081 , n239082 , n239083 , n239084 , n239085 , n239086 , n239087 , n239088 , 
 n239089 , n239090 , n239091 , n239092 , n239093 , n239094 , n239095 , n239096 , n239097 , n239098 , 
 n239099 , n239100 , n239101 , n239102 , n239103 , n239104 , n239105 , n239106 , n239107 , n239108 , 
 n239109 , n239110 , n239111 , n239112 , n239113 , n239114 , n239115 , n239116 , n239117 , n239118 , 
 n239119 , n239120 , n239121 , n239122 , n239123 , n239124 , n239125 , n239126 , n239127 , n239128 , 
 n239129 , n239130 , n239131 , n239132 , n239133 , n239134 , n239135 , n239136 , n239137 , n239138 , 
 n239139 , n239140 , n239141 , n239142 , n239143 , n239144 , n239145 , n239146 , n239147 , n239148 , 
 n239149 , n239150 , n239151 , n239152 , n239153 , n239154 , n239155 , n239156 , n239157 , n239158 , 
 n239159 , n239160 , n239161 , n239162 , n239163 , n239164 , n239165 , n239166 , n239167 , n239168 , 
 n239169 , n239170 , n239171 , n239172 , n239173 , n239174 , n239175 , n239176 , n239177 , n239178 , 
 n239179 , n239180 , n239181 , n239182 , n239183 , n239184 , n239185 , n239186 , n239187 , n239188 , 
 n239189 , n239190 , n239191 , n239192 , n239193 , n239194 , n239195 , n239196 , n239197 , n239198 , 
 n239199 , n239200 , n239201 , n239202 , n239203 , n239204 , n239205 , n239206 , n239207 , n239208 , 
 n239209 , n239210 , n239211 , n239212 , n239213 , n239214 , n239215 , n239216 , n239217 , n239218 , 
 n239219 , n239220 , n239221 , n239222 , n239223 , n239224 , n239225 , n239226 , n239227 , n239228 , 
 n239229 , n239230 , n239231 , n239232 , n239233 , n239234 , n239235 , n239236 , n239237 , n239238 , 
 n239239 , n239240 , n239241 , n239242 , n239243 , n239244 , n239245 , n239246 , n239247 , n239248 , 
 n239249 , n239250 , n239251 , n239252 , n239253 , n239254 , n239255 , n239256 , n239257 , n239258 , 
 n239259 , n239260 , n239261 , n239262 , n239263 , n239264 , n239265 , n239266 , n239267 , n239268 , 
 n239269 , n239270 , n239271 , n239272 , n239273 , n239274 , n239275 , n239276 , n239277 , n239278 , 
 n239279 , n239280 , n239281 , n239282 , n239283 , n239284 , n239285 , n239286 , n239287 , n239288 , 
 n239289 , n239290 , n239291 , n239292 , n239293 , n239294 , n239295 , n239296 , n239297 , n239298 , 
 n239299 , n239300 , n239301 , n239302 , n239303 , n239304 , n239305 , n239306 , n239307 , n239308 , 
 n239309 , n239310 , n239311 , n239312 , n239313 , n239314 , n239315 , n239316 , n239317 , n239318 , 
 n239319 , n239320 , n239321 , n239322 , n239323 , n239324 , n239325 , n239326 , n239327 , n239328 , 
 n239329 , n239330 , n239331 , n239332 , n239333 , n239334 , n239335 , n239336 , n239337 , n239338 , 
 n239339 , n239340 , n239341 , n239342 , n239343 , n239344 , n239345 , n239346 , n239347 , n239348 , 
 n239349 , n239350 , n239351 , n239352 , n239353 , n239354 , n239355 , n239356 , n239357 , n239358 , 
 n239359 , n239360 , n239361 , n239362 , n239363 , n239364 , n239365 , n239366 , n239367 , n239368 , 
 n239369 , n239370 , n239371 , n239372 , n239373 , n239374 , n239375 , n239376 , n239377 , n239378 , 
 n239379 , n239380 , n239381 , n239382 , n239383 , n239384 , n239385 , n239386 , n239387 , n239388 , 
 n239389 , n239390 , n239391 , n239392 , n239393 , n239394 , n239395 , n239396 , n239397 , n239398 , 
 n239399 , n239400 , n239401 , n239402 , n239403 , n239404 , n239405 , n239406 , n239407 , n239408 , 
 n239409 , n239410 , n239411 , n239412 , n239413 , n239414 , n239415 , n239416 , n239417 , n239418 , 
 n239419 , n239420 , n239421 , n239422 , n239423 , n239424 , n239425 , n239426 , n239427 , n239428 , 
 n239429 , n239430 , n239431 , n239432 , n239433 , n239434 , n239435 , n239436 , n239437 , n239438 , 
 n239439 , n239440 , n239441 , n239442 , n239443 , n239444 , n239445 , n239446 , n239447 , n239448 , 
 n239449 , n239450 , n239451 , n239452 , n239453 , n239454 , n239455 , n239456 , n239457 , n239458 , 
 n239459 , n239460 , n239461 , n239462 , n239463 , n239464 , n239465 , n239466 , n239467 , n239468 , 
 n239469 , n239470 , n239471 , n239472 , n239473 , n239474 , n239475 , n239476 , n239477 , n239478 , 
 n239479 , n239480 , n239481 , n239482 , n239483 , n239484 , n239485 , n239486 , n239487 , n239488 , 
 n239489 , n239490 , n239491 , n239492 , n239493 , n239494 , n239495 , n239496 , n239497 , n239498 , 
 n239499 , n239500 , n239501 , n239502 , n239503 , n239504 , n239505 , n239506 , n239507 , n239508 , 
 n239509 , n239510 , n239511 , n239512 , n239513 , n239514 , n239515 , n239516 , n239517 , n239518 , 
 n239519 , n239520 , n239521 , n239522 , n239523 , n239524 , n239525 , n239526 , n239527 , n239528 , 
 n239529 , n239530 , n239531 , n239532 , n239533 , n239534 , n239535 , n239536 , n239537 , n239538 , 
 n239539 , n239540 , n239541 , n239542 , n239543 , n239544 , n239545 , n239546 , n239547 , n239548 , 
 n239549 , n239550 , n239551 , n239552 , n239553 , n239554 , n239555 , n239556 , n239557 , n239558 , 
 n239559 , n239560 , n239561 , n239562 , n239563 , n239564 , n239565 , n239566 , n239567 , n239568 , 
 n239569 , n239570 , n239571 , n239572 , n239573 , n239574 , n239575 , n239576 , n239577 , n239578 , 
 n239579 , n239580 , n239581 , n239582 , n239583 , n239584 , n239585 , n239586 , n239587 , n239588 , 
 n239589 , n239590 , n239591 , n239592 , n239593 , n239594 , n239595 , n239596 , n239597 , n239598 , 
 n239599 , n239600 , n239601 , n239602 , n239603 , n239604 , n239605 , n239606 , n239607 , n239608 , 
 n239609 , n239610 , n239611 , n239612 , n239613 , n239614 , n239615 , n239616 , n239617 , n239618 , 
 n239619 , n239620 , n239621 , n239622 , n239623 , n239624 , n239625 , n239626 , n239627 , n239628 , 
 n239629 , n239630 , n239631 , n239632 , n239633 , n239634 , n239635 , n239636 , n239637 , n239638 , 
 n239639 , n239640 , n239641 , n239642 , n239643 , n239644 , n239645 , n239646 , n239647 , n239648 , 
 n239649 , n239650 , n239651 , n239652 , n239653 , n239654 , n239655 , n239656 , n239657 , n239658 , 
 n239659 , n239660 , n239661 , n239662 , n239663 , n239664 , n239665 , n239666 , n239667 , n239668 , 
 n239669 , n239670 , n239671 , n239672 , n239673 , n239674 , n239675 , n239676 , n239677 , n239678 , 
 n239679 , n239680 , n239681 , n239682 , n239683 , n239684 , n239685 , n239686 , n239687 , n239688 , 
 n239689 , n239690 , n239691 , n239692 , n239693 , n239694 , n239695 , n239696 , n239697 , n239698 , 
 n239699 , n239700 , n239701 , n239702 , n239703 , n239704 , n239705 , n239706 , n239707 , n239708 , 
 n239709 , n239710 , n239711 , n239712 , n239713 , n239714 , n239715 , n239716 , n239717 , n239718 , 
 n239719 , n239720 , n239721 , n239722 , n239723 , n239724 , n239725 , n239726 , n239727 , n239728 , 
 n239729 , n239730 , n239731 , n239732 , n239733 , n239734 , n239735 , n239736 , n239737 , n239738 , 
 n239739 , n239740 , n239741 , n239742 , n239743 , n239744 , n239745 , n239746 , n239747 , n239748 , 
 n239749 , n239750 , n239751 , n239752 , n239753 , n239754 , n239755 , n239756 , n239757 , n239758 , 
 n239759 , n239760 , n239761 , n239762 , n239763 , n239764 , n239765 , n239766 , n239767 , n239768 , 
 n239769 , n239770 , n239771 , n239772 , n239773 , n239774 , n239775 , n239776 , n239777 , n239778 , 
 n239779 , n239780 , n239781 , n239782 , n239783 , n239784 , n239785 , n239786 , n239787 , n239788 , 
 n239789 , n239790 , n239791 , n239792 , n239793 , n239794 , n239795 , n239796 , n239797 , n239798 , 
 n239799 , n239800 , n239801 , n239802 , n239803 , n239804 , n239805 , n239806 , n239807 , n239808 , 
 n239809 , n239810 , n239811 , n239812 , n239813 , n239814 , n239815 , n239816 , n239817 , n239818 , 
 n239819 , n239820 , n239821 , n239822 , n239823 , n239824 , n239825 , n239826 , n239827 , n239828 , 
 n239829 , n239830 , n239831 , n239832 , n239833 , n239834 , n239835 , n239836 , n239837 , n239838 , 
 n239839 , n239840 , n239841 , n239842 , n239843 , n239844 , n239845 , n239846 , n239847 , n239848 , 
 n239849 , n239850 , n239851 , n239852 , n239853 , n239854 , n239855 , n239856 , n239857 , n239858 , 
 n239859 , n239860 , n239861 , n239862 , n239863 , n239864 , n239865 , n239866 , n239867 , n239868 , 
 n239869 , n239870 , n239871 , n239872 , n239873 , n239874 , n239875 , n239876 , n239877 , n239878 , 
 n239879 , n239880 , n239881 , n239882 , n239883 , n239884 , n239885 , n239886 , n239887 , n239888 , 
 n239889 , n239890 , n239891 , n239892 , n239893 , n239894 , n239895 , n239896 , n239897 , n239898 , 
 n239899 , n239900 , n239901 , n239902 , n239903 , n239904 , n239905 , n239906 , n239907 , n239908 , 
 n239909 , n239910 , n239911 , n239912 , n239913 , n239914 , n239915 , n239916 , n239917 , n239918 , 
 n239919 , n239920 , n239921 , n239922 , n239923 , n239924 , n239925 , n239926 , n239927 , n239928 , 
 n239929 , n239930 , n239931 , n239932 , n239933 , n239934 , n239935 , n239936 , n239937 , n239938 , 
 n239939 , n239940 , n239941 , n239942 , n239943 , n239944 , n239945 , n239946 , n239947 , n239948 , 
 n239949 , n239950 , n239951 , n239952 , n239953 , n239954 , n239955 , n239956 , n239957 , n239958 , 
 n239959 , n239960 , n239961 , n239962 , n239963 , n239964 , n239965 , n239966 , n239967 , n239968 , 
 n239969 , n239970 , n239971 , n239972 , n239973 , n239974 , n239975 , n239976 , n239977 , n239978 , 
 n239979 , n239980 , n239981 , n239982 , n239983 , n239984 , n239985 , n239986 , n239987 , n239988 , 
 n239989 , n239990 , n239991 , n239992 , n239993 , n239994 , n239995 , n239996 , n239997 , n239998 , 
 n239999 , n240000 , n240001 , n240002 , n240003 , n240004 , n240005 , n240006 , n240007 , n240008 , 
 n240009 , n240010 , n240011 , n240012 , n240013 , n240014 , n240015 , n240016 , n240017 , n240018 , 
 n240019 , n240020 , n240021 , n240022 , n240023 , n240024 , n240025 , n240026 , n240027 , n240028 , 
 n240029 , n240030 , n240031 , n240032 , n240033 , n240034 , n240035 , n240036 , n240037 , n240038 , 
 n240039 , n240040 , n240041 , n240042 , n240043 , n240044 , n240045 , n240046 , n240047 , n240048 , 
 n240049 , n240050 , n240051 , n240052 , n240053 , n240054 , n240055 , n240056 , n240057 , n240058 , 
 n240059 , n240060 , n240061 , n240062 , n240063 , n240064 , n240065 , n240066 , n240067 , n240068 , 
 n240069 , n240070 , n240071 , n240072 , n240073 , n240074 , n240075 , n240076 , n240077 , n240078 , 
 n240079 , n240080 , n240081 , n240082 , n240083 , n240084 , n240085 , n240086 , n240087 , n240088 , 
 n240089 , n240090 , n240091 , n240092 , n240093 , n240094 , n240095 , n240096 , n240097 , n240098 , 
 n240099 , n240100 , n240101 , n240102 , n240103 , n240104 , n240105 , n240106 , n240107 , n240108 , 
 n240109 , n240110 , n240111 , n240112 , n240113 , n240114 , n240115 , n240116 , n240117 , n240118 , 
 n240119 , n240120 , n240121 , n240122 , n240123 , n240124 , n240125 , n240126 , n240127 , n240128 , 
 n240129 , n240130 , n240131 , n240132 , n240133 , n240134 , n240135 , n240136 , n240137 , n240138 , 
 n240139 , n240140 , n240141 , n240142 , n240143 , n240144 , n240145 , n240146 , n240147 , n240148 , 
 n240149 , n240150 , n240151 , n240152 , n240153 , n240154 , n240155 , n240156 , n240157 , n240158 , 
 n240159 , n240160 , n240161 , n240162 , n240163 , n240164 , n240165 , n240166 , n240167 , n240168 , 
 n240169 , n240170 , n240171 , n240172 , n240173 , n240174 , n240175 , n240176 , n240177 , n240178 , 
 n240179 , n240180 , n240181 , n240182 , n240183 , n240184 , n240185 , n240186 , n240187 , n240188 , 
 n240189 , n240190 , n240191 , n240192 , n240193 , n240194 , n240195 , n240196 , n240197 , n240198 , 
 n240199 , n240200 , n240201 , n240202 , n240203 , n240204 , n240205 , n240206 , n240207 , n240208 , 
 n240209 , n240210 , n240211 , n240212 , n240213 , n240214 , n240215 , n240216 , n240217 , n240218 , 
 n240219 , n240220 , n240221 , n240222 , n240223 , n240224 , n240225 , n240226 , n240227 , n240228 , 
 n240229 , n240230 , n240231 , n240232 , n240233 , n240234 , n240235 , n240236 , n240237 , n240238 , 
 n240239 , n240240 , n240241 , n240242 , n240243 , n240244 , n240245 , n240246 , n240247 , n240248 , 
 n240249 , n240250 , n240251 , n240252 , n240253 , n240254 , n240255 , n240256 , n240257 , n240258 , 
 n240259 , n240260 , n240261 , n240262 , n240263 , n240264 , n240265 , n240266 , n240267 , n240268 , 
 n240269 , n240270 , n240271 , n240272 , n240273 , n240274 , n240275 , n240276 , n240277 , n240278 , 
 n240279 , n240280 , n240281 , n240282 , n240283 , n240284 , n240285 , n240286 , n240287 , n240288 , 
 n240289 , n240290 , n240291 , n240292 , n240293 , n240294 , n240295 , n240296 , n240297 , n240298 , 
 n240299 , n240300 , n240301 , n240302 , n240303 , n240304 , n240305 , n240306 , n240307 , n240308 , 
 n240309 , n240310 , n240311 , n240312 , n240313 , n240314 , n240315 , n240316 , n240317 , n240318 , 
 n240319 , n240320 , n240321 , n240322 , n240323 , n240324 , n240325 , n240326 , n240327 , n240328 , 
 n240329 , n240330 , n240331 , n240332 , n240333 , n240334 , n240335 , n240336 , n240337 , n240338 , 
 n240339 , n240340 , n240341 , n240342 , n240343 , n240344 , n240345 , n240346 , n240347 , n240348 , 
 n240349 , n240350 , n240351 , n240352 , n240353 , n240354 , n240355 , n240356 , n240357 , n240358 , 
 n240359 , n240360 , n240361 , n240362 , n240363 , n240364 , n240365 , n240366 , n240367 , n240368 , 
 n240369 , n240370 , n240371 , n240372 , n240373 , n240374 , n240375 , n240376 , n240377 , n240378 , 
 n240379 , n240380 , n240381 , n240382 , n240383 , n240384 , n240385 , n240386 , n240387 , n240388 , 
 n240389 , n240390 , n240391 , n240392 , n240393 , n240394 , n240395 , n240396 , n240397 , n240398 , 
 n240399 , n240400 , n240401 , n240402 , n240403 , n240404 , n240405 , n240406 , n240407 , n240408 , 
 n240409 , n240410 , n240411 , n240412 , n240413 , n240414 , n240415 , n240416 , n240417 , n240418 , 
 n240419 , n240420 , n240421 , n240422 , n240423 , n240424 , n240425 , n240426 , n240427 , n240428 , 
 n240429 , n240430 , n240431 , n240432 , n240433 , n240434 , n240435 , n240436 , n240437 , n240438 , 
 n240439 , n240440 , n240441 , n240442 , n240443 , n240444 , n240445 , n240446 , n240447 , n240448 , 
 n240449 , n240450 , n240451 , n240452 , n240453 , n240454 , n240455 , n240456 , n240457 , n240458 , 
 n240459 , n240460 , n240461 , n240462 , n240463 , n240464 , n240465 , n240466 , n240467 , n240468 , 
 n240469 , n240470 , n240471 , n240472 , n240473 , n240474 , n240475 , n240476 , n240477 , n240478 , 
 n240479 , n240480 , n240481 , n240482 , n240483 , n240484 , n240485 , n240486 , n240487 , n240488 , 
 n240489 , n240490 , n240491 , n240492 , n240493 , n240494 , n240495 , n240496 , n240497 , n240498 , 
 n240499 , n240500 , n240501 , n240502 , n240503 , n240504 , n240505 , n240506 , n240507 , n240508 , 
 n240509 , n240510 , n240511 , n240512 , n240513 , n240514 , n240515 , n240516 , n240517 , n240518 , 
 n240519 , n240520 , n240521 , n240522 , n240523 , n240524 , n240525 , n240526 , n240527 , n240528 , 
 n240529 , n240530 , n240531 , n240532 , n240533 , n240534 , n240535 , n240536 , n240537 , n240538 , 
 n240539 , n240540 , n240541 , n240542 , n240543 , n240544 , n240545 , n240546 , n240547 , n240548 , 
 n240549 , n240550 , n240551 , n240552 , n240553 , n240554 , n240555 , n240556 , n240557 , n240558 , 
 n240559 , n240560 , n240561 , n240562 , n240563 , n240564 , n240565 , n240566 , n240567 , n240568 , 
 n240569 , n240570 , n240571 , n240572 , n240573 , n240574 , n240575 , n240576 , n240577 , n240578 , 
 n240579 , n240580 , n240581 , n240582 , n240583 , n240584 , n240585 , n240586 , n240587 , n240588 , 
 n240589 , n240590 , n240591 , n240592 , n240593 , n240594 , n240595 , n240596 , n240597 , n240598 , 
 n240599 , n240600 , n240601 , n240602 , n240603 , n240604 , n240605 , n240606 , n240607 , n240608 , 
 n240609 , n240610 , n240611 , n240612 , n240613 , n240614 , n240615 , n240616 , n240617 , n240618 , 
 n240619 , n240620 , n240621 , n240622 , n240623 , n240624 , n240625 , n240626 , n240627 , n240628 , 
 n240629 , n240630 , n240631 , n240632 , n240633 , n240634 , n240635 , n240636 , n240637 , n240638 , 
 n240639 , n240640 , n240641 , n240642 , n240643 , n240644 , n240645 , n240646 , n240647 , n240648 , 
 n240649 , n240650 , n240651 , n240652 , n240653 , n240654 , n240655 , n240656 , n240657 , n240658 , 
 n240659 , n240660 , n240661 , n240662 , n240663 , n240664 , n240665 , n240666 , n240667 , n240668 , 
 n240669 , n240670 , n240671 , n240672 , n240673 , n240674 , n240675 , n240676 , n240677 , n240678 , 
 n240679 , n240680 , n240681 , n240682 , n240683 , n240684 , n240685 , n240686 , n240687 , n240688 , 
 n240689 , n240690 , n240691 , n240692 , n240693 , n240694 , n240695 , n240696 , n240697 , n240698 , 
 n240699 , n240700 , n240701 , n240702 , n240703 , n240704 , n240705 , n240706 , n240707 , n240708 , 
 n240709 , n240710 , n240711 , n240712 , n240713 , n240714 , n240715 , n240716 , n240717 , n240718 , 
 n240719 , n240720 , n240721 , n240722 , n240723 , n240724 , n240725 , n240726 , n240727 , n240728 , 
 n240729 , n240730 , n240731 , n240732 , n240733 , n240734 , n240735 , n240736 , n240737 , n240738 , 
 n240739 , n240740 , n240741 , n240742 , n240743 , n240744 , n240745 , n240746 , n240747 , n240748 , 
 n240749 , n240750 , n240751 , n240752 , n240753 , n240754 , n240755 , n240756 , n240757 , n240758 , 
 n240759 , n240760 , n240761 , n240762 , n240763 , n240764 , n240765 , n240766 , n240767 , n240768 , 
 n240769 , n240770 , n240771 , n240772 , n240773 , n240774 , n240775 , n240776 , n240777 , n240778 , 
 n240779 , n240780 , n240781 , n240782 , n240783 , n240784 , n240785 , n240786 , n240787 , n240788 , 
 n240789 , n240790 , n240791 , n240792 , n240793 , n240794 , n240795 , n240796 , n240797 , n240798 , 
 n240799 , n240800 , n240801 , n240802 , n240803 , n240804 , n240805 , n240806 , n240807 , n240808 , 
 n240809 , n240810 , n240811 , n240812 , n240813 , n240814 , n240815 , n240816 , n240817 , n240818 , 
 n240819 , n240820 , n240821 , n240822 , n240823 , n240824 , n240825 , n240826 , n240827 , n240828 , 
 n240829 , n240830 , n240831 , n240832 , n240833 , n240834 , n240835 , n240836 , n240837 , n240838 , 
 n240839 , n240840 , n240841 , n240842 , n240843 , n240844 , n240845 , n240846 , n240847 , n240848 , 
 n240849 , n240850 , n240851 , n240852 , n240853 , n240854 , n240855 , n240856 , n240857 , n240858 , 
 n240859 , n240860 , n240861 , n240862 , n240863 , n240864 , n240865 , n240866 , n240867 , n240868 , 
 n240869 , n240870 , n240871 , n240872 , n240873 , n240874 , n240875 , n240876 , n240877 , n240878 , 
 n240879 , n240880 , n240881 , n240882 , n240883 , n240884 , n240885 , n240886 , n240887 , n240888 , 
 n240889 , n240890 , n240891 , n240892 , n240893 , n240894 , n240895 , n240896 , n240897 , n240898 , 
 n240899 , n240900 , n240901 , n240902 , n240903 , n240904 , n240905 , n240906 , n240907 , n240908 , 
 n240909 , n240910 , n240911 , n240912 , n240913 , n240914 , n240915 , n240916 , n240917 , n240918 , 
 n240919 , n240920 , n240921 , n240922 , n240923 , n240924 , n240925 , n240926 , n240927 , n240928 , 
 n240929 , n240930 , n240931 , n240932 , n240933 , n240934 , n240935 , n240936 , n240937 , n240938 , 
 n240939 , n240940 , n240941 , n240942 , n240943 , n240944 , n240945 , n240946 , n240947 , n240948 , 
 n240949 , n240950 , n240951 , n240952 , n240953 , n240954 , n240955 , n240956 , n240957 , n240958 , 
 n240959 , n240960 , n240961 , n240962 , n240963 , n240964 , n240965 , n240966 , n240967 , n240968 , 
 n240969 , n240970 , n240971 , n240972 , n240973 , n240974 , n240975 , n240976 , n240977 , n240978 , 
 n240979 , n240980 , n240981 , n240982 , n240983 , n240984 , n240985 , n240986 , n240987 , n240988 , 
 n240989 , n240990 , n240991 , n240992 , n240993 , n240994 , n240995 , n240996 , n240997 , n240998 , 
 n240999 , n241000 , n241001 , n241002 , n241003 , n241004 , n241005 , n241006 , n241007 , n241008 , 
 n241009 , n241010 , n241011 , n241012 , n241013 , n241014 , n241015 , n241016 , n241017 , n241018 , 
 n241019 , n241020 , n241021 , n241022 , n241023 , n241024 , n241025 , n241026 , n241027 , n241028 , 
 n241029 , n241030 , n241031 , n241032 , n241033 , n241034 , n241035 , n241036 , n241037 , n241038 , 
 n241039 , n241040 , n241041 , n241042 , n241043 , n241044 , n241045 , n241046 , n241047 , n241048 , 
 n241049 , n241050 , n241051 , n241052 , n241053 , n241054 , n241055 , n241056 , n241057 , n241058 , 
 n241059 , n241060 , n241061 , n241062 , n241063 , n241064 , n241065 , n241066 , n241067 , n241068 , 
 n241069 , n241070 , n241071 , n241072 , n241073 , n241074 , n241075 , n241076 , n241077 , n241078 , 
 n241079 , n241080 , n241081 , n241082 , n241083 , n241084 , n241085 , n241086 , n241087 , n241088 , 
 n241089 , n241090 , n241091 , n241092 , n241093 , n241094 , n241095 , n241096 , n241097 , n241098 , 
 n241099 , n241100 , n241101 , n241102 , n241103 , n241104 , n241105 , n241106 , n241107 , n241108 , 
 n241109 , n241110 , n241111 , n241112 , n241113 , n241114 , n241115 , n241116 , n241117 , n241118 , 
 n241119 , n241120 , n241121 , n241122 , n241123 , n241124 , n241125 , n241126 , n241127 , n241128 , 
 n241129 , n241130 , n241131 , n241132 , n241133 , n241134 , n241135 , n241136 , n241137 , n241138 , 
 n241139 , n241140 , n241141 , n241142 , n241143 , n241144 , n241145 , n241146 , n241147 , n241148 , 
 n241149 , n241150 , n241151 , n241152 , n241153 , n241154 , n241155 , n241156 , n241157 , n241158 , 
 n241159 , n241160 , n241161 , n241162 , n241163 , n241164 , n241165 , n241166 , n241167 , n241168 , 
 n241169 , n241170 , n241171 , n241172 , n241173 , n241174 , n241175 , n241176 , n241177 , n241178 , 
 n241179 , n241180 , n241181 , n241182 , n241183 , n241184 , n241185 , n241186 , n241187 , n241188 , 
 n241189 , n241190 , n241191 , n241192 , n241193 , n241194 , n241195 , n241196 , n241197 , n241198 , 
 n241199 , n241200 , n241201 , n241202 , n241203 , n241204 , n241205 , n241206 , n241207 , n241208 , 
 n241209 , n241210 , n241211 , n241212 , n241213 , n241214 , n241215 , n241216 , n241217 , n241218 , 
 n241219 , n241220 , n241221 , n241222 , n241223 , n241224 , n241225 , n241226 , n241227 , n241228 , 
 n241229 , n241230 , n241231 , n241232 , n241233 , n241234 , n241235 , n241236 , n241237 , n241238 , 
 n241239 , n241240 , n241241 , n241242 , n241243 , n241244 , n241245 , n241246 , n241247 , n241248 , 
 n241249 , n241250 , n241251 , n241252 , n241253 , n241254 , n241255 , n241256 , n241257 , n241258 , 
 n241259 , n241260 , n241261 , n241262 , n241263 , n241264 , n241265 , n241266 , n241267 , n241268 , 
 n241269 , n241270 , n241271 , n241272 , n241273 , n241274 , n241275 , n241276 , n241277 , n241278 , 
 n241279 , n241280 , n241281 , n241282 , n241283 , n241284 , n241285 , n241286 , n241287 , n241288 , 
 n241289 , n241290 , n241291 , n241292 , n241293 , n241294 , n241295 , n241296 , n241297 , n241298 , 
 n241299 , n241300 , n241301 , n241302 , n241303 , n241304 , n241305 , n241306 , n241307 , n241308 , 
 n241309 , n241310 , n241311 , n241312 , n241313 , n241314 , n241315 , n241316 , n241317 , n241318 , 
 n241319 , n241320 , n241321 , n241322 , n241323 , n241324 , n241325 , n241326 , n241327 , n241328 , 
 n241329 , n241330 , n241331 , n241332 , n241333 , n241334 , n241335 , n241336 , n241337 , n241338 , 
 n241339 , n241340 , n241341 , n241342 , n241343 , n241344 , n241345 , n241346 , n241347 , n241348 , 
 n241349 , n241350 , n241351 , n241352 , n241353 , n241354 , n241355 , n241356 , n241357 , n241358 , 
 n241359 , n241360 , n241361 , n241362 , n241363 , n241364 , n241365 , n241366 , n241367 , n241368 , 
 n241369 , n241370 , n241371 , n241372 , n241373 , n241374 , n241375 , n241376 , n241377 , n241378 , 
 n241379 , n241380 , n241381 , n241382 , n241383 , n241384 , n241385 , n241386 , n241387 , n241388 , 
 n241389 , n241390 , n241391 , n241392 , n241393 , n241394 , n241395 , n241396 , n241397 , n241398 , 
 n241399 , n241400 , n241401 , n241402 , n241403 , n241404 , n241405 , n241406 , n241407 , n241408 , 
 n241409 , n241410 , n241411 , n241412 , n241413 , n241414 , n241415 , n241416 , n241417 , n241418 , 
 n241419 , n241420 , n241421 , n241422 , n241423 , n241424 , n241425 , n241426 , n241427 , n241428 , 
 n241429 , n241430 , n241431 , n241432 , n241433 , n241434 , n241435 , n241436 , n241437 , n241438 , 
 n241439 , n241440 , n241441 , n241442 , n241443 , n241444 , n241445 , n241446 , n241447 , n241448 , 
 n241449 , n241450 , n241451 , n241452 , n241453 , n241454 , n241455 , n241456 , n241457 , n241458 , 
 n241459 , n241460 , n241461 , n241462 , n241463 , n241464 , n241465 , n241466 , n241467 , n241468 , 
 n241469 , n241470 , n241471 , n241472 , n241473 , n241474 , n241475 , n241476 , n241477 , n241478 , 
 n241479 , n241480 , n241481 , n241482 , n241483 , n241484 , n241485 , n241486 , n241487 , n241488 , 
 n241489 , n241490 , n241491 , n241492 , n241493 , n241494 , n241495 , n241496 , n241497 , n241498 , 
 n241499 , n241500 , n241501 , n241502 , n241503 , n241504 , n241505 , n241506 , n241507 , n241508 , 
 n241509 , n241510 , n241511 , n241512 , n241513 , n241514 , n241515 , n241516 , n241517 , n241518 , 
 n241519 , n241520 , n241521 , n241522 , n241523 , n241524 , n241525 , n241526 , n241527 , n241528 , 
 n241529 , n241530 , n241531 , n241532 , n241533 , n241534 , n241535 , n241536 , n241537 , n241538 , 
 n241539 , n241540 , n241541 , n241542 , n241543 , n241544 , n241545 , n241546 , n241547 , n241548 , 
 n241549 , n241550 , n241551 , n241552 , n241553 , n241554 , n241555 , n241556 , n241557 , n241558 , 
 n241559 , n241560 , n241561 , n241562 , n241563 , n241564 , n241565 , n241566 , n241567 , n241568 , 
 n241569 , n241570 , n241571 , n241572 , n241573 , n241574 , n241575 , n241576 , n241577 , n241578 , 
 n241579 , n241580 , n241581 , n241582 , n241583 , n241584 , n241585 , n241586 , n241587 , n241588 , 
 n241589 , n241590 , n241591 , n241592 , n241593 , n241594 , n241595 , n241596 , n241597 , n241598 , 
 n241599 , n241600 , n241601 , n241602 , n241603 , n241604 , n241605 , n241606 , n241607 , n241608 , 
 n241609 , n241610 , n241611 , n241612 , n241613 , n241614 , n241615 , n241616 , n241617 , n241618 , 
 n241619 , n241620 , n241621 , n241622 , n241623 , n241624 , n241625 , n241626 , n241627 , n241628 , 
 n241629 , n241630 , n241631 , n241632 , n241633 , n241634 , n241635 , n241636 , n241637 , n241638 , 
 n241639 , n241640 , n241641 , n241642 , n241643 , n241644 , n241645 , n241646 , n241647 , n241648 , 
 n241649 , n241650 , n241651 , n241652 , n241653 , n241654 , n241655 , n241656 , n241657 , n241658 , 
 n241659 , n241660 , n241661 , n241662 , n241663 , n241664 , n241665 , n241666 , n241667 , n241668 , 
 n241669 , n241670 , n241671 , n241672 , n241673 , n241674 , n241675 , n241676 , n241677 , n241678 , 
 n241679 , n241680 , n241681 , n241682 , n241683 , n241684 , n241685 , n241686 , n241687 , n241688 , 
 n241689 , n241690 , n241691 , n241692 , n241693 , n241694 , n241695 , n241696 , n241697 , n241698 , 
 n241699 , n241700 , n241701 , n241702 , n241703 , n241704 , n241705 , n241706 , n241707 , n241708 , 
 n241709 , n241710 , n241711 , n241712 , n241713 , n241714 , n241715 , n241716 , n241717 , n241718 , 
 n241719 , n241720 , n241721 , n241722 , n241723 , n241724 , n241725 , n241726 , n241727 , n241728 , 
 n241729 , n241730 , n241731 , n241732 , n241733 , n241734 , n241735 , n241736 , n241737 , n241738 , 
 n241739 , n241740 , n241741 , n241742 , n241743 , n241744 , n241745 , n241746 , n241747 , n241748 , 
 n241749 , n241750 , n241751 , n241752 , n241753 , n241754 , n241755 , n241756 , n241757 , n241758 , 
 n241759 , n241760 , n241761 , n241762 , n241763 , n241764 , n241765 , n241766 , n241767 , n241768 , 
 n241769 , n241770 , n241771 , n241772 , n241773 , n241774 , n241775 , n241776 , n241777 , n241778 , 
 n241779 , n241780 , n241781 , n241782 , n241783 , n241784 , n241785 , n241786 , n241787 , n241788 , 
 n241789 , n241790 , n241791 , n241792 , n241793 , n241794 , n241795 , n241796 , n241797 , n241798 , 
 n241799 , n241800 , n241801 , n241802 , n241803 , n241804 , n241805 , n241806 , n241807 , n241808 , 
 n241809 , n241810 , n241811 , n241812 , n241813 , n241814 , n241815 , n241816 , n241817 , n241818 , 
 n241819 , n241820 , n241821 , n241822 , n241823 , n241824 , n241825 , n241826 , n241827 , n241828 , 
 n241829 , n241830 , n241831 , n241832 , n241833 , n241834 , n241835 , n241836 , n241837 , n241838 , 
 n241839 , n241840 , n241841 , n241842 , n241843 , n241844 , n241845 , n241846 , n241847 , n241848 , 
 n241849 , n241850 , n241851 , n241852 , n241853 , n241854 , n241855 , n241856 , n241857 , n241858 , 
 n241859 , n241860 , n241861 , n241862 , n241863 , n241864 , n241865 , n241866 , n241867 , n241868 , 
 n241869 , n241870 , n241871 , n241872 , n241873 , n241874 , n241875 , n241876 , n241877 , n241878 , 
 n241879 , n241880 , n241881 , n241882 , n241883 , n241884 , n241885 , n241886 , n241887 , n241888 , 
 n241889 , n241890 , n241891 , n241892 , n241893 , n241894 , n241895 , n241896 , n241897 , n241898 , 
 n241899 , n241900 , n241901 , n241902 , n241903 , n241904 , n241905 , n241906 , n241907 , n241908 , 
 n241909 , n241910 , n241911 , n241912 , n241913 , n241914 , n241915 , n241916 , n241917 , n241918 , 
 n241919 , n241920 , n241921 , n241922 , n241923 , n241924 , n241925 , n241926 , n241927 , n241928 , 
 n241929 , n241930 , n241931 , n241932 , n241933 , n241934 , n241935 , n241936 , n241937 , n241938 , 
 n241939 , n241940 , n241941 , n241942 , n241943 , n241944 , n241945 , n241946 , n241947 , n241948 , 
 n241949 , n241950 , n241951 , n241952 , n241953 , n241954 , n241955 , n241956 , n241957 , n241958 , 
 n241959 , n241960 , n241961 , n241962 , n241963 , n241964 , n241965 , n241966 , n241967 , n241968 , 
 n241969 , n241970 , n241971 , n241972 , n241973 , n241974 , n241975 , n241976 , n241977 , n241978 , 
 n241979 , n241980 , n241981 , n241982 , n241983 , n241984 , n241985 , n241986 , n241987 , n241988 , 
 n241989 , n241990 , n241991 , n241992 , n241993 , n241994 , n241995 , n241996 , n241997 , n241998 , 
 n241999 , n242000 , n242001 , n242002 , n242003 , n242004 , n242005 , n242006 , n242007 , n242008 , 
 n242009 , n242010 , n242011 , n242012 , n242013 , n242014 , n242015 , n242016 , n242017 , n242018 , 
 n242019 , n242020 , n242021 , n242022 , n242023 , n242024 , n242025 , n242026 , n242027 , n242028 , 
 n242029 , n242030 , n242031 , n242032 , n242033 , n242034 , n242035 , n242036 , n242037 , n242038 , 
 n242039 , n242040 , n242041 , n242042 , n242043 , n242044 , n242045 , n242046 , n242047 , n242048 , 
 n242049 , n242050 , n242051 , n242052 , n242053 , n242054 , n242055 , n242056 , n242057 , n242058 , 
 n242059 , n242060 , n242061 , n242062 , n242063 , n242064 , n242065 , n242066 , n242067 , n242068 , 
 n242069 , n242070 , n242071 , n242072 , n242073 , n242074 , n242075 , n242076 , n242077 , n242078 , 
 n242079 , n242080 , n242081 , n242082 , n242083 , n242084 , n242085 , n242086 , n242087 , n242088 , 
 n242089 , n242090 , n242091 , n242092 , n242093 , n242094 , n242095 , n242096 , n242097 , n242098 , 
 n242099 , n242100 , n242101 , n242102 , n242103 , n242104 , n242105 , n242106 , n242107 , n242108 , 
 n242109 , n242110 , n242111 , n242112 , n242113 , n242114 , n242115 , n242116 , n242117 , n242118 , 
 n242119 , n242120 , n242121 , n242122 , n242123 , n242124 , n242125 , n242126 , n242127 , n242128 , 
 n242129 , n242130 , n242131 , n242132 , n242133 , n242134 , n242135 , n242136 , n242137 , n242138 , 
 n242139 , n242140 , n242141 , n242142 , n242143 , n242144 , n242145 , n242146 , n242147 , n242148 , 
 n242149 , n242150 , n242151 , n242152 , n242153 , n242154 , n242155 , n242156 , n242157 , n242158 , 
 n242159 , n242160 , n242161 , n242162 , n242163 , n242164 , n242165 , n242166 , n242167 , n242168 , 
 n242169 , n242170 , n242171 , n242172 , n242173 , n242174 , n242175 , n242176 , n242177 , n242178 , 
 n242179 , n242180 , n242181 , n242182 , n242183 , n242184 , n242185 , n242186 , n242187 , n242188 , 
 n242189 , n242190 , n242191 , n242192 , n242193 , n242194 , n242195 , n242196 , n242197 , n242198 , 
 n242199 , n242200 , n242201 , n242202 , n242203 , n242204 , n242205 , n242206 , n242207 , n242208 , 
 n242209 , n242210 , n242211 , n242212 , n242213 , n242214 , n242215 , n242216 , n242217 , n242218 , 
 n242219 , n242220 , n242221 , n242222 , n242223 , n242224 , n242225 , n242226 , n242227 , n242228 , 
 n242229 , n242230 , n242231 , n242232 , n242233 , n242234 , n242235 , n242236 , n242237 , n242238 , 
 n242239 , n242240 , n242241 , n242242 , n242243 , n242244 , n242245 , n242246 , n242247 , n242248 , 
 n242249 , n242250 , n242251 , n242252 , n242253 , n242254 , n242255 , n242256 , n242257 , n242258 , 
 n242259 , n242260 , n242261 , n242262 , n242263 , n242264 , n242265 , n242266 , n242267 , n242268 , 
 n242269 , n242270 , n242271 , n242272 , n242273 , n242274 , n242275 , n242276 , n242277 , n242278 , 
 n242279 , n242280 , n242281 , n242282 , n242283 , n242284 , n242285 , n242286 , n242287 , n242288 , 
 n242289 , n242290 , n242291 , n242292 , n242293 , n242294 , n242295 , n242296 , n242297 , n242298 , 
 n242299 , n242300 , n242301 , n242302 , n242303 , n242304 , n242305 , n242306 , n242307 , n242308 , 
 n242309 , n242310 , n242311 , n242312 , n242313 , n242314 , n242315 , n242316 , n242317 , n242318 , 
 n242319 , n242320 , n242321 , n242322 , n242323 , n242324 , n242325 , n242326 , n242327 , n242328 , 
 n242329 , n242330 , n242331 , n242332 , n242333 , n242334 , n242335 , n242336 , n242337 , n242338 , 
 n242339 , n242340 , n242341 , n242342 , n242343 , n242344 , n242345 , n242346 , n242347 , n242348 , 
 n242349 , n242350 , n242351 , n242352 , n242353 , n242354 , n242355 , n242356 , n242357 , n242358 , 
 n242359 , n242360 , n242361 , n242362 , n242363 , n242364 , n242365 , n242366 , n242367 , n242368 , 
 n242369 , n242370 , n242371 , n242372 , n242373 , n242374 , n242375 , n242376 , n242377 , n242378 , 
 n242379 , n242380 , n242381 , n242382 , n242383 , n242384 , n242385 , n242386 , n242387 , n242388 , 
 n242389 , n242390 , n242391 , n242392 , n242393 , n242394 , n242395 , n242396 , n242397 , n242398 , 
 n242399 , n242400 , n242401 , n242402 , n242403 , n242404 , n242405 , n242406 , n242407 , n242408 , 
 n242409 , n242410 , n242411 , n242412 , n242413 , n242414 , n242415 , n242416 , n242417 , n242418 , 
 n242419 , n242420 , n242421 , n242422 , n242423 , n242424 , n242425 , n242426 , n242427 , n242428 , 
 n242429 , n242430 , n242431 , n242432 , n242433 , n242434 , n242435 , n242436 , n242437 , n242438 , 
 n242439 , n242440 , n242441 , n242442 , n242443 , n242444 , n242445 , n242446 , n242447 , n242448 , 
 n242449 , n242450 , n242451 , n242452 , n242453 , n242454 , n242455 , n242456 , n242457 , n242458 , 
 n242459 , n242460 , n242461 , n242462 , n242463 , n242464 , n242465 , n242466 , n242467 , n242468 , 
 n242469 , n242470 , n242471 , n242472 , n242473 , n242474 , n242475 , n242476 , n242477 , n242478 , 
 n242479 , n242480 , n242481 , n242482 , n242483 , n242484 , n242485 , n242486 , n242487 , n242488 , 
 n242489 , n242490 , n242491 , n242492 , n242493 , n242494 , n242495 , n242496 , n242497 , n242498 , 
 n242499 , n242500 , n242501 , n242502 , n242503 , n242504 , n242505 , n242506 , n242507 , n242508 , 
 n242509 , n242510 , n242511 , n242512 , n242513 , n242514 , n242515 , n242516 , n242517 , n242518 , 
 n242519 , n242520 , n242521 , n242522 , n242523 , n242524 , n242525 , n242526 , n242527 , n242528 , 
 n242529 , n242530 , n242531 , n242532 , n242533 , n242534 , n242535 , n242536 , n242537 , n242538 , 
 n242539 , n242540 , n242541 , n242542 , n242543 , n242544 , n242545 , n242546 , n242547 , n242548 , 
 n242549 , n242550 , n242551 , n242552 , n242553 , n242554 , n242555 , n242556 , n242557 , n242558 , 
 n242559 , n242560 , n242561 , n242562 , n242563 , n242564 , n242565 , n242566 , n242567 , n242568 , 
 n242569 , n242570 , n242571 , n242572 , n242573 , n242574 , n242575 , n242576 , n242577 , n242578 , 
 n242579 , n242580 , n242581 , n242582 , n242583 , n242584 , n242585 , n242586 , n242587 , n242588 , 
 n242589 , n242590 , n242591 , n242592 , n242593 , n242594 , n242595 , n242596 , n242597 , n242598 , 
 n242599 , n242600 , n242601 , n242602 , n242603 , n242604 , n242605 , n242606 , n242607 , n242608 , 
 n242609 , n242610 , n242611 , n242612 , n242613 , n242614 , n242615 , n242616 , n242617 , n242618 , 
 n242619 , n242620 , n242621 , n242622 , n242623 , n242624 , n242625 , n242626 , n242627 , n242628 , 
 n242629 , n242630 , n242631 , n242632 , n242633 , n242634 , n242635 , n242636 , n242637 , n242638 , 
 n242639 , n242640 , n242641 , n242642 , n242643 , n242644 , n242645 , n242646 , n242647 , n242648 , 
 n242649 , n242650 , n242651 , n242652 , n242653 , n242654 , n242655 , n242656 , n242657 , n242658 , 
 n242659 , n242660 , n242661 , n242662 , n242663 , n242664 , n242665 , n242666 , n242667 , n242668 , 
 n242669 , n242670 , n242671 , n242672 , n242673 , n242674 , n242675 , n242676 , n242677 , n242678 , 
 n242679 , n242680 , n242681 , n242682 , n242683 , n242684 , n242685 , n242686 , n242687 , n242688 , 
 n242689 , n242690 , n242691 , n242692 , n242693 , n242694 , n242695 , n242696 , n242697 , n242698 , 
 n242699 , n242700 , n242701 , n242702 , n242703 , n242704 , n242705 , n242706 , n242707 , n242708 , 
 n242709 , n242710 , n242711 , n242712 , n242713 , n242714 , n242715 , n242716 , n242717 , n242718 , 
 n242719 , n242720 , n242721 , n242722 , n242723 , n242724 , n242725 , n242726 , n242727 , n242728 , 
 n242729 , n242730 , n242731 , n242732 , n242733 , n242734 , n242735 , n242736 , n242737 , n242738 , 
 n242739 , n242740 , n242741 , n242742 , n242743 , n242744 , n242745 , n242746 , n242747 , n242748 , 
 n242749 , n242750 , n242751 , n242752 , n242753 , n242754 , n242755 , n242756 , n242757 , n242758 , 
 n242759 , n242760 , n242761 , n242762 , n242763 , n242764 , n242765 , n242766 , n242767 , n242768 , 
 n242769 , n242770 , n242771 , n242772 , n242773 , n242774 , n242775 , n242776 , n242777 , n242778 , 
 n242779 , n242780 , n242781 , n242782 , n242783 , n242784 , n242785 , n242786 , n242787 , n242788 , 
 n242789 , n242790 , n242791 , n242792 , n242793 , n242794 , n242795 , n242796 , n242797 , n242798 , 
 n242799 , n242800 , n242801 , n242802 , n242803 , n242804 , n242805 , n242806 , n242807 , n242808 , 
 n242809 , n242810 , n242811 , n242812 , n242813 , n242814 , n242815 , n242816 , n242817 , n242818 , 
 n242819 , n242820 , n242821 , n242822 , n242823 , n242824 , n242825 , n242826 , n242827 , n242828 , 
 n242829 , n242830 , n242831 , n242832 , n242833 , n242834 , n242835 , n242836 , n242837 , n242838 , 
 n242839 , n242840 , n242841 , n242842 , n242843 , n242844 , n242845 , n242846 , n242847 , n242848 , 
 n242849 , n242850 , n242851 , n242852 , n242853 , n242854 , n242855 , n242856 , n242857 , n242858 , 
 n242859 , n242860 , n242861 , n242862 , n242863 , n242864 , n242865 , n242866 , n242867 , n242868 , 
 n242869 , n242870 , n242871 , n242872 , n242873 , n242874 , n242875 , n242876 , n242877 , n242878 , 
 n242879 , n242880 , n242881 , n242882 , n242883 , n242884 , n242885 , n242886 , n242887 , n242888 , 
 n242889 , n242890 , n242891 , n242892 , n242893 , n242894 , n242895 , n242896 , n242897 , n242898 , 
 n242899 , n242900 , n242901 , n242902 , n242903 , n242904 , n242905 , n242906 , n242907 , n242908 , 
 n242909 , n242910 , n242911 , n242912 , n242913 , n242914 , n242915 , n242916 , n242917 , n242918 , 
 n242919 , n242920 , n242921 , n242922 , n242923 , n242924 , n242925 , n242926 , n242927 , n242928 , 
 n242929 , n242930 , n242931 , n242932 , n242933 , n242934 , n242935 , n242936 , n242937 , n242938 , 
 n242939 , n242940 , n242941 , n242942 , n242943 , n242944 , n242945 , n242946 , n242947 , n242948 , 
 n242949 , n242950 , n242951 , n242952 , n242953 , n242954 , n242955 , n242956 , n242957 , n242958 , 
 n242959 , n242960 , n242961 , n242962 , n242963 , n242964 , n242965 , n242966 , n242967 , n242968 , 
 n242969 , n242970 , n242971 , n242972 , n242973 , n242974 , n242975 , n242976 , n242977 , n242978 , 
 n242979 , n242980 , n242981 , n242982 , n242983 , n242984 , n242985 , n242986 , n242987 , n242988 , 
 n242989 , n242990 , n242991 , n242992 , n242993 , n242994 , n242995 , n242996 , n242997 , n242998 , 
 n242999 , n243000 , n243001 , n243002 , n243003 , n243004 , n243005 , n243006 , n243007 , n243008 , 
 n243009 , n243010 , n243011 , n243012 , n243013 , n243014 , n243015 , n243016 , n243017 , n243018 , 
 n243019 , n243020 , n243021 , n243022 , n243023 , n243024 , n243025 , n243026 , n243027 , n243028 , 
 n243029 , n243030 , n243031 , n243032 , n243033 , n243034 , n243035 , n243036 , n243037 , n243038 , 
 n243039 , n243040 , n243041 , n243042 , n243043 , n243044 , n243045 , n243046 , n243047 , n243048 , 
 n243049 , n243050 , n243051 , n243052 , n243053 , n243054 , n243055 , n243056 , n243057 , n243058 , 
 n243059 , n243060 , n243061 , n243062 , n243063 , n243064 , n243065 , n243066 , n243067 , n243068 , 
 n243069 , n243070 , n243071 , n243072 , n243073 , n243074 , n243075 , n243076 , n243077 , n243078 , 
 n243079 , n243080 , n243081 , n243082 , n243083 , n243084 , n243085 , n243086 , n243087 , n243088 , 
 n243089 , n243090 , n243091 , n243092 , n243093 , n243094 , n243095 , n243096 , n243097 , n243098 , 
 n243099 , n243100 , n243101 , n243102 , n243103 , n243104 , n243105 , n243106 , n243107 , n243108 , 
 n243109 , n243110 , n243111 , n243112 , n243113 , n243114 , n243115 , n243116 , n243117 , n243118 , 
 n243119 , n243120 , n243121 , n243122 , n243123 , n243124 , n243125 , n243126 , n243127 , n243128 , 
 n243129 , n243130 , n243131 , n243132 , n243133 , n243134 , n243135 , n243136 , n243137 , n243138 , 
 n243139 , n243140 , n243141 , n243142 , n243143 , n243144 , n243145 , n243146 , n243147 , n243148 , 
 n243149 , n243150 , n243151 , n243152 , n243153 , n243154 , n243155 , n243156 , n243157 , n243158 , 
 n243159 , n243160 , n243161 , n243162 , n243163 , n243164 , n243165 , n243166 , n243167 , n243168 , 
 n243169 , n243170 , n243171 , n243172 , n243173 , n243174 , n243175 , n243176 , n243177 , n243178 , 
 n243179 , n243180 , n243181 , n243182 , n243183 , n243184 , n243185 , n243186 , n243187 , n243188 , 
 n243189 , n243190 , n243191 , n243192 , n243193 , n243194 , n243195 , n243196 , n243197 , n243198 , 
 n243199 , n243200 , n243201 , n243202 , n243203 , n243204 , n243205 , n243206 , n243207 , n243208 , 
 n243209 , n243210 , n243211 , n243212 , n243213 , n243214 , n243215 , n243216 , n243217 , n243218 , 
 n243219 , n243220 , n243221 , n243222 , n243223 , n243224 , n243225 , n243226 , n243227 , n243228 , 
 n243229 , n243230 , n243231 , n243232 , n243233 , n243234 , n243235 , n243236 , n243237 , n243238 , 
 n243239 , n243240 , n243241 , n243242 , n243243 , n243244 , n243245 , n243246 , n243247 , n243248 , 
 n243249 , n243250 , n243251 , n243252 , n243253 , n243254 , n243255 , n243256 , n243257 , n243258 , 
 n243259 , n243260 , n243261 , n243262 , n243263 , n243264 , n243265 , n243266 , n243267 , n243268 , 
 n243269 , n243270 , n243271 , n243272 , n243273 , n243274 , n243275 , n243276 , n243277 , n243278 , 
 n243279 , n243280 , n243281 , n243282 , n243283 , n243284 , n243285 , n243286 , n243287 , n243288 , 
 n243289 , n243290 , n243291 , n243292 , n243293 , n243294 , n243295 , n243296 , n243297 , n243298 , 
 n243299 , n243300 , n243301 , n243302 , n243303 , n243304 , n243305 , n243306 , n243307 , n243308 , 
 n243309 , n243310 , n243311 , n243312 , n243313 , n243314 , n243315 , n243316 , n243317 , n243318 , 
 n243319 , n243320 , n243321 , n243322 , n243323 , n243324 , n243325 , n243326 , n243327 , n243328 , 
 n243329 , n243330 , n243331 , n243332 , n243333 , n243334 , n243335 , n243336 , n243337 , n243338 , 
 n243339 , n243340 , n243341 , n243342 , n243343 , n243344 , n243345 , n243346 , n243347 , n243348 , 
 n243349 , n243350 , n243351 , n243352 , n243353 , n243354 , n243355 , n243356 , n243357 , n243358 , 
 n243359 , n243360 , n243361 , n243362 , n243363 , n243364 , n243365 , n243366 , n243367 , n243368 , 
 n243369 , n243370 , n243371 , n243372 , n243373 , n243374 , n243375 , n243376 , n243377 , n243378 , 
 n243379 , n243380 , n243381 , n243382 , n243383 , n243384 , n243385 , n243386 , n243387 , n243388 , 
 n243389 , n243390 , n243391 , n243392 , n243393 , n243394 , n243395 , n243396 , n243397 , n243398 , 
 n243399 , n243400 , n243401 , n243402 , n243403 , n243404 , n243405 , n243406 , n243407 , n243408 , 
 n243409 , n243410 , n243411 , n243412 , n243413 , n243414 , n243415 , n243416 , n243417 , n243418 , 
 n243419 , n243420 , n243421 , n243422 , n243423 , n243424 , n243425 , n243426 , n243427 , n243428 , 
 n243429 , n243430 , n243431 , n243432 , n243433 , n243434 , n243435 , n243436 , n243437 , n243438 , 
 n243439 , n243440 , n243441 , n243442 , n243443 , n243444 , n243445 , n243446 , n243447 , n243448 , 
 n243449 , n243450 , n243451 , n243452 , n243453 , n243454 , n243455 , n243456 , n243457 , n243458 , 
 n243459 , n243460 , n243461 , n243462 , n243463 , n243464 , n243465 , n243466 , n243467 , n243468 , 
 n243469 , n243470 , n243471 , n243472 , n243473 , n243474 , n243475 , n243476 , n243477 , n243478 , 
 n243479 , n243480 , n243481 , n243482 , n243483 , n243484 , n243485 , n243486 , n243487 , n243488 , 
 n243489 , n243490 , n243491 , n243492 , n243493 , n243494 , n243495 , n243496 , n243497 , n243498 , 
 n243499 , n243500 , n243501 , n243502 , n243503 , n243504 , n243505 , n243506 , n243507 , n243508 , 
 n243509 , n243510 , n243511 , n243512 , n243513 , n243514 , n243515 , n243516 , n243517 , n243518 , 
 n243519 , n243520 , n243521 , n243522 , n243523 , n243524 , n243525 , n243526 , n243527 , n243528 , 
 n243529 , n243530 , n243531 , n243532 , n243533 , n243534 , n243535 , n243536 , n243537 , n243538 , 
 n243539 , n243540 , n243541 , n243542 , n243543 , n243544 , n243545 , n243546 , n243547 , n243548 , 
 n243549 , n243550 , n243551 , n243552 , n243553 , n243554 , n243555 , n243556 , n243557 , n243558 , 
 n243559 , n243560 , n243561 , n243562 , n243563 , n243564 , n243565 , n243566 , n243567 , n243568 , 
 n243569 , n243570 , n243571 , n243572 , n243573 , n243574 , n243575 , n243576 , n243577 , n243578 , 
 n243579 , n243580 , n243581 , n243582 , n243583 , n243584 , n243585 , n243586 , n243587 , n243588 , 
 n243589 , n243590 , n243591 , n243592 , n243593 , n243594 , n243595 , n243596 , n243597 , n243598 , 
 n243599 , n243600 , n243601 , n243602 , n243603 , n243604 , n243605 , n243606 , n243607 , n243608 , 
 n243609 , n243610 , n243611 , n243612 , n243613 , n243614 , n243615 , n243616 , n243617 , n243618 , 
 n243619 , n243620 , n243621 , n243622 , n243623 , n243624 , n243625 , n243626 , n243627 , n243628 , 
 n243629 , n243630 , n243631 , n243632 , n243633 , n243634 , n243635 , n243636 , n243637 , n243638 , 
 n243639 , n243640 , n243641 , n243642 , n243643 , n243644 , n243645 , n243646 , n243647 , n243648 , 
 n243649 , n243650 , n243651 , n243652 , n243653 , n243654 , n243655 , n243656 , n243657 , n243658 , 
 n243659 , n243660 , n243661 , n243662 , n243663 , n243664 , n243665 , n243666 , n243667 , n243668 , 
 n243669 , n243670 , n243671 , n243672 , n243673 , n243674 , n243675 , n243676 , n243677 , n243678 , 
 n243679 , n243680 , n243681 , n243682 , n243683 , n243684 , n243685 , n243686 , n243687 , n243688 , 
 n243689 , n243690 , n243691 , n243692 , n243693 , n243694 , n243695 , n243696 , n243697 , n243698 , 
 n243699 , n243700 , n243701 , n243702 , n243703 , n243704 , n243705 , n243706 , n243707 , n243708 , 
 n243709 , n243710 , n243711 , n243712 , n243713 , n243714 , n243715 , n243716 , n243717 , n243718 , 
 n243719 , n243720 , n243721 , n243722 , n243723 , n243724 , n243725 , n243726 , n243727 , n243728 , 
 n243729 , n243730 , n243731 , n243732 , n243733 , n243734 , n243735 , n243736 , n243737 , n243738 , 
 n243739 , n243740 , n243741 , n243742 , n243743 , n243744 , n243745 , n243746 , n243747 , n243748 , 
 n243749 , n243750 , n243751 , n243752 , n243753 , n243754 , n243755 , n243756 , n243757 , n243758 , 
 n243759 , n243760 , n243761 , n243762 , n243763 , n243764 , n243765 , n243766 , n243767 , n243768 , 
 n243769 , n243770 , n243771 , n243772 , n243773 , n243774 , n243775 , n243776 , n243777 , n243778 , 
 n243779 , n243780 , n243781 , n243782 , n243783 , n243784 , n243785 , n243786 , n243787 , n243788 , 
 n243789 , n243790 , n243791 , n243792 , n243793 , n243794 , n243795 , n243796 , n243797 , n243798 , 
 n243799 , n243800 , n243801 , n243802 , n243803 , n243804 , n243805 , n243806 , n243807 , n243808 , 
 n243809 , n243810 , n243811 , n243812 , n243813 , n243814 , n243815 , n243816 , n243817 , n243818 , 
 n243819 , n243820 , n243821 , n243822 , n243823 , n243824 , n243825 , n243826 , n243827 , n243828 , 
 n243829 , n243830 , n243831 , n243832 , n243833 , n243834 , n243835 , n243836 , n243837 , n243838 , 
 n243839 , n243840 , n243841 , n243842 , n243843 , n243844 , n243845 , n243846 , n243847 , n243848 , 
 n243849 , n243850 , n243851 , n243852 , n243853 , n243854 , n243855 , n243856 , n243857 , n243858 , 
 n243859 , n243860 , n243861 , n243862 , n243863 , n243864 , n243865 , n243866 , n243867 , n243868 , 
 n243869 , n243870 , n243871 , n243872 , n243873 , n243874 , n243875 , n243876 , n243877 , n243878 , 
 n243879 , n243880 , n243881 , n243882 , n243883 , n243884 , n243885 , n243886 , n243887 , n243888 , 
 n243889 , n243890 , n243891 , n243892 , n243893 , n243894 , n243895 , n243896 , n243897 , n243898 , 
 n243899 , n243900 , n243901 , n243902 , n243903 , n243904 , n243905 , n243906 , n243907 , n243908 , 
 n243909 , n243910 , n243911 , n243912 , n243913 , n243914 , n243915 , n243916 , n243917 , n243918 , 
 n243919 , n243920 , n243921 , n243922 , n243923 , n243924 , n243925 , n243926 , n243927 , n243928 , 
 n243929 , n243930 , n243931 , n243932 , n243933 , n243934 , n243935 , n243936 , n243937 , n243938 , 
 n243939 , n243940 , n243941 , n243942 , n243943 , n243944 , n243945 , n243946 , n243947 , n243948 , 
 n243949 , n243950 , n243951 , n243952 , n243953 , n243954 , n243955 , n243956 , n243957 , n243958 , 
 n243959 , n243960 , n243961 , n243962 , n243963 , n243964 , n243965 , n243966 , n243967 , n243968 , 
 n243969 , n243970 , n243971 , n243972 , n243973 , n243974 , n243975 , n243976 , n243977 , n243978 , 
 n243979 , n243980 , n243981 , n243982 , n243983 , n243984 , n243985 , n243986 , n243987 , n243988 , 
 n243989 , n243990 , n243991 , n243992 , n243993 , n243994 , n243995 , n243996 , n243997 , n243998 , 
 n243999 , n244000 , n244001 , n244002 , n244003 , n244004 , n244005 , n244006 , n244007 , n244008 , 
 n244009 , n244010 , n244011 , n244012 , n244013 , n244014 , n244015 , n244016 , n244017 , n244018 , 
 n244019 , n244020 , n244021 , n244022 , n244023 , n244024 , n244025 , n244026 , n244027 , n244028 , 
 n244029 , n244030 , n244031 , n244032 , n244033 , n244034 , n244035 , n244036 , n244037 , n244038 , 
 n244039 , n244040 , n244041 , n244042 , n244043 , n244044 , n244045 , n244046 , n244047 , n244048 , 
 n244049 , n244050 , n244051 , n244052 , n244053 , n244054 , n244055 , n244056 , n244057 , n244058 , 
 n244059 , n244060 , n244061 , n244062 , n244063 , n244064 , n244065 , n244066 , n244067 , n244068 , 
 n244069 , n244070 , n244071 , n244072 , n244073 , n244074 , n244075 , n244076 , n244077 , n244078 , 
 n244079 , n244080 , n244081 , n244082 , n244083 , n244084 , n244085 , n244086 , n244087 , n244088 , 
 n244089 , n244090 , n244091 , n244092 , n244093 , n244094 , n244095 , n244096 , n244097 , n244098 , 
 n244099 , n244100 , n244101 , n244102 , n244103 , n244104 , n244105 , n244106 , n244107 , n244108 , 
 n244109 , n244110 , n244111 , n244112 , n244113 , n244114 , n244115 , n244116 , n244117 , n244118 , 
 n244119 , n244120 , n244121 , n244122 , n244123 , n244124 , n244125 , n244126 , n244127 , n244128 , 
 n244129 , n244130 , n244131 , n244132 , n244133 , n244134 , n244135 , n244136 , n244137 , n244138 , 
 n244139 , n244140 , n244141 , n244142 , n244143 , n244144 , n244145 , n244146 , n244147 , n244148 , 
 n244149 , n244150 , n244151 , n244152 , n244153 , n244154 , n244155 , n244156 , n244157 , n244158 , 
 n244159 , n244160 , n244161 , n244162 , n244163 , n244164 , n244165 , n244166 , n244167 , n244168 , 
 n244169 , n244170 , n244171 , n244172 , n244173 , n244174 , n244175 , n244176 , n244177 , n244178 , 
 n244179 , n244180 , n244181 , n244182 , n244183 , n244184 , n244185 , n244186 , n244187 , n244188 , 
 n244189 , n244190 , n244191 , n244192 , n244193 , n244194 , n244195 , n244196 , n244197 , n244198 , 
 n244199 , n244200 , n244201 , n244202 , n244203 , n244204 , n244205 , n244206 , n244207 , n244208 , 
 n244209 , n244210 , n244211 , n244212 , n244213 , n244214 , n244215 , n244216 , n244217 , n244218 , 
 n244219 , n244220 , n244221 , n244222 , n244223 , n244224 , n244225 , n244226 , n244227 , n244228 , 
 n244229 , n244230 , n244231 , n244232 , n244233 , n244234 , n244235 , n244236 , n244237 , n244238 , 
 n244239 , n244240 , n244241 , n244242 , n244243 , n244244 , n244245 , n244246 , n244247 , n244248 , 
 n244249 , n244250 , n244251 , n244252 , n244253 , n244254 , n244255 , n244256 , n244257 , n244258 , 
 n244259 , n244260 , n244261 , n244262 , n244263 , n244264 , n244265 , n244266 , n244267 , n244268 , 
 n244269 , n244270 , n244271 , n244272 , n244273 , n244274 , n244275 , n244276 , n244277 , n244278 , 
 n244279 , n244280 , n244281 , n244282 , n244283 , n244284 , n244285 , n244286 , n244287 , n244288 , 
 n244289 , n244290 , n244291 , n244292 , n244293 , n244294 , n244295 , n244296 , n244297 , n244298 , 
 n244299 , n244300 , n244301 , n244302 , n244303 , n244304 , n244305 , n244306 , n244307 , n244308 , 
 n244309 , n244310 , n244311 , n244312 , n244313 , n244314 , n244315 , n244316 , n244317 , n244318 , 
 n244319 , n244320 , n244321 , n244322 , n244323 , n244324 , n244325 , n244326 , n244327 , n244328 , 
 n244329 , n244330 , n244331 , n244332 , n244333 , n244334 , n244335 , n244336 , n244337 , n244338 , 
 n244339 , n244340 , n244341 , n244342 , n244343 , n244344 , n244345 , n244346 , n244347 , n244348 , 
 n244349 , n244350 , n244351 , n244352 , n244353 , n244354 , n244355 , n244356 , n244357 , n244358 , 
 n244359 , n244360 , n244361 , n244362 , n244363 , n244364 , n244365 , n244366 , n244367 , n244368 , 
 n244369 , n244370 , n244371 , n244372 , n244373 , n244374 , n244375 , n244376 , n244377 , n244378 , 
 n244379 , n244380 , n244381 , n244382 , n244383 , n244384 , n244385 , n244386 , n244387 , n244388 , 
 n244389 , n244390 , n244391 , n244392 , n244393 , n244394 , n244395 , n244396 , n244397 , n244398 , 
 n244399 , n244400 , n244401 , n244402 , n244403 , n244404 , n244405 , n244406 , n244407 , n244408 , 
 n244409 , n244410 , n244411 , n244412 , n244413 , n244414 , n244415 , n244416 , n244417 , n244418 , 
 n244419 , n244420 , n244421 , n244422 , n244423 , n244424 , n244425 , n244426 , n244427 , n244428 , 
 n244429 , n244430 , n244431 , n244432 , n244433 , n244434 , n244435 , n244436 , n244437 , n244438 , 
 n244439 , n244440 , n244441 , n244442 , n244443 , n244444 , n244445 , n244446 , n244447 , n244448 , 
 n244449 , n244450 , n244451 , n244452 , n244453 , n244454 , n244455 , n244456 , n244457 , n244458 , 
 n244459 , n244460 , n244461 , n244462 , n244463 , n244464 , n244465 , n244466 , n244467 , n244468 , 
 n244469 , n244470 , n244471 , n244472 , n244473 , n244474 , n244475 , n244476 , n244477 , n244478 , 
 n244479 , n244480 , n244481 , n244482 , n244483 , n244484 , n244485 , n244486 , n244487 , n244488 , 
 n244489 , n244490 , n244491 , n244492 , n244493 , n244494 , n244495 , n244496 , n244497 , n244498 , 
 n244499 , n244500 , n244501 , n244502 , n244503 , n244504 , n244505 , n244506 , n244507 , n244508 , 
 n244509 , n244510 , n244511 , n244512 , n244513 , n244514 , n244515 , n244516 , n244517 , n244518 , 
 n244519 , n244520 , n244521 , n244522 , n244523 , n244524 , n244525 , n244526 , n244527 , n244528 , 
 n244529 , n244530 , n244531 , n244532 , n244533 , n244534 , n244535 , n244536 , n244537 , n244538 , 
 n244539 , n244540 , n244541 , n244542 , n244543 , n244544 , n244545 , n244546 , n244547 , n244548 , 
 n244549 , n244550 , n244551 , n244552 , n244553 , n244554 , n244555 , n244556 , n244557 , n244558 , 
 n244559 , n244560 , n244561 , n244562 , n244563 , n244564 , n244565 , n244566 , n244567 , n244568 , 
 n244569 , n244570 , n244571 , n244572 , n244573 , n244574 , n244575 , n244576 , n244577 , n244578 , 
 n244579 , n244580 , n244581 , n244582 , n244583 , n244584 , n244585 , n244586 , n244587 , n244588 , 
 n244589 , n244590 , n244591 , n244592 , n244593 , n244594 , n244595 , n244596 , n244597 , n244598 , 
 n244599 , n244600 , n244601 , n244602 , n244603 , n244604 , n244605 , n244606 , n244607 , n244608 , 
 n244609 , n244610 , n244611 , n244612 , n244613 , n244614 , n244615 , n244616 , n244617 , n244618 , 
 n244619 , n244620 , n244621 , n244622 , n244623 , n244624 , n244625 , n244626 , n244627 , n244628 , 
 n244629 , n244630 , n244631 , n244632 , n244633 , n244634 , n244635 , n244636 , n244637 , n244638 , 
 n244639 , n244640 , n244641 , n244642 , n244643 , n244644 , n244645 , n244646 , n244647 , n244648 , 
 n244649 , n244650 , n244651 , n244652 , n244653 , n244654 , n244655 , n244656 , n244657 , n244658 , 
 n244659 , n244660 , n244661 , n244662 , n244663 , n244664 , n244665 , n244666 , n244667 , n244668 , 
 n244669 , n244670 , n244671 , n244672 , n244673 , n244674 , n244675 , n244676 , n244677 , n244678 , 
 n244679 , n244680 , n244681 , n244682 , n244683 , n244684 , n244685 , n244686 , n244687 , n244688 , 
 n244689 , n244690 , n244691 , n244692 , n244693 , n244694 , n244695 , n244696 , n244697 , n244698 , 
 n244699 , n244700 , n244701 , n244702 , n244703 , n244704 , n244705 , n244706 , n244707 , n244708 , 
 n244709 , n244710 , n244711 , n244712 , n244713 , n244714 , n244715 , n244716 , n244717 , n244718 , 
 n244719 , n244720 , n244721 , n244722 , n244723 , n244724 , n244725 , n244726 , n244727 , n244728 , 
 n244729 , n244730 , n244731 , n244732 , n244733 , n244734 , n244735 , n244736 , n244737 , n244738 , 
 n244739 , n244740 , n244741 , n244742 , n244743 , n244744 , n244745 , n244746 , n244747 , n244748 , 
 n244749 , n244750 , n244751 , n244752 , n244753 , n244754 , n244755 , n244756 , n244757 , n244758 , 
 n244759 , n244760 , n244761 , n244762 , n244763 , n244764 , n244765 , n244766 , n244767 , n244768 , 
 n244769 , n244770 , n244771 , n244772 , n244773 , n244774 , n244775 , n244776 , n244777 , n244778 , 
 n244779 , n244780 , n244781 , n244782 , n244783 , n244784 , n244785 , n244786 , n244787 , n244788 , 
 n244789 , n244790 , n244791 , n244792 , n244793 , n244794 , n244795 , n244796 , n244797 , n244798 , 
 n244799 , n244800 , n244801 , n244802 , n244803 , n244804 , n244805 , n244806 , n244807 , n244808 , 
 n244809 , n244810 , n244811 , n244812 , n244813 , n244814 , n244815 , n244816 , n244817 , n244818 , 
 n244819 , n244820 , n244821 , n244822 , n244823 , n244824 , n244825 , n244826 , n244827 , n244828 , 
 n244829 , n244830 , n244831 , n244832 , n244833 , n244834 , n244835 , n244836 , n244837 , n244838 , 
 n244839 , n244840 , n244841 , n244842 , n244843 , n244844 , n244845 , n244846 , n244847 , n244848 , 
 n244849 , n244850 , n244851 , n244852 , n244853 , n244854 , n244855 , n244856 , n244857 , n244858 , 
 n244859 , n244860 , n244861 , n244862 , n244863 , n244864 , n244865 , n244866 , n244867 , n244868 , 
 n244869 , n244870 , n244871 , n244872 , n244873 , n244874 , n244875 , n244876 , n244877 , n244878 , 
 n244879 , n244880 , n244881 , n244882 , n244883 , n244884 , n244885 , n244886 , n244887 , n244888 , 
 n244889 , n244890 , n244891 , n244892 , n244893 , n244894 , n244895 , n244896 , n244897 , n244898 , 
 n244899 , n244900 , n244901 , n244902 , n244903 , n244904 , n244905 , n244906 , n244907 , n244908 , 
 n244909 , n244910 , n244911 , n244912 , n244913 , n244914 , n244915 , n244916 , n244917 , n244918 , 
 n244919 , n244920 , n244921 , n244922 , n244923 , n244924 , n244925 , n244926 , n244927 , n244928 , 
 n244929 , n244930 , n244931 , n244932 , n244933 , n244934 , n244935 , n244936 , n244937 , n244938 , 
 n244939 , n244940 , n244941 , n244942 , n244943 , n244944 , n244945 , n244946 , n244947 , n244948 , 
 n244949 , n244950 , n244951 , n244952 , n244953 , n244954 , n244955 , n244956 , n244957 , n244958 , 
 n244959 , n244960 , n244961 , n244962 , n244963 , n244964 , n244965 , n244966 , n244967 , n244968 , 
 n244969 , n244970 , n244971 , n244972 , n244973 , n244974 , n244975 , n244976 , n244977 , n244978 , 
 n244979 , n244980 , n244981 , n244982 , n244983 , n244984 , n244985 , n244986 , n244987 , n244988 , 
 n244989 , n244990 , n244991 , n244992 , n244993 , n244994 , n244995 , n244996 , n244997 , n244998 , 
 n244999 , n245000 , n245001 , n245002 , n245003 , n245004 , n245005 , n245006 , n245007 , n245008 , 
 n245009 , n245010 , n245011 , n245012 , n245013 , n245014 , n245015 , n245016 , n245017 , n245018 , 
 n245019 , n245020 , n245021 , n245022 , n245023 , n245024 , n245025 , n245026 , n245027 , n245028 , 
 n245029 , n245030 , n245031 , n245032 , n245033 , n245034 , n245035 , n245036 , n245037 , n245038 , 
 n245039 , n245040 , n245041 , n245042 , n245043 , n245044 , n245045 , n245046 , n245047 , n245048 , 
 n245049 , n245050 , n245051 , n245052 , n245053 , n245054 , n245055 , n245056 , n245057 , n245058 , 
 n245059 , n245060 , n245061 , n245062 , n245063 , n245064 , n245065 , n245066 , n245067 , n245068 , 
 n245069 , n245070 , n245071 , n245072 , n245073 , n245074 , n245075 , n245076 , n245077 , n245078 , 
 n245079 , n245080 , n245081 , n245082 , n245083 , n245084 , n245085 , n245086 , n245087 , n245088 , 
 n245089 , n245090 , n245091 , n245092 , n245093 , n245094 , n245095 , n245096 , n245097 , n245098 , 
 n245099 , n245100 , n245101 , n245102 , n245103 , n245104 , n245105 , n245106 , n245107 , n245108 , 
 n245109 , n245110 , n245111 , n245112 , n245113 , n245114 , n245115 , n245116 , n245117 , n245118 , 
 n245119 , n245120 , n245121 , n245122 , n245123 , n245124 , n245125 , n245126 , n245127 , n245128 , 
 n245129 , n245130 , n245131 , n245132 , n245133 , n245134 , n245135 , n245136 , n245137 , n245138 , 
 n245139 , n245140 , n245141 , n245142 , n245143 , n245144 , n245145 , n245146 , n245147 , n245148 , 
 n245149 , n245150 , n245151 , n245152 , n245153 , n245154 , n245155 , n245156 , n245157 , n245158 , 
 n245159 , n245160 , n245161 , n245162 , n245163 , n245164 , n245165 , n245166 , n245167 , n245168 , 
 n245169 , n245170 , n245171 , n245172 , n245173 , n245174 , n245175 , n245176 , n245177 , n245178 , 
 n245179 , n245180 , n245181 , n245182 , n245183 , n245184 , n245185 , n245186 , n245187 , n245188 , 
 n245189 , n245190 , n245191 , n245192 , n245193 , n245194 , n245195 , n245196 , n245197 , n245198 , 
 n245199 , n245200 , n245201 , n245202 , n245203 , n245204 , n245205 , n245206 , n245207 , n245208 , 
 n245209 , n245210 , n245211 , n245212 , n245213 , n245214 , n245215 , n245216 , n245217 , n245218 , 
 n245219 , n245220 , n245221 , n245222 , n245223 , n245224 , n245225 , n245226 , n245227 , n245228 , 
 n245229 , n245230 , n245231 , n245232 , n245233 , n245234 , n245235 , n245236 , n245237 , n245238 , 
 n245239 , n245240 , n245241 , n245242 , n245243 , n245244 , n245245 , n245246 , n245247 , n245248 , 
 n245249 , n245250 , n245251 , n245252 , n245253 , n245254 , n245255 , n245256 , n245257 , n245258 , 
 n245259 , n245260 , n245261 , n245262 , n245263 , n245264 , n245265 , n245266 , n245267 , n245268 , 
 n245269 , n245270 , n245271 , n245272 , n245273 , n245274 , n245275 , n245276 , n245277 , n245278 , 
 n245279 , n245280 , n245281 , n245282 , n245283 , n245284 , n245285 , n245286 , n245287 , n245288 , 
 n245289 , n245290 , n245291 , n245292 , n245293 , n245294 , n245295 , n245296 , n245297 , n245298 , 
 n245299 , n245300 , n245301 , n245302 , n245303 , n245304 , n245305 , n245306 , n245307 , n245308 , 
 n245309 , n245310 , n245311 , n245312 , n245313 , n245314 , n245315 , n245316 , n245317 , n245318 , 
 n245319 , n245320 , n245321 , n245322 , n245323 , n245324 , n245325 , n245326 , n245327 , n245328 , 
 n245329 , n245330 , n245331 , n245332 , n245333 , n245334 , n245335 , n245336 , n245337 , n245338 , 
 n245339 , n245340 , n245341 , n245342 , n245343 , n245344 , n245345 , n245346 , n245347 , n245348 , 
 n245349 , n245350 , n245351 , n245352 , n245353 , n245354 , n245355 , n245356 , n245357 , n245358 , 
 n245359 , n245360 , n245361 , n245362 , n245363 , n245364 , n245365 , n245366 , n245367 , n245368 , 
 n245369 , n245370 , n245371 , n245372 , n245373 , n245374 , n245375 , n245376 , n245377 , n245378 , 
 n245379 , n245380 , n245381 , n245382 , n245383 , n245384 , n245385 , n245386 , n245387 , n245388 , 
 n245389 , n245390 , n245391 , n245392 , n245393 , n245394 , n245395 , n245396 , n245397 , n245398 , 
 n245399 , n245400 , n245401 , n245402 , n245403 , n245404 , n245405 , n245406 , n245407 , n245408 , 
 n245409 , n245410 , n245411 , n245412 , n245413 , n245414 , n245415 , n245416 , n245417 , n245418 , 
 n245419 , n245420 , n245421 , n245422 , n245423 , n245424 , n245425 , n245426 , n245427 , n245428 , 
 n245429 , n245430 , n245431 , n245432 , n245433 , n245434 , n245435 , n245436 , n245437 , n245438 , 
 n245439 , n245440 , n245441 , n245442 , n245443 , n245444 , n245445 , n245446 , n245447 , n245448 , 
 n245449 , n245450 , n245451 , n245452 , n245453 , n245454 , n245455 , n245456 , n245457 , n245458 , 
 n245459 , n245460 , n245461 , n245462 , n245463 , n245464 , n245465 , n245466 , n245467 , n245468 , 
 n245469 , n245470 , n245471 , n245472 , n245473 , n245474 , n245475 , n245476 , n245477 , n245478 , 
 n245479 , n245480 , n245481 , n245482 , n245483 , n245484 , n245485 , n245486 , n245487 , n245488 , 
 n245489 , n245490 , n245491 , n245492 , n245493 , n245494 , n245495 , n245496 , n245497 , n245498 , 
 n245499 , n245500 , n245501 , n245502 , n245503 , n245504 , n245505 , n245506 , n245507 , n245508 , 
 n245509 , n245510 , n245511 , n245512 , n245513 , n245514 , n245515 , n245516 , n245517 , n245518 , 
 n245519 , n245520 , n245521 , n245522 , n245523 , n245524 , n245525 , n245526 , n245527 , n245528 , 
 n245529 , n245530 , n245531 , n245532 , n245533 , n245534 , n245535 , n245536 , n245537 , n245538 , 
 n245539 , n245540 , n245541 , n245542 , n245543 , n245544 , n245545 , n245546 , n245547 , n245548 , 
 n245549 , n245550 , n245551 , n245552 , n245553 , n245554 , n245555 , n245556 , n245557 , n245558 , 
 n245559 , n245560 , n245561 , n245562 , n245563 , n245564 , n245565 , n245566 , n245567 , n245568 , 
 n245569 , n245570 , n245571 , n245572 , n245573 , n245574 , n245575 , n245576 , n245577 , n245578 , 
 n245579 , n245580 , n245581 , n245582 , n245583 , n245584 , n245585 , n245586 , n245587 , n245588 , 
 n245589 , n245590 , n245591 , n245592 , n245593 , n245594 , n245595 , n245596 , n245597 , n245598 , 
 n245599 , n245600 , n245601 , n245602 , n245603 , n245604 , n245605 , n245606 , n245607 , n245608 , 
 n245609 , n245610 , n245611 , n245612 , n245613 , n245614 , n245615 , n245616 , n245617 , n245618 , 
 n245619 , n245620 , n245621 , n245622 , n245623 , n245624 , n245625 , n245626 , n245627 , n245628 , 
 n245629 , n245630 , n245631 , n245632 , n245633 , n245634 , n245635 , n245636 , n245637 , n245638 , 
 n245639 , n245640 , n245641 , n245642 , n245643 , n245644 , n245645 , n245646 , n245647 , n245648 , 
 n245649 , n245650 , n245651 , n245652 , n245653 , n245654 , n245655 , n245656 , n245657 , n245658 , 
 n245659 , n245660 , n245661 , n245662 , n245663 , n245664 , n245665 , n245666 , n245667 , n245668 , 
 n245669 , n245670 , n245671 , n245672 , n245673 , n245674 , n245675 , n245676 , n245677 , n245678 , 
 n245679 , n245680 , n245681 , n245682 , n245683 , n245684 , n245685 , n245686 , n245687 , n245688 , 
 n245689 , n245690 , n245691 , n245692 , n245693 , n245694 , n245695 , n245696 , n245697 , n245698 , 
 n245699 , n245700 , n245701 , n245702 , n245703 , n245704 , n245705 , n245706 , n245707 , n245708 , 
 n245709 , n245710 , n245711 , n245712 , n245713 , n245714 , n245715 , n245716 , n245717 , n245718 , 
 n245719 , n245720 , n245721 , n245722 , n245723 , n245724 , n245725 , n245726 , n245727 , n245728 , 
 n245729 , n245730 , n245731 , n245732 , n245733 , n245734 , n245735 , n245736 , n245737 , n245738 , 
 n245739 , n245740 , n245741 , n245742 , n245743 , n245744 , n245745 , n245746 , n245747 , n245748 , 
 n245749 , n245750 , n245751 , n245752 , n245753 , n245754 , n245755 , n245756 , n245757 , n245758 , 
 n245759 , n245760 , n245761 , n245762 , n245763 , n245764 , n245765 , n245766 , n245767 , n245768 , 
 n245769 , n245770 , n245771 , n245772 , n245773 , n245774 , n245775 , n245776 , n245777 , n245778 , 
 n245779 , n245780 , n245781 , n245782 , n245783 , n245784 , n245785 , n245786 , n245787 , n245788 , 
 n245789 , n245790 , n245791 , n245792 , n245793 , n245794 , n245795 , n245796 , n245797 , n245798 , 
 n245799 , n245800 , n245801 , n245802 , n245803 , n245804 , n245805 , n245806 , n245807 , n245808 , 
 n245809 , n245810 , n245811 , n245812 , n245813 , n245814 , n245815 , n245816 , n245817 , n245818 , 
 n245819 , n245820 , n245821 , n245822 , n245823 , n245824 , n245825 , n245826 , n245827 , n245828 , 
 n245829 , n245830 , n245831 , n245832 , n245833 , n245834 , n245835 , n245836 , n245837 , n245838 , 
 n245839 , n245840 , n245841 , n245842 , n245843 , n245844 , n245845 , n245846 , n245847 , n245848 , 
 n245849 , n245850 , n245851 , n245852 , n245853 , n245854 , n245855 , n245856 , n245857 , n245858 , 
 n245859 , n245860 , n245861 , n245862 , n245863 , n245864 , n245865 , n245866 , n245867 , n245868 , 
 n245869 , n245870 , n245871 , n245872 , n245873 , n245874 , n245875 , n245876 , n245877 , n245878 , 
 n245879 , n245880 , n245881 , n245882 , n245883 , n245884 , n245885 , n245886 , n245887 , n245888 , 
 n245889 , n245890 , n245891 , n245892 , n245893 , n245894 , n245895 , n245896 , n245897 , n245898 , 
 n245899 , n245900 , n245901 , n245902 , n245903 , n245904 , n245905 , n245906 , n245907 , n245908 , 
 n245909 , n245910 , n245911 , n245912 , n245913 , n245914 , n245915 , n245916 , n245917 , n245918 , 
 n245919 , n245920 , n245921 , n245922 , n245923 , n245924 , n245925 , n245926 , n245927 , n245928 , 
 n245929 , n245930 , n245931 , n245932 , n245933 , n245934 , n245935 , n245936 , n245937 , n245938 , 
 n245939 , n245940 , n245941 , n245942 , n245943 , n245944 , n245945 , n245946 , n245947 , n245948 , 
 n245949 , n245950 , n245951 , n245952 , n245953 , n245954 , n245955 , n245956 , n245957 , n245958 , 
 n245959 , n245960 , n245961 , n245962 , n245963 , n245964 , n245965 , n245966 , n245967 , n245968 , 
 n245969 , n245970 , n245971 , n245972 , n245973 , n245974 , n245975 , n245976 , n245977 , n245978 , 
 n245979 , n245980 , n245981 , n245982 , n245983 , n245984 , n245985 , n245986 , n245987 , n245988 , 
 n245989 , n245990 , n245991 , n245992 , n245993 , n245994 , n245995 , n245996 , n245997 , n245998 , 
 n245999 , n246000 , n246001 , n246002 , n246003 , n246004 , n246005 , n246006 , n246007 , n246008 , 
 n246009 , n246010 , n246011 , n246012 , n246013 , n246014 , n246015 , n246016 , n246017 , n246018 , 
 n246019 , n246020 , n246021 , n246022 , n246023 , n246024 , n246025 , n246026 , n246027 , n246028 , 
 n246029 , n246030 , n246031 , n246032 , n246033 , n246034 , n246035 , n246036 , n246037 , n246038 , 
 n246039 , n246040 , n246041 , n246042 , n246043 , n246044 , n246045 , n246046 , n246047 , n246048 , 
 n246049 , n246050 , n246051 , n246052 , n246053 , n246054 , n246055 , n246056 , n246057 , n246058 , 
 n246059 , n246060 , n246061 , n246062 , n246063 , n246064 , n246065 , n246066 , n246067 , n246068 , 
 n246069 , n246070 , n246071 , n246072 , n246073 , n246074 , n246075 , n246076 , n246077 , n246078 , 
 n246079 , n246080 , n246081 , n246082 , n246083 , n246084 , n246085 , n246086 , n246087 , n246088 , 
 n246089 , n246090 , n246091 , n246092 , n246093 , n246094 , n246095 , n246096 , n246097 , n246098 , 
 n246099 , n246100 , n246101 , n246102 , n246103 , n246104 , n246105 , n246106 , n246107 , n246108 , 
 n246109 , n246110 , n246111 , n246112 , n246113 , n246114 , n246115 , n246116 , n246117 , n246118 , 
 n246119 , n246120 , n246121 , n246122 , n246123 , n246124 , n246125 , n246126 , n246127 , n246128 , 
 n246129 , n246130 , n246131 , n246132 , n246133 , n246134 , n246135 , n246136 , n246137 , n246138 , 
 n246139 , n246140 , n246141 , n246142 , n246143 , n246144 , n246145 , n246146 , n246147 , n246148 , 
 n246149 , n246150 , n246151 , n246152 , n246153 , n246154 , n246155 , n246156 , n246157 , n246158 , 
 n246159 , n246160 , n246161 , n246162 , n246163 , n246164 , n246165 , n246166 , n246167 , n246168 , 
 n246169 , n246170 , n246171 , n246172 , n246173 , n246174 , n246175 , n246176 , n246177 , n246178 , 
 n246179 , n246180 , n246181 , n246182 , n246183 , n246184 , n246185 , n246186 , n246187 , n246188 , 
 n246189 , n246190 , n246191 , n246192 , n246193 , n246194 , n246195 , n246196 , n246197 , n246198 , 
 n246199 , n246200 , n246201 , n246202 , n246203 , n246204 , n246205 , n246206 , n246207 , n246208 , 
 n246209 , n246210 , n246211 , n246212 , n246213 , n246214 , n246215 , n246216 , n246217 , n246218 , 
 n246219 , n246220 , n246221 , n246222 , n246223 , n246224 , n246225 , n246226 , n246227 , n246228 , 
 n246229 , n246230 , n246231 , n246232 , n246233 , n246234 , n246235 , n246236 , n246237 , n246238 , 
 n246239 , n246240 , n246241 , n246242 , n246243 , n246244 , n246245 , n246246 , n246247 , n246248 , 
 n246249 , n246250 , n246251 , n246252 , n246253 , n246254 , n246255 , n246256 , n246257 , n246258 , 
 n246259 , n246260 , n246261 , n246262 , n246263 , n246264 , n246265 , n246266 , n246267 , n246268 , 
 n246269 , n246270 , n246271 , n246272 , n246273 , n246274 , n246275 , n246276 , n246277 , n246278 , 
 n246279 , n246280 , n246281 , n246282 , n246283 , n246284 , n246285 , n246286 , n246287 , n246288 , 
 n246289 , n246290 , n246291 , n246292 , n246293 , n246294 , n246295 , n246296 , n246297 , n246298 , 
 n246299 , n246300 , n246301 , n246302 , n246303 , n246304 , n246305 , n246306 , n246307 , n246308 , 
 n246309 , n246310 , n246311 , n246312 , n246313 , n246314 , n246315 , n246316 , n246317 , n246318 , 
 n246319 , n246320 , n246321 , n246322 , n246323 , n246324 , n246325 , n246326 , n246327 , n246328 , 
 n246329 , n246330 , n246331 , n246332 , n246333 , n246334 , n246335 , n246336 , n246337 , n246338 , 
 n246339 , n246340 , n246341 , n246342 , n246343 , n246344 , n246345 , n246346 , n246347 , n246348 , 
 n246349 , n246350 , n246351 , n246352 , n246353 , n246354 , n246355 , n246356 , n246357 , n246358 , 
 n246359 , n246360 , n246361 , n246362 , n246363 , n246364 , n246365 , n246366 , n246367 , n246368 , 
 n246369 , n246370 , n246371 , n246372 , n246373 , n246374 , n246375 , n246376 , n246377 , n246378 , 
 n246379 , n246380 , n246381 , n246382 , n246383 , n246384 , n246385 , n246386 , n246387 , n246388 , 
 n246389 , n246390 , n246391 , n246392 , n246393 , n246394 , n246395 , n246396 , n246397 , n246398 , 
 n246399 , n246400 , n246401 , n246402 , n246403 , n246404 , n246405 , n246406 , n246407 , n246408 , 
 n246409 , n246410 , n246411 , n246412 , n246413 , n246414 , n246415 , n246416 , n246417 , n246418 , 
 n246419 , n246420 , n246421 , n246422 , n246423 , n246424 , n246425 , n246426 , n246427 , n246428 , 
 n246429 , n246430 , n246431 , n246432 , n246433 , n246434 , n246435 , n246436 , n246437 , n246438 , 
 n246439 , n246440 , n246441 , n246442 , n246443 , n246444 , n246445 , n246446 , n246447 , n246448 , 
 n246449 , n246450 , n246451 , n246452 , n246453 , n246454 , n246455 , n246456 , n246457 , n246458 , 
 n246459 , n246460 , n246461 , n246462 , n246463 , n246464 , n246465 , n246466 , n246467 , n246468 , 
 n246469 , n246470 , n246471 , n246472 , n246473 , n246474 , n246475 , n246476 , n246477 , n246478 , 
 n246479 , n246480 , n246481 , n246482 , n246483 , n246484 , n246485 , n246486 , n246487 , n246488 , 
 n246489 , n246490 , n246491 , n246492 , n246493 , n246494 , n246495 , n246496 , n246497 , n246498 , 
 n246499 , n246500 , n246501 , n246502 , n246503 , n246504 , n246505 , n246506 , n246507 , n246508 , 
 n246509 , n246510 , n246511 , n246512 , n246513 , n246514 , n246515 , n246516 , n246517 , n246518 , 
 n246519 , n246520 , n246521 , n246522 , n246523 , n246524 , n246525 , n246526 , n246527 , n246528 , 
 n246529 , n246530 , n246531 , n246532 , n246533 , n246534 , n246535 , n246536 , n246537 , n246538 , 
 n246539 , n246540 , n246541 , n246542 , n246543 , n246544 , n246545 , n246546 , n246547 , n246548 , 
 n246549 , n246550 , n246551 , n246552 , n246553 , n246554 , n246555 , n246556 , n246557 , n246558 , 
 n246559 , n246560 , n246561 , n246562 , n246563 , n246564 , n246565 , n246566 , n246567 , n246568 , 
 n246569 , n246570 , n246571 , n246572 , n246573 , n246574 , n246575 , n246576 , n246577 , n246578 , 
 n246579 , n246580 , n246581 , n246582 , n246583 , n246584 , n246585 , n246586 , n246587 , n246588 , 
 n246589 , n246590 , n246591 , n246592 , n246593 , n246594 , n246595 , n246596 , n246597 , n246598 , 
 n246599 , n246600 , n246601 , n246602 , n246603 , n246604 , n246605 , n246606 , n246607 , n246608 , 
 n246609 , n246610 , n246611 , n246612 , n246613 , n246614 , n246615 , n246616 , n246617 , n246618 , 
 n246619 , n246620 , n246621 , n246622 , n246623 , n246624 , n246625 , n246626 , n246627 , n246628 , 
 n246629 , n246630 , n246631 , n246632 , n246633 , n246634 , n246635 , n246636 , n246637 , n246638 , 
 n246639 , n246640 , n246641 , n246642 , n246643 , n246644 , n246645 , n246646 , n246647 , n246648 , 
 n246649 , n246650 , n246651 , n246652 , n246653 , n246654 , n246655 , n246656 , n246657 , n246658 , 
 n246659 , n246660 , n246661 , n246662 , n246663 , n246664 , n246665 , n246666 , n246667 , n246668 , 
 n246669 , n246670 , n246671 , n246672 , n246673 , n246674 , n246675 , n246676 , n246677 , n246678 , 
 n246679 , n246680 , n246681 , n246682 , n246683 , n246684 , n246685 , n246686 , n246687 , n246688 , 
 n246689 , n246690 , n246691 , n246692 , n246693 , n246694 , n246695 , n246696 , n246697 , n246698 , 
 n246699 , n246700 , n246701 , n246702 , n246703 , n246704 , n246705 , n246706 , n246707 , n246708 , 
 n246709 , n246710 , n246711 , n246712 , n246713 , n246714 , n246715 , n246716 , n246717 , n246718 , 
 n246719 , n246720 , n246721 , n246722 , n246723 , n246724 , n246725 , n246726 , n246727 , n246728 , 
 n246729 , n246730 , n246731 , n246732 , n246733 , n246734 , n246735 , n246736 , n246737 , n246738 , 
 n246739 , n246740 , n246741 , n246742 , n246743 , n246744 , n246745 , n246746 , n246747 , n246748 , 
 n246749 , n246750 , n246751 , n246752 , n246753 , n246754 , n246755 , n246756 , n246757 , n246758 , 
 n246759 , n246760 , n246761 , n246762 , n246763 , n246764 , n246765 , n246766 , n246767 , n246768 , 
 n246769 , n246770 , n246771 , n246772 , n246773 , n246774 , n246775 , n246776 , n246777 , n246778 , 
 n246779 , n246780 , n246781 , n246782 , n246783 , n246784 , n246785 , n246786 , n246787 , n246788 , 
 n246789 , n246790 , n246791 , n246792 , n246793 , n246794 , n246795 , n246796 , n246797 , n246798 , 
 n246799 , n246800 , n246801 , n246802 , n246803 , n246804 , n246805 , n246806 , n246807 , n246808 , 
 n246809 , n246810 , n246811 , n246812 , n246813 , n246814 , n246815 , n246816 , n246817 , n246818 , 
 n246819 , n246820 , n246821 , n246822 , n246823 , n246824 , n246825 , n246826 , n246827 , n246828 , 
 n246829 , n246830 , n246831 , n246832 , n246833 , n246834 , n246835 , n246836 , n246837 , n246838 , 
 n246839 , n246840 , n246841 , n246842 , n246843 , n246844 , n246845 , n246846 , n246847 , n246848 , 
 n246849 , n246850 , n246851 , n246852 , n246853 , n246854 , n246855 , n246856 , n246857 , n246858 , 
 n246859 , n246860 , n246861 , n246862 , n246863 , n246864 , n246865 , n246866 , n246867 , n246868 , 
 n246869 , n246870 , n246871 , n246872 , n246873 , n246874 , n246875 , n246876 , n246877 , n246878 , 
 n246879 , n246880 , n246881 , n246882 , n246883 , n246884 , n246885 , n246886 , n246887 , n246888 , 
 n246889 , n246890 , n246891 , n246892 , n246893 , n246894 , n246895 , n246896 , n246897 , n246898 , 
 n246899 , n246900 , n246901 , n246902 , n246903 , n246904 , n246905 , n246906 , n246907 , n246908 , 
 n246909 , n246910 , n246911 , n246912 , n246913 , n246914 , n246915 , n246916 , n246917 , n246918 , 
 n246919 , n246920 , n246921 , n246922 , n246923 , n246924 , n246925 , n246926 , n246927 , n246928 , 
 n246929 , n246930 , n246931 , n246932 , n246933 , n246934 , n246935 , n246936 , n246937 , n246938 , 
 n246939 , n246940 , n246941 , n246942 , n246943 , n246944 , n246945 , n246946 , n246947 , n246948 , 
 n246949 , n246950 , n246951 , n246952 , n246953 , n246954 , n246955 , n246956 , n246957 , n246958 , 
 n246959 , n246960 , n246961 , n246962 , n246963 , n246964 , n246965 , n246966 , n246967 , n246968 , 
 n246969 , n246970 , n246971 , n246972 , n246973 , n246974 , n246975 , n246976 , n246977 , n246978 , 
 n246979 , n246980 , n246981 , n246982 , n246983 , n246984 , n246985 , n246986 , n246987 , n246988 , 
 n246989 , n246990 , n246991 , n246992 , n246993 , n246994 , n246995 , n246996 , n246997 , n246998 , 
 n246999 , n247000 , n247001 , n247002 , n247003 , n247004 , n247005 , n247006 , n247007 , n247008 , 
 n247009 , n247010 , n247011 , n247012 , n247013 , n247014 , n247015 , n247016 , n247017 , n247018 , 
 n247019 , n247020 , n247021 , n247022 , n247023 , n247024 , n247025 , n247026 , n247027 , n247028 , 
 n247029 , n247030 , n247031 , n247032 , n247033 , n247034 , n247035 , n247036 , n247037 , n247038 , 
 n247039 , n247040 , n247041 , n247042 , n247043 , n247044 , n247045 , n247046 , n247047 , n247048 , 
 n247049 , n247050 , n247051 , n247052 , n247053 , n247054 , n247055 , n247056 , n247057 , n247058 , 
 n247059 , n247060 , n247061 , n247062 , n247063 , n247064 , n247065 , n247066 , n247067 , n247068 , 
 n247069 , n247070 , n247071 , n247072 , n247073 , n247074 , n247075 , n247076 , n247077 , n247078 , 
 n247079 , n247080 , n247081 , n247082 , n247083 , n247084 , n247085 , n247086 , n247087 , n247088 , 
 n247089 , n247090 , n247091 , n247092 , n247093 , n247094 , n247095 , n247096 , n247097 , n247098 , 
 n247099 , n247100 , n247101 , n247102 , n247103 , n247104 , n247105 , n247106 , n247107 , n247108 , 
 n247109 , n247110 , n247111 , n247112 , n247113 , n247114 , n247115 , n247116 , n247117 , n247118 , 
 n247119 , n247120 , n247121 , n247122 , n247123 , n247124 , n247125 , n247126 , n247127 , n247128 , 
 n247129 , n247130 , n247131 , n247132 , n247133 , n247134 , n247135 , n247136 , n247137 , n247138 , 
 n247139 , n247140 , n247141 , n247142 , n247143 , n247144 , n247145 , n247146 , n247147 , n247148 , 
 n247149 , n247150 , n247151 , n247152 , n247153 , n247154 , n247155 , n247156 , n247157 , n247158 , 
 n247159 , n247160 , n247161 , n247162 , n247163 , n247164 , n247165 , n247166 , n247167 , n247168 , 
 n247169 , n247170 , n247171 , n247172 , n247173 , n247174 , n247175 , n247176 , n247177 , n247178 , 
 n247179 , n247180 , n247181 , n247182 , n247183 , n247184 , n247185 , n247186 , n247187 , n247188 , 
 n247189 , n247190 , n247191 , n247192 , n247193 , n247194 , n247195 , n247196 , n247197 , n247198 , 
 n247199 , n247200 , n247201 , n247202 , n247203 , n247204 , n247205 , n247206 , n247207 , n247208 , 
 n247209 , n247210 , n247211 , n247212 , n247213 , n247214 , n247215 , n247216 , n247217 , n247218 , 
 n247219 , n247220 , n247221 , n247222 , n247223 , n247224 , n247225 , n247226 , n247227 , n247228 , 
 n247229 , n247230 , n247231 , n247232 , n247233 , n247234 , n247235 , n247236 , n247237 , n247238 , 
 n247239 , n247240 , n247241 , n247242 , n247243 , n247244 , n247245 , n247246 , n247247 , n247248 , 
 n247249 , n247250 , n247251 , n247252 , n247253 , n247254 , n247255 , n247256 , n247257 , n247258 , 
 n247259 , n247260 , n247261 , n247262 , n247263 , n247264 , n247265 , n247266 , n247267 , n247268 , 
 n247269 , n247270 , n247271 , n247272 , n247273 , n247274 , n247275 , n247276 , n247277 , n247278 , 
 n247279 , n247280 , n247281 , n247282 , n247283 , n247284 , n247285 , n247286 , n247287 , n247288 , 
 n247289 , n247290 , n247291 , n247292 , n247293 , n247294 , n247295 , n247296 , n247297 , n247298 , 
 n247299 , n247300 , n247301 , n247302 , n247303 , n247304 , n247305 , n247306 , n247307 , n247308 , 
 n247309 , n247310 , n247311 , n247312 , n247313 , n247314 , n247315 , n247316 , n247317 , n247318 , 
 n247319 , n247320 , n247321 , n247322 , n247323 , n247324 , n247325 , n247326 , n247327 , n247328 , 
 n247329 , n247330 , n247331 , n247332 , n247333 , n247334 , n247335 , n247336 , n247337 , n247338 , 
 n247339 , n247340 , n247341 , n247342 , n247343 , n247344 , n247345 , n247346 , n247347 , n247348 , 
 n247349 , n247350 , n247351 , n247352 , n247353 , n247354 , n247355 , n247356 , n247357 , n247358 , 
 n247359 , n247360 , n247361 , n247362 , n247363 , n247364 , n247365 , n247366 , n247367 , n247368 , 
 n247369 , n247370 , n247371 , n247372 , n247373 , n247374 , n247375 , n247376 , n247377 , n247378 , 
 n247379 , n247380 , n247381 , n247382 , n247383 , n247384 , n247385 , n247386 , n247387 , n247388 , 
 n247389 , n247390 , n247391 , n247392 , n247393 , n247394 , n247395 , n247396 , n247397 , n247398 , 
 n247399 , n247400 , n247401 , n247402 , n247403 , n247404 , n247405 , n247406 , n247407 , n247408 , 
 n247409 , n247410 , n247411 , n247412 , n247413 , n247414 , n247415 , n247416 , n247417 , n247418 , 
 n247419 , n247420 , n247421 , n247422 , n247423 , n247424 , n247425 , n247426 , n247427 , n247428 , 
 n247429 , n247430 , n247431 , n247432 , n247433 , n247434 , n247435 , n247436 , n247437 , n247438 , 
 n247439 , n247440 , n247441 , n247442 , n247443 , n247444 , n247445 , n247446 , n247447 , n247448 , 
 n247449 , n247450 , n247451 , n247452 , n247453 , n247454 , n247455 , n247456 , n247457 , n247458 , 
 n247459 , n247460 , n247461 , n247462 , n247463 , n247464 , n247465 , n247466 , n247467 , n247468 , 
 n247469 , n247470 , n247471 , n247472 , n247473 , n247474 , n247475 , n247476 , n247477 , n247478 , 
 n247479 , n247480 , n247481 , n247482 , n247483 , n247484 , n247485 , n247486 , n247487 , n247488 , 
 n247489 , n247490 , n247491 , n247492 , n247493 , n247494 , n247495 , n247496 , n247497 , n247498 , 
 n247499 , n247500 , n247501 , n247502 , n247503 , n247504 , n247505 , n247506 , n247507 , n247508 , 
 n247509 , n247510 , n247511 , n247512 , n247513 , n247514 , n247515 , n247516 , n247517 , n247518 , 
 n247519 , n247520 , n247521 , n247522 , n247523 , n247524 , n247525 , n247526 , n247527 , n247528 , 
 n247529 , n247530 , n247531 , n247532 , n247533 , n247534 , n247535 , n247536 , n247537 , n247538 , 
 n247539 , n247540 , n247541 , n247542 , n247543 , n247544 , n247545 , n247546 , n247547 , n247548 , 
 n247549 , n247550 , n247551 , n247552 , n247553 , n247554 , n247555 , n247556 , n247557 , n247558 , 
 n247559 , n247560 , n247561 , n247562 , n247563 , n247564 , n247565 , n247566 , n247567 , n247568 , 
 n247569 , n247570 , n247571 , n247572 , n247573 , n247574 , n247575 , n247576 , n247577 , n247578 , 
 n247579 , n247580 , n247581 , n247582 , n247583 , n247584 , n247585 , n247586 , n247587 , n247588 , 
 n247589 , n247590 , n247591 , n247592 , n247593 , n247594 , n247595 , n247596 , n247597 , n247598 , 
 n247599 , n247600 , n247601 , n247602 , n247603 , n247604 , n247605 , n247606 , n247607 , n247608 , 
 n247609 , n247610 , n247611 , n247612 , n247613 , n247614 , n247615 , n247616 , n247617 , n247618 , 
 n247619 , n247620 , n247621 , n247622 , n247623 , n247624 , n247625 , n247626 , n247627 , n247628 , 
 n247629 , n247630 , n247631 , n247632 , n247633 , n247634 , n247635 , n247636 , n247637 , n247638 , 
 n247639 , n247640 , n247641 , n247642 , n247643 , n247644 , n247645 , n247646 , n247647 , n247648 , 
 n247649 , n247650 , n247651 , n247652 , n247653 , n247654 , n247655 , n247656 , n247657 , n247658 , 
 n247659 , n247660 , n247661 , n247662 , n247663 , n247664 , n247665 , n247666 , n247667 , n247668 , 
 n247669 , n247670 , n247671 , n247672 , n247673 , n247674 , n247675 , n247676 , n247677 , n247678 , 
 n247679 , n247680 , n247681 , n247682 , n247683 , n247684 , n247685 , n247686 , n247687 , n247688 , 
 n247689 , n247690 , n247691 , n247692 , n247693 , n247694 , n247695 , n247696 , n247697 , n247698 , 
 n247699 , n247700 , n247701 , n247702 , n247703 , n247704 , n247705 , n247706 , n247707 , n247708 , 
 n247709 , n247710 , n247711 , n247712 , n247713 , n247714 , n247715 , n247716 , n247717 , n247718 , 
 n247719 , n247720 , n247721 , n247722 , n247723 , n247724 , n247725 , n247726 , n247727 , n247728 , 
 n247729 , n247730 , n247731 , n247732 , n247733 , n247734 , n247735 , n247736 , n247737 , n247738 , 
 n247739 , n247740 , n247741 , n247742 , n247743 , n247744 , n247745 , n247746 , n247747 , n247748 , 
 n247749 , n247750 , n247751 , n247752 , n247753 , n247754 , n247755 , n247756 , n247757 , n247758 , 
 n247759 , n247760 , n247761 , n247762 , n247763 , n247764 , n247765 , n247766 , n247767 , n247768 , 
 n247769 , n247770 , n247771 , n247772 , n247773 , n247774 , n247775 , n247776 , n247777 , n247778 , 
 n247779 , n247780 , n247781 , n247782 , n247783 , n247784 , n247785 , n247786 , n247787 , n247788 , 
 n247789 , n247790 , n247791 , n247792 , n247793 , n247794 , n247795 , n247796 , n247797 , n247798 , 
 n247799 , n247800 , n247801 , n247802 , n247803 , n247804 , n247805 , n247806 , n247807 , n247808 , 
 n247809 , n247810 , n247811 , n247812 , n247813 , n247814 , n247815 , n247816 , n247817 , n247818 , 
 n247819 , n247820 , n247821 , n247822 , n247823 , n247824 , n247825 , n247826 , n247827 , n247828 , 
 n247829 , n247830 , n247831 , n247832 , n247833 , n247834 , n247835 , n247836 , n247837 , n247838 , 
 n247839 , n247840 , n247841 , n247842 , n247843 , n247844 , n247845 , n247846 , n247847 , n247848 , 
 n247849 , n247850 , n247851 , n247852 , n247853 , n247854 , n247855 , n247856 , n247857 , n247858 , 
 n247859 , n247860 , n247861 , n247862 , n247863 , n247864 , n247865 , n247866 , n247867 , n247868 , 
 n247869 , n247870 , n247871 , n247872 , n247873 , n247874 , n247875 , n247876 , n247877 , n247878 , 
 n247879 , n247880 , n247881 , n247882 , n247883 , n247884 , n247885 , n247886 , n247887 , n247888 , 
 n247889 , n247890 , n247891 , n247892 , n247893 , n247894 , n247895 , n247896 , n247897 , n247898 , 
 n247899 , n247900 , n247901 , n247902 , n247903 , n247904 , n247905 , n247906 , n247907 , n247908 , 
 n247909 , n247910 , n247911 , n247912 , n247913 , n247914 , n247915 , n247916 , n247917 , n247918 , 
 n247919 , n247920 , n247921 , n247922 , n247923 , n247924 , n247925 , n247926 , n247927 , n247928 , 
 n247929 , n247930 , n247931 , n247932 , n247933 , n247934 , n247935 , n247936 , n247937 , n247938 , 
 n247939 , n247940 , n247941 , n247942 , n247943 , n247944 , n247945 , n247946 , n247947 , n247948 , 
 n247949 , n247950 , n247951 , n247952 , n247953 , n247954 , n247955 , n247956 , n247957 , n247958 , 
 n247959 , n247960 , n247961 , n247962 , n247963 , n247964 , n247965 , n247966 , n247967 , n247968 , 
 n247969 , n247970 , n247971 , n247972 , n247973 , n247974 , n247975 , n247976 , n247977 , n247978 , 
 n247979 , n247980 , n247981 , n247982 , n247983 , n247984 , n247985 , n247986 , n247987 , n247988 , 
 n247989 , n247990 , n247991 , n247992 , n247993 , n247994 , n247995 , n247996 , n247997 , n247998 , 
 n247999 , n248000 , n248001 , n248002 , n248003 , n248004 , n248005 , n248006 , n248007 , n248008 , 
 n248009 , n248010 , n248011 , n248012 , n248013 , n248014 , n248015 , n248016 , n248017 , n248018 , 
 n248019 , n248020 , n248021 , n248022 , n248023 , n248024 , n248025 , n248026 , n248027 , n248028 , 
 n248029 , n248030 , n248031 , n248032 , n248033 , n248034 , n248035 , n248036 , n248037 , n248038 , 
 n248039 , n248040 , n248041 , n248042 , n248043 , n248044 , n248045 , n248046 , n248047 , n248048 , 
 n248049 , n248050 , n248051 , n248052 , n248053 , n248054 , n248055 , n248056 , n248057 , n248058 , 
 n248059 , n248060 , n248061 , n248062 , n248063 , n248064 , n248065 , n248066 , n248067 , n248068 , 
 n248069 , n248070 , n248071 , n248072 , n248073 , n248074 , n248075 , n248076 , n248077 , n248078 , 
 n248079 , n248080 , n248081 , n248082 , n248083 , n248084 , n248085 , n248086 , n248087 , n248088 , 
 n248089 , n248090 , n248091 , n248092 , n248093 , n248094 , n248095 , n248096 , n248097 , n248098 , 
 n248099 , n248100 , n248101 , n248102 , n248103 , n248104 , n248105 , n248106 , n248107 , n248108 , 
 n248109 , n248110 , n248111 , n248112 , n248113 , n248114 , n248115 , n248116 , n248117 , n248118 , 
 n248119 , n248120 , n248121 , n248122 , n248123 , n248124 , n248125 , n248126 , n248127 , n248128 , 
 n248129 , n248130 , n248131 , n248132 , n248133 , n248134 , n248135 , n248136 , n248137 , n248138 , 
 n248139 , n248140 , n248141 , n248142 , n248143 , n248144 , n248145 , n248146 , n248147 , n248148 , 
 n248149 , n248150 , n248151 , n248152 , n248153 , n248154 , n248155 , n248156 , n248157 , n248158 , 
 n248159 , n248160 , n248161 , n248162 , n248163 , n248164 , n248165 , n248166 , n248167 , n248168 , 
 n248169 , n248170 , n248171 , n248172 , n248173 , n248174 , n248175 , n248176 , n248177 , n248178 , 
 n248179 , n248180 , n248181 , n248182 , n248183 , n248184 , n248185 , n248186 , n248187 , n248188 , 
 n248189 , n248190 , n248191 , n248192 , n248193 , n248194 , n248195 , n248196 , n248197 , n248198 , 
 n248199 , n248200 , n248201 , n248202 , n248203 , n248204 , n248205 , n248206 , n248207 , n248208 , 
 n248209 , n248210 , n248211 , n248212 , n248213 , n248214 , n248215 , n248216 , n248217 , n248218 , 
 n248219 , n248220 , n248221 , n248222 , n248223 , n248224 , n248225 , n248226 , n248227 , n248228 , 
 n248229 , n248230 , n248231 , n248232 , n248233 , n248234 , n248235 , n248236 , n248237 , n248238 , 
 n248239 , n248240 , n248241 , n248242 , n248243 , n248244 , n248245 , n248246 , n248247 , n248248 , 
 n248249 , n248250 , n248251 , n248252 , n248253 , n248254 , n248255 , n248256 , n248257 , n248258 , 
 n248259 , n248260 , n248261 , n248262 , n248263 , n248264 , n248265 , n248266 , n248267 , n248268 , 
 n248269 , n248270 , n248271 , n248272 , n248273 , n248274 , n248275 , n248276 , n248277 , n248278 , 
 n248279 , n248280 , n248281 , n248282 , n248283 , n248284 , n248285 , n248286 , n248287 , n248288 , 
 n248289 , n248290 , n248291 , n248292 , n248293 , n248294 , n248295 , n248296 , n248297 , n248298 , 
 n248299 , n248300 , n248301 , n248302 , n248303 , n248304 , n248305 , n248306 , n248307 , n248308 , 
 n248309 , n248310 , n248311 , n248312 , n248313 , n248314 , n248315 , n248316 , n248317 , n248318 , 
 n248319 , n248320 , n248321 , n248322 , n248323 , n248324 , n248325 , n248326 , n248327 , n248328 , 
 n248329 , n248330 , n248331 , n248332 , n248333 , n248334 , n248335 , n248336 , n248337 , n248338 , 
 n248339 , n248340 , n248341 , n248342 , n248343 , n248344 , n248345 , n248346 , n248347 , n248348 , 
 n248349 , n248350 , n248351 , n248352 , n248353 , n248354 , n248355 , n248356 , n248357 , n248358 , 
 n248359 , n248360 , n248361 , n248362 , n248363 , n248364 , n248365 , n248366 , n248367 , n248368 , 
 n248369 , n248370 , n248371 , n248372 , n248373 , n248374 , n248375 , n248376 , n248377 , n248378 , 
 n248379 , n248380 , n248381 , n248382 , n248383 , n248384 , n248385 , n248386 , n248387 , n248388 , 
 n248389 , n248390 , n248391 , n248392 , n248393 , n248394 , n248395 , n248396 , n248397 , n248398 , 
 n248399 , n248400 , n248401 , n248402 , n248403 , n248404 , n248405 , n248406 , n248407 , n248408 , 
 n248409 , n248410 , n248411 , n248412 , n248413 , n248414 , n248415 , n248416 , n248417 , n248418 , 
 n248419 , n248420 , n248421 , n248422 , n248423 , n248424 , n248425 , n248426 , n248427 , n248428 , 
 n248429 , n248430 , n248431 , n248432 , n248433 , n248434 , n248435 , n248436 , n248437 , n248438 , 
 n248439 , n248440 , n248441 , n248442 , n248443 , n248444 , n248445 , n248446 , n248447 , n248448 , 
 n248449 , n248450 , n248451 , n248452 , n248453 , n248454 , n248455 , n248456 , n248457 , n248458 , 
 n248459 , n248460 , n248461 , n248462 , n248463 , n248464 , n248465 , n248466 , n248467 , n248468 , 
 n248469 , n248470 , n248471 , n248472 , n248473 , n248474 , n248475 , n248476 , n248477 , n248478 , 
 n248479 , n248480 , n248481 , n248482 , n248483 , n248484 , n248485 , n248486 , n248487 , n248488 , 
 n248489 , n248490 , n248491 , n248492 , n248493 , n248494 , n248495 , n248496 , n248497 , n248498 , 
 n248499 , n248500 , n248501 , n248502 , n248503 , n248504 , n248505 , n248506 , n248507 , n248508 , 
 n248509 , n248510 , n248511 , n248512 , n248513 , n248514 , n248515 , n248516 , n248517 , n248518 , 
 n248519 , n248520 , n248521 , n248522 , n248523 , n248524 , n248525 , n248526 , n248527 , n248528 , 
 n248529 , n248530 , n248531 , n248532 , n248533 , n248534 , n248535 , n248536 , n248537 , n248538 , 
 n248539 , n248540 , n248541 , n248542 , n248543 , n248544 , n248545 , n248546 , n248547 , n248548 , 
 n248549 , n248550 , n248551 , n248552 , n248553 , n248554 , n248555 , n248556 , n248557 , n248558 , 
 n248559 , n248560 , n248561 , n248562 , n248563 , n248564 , n248565 , n248566 , n248567 , n248568 , 
 n248569 , n248570 , n248571 , n248572 , n248573 , n248574 , n248575 , n248576 , n248577 , n248578 , 
 n248579 , n248580 , n248581 , n248582 , n248583 , n248584 , n248585 , n248586 , n248587 , n248588 , 
 n248589 , n248590 , n248591 , n248592 , n248593 , n248594 , n248595 , n248596 , n248597 , n248598 , 
 n248599 , n248600 , n248601 , n248602 , n248603 , n248604 , n248605 , n248606 , n248607 , n248608 , 
 n248609 , n248610 , n248611 , n248612 , n248613 , n248614 , n248615 , n248616 , n248617 , n248618 , 
 n248619 , n248620 , n248621 , n248622 , n248623 , n248624 , n248625 , n248626 , n248627 , n248628 , 
 n248629 , n248630 , n248631 , n248632 , n248633 , n248634 , n248635 , n248636 , n248637 , n248638 , 
 n248639 , n248640 , n248641 , n248642 , n248643 , n248644 , n248645 , n248646 , n248647 , n248648 , 
 n248649 , n248650 , n248651 , n248652 , n248653 , n248654 , n248655 , n248656 , n248657 , n248658 , 
 n248659 , n248660 , n248661 , n248662 , n248663 , n248664 , n248665 , n248666 , n248667 , n248668 , 
 n248669 , n248670 , n248671 , n248672 , n248673 , n248674 , n248675 , n248676 , n248677 , n248678 , 
 n248679 , n248680 , n248681 , n248682 , n248683 , n248684 , n248685 , n248686 , n248687 , n248688 , 
 n248689 , n248690 , n248691 , n248692 , n248693 , n248694 , n248695 , n248696 , n248697 , n248698 , 
 n248699 , n248700 , n248701 , n248702 , n248703 , n248704 , n248705 , n248706 , n248707 , n248708 , 
 n248709 , n248710 , n248711 , n248712 , n248713 , n248714 , n248715 , n248716 , n248717 , n248718 , 
 n248719 , n248720 , n248721 , n248722 , n248723 , n248724 , n248725 , n248726 , n248727 , n248728 , 
 n248729 , n248730 , n248731 , n248732 , n248733 , n248734 , n248735 , n248736 , n248737 , n248738 , 
 n248739 , n248740 , n248741 , n248742 , n248743 , n248744 , n248745 , n248746 , n248747 , n248748 , 
 n248749 , n248750 , n248751 , n248752 , n248753 , n248754 , n248755 , n248756 , n248757 , n248758 , 
 n248759 , n248760 , n248761 , n248762 , n248763 , n248764 , n248765 , n248766 , n248767 , n248768 , 
 n248769 , n248770 , n248771 , n248772 , n248773 , n248774 , n248775 , n248776 , n248777 , n248778 , 
 n248779 , n248780 , n248781 , n248782 , n248783 , n248784 , n248785 , n248786 , n248787 , n248788 , 
 n248789 , n248790 , n248791 , n248792 , n248793 , n248794 , n248795 , n248796 , n248797 , n248798 , 
 n248799 , n248800 , n248801 , n248802 , n248803 , n248804 , n248805 , n248806 , n248807 , n248808 , 
 n248809 , n248810 , n248811 , n248812 , n248813 , n248814 , n248815 , n248816 , n248817 , n248818 , 
 n248819 , n248820 , n248821 , n248822 , n248823 , n248824 , n248825 , n248826 , n248827 , n248828 , 
 n248829 , n248830 , n248831 , n248832 , n248833 , n248834 , n248835 , n248836 , n248837 , n248838 , 
 n248839 , n248840 , n248841 , n248842 , n248843 , n248844 , n248845 , n248846 , n248847 , n248848 , 
 n248849 , n248850 , n248851 , n248852 , n248853 , n248854 , n248855 , n248856 , n248857 , n248858 , 
 n248859 , n248860 , n248861 , n248862 , n248863 , n248864 , n248865 , n248866 , n248867 , n248868 , 
 n248869 , n248870 , n248871 , n248872 , n248873 , n248874 , n248875 , n248876 , n248877 , n248878 , 
 n248879 , n248880 , n248881 , n248882 , n248883 , n248884 , n248885 , n248886 , n248887 , n248888 , 
 n248889 , n248890 , n248891 , n248892 , n248893 , n248894 , n248895 , n248896 , n248897 , n248898 , 
 n248899 , n248900 , n248901 , n248902 , n248903 , n248904 , n248905 , n248906 , n248907 , n248908 , 
 n248909 , n248910 , n248911 , n248912 , n248913 , n248914 , n248915 , n248916 , n248917 , n248918 , 
 n248919 , n248920 , n248921 , n248922 , n248923 , n248924 , n248925 , n248926 , n248927 , n248928 , 
 n248929 , n248930 , n248931 , n248932 , n248933 , n248934 , n248935 , n248936 , n248937 , n248938 , 
 n248939 , n248940 , n248941 , n248942 , n248943 , n248944 , n248945 , n248946 , n248947 , n248948 , 
 n248949 , n248950 , n248951 , n248952 , n248953 , n248954 , n248955 , n248956 , n248957 , n248958 , 
 n248959 , n248960 , n248961 , n248962 , n248963 , n248964 , n248965 , n248966 , n248967 , n248968 , 
 n248969 , n248970 , n248971 , n248972 , n248973 , n248974 , n248975 , n248976 , n248977 , n248978 , 
 n248979 , n248980 , n248981 , n248982 , n248983 , n248984 , n248985 , n248986 , n248987 , n248988 , 
 n248989 , n248990 , n248991 , n248992 , n248993 , n248994 , n248995 , n248996 , n248997 , n248998 , 
 n248999 , n249000 , n249001 , n249002 , n249003 , n249004 , n249005 , n249006 , n249007 , n249008 , 
 n249009 , n249010 , n249011 , n249012 , n249013 , n249014 , n249015 , n249016 , n249017 , n249018 , 
 n249019 , n249020 , n249021 , n249022 , n249023 , n249024 , n249025 , n249026 , n249027 , n249028 , 
 n249029 , n249030 , n249031 , n249032 , n249033 , n249034 , n249035 , n249036 , n249037 , n249038 , 
 n249039 , n249040 , n249041 , n249042 , n249043 , n249044 , n249045 , n249046 , n249047 , n249048 , 
 n249049 , n249050 , n249051 , n249052 , n249053 , n249054 , n249055 , n249056 , n249057 , n249058 , 
 n249059 , n249060 , n249061 , n249062 , n249063 , n249064 , n249065 , n249066 , n249067 , n249068 , 
 n249069 , n249070 , n249071 , n249072 , n249073 , n249074 , n249075 , n249076 , n249077 , n249078 , 
 n249079 , n249080 , n249081 , n249082 , n249083 , n249084 , n249085 , n249086 , n249087 , n249088 , 
 n249089 , n249090 , n249091 , n249092 , n249093 , n249094 , n249095 , n249096 , n249097 , n249098 , 
 n249099 , n249100 , n249101 , n249102 , n249103 , n249104 , n249105 , n249106 , n249107 , n249108 , 
 n249109 , n249110 , n249111 , n249112 , n249113 , n249114 , n249115 , n249116 , n249117 , n249118 , 
 n249119 , n249120 , n249121 , n249122 , n249123 , n249124 , n249125 , n249126 , n249127 , n249128 , 
 n249129 , n249130 , n249131 , n249132 , n249133 , n249134 , n249135 , n249136 , n249137 , n249138 , 
 n249139 , n249140 , n249141 , n249142 , n249143 , n249144 , n249145 , n249146 , n249147 , n249148 , 
 n249149 , n249150 , n249151 , n249152 , n249153 , n249154 , n249155 , n249156 , n249157 , n249158 , 
 n249159 , n249160 , n249161 , n249162 , n249163 , n249164 , n249165 , n249166 , n249167 , n249168 , 
 n249169 , n249170 , n249171 , n249172 , n249173 , n249174 , n249175 , n249176 , n249177 , n249178 , 
 n249179 , n249180 , n249181 , n249182 , n249183 , n249184 , n249185 , n249186 , n249187 , n249188 , 
 n249189 , n249190 , n249191 , n249192 , n249193 , n249194 , n249195 , n249196 , n249197 , n249198 , 
 n249199 , n249200 , n249201 , n249202 , n249203 , n249204 , n249205 , n249206 , n249207 , n249208 , 
 n249209 , n249210 , n249211 , n249212 , n249213 , n249214 , n249215 , n249216 , n249217 , n249218 , 
 n249219 , n249220 , n249221 , n249222 , n249223 , n249224 , n249225 , n249226 , n249227 , n249228 , 
 n249229 , n249230 , n249231 , n249232 , n249233 , n249234 , n249235 , n249236 , n249237 , n249238 , 
 n249239 , n249240 , n249241 , n249242 , n249243 , n249244 , n249245 , n249246 , n249247 , n249248 , 
 n249249 , n249250 , n249251 , n249252 , n249253 , n249254 , n249255 , n249256 , n249257 , n249258 , 
 n249259 , n249260 , n249261 , n249262 , n249263 , n249264 , n249265 , n249266 , n249267 , n249268 , 
 n249269 , n249270 , n249271 , n249272 , n249273 , n249274 , n249275 , n249276 , n249277 , n249278 , 
 n249279 , n249280 , n249281 , n249282 , n249283 , n249284 , n249285 , n249286 , n249287 , n249288 , 
 n249289 , n249290 , n249291 , n249292 , n249293 , n249294 , n249295 , n249296 , n249297 , n249298 , 
 n249299 , n249300 , n249301 , n249302 , n249303 , n249304 , n249305 , n249306 , n249307 , n249308 , 
 n249309 , n249310 , n249311 , n249312 , n249313 , n249314 , n249315 , n249316 , n249317 , n249318 , 
 n249319 , n249320 , n249321 , n249322 , n249323 , n249324 , n249325 , n249326 , n249327 , n249328 , 
 n249329 , n249330 , n249331 , n249332 , n249333 , n249334 , n249335 , n249336 , n249337 , n249338 , 
 n249339 , n249340 , n249341 , n249342 , n249343 , n249344 , n249345 , n249346 , n249347 , n249348 , 
 n249349 , n249350 , n249351 , n249352 , n249353 , n249354 , n249355 , n249356 , n249357 , n249358 , 
 n249359 , n249360 , n249361 , n249362 , n249363 , n249364 , n249365 , n249366 , n249367 , n249368 , 
 n249369 , n249370 , n249371 , n249372 , n249373 , n249374 , n249375 , n249376 , n249377 , n249378 , 
 n249379 , n249380 , n249381 , n249382 , n249383 , n249384 , n249385 , n249386 , n249387 , n249388 , 
 n249389 , n249390 , n249391 , n249392 , n249393 , n249394 , n249395 , n249396 , n249397 , n249398 , 
 n249399 , n249400 , n249401 , n249402 , n249403 , n249404 , n249405 , n249406 , n249407 , n249408 , 
 n249409 , n249410 , n249411 , n249412 , n249413 , n249414 , n249415 , n249416 , n249417 , n249418 , 
 n249419 , n249420 , n249421 , n249422 , n249423 , n249424 , n249425 , n249426 , n249427 , n249428 , 
 n249429 , n249430 , n249431 , n249432 , n249433 , n249434 , n249435 , n249436 , n249437 , n249438 , 
 n249439 , n249440 , n249441 , n249442 , n249443 , n249444 , n249445 , n249446 , n249447 , n249448 , 
 n249449 , n249450 , n249451 , n249452 , n249453 , n249454 , n249455 , n249456 , n249457 , n249458 , 
 n249459 , n249460 , n249461 , n249462 , n249463 , n249464 , n249465 , n249466 , n249467 , n249468 , 
 n249469 , n249470 , n249471 , n249472 , n249473 , n249474 , n249475 , n249476 , n249477 , n249478 , 
 n249479 , n249480 , n249481 , n249482 , n249483 , n249484 , n249485 , n249486 , n249487 , n249488 , 
 n249489 , n249490 , n249491 , n249492 , n249493 , n249494 , n249495 , n249496 , n249497 , n249498 , 
 n249499 , n249500 , n249501 , n249502 , n249503 , n249504 , n249505 , n249506 , n249507 , n249508 , 
 n249509 , n249510 , n249511 , n249512 , n249513 , n249514 , n249515 , n249516 , n249517 , n249518 , 
 n249519 , n249520 , n249521 , n249522 , n249523 , n249524 , n249525 , n249526 , n249527 , n249528 , 
 n249529 , n249530 , n249531 , n249532 , n249533 , n249534 , n249535 , n249536 , n249537 , n249538 , 
 n249539 , n249540 , n249541 , n249542 , n249543 , n249544 , n249545 , n249546 , n249547 , n249548 , 
 n249549 , n249550 , n249551 , n249552 , n249553 , n249554 , n249555 , n249556 , n249557 , n249558 , 
 n249559 , n249560 , n249561 , n249562 , n249563 , n249564 , n249565 , n249566 , n249567 , n249568 , 
 n249569 , n249570 , n249571 , n249572 , n249573 , n249574 , n249575 , n249576 , n249577 , n249578 , 
 n249579 , n249580 , n249581 , n249582 , n249583 , n249584 , n249585 , n249586 , n249587 , n249588 , 
 n249589 , n249590 , n249591 , n249592 , n249593 , n249594 , n249595 , n249596 , n249597 , n249598 , 
 n249599 , n249600 , n249601 , n249602 , n249603 , n249604 , n249605 , n249606 , n249607 , n249608 , 
 n249609 , n249610 , n249611 , n249612 , n249613 , n249614 , n249615 , n249616 , n249617 , n249618 , 
 n249619 , n249620 , n249621 , n249622 , n249623 , n249624 , n249625 , n249626 , n249627 , n249628 , 
 n249629 , n249630 , n249631 , n249632 , n249633 , n249634 , n249635 , n249636 , n249637 , n249638 , 
 n249639 , n249640 , n249641 , n249642 , n249643 , n249644 , n249645 , n249646 , n249647 , n249648 , 
 n249649 , n249650 , n249651 , n249652 , n249653 , n249654 , n249655 , n249656 , n249657 , n249658 , 
 n249659 , n249660 , n249661 , n249662 , n249663 , n249664 , n249665 , n249666 , n249667 , n249668 , 
 n249669 , n249670 , n249671 , n249672 , n249673 , n249674 , n249675 , n249676 , n249677 , n249678 , 
 n249679 , n249680 , n249681 , n249682 , n249683 , n249684 , n249685 , n249686 , n249687 , n249688 , 
 n249689 , n249690 , n249691 , n249692 , n249693 , n249694 , n249695 , n249696 , n249697 , n249698 , 
 n249699 , n249700 , n249701 , n249702 , n249703 , n249704 , n249705 , n249706 , n249707 , n249708 , 
 n249709 , n249710 , n249711 , n249712 , n249713 , n249714 , n249715 , n249716 , n249717 , n249718 , 
 n249719 , n249720 , n249721 , n249722 , n249723 , n249724 , n249725 , n249726 , n249727 , n249728 , 
 n249729 , n249730 , n249731 , n249732 , n249733 , n249734 , n249735 , n249736 , n249737 , n249738 , 
 n249739 , n249740 , n249741 , n249742 , n249743 , n249744 , n249745 , n249746 , n249747 , n249748 , 
 n249749 , n249750 , n249751 , n249752 , n249753 , n249754 , n249755 , n249756 , n249757 , n249758 , 
 n249759 , n249760 , n249761 , n249762 , n249763 , n249764 , n249765 , n249766 , n249767 , n249768 , 
 n249769 , n249770 , n249771 , n249772 , n249773 , n249774 , n249775 , n249776 , n249777 , n249778 , 
 n249779 , n249780 , n249781 , n249782 , n249783 , n249784 , n249785 , n249786 , n249787 , n249788 , 
 n249789 , n249790 , n249791 , n249792 , n249793 , n249794 , n249795 , n249796 , n249797 , n249798 , 
 n249799 , n249800 , n249801 , n249802 , n249803 , n249804 , n249805 , n249806 , n249807 , n249808 , 
 n249809 , n249810 , n249811 , n249812 , n249813 , n249814 , n249815 , n249816 , n249817 , n249818 , 
 n249819 , n249820 , n249821 , n249822 , n249823 , n249824 , n249825 , n249826 , n249827 , n249828 , 
 n249829 , n249830 , n249831 , n249832 , n249833 , n249834 , n249835 , n249836 , n249837 , n249838 , 
 n249839 , n249840 , n249841 , n249842 , n249843 , n249844 , n249845 , n249846 , n249847 , n249848 , 
 n249849 , n249850 , n249851 , n249852 , n249853 , n249854 , n249855 , n249856 , n249857 , n249858 , 
 n249859 , n249860 , n249861 , n249862 , n249863 , n249864 , n249865 , n249866 , n249867 , n249868 , 
 n249869 , n249870 , n249871 , n249872 , n249873 , n249874 , n249875 , n249876 , n249877 , n249878 , 
 n249879 , n249880 , n249881 , n249882 , n249883 , n249884 , n249885 , n249886 , n249887 , n249888 , 
 n249889 , n249890 , n249891 , n249892 , n249893 , n249894 , n249895 , n249896 , n249897 , n249898 , 
 n249899 , n249900 , n249901 , n249902 , n249903 , n249904 , n249905 , n249906 , n249907 , n249908 , 
 n249909 , n249910 , n249911 , n249912 , n249913 , n249914 , n249915 , n249916 , n249917 , n249918 , 
 n249919 , n249920 , n249921 , n249922 , n249923 , n249924 , n249925 , n249926 , n249927 , n249928 , 
 n249929 , n249930 , n249931 , n249932 , n249933 , n249934 , n249935 , n249936 , n249937 , n249938 , 
 n249939 , n249940 , n249941 , n249942 , n249943 , n249944 , n249945 , n249946 , n249947 , n249948 , 
 n249949 , n249950 , n249951 , n249952 , n249953 , n249954 , n249955 , n249956 , n249957 , n249958 , 
 n249959 , n249960 , n249961 , n249962 , n249963 , n249964 , n249965 , n249966 , n249967 , n249968 , 
 n249969 , n249970 , n249971 , n249972 , n249973 , n249974 , n249975 , n249976 , n249977 , n249978 , 
 n249979 , n249980 , n249981 , n249982 , n249983 , n249984 , n249985 , n249986 , n249987 , n249988 , 
 n249989 , n249990 , n249991 , n249992 , n249993 , n249994 , n249995 , n249996 , n249997 , n249998 , 
 n249999 , n250000 , n250001 , n250002 , n250003 , n250004 , n250005 , n250006 , n250007 , n250008 , 
 n250009 , n250010 , n250011 , n250012 , n250013 , n250014 , n250015 , n250016 , n250017 , n250018 , 
 n250019 , n250020 , n250021 , n250022 , n250023 , n250024 , n250025 , n250026 , n250027 , n250028 , 
 n250029 , n250030 , n250031 , n250032 , n250033 , n250034 , n250035 , n250036 , n250037 , n250038 , 
 n250039 , n250040 , n250041 , n250042 , n250043 , n250044 , n250045 , n250046 , n250047 , n250048 , 
 n250049 , n250050 , n250051 , n250052 , n250053 , n250054 , n250055 , n250056 , n250057 , n250058 , 
 n250059 , n250060 , n250061 , n250062 , n250063 , n250064 , n250065 , n250066 , n250067 , n250068 , 
 n250069 , n250070 , n250071 , n250072 , n250073 , n250074 , n250075 , n250076 , n250077 , n250078 , 
 n250079 , n250080 , n250081 , n250082 , n250083 , n250084 , n250085 , n250086 , n250087 , n250088 , 
 n250089 , n250090 , n250091 , n250092 , n250093 , n250094 , n250095 , n250096 , n250097 , n250098 , 
 n250099 , n250100 , n250101 , n250102 , n250103 , n250104 , n250105 , n250106 , n250107 , n250108 , 
 n250109 , n250110 , n250111 , n250112 , n250113 , n250114 , n250115 , n250116 , n250117 , n250118 , 
 n250119 , n250120 , n250121 , n250122 , n250123 , n250124 , n250125 , n250126 , n250127 , n250128 , 
 n250129 , n250130 , n250131 , n250132 , n250133 , n250134 , n250135 , n250136 , n250137 , n250138 , 
 n250139 , n250140 , n250141 , n250142 , n250143 , n250144 , n250145 , n250146 , n250147 , n250148 , 
 n250149 , n250150 , n250151 , n250152 , n250153 , n250154 , n250155 , n250156 , n250157 , n250158 , 
 n250159 , n250160 , n250161 , n250162 , n250163 , n250164 , n250165 , n250166 , n250167 , n250168 , 
 n250169 , n250170 , n250171 , n250172 , n250173 , n250174 , n250175 , n250176 , n250177 , n250178 , 
 n250179 , n250180 , n250181 , n250182 , n250183 , n250184 , n250185 , n250186 , n250187 , n250188 , 
 n250189 , n250190 , n250191 , n250192 , n250193 , n250194 , n250195 , n250196 , n250197 , n250198 , 
 n250199 , n250200 , n250201 , n250202 , n250203 , n250204 , n250205 , n250206 , n250207 , n250208 , 
 n250209 , n250210 , n250211 , n250212 , n250213 , n250214 , n250215 , n250216 , n250217 , n250218 , 
 n250219 , n250220 , n250221 , n250222 , n250223 , n250224 , n250225 , n250226 , n250227 , n250228 , 
 n250229 , n250230 , n250231 , n250232 , n250233 , n250234 , n250235 , n250236 , n250237 , n250238 , 
 n250239 , n250240 , n250241 , n250242 , n250243 , n250244 , n250245 , n250246 , n250247 , n250248 , 
 n250249 , n250250 , n250251 , n250252 , n250253 , n250254 , n250255 , n250256 , n250257 , n250258 , 
 n250259 , n250260 , n250261 , n250262 , n250263 , n250264 , n250265 , n250266 , n250267 , n250268 , 
 n250269 , n250270 , n250271 , n250272 , n250273 , n250274 , n250275 , n250276 , n250277 , n250278 , 
 n250279 , n250280 , n250281 , n250282 , n250283 , n250284 , n250285 , n250286 , n250287 , n250288 , 
 n250289 , n250290 , n250291 , n250292 , n250293 , n250294 , n250295 , n250296 , n250297 , n250298 , 
 n250299 , C0n , C0 ;
buf ( n768 , n0 );
buf ( n769 , n1 );
buf ( n770 , n2 );
buf ( n771 , n3 );
buf ( n772 , n4 );
buf ( n773 , n5 );
buf ( n774 , n6 );
buf ( n775 , n7 );
buf ( n776 , n8 );
buf ( n777 , n9 );
buf ( n778 , n10 );
buf ( n779 , n11 );
buf ( n780 , n12 );
buf ( n781 , n13 );
buf ( n782 , n14 );
buf ( n783 , n15 );
buf ( n784 , n16 );
buf ( n785 , n17 );
buf ( n786 , n18 );
buf ( n787 , n19 );
buf ( n788 , n20 );
buf ( n789 , n21 );
buf ( n790 , n22 );
buf ( n791 , n23 );
buf ( n792 , n24 );
buf ( n793 , n25 );
buf ( n794 , n26 );
buf ( n795 , n27 );
buf ( n796 , n28 );
buf ( n797 , n29 );
buf ( n798 , n30 );
buf ( n799 , n31 );
buf ( n800 , n32 );
buf ( n801 , n33 );
buf ( n802 , n34 );
buf ( n803 , n35 );
buf ( n804 , n36 );
buf ( n805 , n37 );
buf ( n806 , n38 );
buf ( n807 , n39 );
buf ( n808 , n40 );
buf ( n809 , n41 );
buf ( n810 , n42 );
buf ( n811 , n43 );
buf ( n812 , n44 );
buf ( n813 , n45 );
buf ( n814 , n46 );
buf ( n815 , n47 );
buf ( n816 , n48 );
buf ( n817 , n49 );
buf ( n818 , n50 );
buf ( n819 , n51 );
buf ( n820 , n52 );
buf ( n821 , n53 );
buf ( n822 , n54 );
buf ( n823 , n55 );
buf ( n824 , n56 );
buf ( n825 , n57 );
buf ( n826 , n58 );
buf ( n827 , n59 );
buf ( n828 , n60 );
buf ( n829 , n61 );
buf ( n830 , n62 );
buf ( n831 , n63 );
buf ( n832 , n64 );
buf ( n833 , n65 );
buf ( n834 , n66 );
buf ( n835 , n67 );
buf ( n836 , n68 );
buf ( n837 , n69 );
buf ( n838 , n70 );
buf ( n839 , n71 );
buf ( n840 , n72 );
buf ( n841 , n73 );
buf ( n842 , n74 );
buf ( n843 , n75 );
buf ( n844 , n76 );
buf ( n845 , n77 );
buf ( n846 , n78 );
buf ( n847 , n79 );
buf ( n848 , n80 );
buf ( n849 , n81 );
buf ( n850 , n82 );
buf ( n851 , n83 );
buf ( n852 , n84 );
buf ( n853 , n85 );
buf ( n854 , n86 );
buf ( n855 , n87 );
buf ( n856 , n88 );
buf ( n857 , n89 );
buf ( n858 , n90 );
buf ( n859 , n91 );
buf ( n860 , n92 );
buf ( n861 , n93 );
buf ( n862 , n94 );
buf ( n863 , n95 );
buf ( n864 , n96 );
buf ( n865 , n97 );
buf ( n866 , n98 );
buf ( n867 , n99 );
buf ( n868 , n100 );
buf ( n869 , n101 );
buf ( n870 , n102 );
buf ( n871 , n103 );
buf ( n872 , n104 );
buf ( n873 , n105 );
buf ( n874 , n106 );
buf ( n875 , n107 );
buf ( n876 , n108 );
buf ( n877 , n109 );
buf ( n878 , n110 );
buf ( n879 , n111 );
buf ( n880 , n112 );
buf ( n881 , n113 );
buf ( n882 , n114 );
buf ( n883 , n115 );
buf ( n884 , n116 );
buf ( n885 , n117 );
buf ( n886 , n118 );
buf ( n887 , n119 );
buf ( n888 , n120 );
buf ( n889 , n121 );
buf ( n890 , n122 );
buf ( n891 , n123 );
buf ( n892 , n124 );
buf ( n893 , n125 );
buf ( n894 , n126 );
buf ( n895 , n127 );
buf ( n128 , n896 );
buf ( n129 , n897 );
buf ( n130 , n898 );
buf ( n131 , n899 );
buf ( n132 , n900 );
buf ( n133 , n901 );
buf ( n134 , n902 );
buf ( n135 , n903 );
buf ( n136 , n904 );
buf ( n137 , n905 );
buf ( n138 , n906 );
buf ( n139 , n907 );
buf ( n140 , n908 );
buf ( n141 , n909 );
buf ( n142 , n910 );
buf ( n143 , n911 );
buf ( n144 , n912 );
buf ( n145 , n913 );
buf ( n146 , n914 );
buf ( n147 , n915 );
buf ( n148 , n916 );
buf ( n149 , n917 );
buf ( n150 , n918 );
buf ( n151 , n919 );
buf ( n152 , n920 );
buf ( n153 , n921 );
buf ( n154 , n922 );
buf ( n155 , n923 );
buf ( n156 , n924 );
buf ( n157 , n925 );
buf ( n158 , n926 );
buf ( n159 , n927 );
buf ( n160 , n928 );
buf ( n161 , n929 );
buf ( n162 , n930 );
buf ( n163 , n931 );
buf ( n164 , n932 );
buf ( n165 , n933 );
buf ( n166 , n934 );
buf ( n167 , n935 );
buf ( n168 , n936 );
buf ( n169 , n937 );
buf ( n170 , n938 );
buf ( n171 , n939 );
buf ( n172 , n940 );
buf ( n173 , n941 );
buf ( n174 , n942 );
buf ( n175 , n943 );
buf ( n176 , n944 );
buf ( n177 , n945 );
buf ( n178 , n946 );
buf ( n179 , n947 );
buf ( n180 , n948 );
buf ( n181 , n949 );
buf ( n182 , n950 );
buf ( n183 , n951 );
buf ( n184 , n952 );
buf ( n185 , n953 );
buf ( n186 , n954 );
buf ( n187 , n955 );
buf ( n188 , n956 );
buf ( n189 , n957 );
buf ( n190 , n958 );
buf ( n191 , n959 );
buf ( n192 , n960 );
buf ( n193 , n961 );
buf ( n194 , n962 );
buf ( n195 , n963 );
buf ( n196 , n964 );
buf ( n197 , n965 );
buf ( n198 , n966 );
buf ( n199 , n967 );
buf ( n200 , n968 );
buf ( n201 , n969 );
buf ( n202 , n970 );
buf ( n203 , n971 );
buf ( n204 , n972 );
buf ( n205 , n973 );
buf ( n206 , n974 );
buf ( n207 , n975 );
buf ( n208 , n976 );
buf ( n209 , n977 );
buf ( n210 , n978 );
buf ( n211 , n979 );
buf ( n212 , n980 );
buf ( n213 , n981 );
buf ( n214 , n982 );
buf ( n215 , n983 );
buf ( n216 , n984 );
buf ( n217 , n985 );
buf ( n218 , n986 );
buf ( n219 , n987 );
buf ( n220 , n988 );
buf ( n221 , n989 );
buf ( n222 , n990 );
buf ( n223 , n991 );
buf ( n224 , n992 );
buf ( n225 , n993 );
buf ( n226 , n994 );
buf ( n227 , n995 );
buf ( n228 , n996 );
buf ( n229 , n997 );
buf ( n230 , n998 );
buf ( n231 , n999 );
buf ( n232 , n1000 );
buf ( n233 , n1001 );
buf ( n234 , n1002 );
buf ( n235 , n1003 );
buf ( n236 , n1004 );
buf ( n237 , n1005 );
buf ( n238 , n1006 );
buf ( n239 , n1007 );
buf ( n240 , n1008 );
buf ( n241 , n1009 );
buf ( n242 , n1010 );
buf ( n243 , n1011 );
buf ( n244 , n1012 );
buf ( n245 , n1013 );
buf ( n246 , n1014 );
buf ( n247 , n1015 );
buf ( n248 , n1016 );
buf ( n249 , n1017 );
buf ( n250 , n1018 );
buf ( n251 , n1019 );
buf ( n252 , n1020 );
buf ( n253 , n1021 );
buf ( n254 , n1022 );
buf ( n255 , n1023 );
buf ( n256 , n1024 );
buf ( n257 , n1025 );
buf ( n258 , n1026 );
buf ( n259 , n1027 );
buf ( n260 , n1028 );
buf ( n261 , n1029 );
buf ( n262 , n1030 );
buf ( n263 , n1031 );
buf ( n264 , n1032 );
buf ( n265 , n1033 );
buf ( n266 , n1034 );
buf ( n267 , n1035 );
buf ( n268 , n1036 );
buf ( n269 , n1037 );
buf ( n270 , n1038 );
buf ( n271 , n1039 );
buf ( n272 , n1040 );
buf ( n273 , n1041 );
buf ( n274 , n1042 );
buf ( n275 , n1043 );
buf ( n276 , n1044 );
buf ( n277 , n1045 );
buf ( n278 , n1046 );
buf ( n279 , n1047 );
buf ( n280 , n1048 );
buf ( n281 , n1049 );
buf ( n282 , n1050 );
buf ( n283 , n1051 );
buf ( n284 , n1052 );
buf ( n285 , n1053 );
buf ( n286 , n1054 );
buf ( n287 , n1055 );
buf ( n288 , n1056 );
buf ( n289 , n1057 );
buf ( n290 , n1058 );
buf ( n291 , n1059 );
buf ( n292 , n1060 );
buf ( n293 , n1061 );
buf ( n294 , n1062 );
buf ( n295 , n1063 );
buf ( n296 , n1064 );
buf ( n297 , n1065 );
buf ( n298 , n1066 );
buf ( n299 , n1067 );
buf ( n300 , n1068 );
buf ( n301 , n1069 );
buf ( n302 , n1070 );
buf ( n303 , n1071 );
buf ( n304 , n1072 );
buf ( n305 , n1073 );
buf ( n306 , n1074 );
buf ( n307 , n1075 );
buf ( n308 , n1076 );
buf ( n309 , n1077 );
buf ( n310 , n1078 );
buf ( n311 , n1079 );
buf ( n312 , n1080 );
buf ( n313 , n1081 );
buf ( n314 , n1082 );
buf ( n315 , n1083 );
buf ( n316 , n1084 );
buf ( n317 , n1085 );
buf ( n318 , n1086 );
buf ( n319 , n1087 );
buf ( n320 , n1088 );
buf ( n321 , n1089 );
buf ( n322 , n1090 );
buf ( n323 , n1091 );
buf ( n324 , n1092 );
buf ( n325 , n1093 );
buf ( n326 , n1094 );
buf ( n327 , n1095 );
buf ( n328 , n1096 );
buf ( n329 , n1097 );
buf ( n330 , n1098 );
buf ( n331 , n1099 );
buf ( n332 , n1100 );
buf ( n333 , n1101 );
buf ( n334 , n1102 );
buf ( n335 , n1103 );
buf ( n336 , n1104 );
buf ( n337 , n1105 );
buf ( n338 , n1106 );
buf ( n339 , n1107 );
buf ( n340 , n1108 );
buf ( n341 , n1109 );
buf ( n342 , n1110 );
buf ( n343 , n1111 );
buf ( n344 , n1112 );
buf ( n345 , n1113 );
buf ( n346 , n1114 );
buf ( n347 , n1115 );
buf ( n348 , n1116 );
buf ( n349 , n1117 );
buf ( n350 , n1118 );
buf ( n351 , n1119 );
buf ( n352 , n1120 );
buf ( n353 , n1121 );
buf ( n354 , n1122 );
buf ( n355 , n1123 );
buf ( n356 , n1124 );
buf ( n357 , n1125 );
buf ( n358 , n1126 );
buf ( n359 , n1127 );
buf ( n360 , n1128 );
buf ( n361 , n1129 );
buf ( n362 , n1130 );
buf ( n363 , n1131 );
buf ( n364 , n1132 );
buf ( n365 , n1133 );
buf ( n366 , n1134 );
buf ( n367 , n1135 );
buf ( n368 , n1136 );
buf ( n369 , n1137 );
buf ( n370 , n1138 );
buf ( n371 , n1139 );
buf ( n372 , n1140 );
buf ( n373 , n1141 );
buf ( n374 , n1142 );
buf ( n375 , n1143 );
buf ( n376 , n1144 );
buf ( n377 , n1145 );
buf ( n378 , n1146 );
buf ( n379 , n1147 );
buf ( n380 , n1148 );
buf ( n381 , n1149 );
buf ( n382 , n1150 );
buf ( n383 , n1151 );
buf ( n896 , n209979 );
buf ( n897 , n209983 );
buf ( n898 , n250076 );
buf ( n899 , n209987 );
buf ( n900 , n209999 );
buf ( n901 , n210005 );
buf ( n902 , n210393 );
buf ( n903 , n210032 );
buf ( n904 , n210020 );
buf ( n905 , n210379 );
buf ( n906 , n210384 );
buf ( n907 , n210385 );
buf ( n908 , n210386 );
buf ( n909 , n210382 );
buf ( n910 , n210383 );
buf ( n911 , n210116 );
buf ( n912 , n210387 );
buf ( n913 , n210388 );
buf ( n914 , n210389 );
buf ( n915 , n210122 );
buf ( n916 , n210391 );
buf ( n917 , n210392 );
buf ( n918 , n250148 );
buf ( n919 , n210141 );
buf ( n920 , n210381 );
buf ( n921 , n210110 );
buf ( n922 , n210104 );
buf ( n923 , n210147 );
buf ( n924 , n210380 );
buf ( n925 , n210135 );
buf ( n926 , n210156 );
buf ( n927 , n210173 );
buf ( n928 , n210167 );
buf ( n929 , n250279 );
buf ( n930 , n210185 );
buf ( n931 , n210201 );
buf ( n932 , n210390 );
buf ( n933 , n249932 );
buf ( n934 , n210208 );
buf ( n935 , n210239 );
buf ( n936 , n250191 );
buf ( n937 , n249936 );
buf ( n938 , n210233 );
buf ( n939 , n250205 );
buf ( n940 , n210220 );
buf ( n941 , n210245 );
buf ( n942 , n210254 );
buf ( n943 , n210260 );
buf ( n944 , n210272 );
buf ( n945 , n210278 );
buf ( n946 , n210286 );
buf ( n947 , n210304 );
buf ( n948 , n210298 );
buf ( n949 , n210310 );
buf ( n950 , n210318 );
buf ( n951 , n210324 );
buf ( n952 , n210326 );
buf ( n953 , n210332 );
buf ( n954 , n210338 );
buf ( n955 , n210344 );
buf ( n956 , n250242 );
buf ( n957 , n210350 );
buf ( n958 , n210357 );
buf ( n959 , n250273 );
buf ( n960 , n250256 );
buf ( n961 , n212114 );
buf ( n962 , n250225 );
buf ( n963 , n212990 );
buf ( n964 , n212146 );
buf ( n965 , n212901 );
buf ( n966 , n250162 );
buf ( n967 , n212994 );
buf ( n968 , n250215 );
buf ( n969 , n212998 );
buf ( n970 , n213002 );
buf ( n971 , n213014 );
buf ( n972 , n213018 );
buf ( n973 , n213022 );
buf ( n974 , n213026 );
buf ( n975 , n213030 );
buf ( n976 , n212962 );
buf ( n977 , n212986 );
buf ( n978 , n212966 );
buf ( n979 , n212914 );
buf ( n980 , n212918 );
buf ( n981 , n250120 );
buf ( n982 , n212978 );
buf ( n983 , n250285 );
buf ( n984 , n212922 );
buf ( n985 , n212958 );
buf ( n986 , n212974 );
buf ( n987 , n212934 );
buf ( n988 , n250172 );
buf ( n989 , n212938 );
buf ( n990 , n212942 );
buf ( n991 , n212406 );
buf ( n992 , n212982 );
buf ( n993 , n212910 );
buf ( n994 , n250199 );
buf ( n995 , n212946 );
buf ( n996 , n212926 );
buf ( n997 , n212970 );
buf ( n998 , n213034 );
buf ( n999 , n212450 );
buf ( n1000 , n213010 );
buf ( n1001 , n212954 );
buf ( n1002 , n212930 );
buf ( n1003 , n212505 );
buf ( n1004 , n250100 );
buf ( n1005 , n212476 );
buf ( n1006 , n212525 );
buf ( n1007 , n212566 );
buf ( n1008 , n212551 );
buf ( n1009 , n212580 );
buf ( n1010 , n212599 );
buf ( n1011 , n212642 );
buf ( n1012 , n212628 );
buf ( n1013 , n212656 );
buf ( n1014 , n212682 );
buf ( n1015 , n212696 );
buf ( n1016 , n212699 );
buf ( n1017 , n212702 );
buf ( n1018 , n212705 );
buf ( n1019 , n212708 );
buf ( n1020 , n212711 );
buf ( n1021 , n212726 );
buf ( n1022 , n212748 );
buf ( n1023 , n250284 );
buf ( n1024 , n249984 );
buf ( n1025 , n249339 );
buf ( n1026 , n249362 );
buf ( n1027 , n249027 );
buf ( n1028 , n248773 );
buf ( n1029 , n250004 );
buf ( n1030 , n250083 );
buf ( n1031 , n249384 );
buf ( n1032 , n250050 );
buf ( n1033 , n248855 );
buf ( n1034 , n249192 );
buf ( n1035 , n249050 );
buf ( n1036 , n249168 );
buf ( n1037 , n249970 );
buf ( n1038 , n248894 );
buf ( n1039 , n249182 );
buf ( n1040 , n248926 );
buf ( n1041 , n249131 );
buf ( n1042 , n249147 );
buf ( n1043 , n248937 );
buf ( n1044 , n249116 );
buf ( n1045 , n248905 );
buf ( n1046 , n250272 );
buf ( n1047 , n248788 );
buf ( n1048 , n249921 );
buf ( n1049 , n249096 );
buf ( n1050 , n249938 );
buf ( n1051 , n250299 );
buf ( n1052 , n248955 );
buf ( n1053 , n248967 );
buf ( n1054 , n249937 );
buf ( n1055 , n249083 );
buf ( n1056 , n249069 );
buf ( n1057 , n250014 );
buf ( n1058 , n249211 );
buf ( n1059 , n249223 );
buf ( n1060 , n249234 );
buf ( n1061 , n249454 );
buf ( n1062 , n248818 );
buf ( n1063 , n249240 );
buf ( n1064 , n248987 );
buf ( n1065 , n249250 );
buf ( n1066 , n249001 );
buf ( n1067 , n249260 );
buf ( n1068 , n249448 );
buf ( n1069 , n249279 );
buf ( n1070 , n249886 );
buf ( n1071 , n249442 );
buf ( n1072 , n249480 );
buf ( n1073 , n249429 );
buf ( n1074 , n250266 );
buf ( n1075 , n249306 );
buf ( n1076 , n249409 );
buf ( n1077 , n250252 );
buf ( n1078 , n249943 );
buf ( n1079 , n249487 );
buf ( n1080 , n249403 );
buf ( n1081 , n249944 );
buf ( n1082 , n249518 );
buf ( n1083 , n249524 );
buf ( n1084 , n249505 );
buf ( n1085 , n249530 );
buf ( n1086 , n249474 );
buf ( n1087 , n249536 );
buf ( n1088 , n249549 );
buf ( n1089 , n250089 );
buf ( n1090 , n249566 );
buf ( n1091 , n249589 );
buf ( n1092 , n249583 );
buf ( n1093 , n250071 );
buf ( n1094 , n249603 );
buf ( n1095 , n250029 );
buf ( n1096 , n249618 );
buf ( n1097 , n249637 );
buf ( n1098 , n249630 );
buf ( n1099 , n249645 );
buf ( n1100 , n250034 );
buf ( n1101 , n249880 );
buf ( n1102 , n249659 );
buf ( n1103 , n249673 );
buf ( n1104 , n250039 );
buf ( n1105 , n250114 );
buf ( n1106 , n249883 );
buf ( n1107 , n249884 );
buf ( n1108 , n249686 );
buf ( n1109 , n250180 );
buf ( n1110 , n249887 );
buf ( n1111 , n250061 );
buf ( n1112 , n250154 );
buf ( n1113 , n250132 );
buf ( n1114 , n249891 );
buf ( n1115 , n249892 );
buf ( n1116 , n250141 );
buf ( n1117 , n249893 );
buf ( n1118 , n249895 );
buf ( n1119 , n249896 );
buf ( n1120 , n249897 );
buf ( n1121 , n249903 );
buf ( n1122 , n250280 );
buf ( n1123 , n249909 );
buf ( n1124 , n250019 );
buf ( n1125 , n249912 );
buf ( n1126 , n250236 );
buf ( n1127 , n249913 );
buf ( n1128 , n249920 );
buf ( n1129 , n249923 );
buf ( n1130 , n249925 );
buf ( n1131 , n249924 );
buf ( n1132 , n249888 );
buf ( n1133 , n249748 );
buf ( n1134 , n250108 );
buf ( n1135 , n249767 );
buf ( n1136 , n249778 );
buf ( n1137 , n249791 );
buf ( n1138 , n249945 );
buf ( n1139 , n249812 );
buf ( n1140 , n249822 );
buf ( n1141 , n249829 );
buf ( n1142 , n249838 );
buf ( n1143 , n249847 );
buf ( n1144 , n249853 );
buf ( n1145 , n249855 );
buf ( n1146 , n249857 );
buf ( n1147 , n249864 );
buf ( n1148 , n249866 );
buf ( n1149 , n249868 );
buf ( n1150 , n249870 );
buf ( n1151 , n248193 );
not ( n168462 , n831 );
not ( n168463 , n168462 );
buf ( n168464 , n799 );
not ( n168465 , n168464 );
buf ( n168466 , n168465 );
buf ( n168467 , n168466 );
not ( n168468 , n168467 );
not ( n168469 , n831 );
nand ( n168470 , n168469 , n830 );
not ( n168471 , n168470 );
buf ( n168472 , n168471 );
not ( n168473 , n168472 );
or ( n168474 , n168468 , n168473 );
buf ( n168475 , n798 );
buf ( n168476 , n830 );
xor ( n168477 , n168475 , n168476 );
buf ( n168478 , n168477 );
buf ( n168479 , n168478 );
buf ( n168480 , n831 );
nand ( n168481 , n168479 , n168480 );
buf ( n168482 , n168481 );
buf ( n168483 , n168482 );
nand ( n168484 , n168474 , n168483 );
buf ( n168485 , n168484 );
not ( n168486 , n168485 );
buf ( n168487 , n799 );
buf ( n168488 , n831 );
nand ( n168489 , n168487 , n168488 );
buf ( n168490 , n168489 );
buf ( n168491 , n168490 );
not ( n168492 , n168491 );
buf ( n168493 , n168492 );
and ( n168494 , n168493 , n895 );
buf ( n168495 , n894 );
buf ( n168496 , n168490 );
buf ( n168497 , n830 );
and ( n168498 , n168496 , n168497 );
buf ( n168499 , n168498 );
buf ( n168500 , n168499 );
xor ( n168501 , n168495 , n168500 );
buf ( n168502 , n168501 );
not ( n168503 , n168502 );
and ( n168504 , n168494 , n168503 );
not ( n168505 , n168494 );
and ( n168506 , n168505 , n168502 );
nor ( n168507 , n168504 , n168506 );
xor ( n168508 , n168486 , n168507 );
not ( n168509 , n168508 );
or ( n168510 , n168463 , n168509 );
nand ( n168511 , n168493 , n863 );
buf ( n168512 , n862 );
buf ( n168513 , n168499 );
xor ( n168514 , n168512 , n168513 );
buf ( n168515 , n168514 );
buf ( n168516 , n168515 );
not ( n168517 , n168516 );
buf ( n168518 , n168517 );
xor ( n168519 , n168511 , n168518 );
xor ( n168520 , n168519 , n168485 );
nand ( n168521 , n168520 , n831 );
nand ( n168522 , n168510 , n168521 );
buf ( n168523 , n168522 );
buf ( n168524 , n832 );
buf ( n168525 , n801 );
buf ( n168526 , n802 );
xor ( n168527 , n168525 , n168526 );
buf ( n168528 , n168527 );
buf ( n168529 , n168528 );
buf ( n168530 , n799 );
and ( n168531 , n168529 , n168530 );
buf ( n168532 , n168531 );
buf ( n168533 , n168532 );
buf ( n168534 , n772 );
buf ( n168535 , n828 );
xor ( n168536 , n168534 , n168535 );
buf ( n168537 , n168536 );
buf ( n168538 , n168537 );
not ( n168539 , n168538 );
buf ( n168540 , n829 );
buf ( n168541 , n830 );
xnor ( n168542 , n168540 , n168541 );
buf ( n168543 , n168542 );
buf ( n168544 , n828 );
buf ( n168545 , n829 );
xor ( n168546 , n168544 , n168545 );
buf ( n168547 , n168546 );
nand ( n168548 , n168543 , n168547 );
not ( n168549 , n168548 );
buf ( n168550 , n168549 );
not ( n168551 , n168550 );
or ( n168552 , n168539 , n168551 );
buf ( n168553 , n829 );
buf ( n168554 , n830 );
xor ( n168555 , n168553 , n168554 );
buf ( n168556 , n168555 );
buf ( n168557 , n168556 );
buf ( n168558 , n168557 );
buf ( n168559 , n168558 );
buf ( n168560 , n168559 );
buf ( n168561 , n771 );
buf ( n168562 , n828 );
xor ( n168563 , n168561 , n168562 );
buf ( n168564 , n168563 );
buf ( n168565 , n168564 );
nand ( n168566 , n168560 , n168565 );
buf ( n168567 , n168566 );
buf ( n168568 , n168567 );
nand ( n168569 , n168552 , n168568 );
buf ( n168570 , n168569 );
buf ( n168571 , n168570 );
xor ( n168572 , n168533 , n168571 );
buf ( n168573 , n770 );
buf ( n168574 , n830 );
xor ( n168575 , n168573 , n168574 );
buf ( n168576 , n168575 );
buf ( n168577 , n168576 );
not ( n168578 , n168577 );
buf ( n168579 , n168471 );
not ( n168580 , n168579 );
or ( n168581 , n168578 , n168580 );
buf ( n168582 , n769 );
buf ( n168583 , n830 );
xor ( n168584 , n168582 , n168583 );
buf ( n168585 , n168584 );
buf ( n168586 , n168585 );
buf ( n168587 , n831 );
nand ( n168588 , n168586 , n168587 );
buf ( n168589 , n168588 );
buf ( n168590 , n168589 );
nand ( n168591 , n168581 , n168590 );
buf ( n168592 , n168591 );
buf ( n168593 , n168592 );
xor ( n168594 , n168572 , n168593 );
buf ( n168595 , n168594 );
buf ( n168596 , n168595 );
buf ( n168597 , n792 );
buf ( n168598 , n808 );
xor ( n168599 , n168597 , n168598 );
buf ( n168600 , n168599 );
buf ( n168601 , n168600 );
not ( n168602 , n168601 );
buf ( n168603 , n809 );
buf ( n168604 , n810 );
xor ( n168605 , n168603 , n168604 );
buf ( n168606 , n168605 );
not ( n168607 , n168606 );
buf ( n168608 , n168607 );
xor ( n168609 , n809 , n808 );
buf ( n168610 , n168609 );
nand ( n168611 , n168608 , n168610 );
buf ( n168612 , n168611 );
buf ( n168613 , n168612 );
not ( n168614 , n168613 );
buf ( n168615 , n168614 );
buf ( n168616 , n168615 );
not ( n168617 , n168616 );
or ( n168618 , n168602 , n168617 );
buf ( n168619 , n168606 );
buf ( n168620 , n168619 );
buf ( n168621 , n791 );
buf ( n168622 , n808 );
xor ( n168623 , n168621 , n168622 );
buf ( n168624 , n168623 );
buf ( n168625 , n168624 );
nand ( n168626 , n168620 , n168625 );
buf ( n168627 , n168626 );
buf ( n168628 , n168627 );
nand ( n168629 , n168618 , n168628 );
buf ( n168630 , n168629 );
not ( n168631 , n780 );
and ( n168632 , n820 , n168631 );
not ( n168633 , n820 );
and ( n168634 , n168633 , n780 );
or ( n168635 , n168632 , n168634 );
not ( n168636 , n168635 );
buf ( n168637 , n821 );
not ( n168638 , n168637 );
buf ( n168639 , n822 );
nand ( n168640 , n168638 , n168639 );
buf ( n168641 , n168640 );
xor ( n168642 , n821 , n820 );
buf ( n168643 , n822 );
not ( n168644 , n168643 );
buf ( n168645 , n821 );
nand ( n168646 , n168644 , n168645 );
buf ( n168647 , n168646 );
and ( n168648 , n168641 , n168642 , n168647 );
not ( n168649 , n168648 );
or ( n168650 , n168636 , n168649 );
buf ( n168651 , n779 );
buf ( n168652 , n820 );
xor ( n168653 , n168651 , n168652 );
buf ( n168654 , n168653 );
xor ( n168655 , n821 , n822 );
buf ( n168656 , n168655 );
nand ( n168657 , n168654 , n168656 );
nand ( n168658 , n168650 , n168657 );
xor ( n168659 , n168630 , n168658 );
not ( n168660 , n826 );
nand ( n168661 , n168660 , n827 );
not ( n168662 , n827 );
nand ( n168663 , n168662 , n826 );
nand ( n168664 , n168661 , n168663 );
xnor ( n168665 , n828 , n827 );
and ( n168666 , n168664 , n168665 );
not ( n168667 , n168666 );
buf ( n168668 , n168667 );
buf ( n168669 , n774 );
buf ( n168670 , n826 );
xor ( n168671 , n168669 , n168670 );
buf ( n168672 , n168671 );
buf ( n168673 , n168672 );
not ( n168674 , n168673 );
buf ( n168675 , n168674 );
buf ( n168676 , n168675 );
or ( n168677 , n168668 , n168676 );
buf ( n168678 , n827 );
buf ( n168679 , n828 );
xor ( n168680 , n168678 , n168679 );
buf ( n168681 , n168680 );
buf ( n168682 , n168681 );
buf ( n168683 , n168682 );
buf ( n168684 , n168683 );
buf ( n168685 , n168684 );
xor ( n1217 , n826 , n773 );
buf ( n168687 , n1217 );
nand ( n1219 , n168685 , n168687 );
buf ( n168689 , n1219 );
buf ( n168690 , n168689 );
nand ( n1222 , n168677 , n168690 );
buf ( n168692 , n1222 );
xor ( n1224 , n168659 , n168692 );
buf ( n168694 , n1224 );
xor ( n1226 , n168596 , n168694 );
buf ( n168696 , n794 );
buf ( n168697 , n806 );
xor ( n1229 , n168696 , n168697 );
buf ( n168699 , n1229 );
buf ( n168700 , n168699 );
not ( n1232 , n168700 );
xor ( n1233 , n807 , n808 );
not ( n1234 , n1233 );
buf ( n168704 , n1234 );
and ( n1236 , n806 , n807 );
nor ( n1237 , n806 , n807 );
nor ( n1238 , n1236 , n1237 );
buf ( n168708 , n1238 );
nand ( n1240 , n168704 , n168708 );
buf ( n168710 , n1240 );
buf ( n168711 , n168710 );
not ( n1243 , n168711 );
buf ( n168713 , n1243 );
buf ( n168714 , n168713 );
not ( n1246 , n168714 );
or ( n1247 , n1232 , n1246 );
buf ( n168717 , n1234 );
not ( n1249 , n168717 );
buf ( n168719 , n1249 );
buf ( n168720 , n168719 );
buf ( n168721 , n793 );
buf ( n168722 , n806 );
xor ( n1254 , n168721 , n168722 );
buf ( n168724 , n1254 );
buf ( n168725 , n168724 );
nand ( n1257 , n168720 , n168725 );
buf ( n168727 , n1257 );
buf ( n168728 , n168727 );
nand ( n1260 , n1247 , n168728 );
buf ( n168730 , n1260 );
not ( n1262 , n168730 );
not ( n1263 , n1262 );
buf ( n168733 , n796 );
buf ( n168734 , n804 );
xor ( n1266 , n168733 , n168734 );
buf ( n168736 , n1266 );
buf ( n168737 , n168736 );
not ( n1269 , n168737 );
xnor ( n1270 , n804 , n805 );
buf ( n168740 , n805 );
buf ( n168741 , n806 );
xor ( n1273 , n168740 , n168741 );
buf ( n168743 , n1273 );
nor ( n1275 , n1270 , n168743 );
buf ( n168745 , n1275 );
not ( n1277 , n168745 );
buf ( n168747 , n1277 );
buf ( n168748 , n168747 );
not ( n1280 , n168748 );
buf ( n168750 , n1280 );
buf ( n168751 , n168750 );
not ( n1283 , n168751 );
or ( n1284 , n1269 , n1283 );
buf ( n168754 , n168743 );
not ( n1286 , n168754 );
buf ( n168756 , n1286 );
buf ( n168757 , n168756 );
not ( n1289 , n168757 );
buf ( n168759 , n1289 );
buf ( n168760 , n168759 );
buf ( n168761 , n795 );
buf ( n168762 , n804 );
xor ( n1294 , n168761 , n168762 );
buf ( n168764 , n1294 );
buf ( n168765 , n168764 );
nand ( n1297 , n168760 , n168765 );
buf ( n168767 , n1297 );
buf ( n168768 , n168767 );
nand ( n1300 , n1284 , n168768 );
buf ( n168770 , n1300 );
not ( n1302 , n168770 );
or ( n1303 , n1263 , n1302 );
not ( n1304 , n168770 );
nand ( n1305 , n1304 , n168730 );
nand ( n1306 , n1303 , n1305 );
buf ( n168776 , n782 );
buf ( n168777 , n818 );
xor ( n1309 , n168776 , n168777 );
buf ( n168779 , n1309 );
buf ( n168780 , n168779 );
not ( n1312 , n168780 );
or ( n1313 , n818 , n819 );
nand ( n1314 , n818 , n819 );
nand ( n1315 , n1313 , n1314 );
buf ( n168785 , n819 );
buf ( n168786 , n820 );
xor ( n1318 , n168785 , n168786 );
buf ( n168788 , n1318 );
nor ( n1320 , n1315 , n168788 );
buf ( n1321 , n1320 );
buf ( n168791 , n1321 );
not ( n1323 , n168791 );
buf ( n168793 , n1323 );
buf ( n168794 , n168793 );
not ( n1326 , n168794 );
buf ( n168796 , n1326 );
buf ( n168797 , n168796 );
not ( n1329 , n168797 );
or ( n1330 , n1312 , n1329 );
buf ( n168800 , n819 );
buf ( n168801 , n820 );
xor ( n1333 , n168800 , n168801 );
buf ( n168803 , n1333 );
buf ( n168804 , n168803 );
buf ( n1336 , n168804 );
buf ( n168806 , n1336 );
buf ( n168807 , n168806 );
xor ( n1339 , n818 , n781 );
buf ( n168809 , n1339 );
nand ( n1341 , n168807 , n168809 );
buf ( n168811 , n1341 );
buf ( n168812 , n168811 );
nand ( n1344 , n1330 , n168812 );
buf ( n168814 , n1344 );
and ( n1346 , n1306 , n168814 );
not ( n1347 , n1306 );
not ( n1348 , n168814 );
and ( n1349 , n1347 , n1348 );
nor ( n1350 , n1346 , n1349 );
buf ( n168820 , n1350 );
xor ( n1352 , n1226 , n168820 );
buf ( n168822 , n1352 );
buf ( n168823 , n168822 );
buf ( n168824 , n797 );
buf ( n168825 , n804 );
xor ( n1357 , n168824 , n168825 );
buf ( n168827 , n1357 );
buf ( n168828 , n168827 );
not ( n1360 , n168828 );
buf ( n168830 , n168747 );
not ( n1362 , n168830 );
buf ( n168832 , n1362 );
buf ( n168833 , n168832 );
not ( n1365 , n168833 );
or ( n1366 , n1360 , n1365 );
buf ( n168836 , n168756 );
not ( n1368 , n168836 );
buf ( n168838 , n1368 );
buf ( n168839 , n168838 );
buf ( n168840 , n168736 );
nand ( n1372 , n168839 , n168840 );
buf ( n168842 , n1372 );
buf ( n168843 , n168842 );
nand ( n1375 , n1366 , n168843 );
buf ( n168845 , n1375 );
buf ( n168846 , n168845 );
buf ( n168847 , n799 );
buf ( n168848 , n802 );
xor ( n1380 , n168847 , n168848 );
buf ( n168850 , n1380 );
buf ( n168851 , n168850 );
not ( n1383 , n168851 );
xnor ( n1384 , n802 , n803 );
buf ( n168854 , n803 );
buf ( n168855 , n804 );
xor ( n1387 , n168854 , n168855 );
buf ( n168857 , n1387 );
nor ( n1389 , n1384 , n168857 );
buf ( n168859 , n1389 );
buf ( n1391 , n168859 );
buf ( n168861 , n1391 );
buf ( n168862 , n168861 );
not ( n1394 , n168862 );
or ( n1395 , n1383 , n1394 );
buf ( n168865 , n168857 );
buf ( n1397 , n168865 );
buf ( n168867 , n1397 );
buf ( n168868 , n168867 );
buf ( n1400 , n168868 );
buf ( n168870 , n1400 );
buf ( n168871 , n168870 );
buf ( n168872 , n798 );
buf ( n168873 , n802 );
xor ( n1405 , n168872 , n168873 );
buf ( n168875 , n1405 );
buf ( n168876 , n168875 );
nand ( n1408 , n168871 , n168876 );
buf ( n168878 , n1408 );
buf ( n168879 , n168878 );
nand ( n1411 , n1395 , n168879 );
buf ( n168881 , n1411 );
buf ( n168882 , n168881 );
and ( n1414 , n168846 , n168882 );
not ( n1415 , n168846 );
buf ( n168885 , n168881 );
not ( n1417 , n168885 );
buf ( n168887 , n1417 );
buf ( n168888 , n168887 );
and ( n1420 , n1415 , n168888 );
nor ( n1421 , n1414 , n1420 );
buf ( n168891 , n1421 );
buf ( n168892 , n168891 );
buf ( n168893 , n771 );
buf ( n168894 , n830 );
xor ( n1426 , n168893 , n168894 );
buf ( n168896 , n1426 );
not ( n1428 , n168896 );
not ( n1429 , n168471 );
or ( n1430 , n1428 , n1429 );
buf ( n168900 , n168576 );
buf ( n168901 , n831 );
nand ( n1433 , n168900 , n168901 );
buf ( n168903 , n1433 );
nand ( n1435 , n1430 , n168903 );
buf ( n168905 , n799 );
buf ( n168906 , n803 );
or ( n1438 , n168905 , n168906 );
buf ( n168908 , n804 );
nand ( n1440 , n1438 , n168908 );
buf ( n168910 , n1440 );
buf ( n168911 , n168910 );
buf ( n168912 , n799 );
buf ( n168913 , n803 );
nand ( n1445 , n168912 , n168913 );
buf ( n168915 , n1445 );
buf ( n168916 , n168915 );
buf ( n168917 , n802 );
nand ( n1449 , n168911 , n168916 , n168917 );
buf ( n168919 , n1449 );
buf ( n168920 , n168919 );
not ( n1452 , n168920 );
buf ( n168922 , n1452 );
and ( n1454 , n1435 , n168922 );
not ( n1455 , n1435 );
and ( n1456 , n1455 , n168919 );
nor ( n1457 , n1454 , n1456 );
buf ( n1458 , n1457 );
buf ( n168928 , n1458 );
xor ( n1460 , n168892 , n168928 );
buf ( n168930 , n1460 );
buf ( n168931 , n168930 );
not ( n1463 , n168931 );
buf ( n168933 , n772 );
buf ( n168934 , n830 );
xor ( n1466 , n168933 , n168934 );
buf ( n168936 , n1466 );
buf ( n168937 , n168936 );
not ( n1469 , n168937 );
nand ( n1470 , n168469 , n830 );
not ( n1471 , n1470 );
buf ( n168941 , n1471 );
not ( n1473 , n168941 );
or ( n1474 , n1469 , n1473 );
buf ( n168944 , n168896 );
buf ( n168945 , n831 );
nand ( n1477 , n168944 , n168945 );
buf ( n168947 , n1477 );
buf ( n168948 , n168947 );
nand ( n1480 , n1474 , n168948 );
buf ( n168950 , n1480 );
buf ( n168951 , n792 );
buf ( n168952 , n810 );
xor ( n1484 , n168951 , n168952 );
buf ( n168954 , n1484 );
buf ( n168955 , n168954 );
not ( n1487 , n168955 );
not ( n1488 , n810 );
nand ( n1489 , n1488 , n811 );
not ( n1490 , n1489 );
buf ( n168960 , n811 );
not ( n1492 , n168960 );
buf ( n168962 , n810 );
nand ( n1494 , n1492 , n168962 );
buf ( n168964 , n1494 );
not ( n1496 , n168964 );
or ( n1497 , n1490 , n1496 );
buf ( n168967 , n811 );
buf ( n168968 , n812 );
xor ( n1500 , n168967 , n168968 );
buf ( n168970 , n1500 );
buf ( n168971 , n168970 );
not ( n1503 , n168971 );
buf ( n168973 , n1503 );
nand ( n1505 , n1497 , n168973 );
buf ( n168975 , n1505 );
buf ( n1507 , n168975 );
buf ( n168977 , n1507 );
buf ( n168978 , n168977 );
not ( n1510 , n168978 );
buf ( n168980 , n1510 );
buf ( n168981 , n168980 );
not ( n1513 , n168981 );
or ( n1514 , n1487 , n1513 );
buf ( n168984 , n168973 );
buf ( n1516 , n168984 );
buf ( n168986 , n1516 );
buf ( n168987 , n168986 );
not ( n1519 , n168987 );
buf ( n168989 , n1519 );
buf ( n168990 , n168989 );
buf ( n168991 , n791 );
buf ( n168992 , n810 );
xor ( n1524 , n168991 , n168992 );
buf ( n168994 , n1524 );
buf ( n168995 , n168994 );
nand ( n1527 , n168990 , n168995 );
buf ( n168997 , n1527 );
buf ( n168998 , n168997 );
nand ( n1530 , n1514 , n168998 );
buf ( n169000 , n1530 );
xor ( n1532 , n168950 , n169000 );
xor ( n1533 , n813 , n814 );
buf ( n1534 , n1533 );
buf ( n1535 , n1534 );
not ( n1536 , n1535 );
buf ( n169006 , n789 );
buf ( n169007 , n812 );
xor ( n1539 , n169006 , n169007 );
buf ( n169009 , n1539 );
buf ( n169010 , n169009 );
not ( n1542 , n169010 );
buf ( n169012 , n1542 );
or ( n1544 , n1536 , n169012 );
not ( n1545 , n812 );
not ( n1546 , n1545 );
nand ( n1547 , n813 , n814 );
not ( n1548 , n1547 );
not ( n1549 , n1548 );
or ( n1550 , n1546 , n1549 );
nor ( n1551 , n813 , n814 );
nand ( n1552 , n1551 , n812 );
nand ( n1553 , n1550 , n1552 );
not ( n1554 , n1553 );
not ( n1555 , n1554 );
buf ( n169025 , n790 );
buf ( n169026 , n812 );
xor ( n1558 , n169025 , n169026 );
buf ( n169028 , n1558 );
nand ( n1560 , n1555 , n169028 );
nand ( n1561 , n1544 , n1560 );
xor ( n1562 , n1532 , n1561 );
buf ( n169032 , n1562 );
not ( n1564 , n169032 );
buf ( n169034 , n798 );
buf ( n169035 , n804 );
xor ( n1567 , n169034 , n169035 );
buf ( n169037 , n1567 );
buf ( n169038 , n169037 );
not ( n1570 , n169038 );
xor ( n1571 , n806 , n805 );
and ( n1572 , n804 , n805 );
not ( n1573 , n804 );
not ( n1574 , n805 );
and ( n1575 , n1573 , n1574 );
nor ( n1576 , n1572 , n1575 );
not ( n1577 , n1576 );
nor ( n1578 , n1571 , n1577 );
buf ( n169048 , n1578 );
not ( n1580 , n169048 );
or ( n1581 , n1570 , n1580 );
buf ( n169051 , n168759 );
buf ( n169052 , n168827 );
nand ( n1584 , n169051 , n169052 );
buf ( n169054 , n1584 );
buf ( n169055 , n169054 );
nand ( n1587 , n1581 , n169055 );
buf ( n169057 , n1587 );
buf ( n169058 , n784 );
buf ( n169059 , n818 );
xor ( n1591 , n169058 , n169059 );
buf ( n169061 , n1591 );
buf ( n169062 , n169061 );
not ( n1594 , n169062 );
buf ( n169064 , n1321 );
not ( n1596 , n169064 );
or ( n1597 , n1594 , n1596 );
buf ( n169067 , n168806 );
buf ( n169068 , n783 );
buf ( n169069 , n818 );
xor ( n1601 , n169068 , n169069 );
buf ( n169071 , n1601 );
buf ( n169072 , n169071 );
nand ( n1604 , n169067 , n169072 );
buf ( n169074 , n1604 );
buf ( n169075 , n169074 );
nand ( n1607 , n1597 , n169075 );
buf ( n169077 , n1607 );
xor ( n1609 , n169057 , n169077 );
buf ( n169079 , n168681 );
buf ( n1611 , n169079 );
buf ( n169081 , n1611 );
not ( n1613 , n169081 );
xor ( n1614 , n826 , n775 );
not ( n1615 , n1614 );
or ( n1616 , n1613 , n1615 );
not ( n1617 , n168663 );
not ( n1618 , n168661 );
or ( n1619 , n1617 , n1618 );
nand ( n1620 , n1619 , n168665 );
not ( n1621 , n1620 );
buf ( n169091 , n1621 );
not ( n1623 , n169091 );
buf ( n169093 , n1623 );
buf ( n169094 , n776 );
buf ( n169095 , n826 );
xnor ( n1627 , n169094 , n169095 );
buf ( n169097 , n1627 );
or ( n1629 , n169093 , n169097 );
nand ( n1630 , n1616 , n1629 );
xor ( n1631 , n1609 , n1630 );
buf ( n169101 , n1631 );
not ( n1633 , n169101 );
or ( n1634 , n1564 , n1633 );
not ( n1635 , n1631 );
not ( n1636 , n1635 );
not ( n1637 , n1562 );
not ( n1638 , n1637 );
or ( n1639 , n1636 , n1638 );
buf ( n169109 , n168867 );
buf ( n169110 , n799 );
and ( n1642 , n169109 , n169110 );
buf ( n169112 , n1642 );
buf ( n169113 , n168549 );
buf ( n169114 , n774 );
buf ( n169115 , n828 );
xor ( n1647 , n169114 , n169115 );
buf ( n169117 , n1647 );
buf ( n169118 , n169117 );
and ( n1650 , n169113 , n169118 );
buf ( n169120 , n168559 );
buf ( n169121 , n773 );
buf ( n169122 , n828 );
xor ( n1654 , n169121 , n169122 );
buf ( n169124 , n1654 );
buf ( n169125 , n169124 );
and ( n1657 , n169120 , n169125 );
nor ( n1658 , n1650 , n1657 );
buf ( n169128 , n1658 );
not ( n1660 , n169128 );
xor ( n1661 , n169112 , n1660 );
buf ( n169131 , n778 );
buf ( n169132 , n824 );
xor ( n1664 , n169131 , n169132 );
buf ( n169134 , n1664 );
buf ( n169135 , n169134 );
not ( n1667 , n169135 );
and ( n1668 , n825 , n824 );
not ( n1669 , n825 );
not ( n1670 , n824 );
and ( n1671 , n1669 , n1670 );
nor ( n1672 , n1668 , n1671 );
not ( n1673 , n826 );
and ( n1674 , n825 , n1673 );
not ( n1675 , n825 );
and ( n1676 , n1675 , n826 );
nor ( n1677 , n1674 , n1676 );
nand ( n1678 , n1672 , n1677 );
not ( n1679 , n1678 );
buf ( n169149 , n1679 );
not ( n1681 , n169149 );
buf ( n169151 , n1681 );
buf ( n169152 , n169151 );
not ( n1684 , n169152 );
buf ( n169154 , n1684 );
buf ( n169155 , n169154 );
not ( n1687 , n169155 );
or ( n1688 , n1667 , n1687 );
buf ( n169158 , n777 );
buf ( n169159 , n824 );
xor ( n1691 , n169158 , n169159 );
buf ( n169161 , n1691 );
buf ( n169162 , n169161 );
buf ( n169163 , n825 );
buf ( n169164 , n826 );
xnor ( n1696 , n169163 , n169164 );
buf ( n169166 , n1696 );
buf ( n169167 , n169166 );
not ( n1699 , n169167 );
buf ( n169169 , n1699 );
buf ( n169170 , n169169 );
nand ( n1702 , n169162 , n169170 );
buf ( n169172 , n1702 );
buf ( n169173 , n169172 );
nand ( n1705 , n1688 , n169173 );
buf ( n169175 , n1705 );
xnor ( n1707 , n1661 , n169175 );
not ( n1708 , n1707 );
nand ( n1709 , n1639 , n1708 );
buf ( n169179 , n1709 );
nand ( n1711 , n1634 , n169179 );
buf ( n169181 , n1711 );
buf ( n169182 , n169181 );
not ( n1714 , n169182 );
or ( n1715 , n1463 , n1714 );
buf ( n169185 , n169181 );
buf ( n169186 , n168930 );
or ( n1718 , n169185 , n169186 );
buf ( n169188 , n799 );
buf ( n169189 , n805 );
or ( n1721 , n169188 , n169189 );
buf ( n169191 , n806 );
nand ( n1723 , n1721 , n169191 );
buf ( n169193 , n1723 );
buf ( n169194 , n169193 );
buf ( n169195 , n799 );
buf ( n169196 , n805 );
nand ( n1728 , n169195 , n169196 );
buf ( n169198 , n1728 );
buf ( n169199 , n169198 );
buf ( n169200 , n804 );
and ( n1732 , n169194 , n169199 , n169200 );
buf ( n169202 , n1732 );
buf ( n169203 , n169202 );
buf ( n169204 , n775 );
buf ( n169205 , n828 );
xor ( n1737 , n169204 , n169205 );
buf ( n169207 , n1737 );
buf ( n169208 , n169207 );
not ( n1740 , n169208 );
nand ( n1741 , n168543 , n168547 );
not ( n1742 , n1741 );
buf ( n169212 , n1742 );
not ( n1744 , n169212 );
or ( n1745 , n1740 , n1744 );
buf ( n169215 , n168559 );
buf ( n169216 , n169117 );
nand ( n1748 , n169215 , n169216 );
buf ( n169218 , n1748 );
buf ( n169219 , n169218 );
nand ( n1751 , n1745 , n169219 );
buf ( n169221 , n1751 );
buf ( n169222 , n169221 );
nand ( n1754 , n169203 , n169222 );
buf ( n169224 , n1754 );
buf ( n169225 , n169224 );
not ( n1757 , n169225 );
buf ( n169227 , n1757 );
buf ( n169228 , n169227 );
not ( n1760 , n169228 );
buf ( n169230 , n789 );
buf ( n169231 , n814 );
xor ( n1763 , n169230 , n169231 );
buf ( n169233 , n1763 );
buf ( n169234 , n169233 );
not ( n1766 , n169234 );
xnor ( n1767 , n814 , n815 );
xor ( n1768 , n815 , n816 );
nor ( n1769 , n1767 , n1768 );
buf ( n169239 , n1769 );
buf ( n1771 , n169239 );
buf ( n169241 , n1771 );
buf ( n169242 , n169241 );
not ( n1774 , n169242 );
or ( n1775 , n1766 , n1774 );
buf ( n169245 , n1768 );
buf ( n1777 , n169245 );
buf ( n169247 , n1777 );
buf ( n169248 , n169247 );
buf ( n1780 , n169248 );
buf ( n169250 , n1780 );
buf ( n169251 , n169250 );
buf ( n169252 , n788 );
buf ( n169253 , n814 );
xor ( n1785 , n169252 , n169253 );
buf ( n169255 , n1785 );
buf ( n169256 , n169255 );
nand ( n1788 , n169251 , n169256 );
buf ( n169258 , n1788 );
buf ( n169259 , n169258 );
nand ( n1791 , n1775 , n169259 );
buf ( n169261 , n1791 );
buf ( n169262 , n169261 );
not ( n1794 , n169262 );
buf ( n169264 , n779 );
buf ( n169265 , n824 );
xor ( n1797 , n169264 , n169265 );
buf ( n169267 , n1797 );
buf ( n169268 , n169267 );
not ( n1800 , n169268 );
and ( n1801 , n825 , n1673 );
not ( n1802 , n825 );
and ( n1803 , n1802 , n826 );
nor ( n1804 , n1801 , n1803 );
nand ( n1805 , n1804 , n1672 );
not ( n1806 , n1805 );
buf ( n169276 , n1806 );
not ( n1808 , n169276 );
or ( n1809 , n1800 , n1808 );
buf ( n169279 , n169134 );
buf ( n169280 , n169169 );
nand ( n1812 , n169279 , n169280 );
buf ( n169282 , n1812 );
buf ( n169283 , n169282 );
nand ( n1815 , n1809 , n169283 );
buf ( n169285 , n1815 );
buf ( n169286 , n169285 );
not ( n1818 , n169286 );
or ( n1819 , n1794 , n1818 );
buf ( n169289 , n169261 );
not ( n1821 , n169289 );
buf ( n169291 , n1821 );
buf ( n169292 , n169291 );
not ( n1824 , n169292 );
buf ( n169294 , n169285 );
not ( n1826 , n169294 );
buf ( n169296 , n1826 );
buf ( n169297 , n169296 );
not ( n1829 , n169297 );
or ( n1830 , n1824 , n1829 );
buf ( n169300 , n787 );
buf ( n169301 , n816 );
xor ( n1833 , n169300 , n169301 );
buf ( n169303 , n1833 );
buf ( n169304 , n169303 );
not ( n1836 , n169304 );
xnor ( n1837 , n817 , n816 );
buf ( n169307 , n817 );
buf ( n169308 , n818 );
xor ( n1840 , n169307 , n169308 );
buf ( n169310 , n1840 );
nor ( n1842 , n1837 , n169310 );
buf ( n169312 , n1842 );
buf ( n1844 , n169312 );
buf ( n169314 , n1844 );
buf ( n169315 , n169314 );
not ( n1847 , n169315 );
or ( n1848 , n1836 , n1847 );
buf ( n169318 , n169310 );
buf ( n1850 , n169318 );
buf ( n169320 , n1850 );
buf ( n169321 , n169320 );
buf ( n169322 , n786 );
buf ( n169323 , n816 );
xor ( n1855 , n169322 , n169323 );
buf ( n169325 , n1855 );
buf ( n169326 , n169325 );
nand ( n1858 , n169321 , n169326 );
buf ( n169328 , n1858 );
buf ( n169329 , n169328 );
nand ( n1861 , n1848 , n169329 );
buf ( n169331 , n1861 );
buf ( n169332 , n169331 );
nand ( n1864 , n1830 , n169332 );
buf ( n169334 , n1864 );
buf ( n169335 , n169334 );
nand ( n1867 , n1819 , n169335 );
buf ( n169337 , n1867 );
buf ( n169338 , n169337 );
not ( n1870 , n169338 );
or ( n1871 , n1760 , n1870 );
buf ( n169341 , n169224 );
not ( n1873 , n169341 );
buf ( n169343 , n169337 );
not ( n1875 , n169343 );
buf ( n169345 , n1875 );
buf ( n169346 , n169345 );
not ( n1878 , n169346 );
or ( n1879 , n1873 , n1878 );
buf ( n169349 , n793 );
buf ( n169350 , n810 );
xor ( n1882 , n169349 , n169350 );
buf ( n169352 , n1882 );
buf ( n169353 , n169352 );
not ( n1885 , n169353 );
buf ( n169355 , n168980 );
not ( n1887 , n169355 );
or ( n1888 , n1885 , n1887 );
buf ( n169358 , n168989 );
buf ( n169359 , n168954 );
nand ( n1891 , n169358 , n169359 );
buf ( n169361 , n1891 );
buf ( n169362 , n169361 );
nand ( n1894 , n1888 , n169362 );
buf ( n169364 , n1894 );
buf ( n169365 , n169364 );
buf ( n169366 , n791 );
buf ( n169367 , n812 );
xor ( n1899 , n169366 , n169367 );
buf ( n169369 , n1899 );
buf ( n169370 , n169369 );
not ( n1902 , n169370 );
not ( n1903 , n1545 );
not ( n1904 , n1548 );
or ( n1905 , n1903 , n1904 );
nand ( n1906 , n1905 , n1552 );
buf ( n1907 , n1906 );
buf ( n169377 , n1907 );
not ( n1909 , n169377 );
or ( n1910 , n1902 , n1909 );
buf ( n169380 , n1535 );
buf ( n169381 , n169028 );
nand ( n1913 , n169380 , n169381 );
buf ( n169383 , n1913 );
buf ( n169384 , n169383 );
nand ( n1916 , n1910 , n169384 );
buf ( n169386 , n1916 );
buf ( n169387 , n169386 );
xor ( n1919 , n169365 , n169387 );
buf ( n169389 , n781 );
buf ( n169390 , n822 );
xor ( n1922 , n169389 , n169390 );
buf ( n169392 , n1922 );
buf ( n169393 , n169392 );
not ( n1925 , n169393 );
and ( n1926 , n823 , n822 );
not ( n1927 , n823 );
not ( n1928 , n822 );
and ( n1929 , n1927 , n1928 );
nor ( n1930 , n1926 , n1929 );
buf ( n169400 , n1930 );
not ( n1932 , n169400 );
buf ( n169402 , n1932 );
buf ( n169403 , n823 );
buf ( n169404 , n824 );
xor ( n1936 , n169403 , n169404 );
buf ( n169406 , n1936 );
nor ( n1938 , n169402 , n169406 );
buf ( n1939 , n1938 );
buf ( n169409 , n1939 );
buf ( n1941 , n169409 );
buf ( n169411 , n1941 );
buf ( n169412 , n169411 );
not ( n1944 , n169412 );
or ( n1945 , n1925 , n1944 );
buf ( n169415 , n169406 );
buf ( n1947 , n169415 );
buf ( n169417 , n1947 );
buf ( n169418 , n169417 );
not ( n1950 , n169418 );
buf ( n169420 , n1950 );
buf ( n169421 , n169420 );
not ( n1953 , n169421 );
buf ( n169423 , n1953 );
buf ( n169424 , n169423 );
buf ( n169425 , n780 );
buf ( n169426 , n822 );
xor ( n1958 , n169425 , n169426 );
buf ( n169428 , n1958 );
buf ( n169429 , n169428 );
nand ( n1961 , n169424 , n169429 );
buf ( n169431 , n1961 );
buf ( n169432 , n169431 );
nand ( n1964 , n1945 , n169432 );
buf ( n169434 , n1964 );
buf ( n169435 , n169434 );
and ( n1967 , n1919 , n169435 );
and ( n1968 , n169365 , n169387 );
or ( n1969 , n1967 , n1968 );
buf ( n169439 , n1969 );
buf ( n169440 , n169439 );
nand ( n1972 , n1879 , n169440 );
buf ( n169442 , n1972 );
buf ( n169443 , n169442 );
nand ( n1975 , n1871 , n169443 );
buf ( n169445 , n1975 );
buf ( n169446 , n169445 );
nand ( n1978 , n1718 , n169446 );
buf ( n169448 , n1978 );
buf ( n169449 , n169448 );
nand ( n1981 , n1715 , n169449 );
buf ( n169451 , n1981 );
buf ( n169452 , n169451 );
xor ( n1984 , n168823 , n169452 );
not ( n1985 , n169175 );
not ( n1986 , n169112 );
or ( n1987 , n1985 , n1986 );
buf ( n1988 , n169128 );
buf ( n169458 , n169175 );
buf ( n169459 , n169112 );
nor ( n1991 , n169458 , n169459 );
buf ( n169461 , n1991 );
or ( n1993 , n1988 , n169461 );
nand ( n1994 , n1987 , n1993 );
xor ( n1995 , n168950 , n169000 );
and ( n1996 , n1995 , n1561 );
and ( n1997 , n168950 , n169000 );
or ( n1998 , n1996 , n1997 );
xor ( n1999 , n1994 , n1998 );
not ( n2000 , n169428 );
not ( n2001 , n169411 );
or ( n2002 , n2000 , n2001 );
buf ( n169472 , n169423 );
buf ( n169473 , n779 );
buf ( n169474 , n822 );
xor ( n2006 , n169473 , n169474 );
buf ( n169476 , n2006 );
buf ( n169477 , n169476 );
nand ( n2009 , n169472 , n169477 );
buf ( n169479 , n2009 );
nand ( n2011 , n2002 , n169479 );
not ( n2012 , n169255 );
not ( n2013 , n169241 );
or ( n2014 , n2012 , n2013 );
buf ( n169484 , n169250 );
buf ( n169485 , n787 );
buf ( n169486 , n814 );
xor ( n2018 , n169485 , n169486 );
buf ( n169488 , n2018 );
buf ( n169489 , n169488 );
nand ( n2021 , n169484 , n169489 );
buf ( n169491 , n2021 );
nand ( n2023 , n2014 , n169491 );
buf ( n2024 , n2023 );
nand ( n2025 , n2011 , n2024 );
or ( n2026 , n2024 , n2011 );
buf ( n169496 , n169325 );
not ( n2028 , n169496 );
buf ( n169498 , n169314 );
not ( n2030 , n169498 );
or ( n2031 , n2028 , n2030 );
buf ( n169501 , n169320 );
buf ( n169502 , n785 );
buf ( n169503 , n816 );
xor ( n2035 , n169502 , n169503 );
buf ( n169505 , n2035 );
buf ( n169506 , n169505 );
nand ( n2038 , n169501 , n169506 );
buf ( n169508 , n2038 );
buf ( n169509 , n169508 );
nand ( n2041 , n2031 , n169509 );
buf ( n169511 , n2041 );
nand ( n2043 , n2026 , n169511 );
nand ( n2044 , n2025 , n2043 );
xor ( n2045 , n1999 , n2044 );
buf ( n169515 , n2045 );
not ( n2047 , n831 );
and ( n2048 , n2047 , n830 );
not ( n2049 , n2048 );
buf ( n169519 , n773 );
buf ( n169520 , n830 );
xor ( n2052 , n169519 , n169520 );
buf ( n169522 , n2052 );
not ( n2054 , n169522 );
or ( n2055 , n2049 , n2054 );
buf ( n169525 , n168936 );
buf ( n169526 , n831 );
nand ( n2058 , n169525 , n169526 );
buf ( n169528 , n2058 );
nand ( n2060 , n2055 , n169528 );
not ( n2061 , n2060 );
buf ( n169531 , n2061 );
not ( n2063 , n169531 );
buf ( n169533 , n795 );
buf ( n169534 , n808 );
xor ( n2066 , n169533 , n169534 );
buf ( n169536 , n2066 );
buf ( n169537 , n169536 );
not ( n2069 , n169537 );
buf ( n169539 , n168607 );
buf ( n169540 , n168609 );
nand ( n2072 , n169539 , n169540 );
buf ( n169542 , n2072 );
buf ( n169543 , n169542 );
not ( n2075 , n169543 );
buf ( n169545 , n2075 );
buf ( n169546 , n169545 );
not ( n2078 , n169546 );
or ( n2079 , n2069 , n2078 );
buf ( n169549 , n794 );
buf ( n169550 , n808 );
xor ( n2082 , n169549 , n169550 );
buf ( n169552 , n2082 );
buf ( n169553 , n169552 );
buf ( n169554 , n168619 );
nand ( n2086 , n169553 , n169554 );
buf ( n169556 , n2086 );
buf ( n169557 , n169556 );
nand ( n2089 , n2079 , n169557 );
buf ( n169559 , n2089 );
not ( n2091 , n169559 );
buf ( n169561 , n2091 );
not ( n2093 , n169561 );
or ( n2094 , n2063 , n2093 );
buf ( n169564 , n783 );
buf ( n169565 , n820 );
xor ( n2097 , n169564 , n169565 );
buf ( n169567 , n2097 );
buf ( n169568 , n169567 );
not ( n2100 , n169568 );
not ( n2101 , n820 );
nor ( n2102 , n821 , n822 );
not ( n2103 , n2102 );
or ( n2104 , n2101 , n2103 );
not ( n2105 , n820 );
nand ( n2106 , n2105 , n821 , n822 );
nand ( n2107 , n2104 , n2106 );
buf ( n2108 , n2107 );
buf ( n169578 , n2108 );
not ( n2110 , n169578 );
or ( n2111 , n2100 , n2110 );
buf ( n169581 , n168656 );
buf ( n169582 , n782 );
buf ( n169583 , n820 );
xor ( n2115 , n169582 , n169583 );
buf ( n169585 , n2115 );
buf ( n169586 , n169585 );
nand ( n2118 , n169581 , n169586 );
buf ( n169588 , n2118 );
buf ( n169589 , n169588 );
nand ( n2121 , n2111 , n169589 );
buf ( n169591 , n2121 );
buf ( n169592 , n169591 );
nand ( n2124 , n2094 , n169592 );
buf ( n169594 , n2124 );
buf ( n169595 , n169594 );
buf ( n169596 , n2061 );
not ( n2128 , n169596 );
buf ( n169598 , n169559 );
nand ( n2130 , n2128 , n169598 );
buf ( n169600 , n2130 );
buf ( n169601 , n169600 );
nand ( n2133 , n169595 , n169601 );
buf ( n169603 , n2133 );
buf ( n169604 , n169603 );
buf ( n169605 , n799 );
buf ( n169606 , n804 );
xor ( n2138 , n169605 , n169606 );
buf ( n169608 , n2138 );
buf ( n169609 , n169608 );
not ( n2141 , n169609 );
buf ( n169611 , n168832 );
not ( n2143 , n169611 );
or ( n2144 , n2141 , n2143 );
buf ( n169614 , n168838 );
buf ( n169615 , n169037 );
nand ( n2147 , n169614 , n169615 );
buf ( n169617 , n2147 );
buf ( n169618 , n169617 );
nand ( n2150 , n2144 , n169618 );
buf ( n169620 , n2150 );
buf ( n169621 , n169620 );
not ( n2153 , n169621 );
buf ( n169623 , n797 );
buf ( n169624 , n806 );
xor ( n2156 , n169623 , n169624 );
buf ( n169626 , n2156 );
buf ( n169627 , n169626 );
not ( n2159 , n169627 );
buf ( n169629 , n1234 );
buf ( n169630 , n1238 );
nand ( n2162 , n169629 , n169630 );
buf ( n169632 , n2162 );
buf ( n169633 , n169632 );
not ( n2165 , n169633 );
buf ( n169635 , n2165 );
buf ( n169636 , n169635 );
not ( n2168 , n169636 );
or ( n2169 , n2159 , n2168 );
buf ( n169639 , n1234 );
not ( n2171 , n169639 );
buf ( n169641 , n2171 );
buf ( n169642 , n169641 );
buf ( n169643 , n796 );
buf ( n169644 , n806 );
xor ( n2176 , n169643 , n169644 );
buf ( n169646 , n2176 );
buf ( n169647 , n169646 );
nand ( n2179 , n169642 , n169647 );
buf ( n169649 , n2179 );
buf ( n169650 , n169649 );
nand ( n2182 , n2169 , n169650 );
buf ( n169652 , n2182 );
buf ( n169653 , n169652 );
not ( n2185 , n169653 );
or ( n2186 , n2153 , n2185 );
buf ( n169656 , n169620 );
not ( n2188 , n169656 );
buf ( n169658 , n2188 );
buf ( n169659 , n169658 );
not ( n2191 , n169659 );
buf ( n169661 , n169652 );
not ( n2193 , n169661 );
buf ( n169663 , n2193 );
buf ( n169664 , n169663 );
not ( n2196 , n169664 );
or ( n2197 , n2191 , n2196 );
not ( n2198 , n168661 );
not ( n2199 , n168663 );
or ( n2200 , n2198 , n2199 );
xnor ( n2201 , n828 , n827 );
nand ( n2202 , n2200 , n2201 );
buf ( n169672 , n2202 );
not ( n2204 , n169672 );
buf ( n169674 , n2204 );
not ( n2206 , n169674 );
xor ( n2207 , n777 , n826 );
not ( n2208 , n2207 );
or ( n2209 , n2206 , n2208 );
buf ( n169679 , n168684 );
not ( n2211 , n169679 );
buf ( n169681 , n2211 );
or ( n2213 , n169097 , n169681 );
nand ( n2214 , n2209 , n2213 );
buf ( n169684 , n2214 );
nand ( n2216 , n2197 , n169684 );
buf ( n169686 , n2216 );
buf ( n169687 , n169686 );
nand ( n2219 , n2186 , n169687 );
buf ( n169689 , n2219 );
buf ( n169690 , n169689 );
xor ( n2222 , n169604 , n169690 );
buf ( n169692 , n2011 );
not ( n2224 , n169692 );
not ( n2225 , n2023 );
buf ( n169695 , n2225 );
not ( n2227 , n169695 );
buf ( n169697 , n169511 );
not ( n2229 , n169697 );
and ( n2230 , n2227 , n2229 );
buf ( n169700 , n169511 );
buf ( n169701 , n2225 );
and ( n2233 , n169700 , n169701 );
nor ( n2234 , n2230 , n2233 );
buf ( n169704 , n2234 );
buf ( n169705 , n169704 );
not ( n2237 , n169705 );
or ( n2238 , n2224 , n2237 );
buf ( n169708 , n169704 );
buf ( n169709 , n2011 );
or ( n2241 , n169708 , n169709 );
nand ( n2242 , n2238 , n2241 );
buf ( n169712 , n2242 );
buf ( n169713 , n169712 );
and ( n2245 , n2222 , n169713 );
and ( n2246 , n169604 , n169690 );
or ( n2247 , n2245 , n2246 );
buf ( n169717 , n2247 );
buf ( n169718 , n169717 );
xor ( n2250 , n169515 , n169718 );
buf ( n2251 , n2107 );
not ( n2252 , n2251 );
not ( n2253 , n169585 );
or ( n2254 , n2252 , n2253 );
buf ( n169724 , n168655 );
buf ( n169725 , n781 );
buf ( n169726 , n820 );
xor ( n2258 , n169725 , n169726 );
buf ( n169728 , n2258 );
buf ( n169729 , n169728 );
nand ( n2261 , n169724 , n169729 );
buf ( n169731 , n2261 );
nand ( n2263 , n2254 , n169731 );
buf ( n169733 , n2263 );
buf ( n169734 , n169552 );
not ( n2266 , n169734 );
buf ( n169736 , n169545 );
not ( n2268 , n169736 );
or ( n2269 , n2266 , n2268 );
buf ( n169739 , n168619 );
buf ( n169740 , n793 );
buf ( n169741 , n808 );
xor ( n2273 , n169740 , n169741 );
buf ( n169743 , n2273 );
buf ( n169744 , n169743 );
nand ( n2276 , n169739 , n169744 );
buf ( n169746 , n2276 );
buf ( n169747 , n169746 );
nand ( n2279 , n2269 , n169747 );
buf ( n169749 , n2279 );
buf ( n169750 , n169749 );
or ( n2282 , n169733 , n169750 );
buf ( n169752 , n169646 );
not ( n2284 , n169752 );
buf ( n169754 , n168713 );
not ( n2286 , n169754 );
or ( n2287 , n2284 , n2286 );
buf ( n169757 , n168719 );
buf ( n2289 , n169757 );
buf ( n169759 , n2289 );
buf ( n169760 , n169759 );
buf ( n169761 , n795 );
buf ( n169762 , n806 );
xor ( n2294 , n169761 , n169762 );
buf ( n169764 , n2294 );
buf ( n169765 , n169764 );
nand ( n2297 , n169760 , n169765 );
buf ( n169767 , n2297 );
buf ( n169768 , n169767 );
nand ( n2300 , n2287 , n169768 );
buf ( n169770 , n2300 );
buf ( n169771 , n169770 );
nand ( n2303 , n2282 , n169771 );
buf ( n169773 , n2303 );
buf ( n169774 , n169773 );
buf ( n169775 , n2263 );
buf ( n169776 , n169749 );
nand ( n2308 , n169775 , n169776 );
buf ( n169778 , n2308 );
buf ( n169779 , n169778 );
nand ( n2311 , n169774 , n169779 );
buf ( n169781 , n2311 );
buf ( n169782 , n169781 );
xor ( n2314 , n169057 , n169077 );
and ( n2315 , n2314 , n1630 );
and ( n2316 , n169057 , n169077 );
or ( n2317 , n2315 , n2316 );
buf ( n169787 , n2317 );
xor ( n2319 , n169782 , n169787 );
buf ( n169789 , n169161 );
not ( n2321 , n169789 );
buf ( n169791 , n1679 );
buf ( n2323 , n169791 );
buf ( n169793 , n2323 );
buf ( n169794 , n169793 );
not ( n2326 , n169794 );
or ( n2327 , n2321 , n2326 );
buf ( n169797 , n169166 );
buf ( n2329 , n169797 );
buf ( n169799 , n2329 );
buf ( n169800 , n169799 );
not ( n2332 , n169800 );
buf ( n169802 , n2332 );
buf ( n169803 , n169802 );
buf ( n169804 , n776 );
buf ( n169805 , n824 );
xor ( n2337 , n169804 , n169805 );
buf ( n169807 , n2337 );
buf ( n169808 , n169807 );
nand ( n2340 , n169803 , n169808 );
buf ( n169810 , n2340 );
buf ( n169811 , n169810 );
nand ( n2343 , n2327 , n169811 );
buf ( n169813 , n2343 );
buf ( n169814 , n169813 );
buf ( n169815 , n169124 );
not ( n2347 , n169815 );
buf ( n169817 , n1742 );
not ( n2349 , n169817 );
or ( n2350 , n2347 , n2349 );
buf ( n169820 , n168559 );
buf ( n169821 , n168537 );
nand ( n2353 , n169820 , n169821 );
buf ( n169823 , n2353 );
buf ( n169824 , n169823 );
nand ( n2356 , n2350 , n169824 );
buf ( n169826 , n2356 );
buf ( n169827 , n169826 );
xor ( n2359 , n169814 , n169827 );
buf ( n169829 , n169505 );
not ( n2361 , n169829 );
buf ( n169831 , n1842 );
buf ( n2363 , n169831 );
buf ( n169833 , n2363 );
buf ( n169834 , n169833 );
buf ( n2366 , n169834 );
buf ( n169836 , n2366 );
buf ( n169837 , n169836 );
not ( n2369 , n169837 );
or ( n2370 , n2361 , n2369 );
buf ( n169840 , n169310 );
buf ( n2372 , n169840 );
buf ( n169842 , n2372 );
buf ( n169843 , n169842 );
buf ( n2375 , n169843 );
buf ( n169845 , n2375 );
buf ( n169846 , n169845 );
buf ( n169847 , n784 );
buf ( n169848 , n816 );
xor ( n2380 , n169847 , n169848 );
buf ( n169850 , n2380 );
buf ( n169851 , n169850 );
nand ( n2383 , n169846 , n169851 );
buf ( n169853 , n2383 );
buf ( n169854 , n169853 );
nand ( n2386 , n2370 , n169854 );
buf ( n169856 , n2386 );
buf ( n169857 , n169856 );
xor ( n2389 , n2359 , n169857 );
buf ( n169859 , n2389 );
buf ( n169860 , n169859 );
xor ( n2392 , n2319 , n169860 );
buf ( n169862 , n2392 );
buf ( n169863 , n169862 );
and ( n2395 , n2250 , n169863 );
and ( n2396 , n169515 , n169718 );
or ( n2397 , n2395 , n2396 );
buf ( n169867 , n2397 );
buf ( n169868 , n169867 );
xor ( n2400 , n1984 , n169868 );
buf ( n169870 , n2400 );
buf ( n169871 , n169870 );
xor ( n2403 , n169515 , n169718 );
xor ( n2404 , n2403 , n169863 );
buf ( n169874 , n2404 );
buf ( n169875 , n169874 );
not ( n2407 , n169875 );
xor ( n2408 , n168930 , n169445 );
xnor ( n2409 , n2408 , n169181 );
buf ( n169879 , n2409 );
nand ( n2411 , n2407 , n169879 );
buf ( n169881 , n2411 );
buf ( n169882 , n169881 );
not ( n2414 , n169882 );
buf ( n169884 , n169476 );
not ( n2416 , n169884 );
xnor ( n2417 , n822 , n823 );
nor ( n2418 , n2417 , n169406 );
buf ( n169888 , n2418 );
not ( n2420 , n169888 );
or ( n2421 , n2416 , n2420 );
buf ( n169891 , n169417 );
buf ( n169892 , n778 );
buf ( n169893 , n822 );
xor ( n2425 , n169892 , n169893 );
buf ( n169895 , n2425 );
buf ( n169896 , n169895 );
nand ( n2428 , n169891 , n169896 );
buf ( n169898 , n2428 );
buf ( n169899 , n169898 );
nand ( n2431 , n2421 , n169899 );
buf ( n169901 , n2431 );
buf ( n169902 , n169901 );
buf ( n169903 , n169009 );
not ( n2435 , n169903 );
buf ( n169905 , n1907 );
not ( n2437 , n169905 );
or ( n2438 , n2435 , n2437 );
buf ( n169908 , n1534 );
xor ( n2440 , n812 , n788 );
buf ( n169910 , n2440 );
nand ( n2442 , n169908 , n169910 );
buf ( n169912 , n2442 );
buf ( n169913 , n169912 );
nand ( n2445 , n2438 , n169913 );
buf ( n169915 , n2445 );
buf ( n169916 , n169915 );
xor ( n2448 , n169902 , n169916 );
buf ( n169918 , n169488 );
not ( n2450 , n169918 );
buf ( n169920 , n169241 );
buf ( n2452 , n169920 );
buf ( n169922 , n2452 );
buf ( n169923 , n169922 );
not ( n2455 , n169923 );
or ( n2456 , n2450 , n2455 );
buf ( n169926 , n169247 );
not ( n2458 , n169926 );
buf ( n169928 , n2458 );
buf ( n169929 , n169928 );
not ( n2461 , n169929 );
buf ( n169931 , n2461 );
buf ( n169932 , n169931 );
buf ( n169933 , n786 );
buf ( n169934 , n814 );
xor ( n2466 , n169933 , n169934 );
buf ( n169936 , n2466 );
buf ( n169937 , n169936 );
nand ( n2469 , n169932 , n169937 );
buf ( n169939 , n2469 );
buf ( n169940 , n169939 );
nand ( n2472 , n2456 , n169940 );
buf ( n169942 , n2472 );
buf ( n169943 , n169942 );
xor ( n2475 , n2448 , n169943 );
buf ( n169945 , n2475 );
buf ( n169946 , n169945 );
buf ( n169947 , n168994 );
not ( n2479 , n169947 );
buf ( n169949 , n168977 );
not ( n2481 , n169949 );
buf ( n169951 , n2481 );
buf ( n169952 , n169951 );
not ( n2484 , n169952 );
or ( n2485 , n2479 , n2484 );
buf ( n169955 , n168973 );
not ( n2487 , n169955 );
buf ( n169957 , n2487 );
buf ( n169958 , n169957 );
xor ( n2490 , n810 , n790 );
buf ( n169960 , n2490 );
nand ( n2492 , n169958 , n169960 );
buf ( n169962 , n2492 );
buf ( n169963 , n169962 );
nand ( n2495 , n2485 , n169963 );
buf ( n169965 , n2495 );
buf ( n169966 , n169965 );
buf ( n169967 , n1614 );
not ( n2499 , n169967 );
buf ( n169969 , n1621 );
not ( n2501 , n169969 );
or ( n2502 , n2499 , n2501 );
buf ( n169972 , n169081 );
buf ( n169973 , n168672 );
nand ( n2505 , n169972 , n169973 );
buf ( n169975 , n2505 );
buf ( n169976 , n169975 );
nand ( n2508 , n2502 , n169976 );
buf ( n169978 , n2508 );
buf ( n169979 , n169978 );
xor ( n2511 , n169966 , n169979 );
not ( n2512 , n168655 );
not ( n2513 , n2512 );
not ( n2514 , n2513 );
not ( n2515 , n168635 );
or ( n2516 , n2514 , n2515 );
buf ( n169986 , n2108 );
not ( n2518 , n169986 );
buf ( n169988 , n2518 );
buf ( n169989 , n169988 );
buf ( n2521 , n169989 );
buf ( n169991 , n2521 );
buf ( n169992 , n169728 );
not ( n2524 , n169992 );
buf ( n169994 , n2524 );
or ( n2526 , n169991 , n169994 );
nand ( n2527 , n2516 , n2526 );
buf ( n169997 , n2527 );
xor ( n2529 , n2511 , n169997 );
buf ( n169999 , n2529 );
buf ( n170000 , n169999 );
xor ( n2532 , n169946 , n170000 );
buf ( n170002 , n169764 );
not ( n2534 , n170002 );
buf ( n170004 , n168713 );
not ( n2536 , n170004 );
or ( n2537 , n2534 , n2536 );
buf ( n170007 , n169759 );
buf ( n170008 , n168699 );
nand ( n2540 , n170007 , n170008 );
buf ( n170010 , n2540 );
buf ( n170011 , n170010 );
nand ( n2543 , n2537 , n170011 );
buf ( n170013 , n2543 );
buf ( n170014 , n170013 );
buf ( n170015 , n169743 );
not ( n2547 , n170015 );
buf ( n170017 , n169545 );
buf ( n2549 , n170017 );
buf ( n170019 , n2549 );
buf ( n170020 , n170019 );
not ( n2552 , n170020 );
or ( n2553 , n2547 , n2552 );
buf ( n2554 , n168619 );
buf ( n170024 , n2554 );
buf ( n170025 , n168600 );
nand ( n2557 , n170024 , n170025 );
buf ( n170027 , n2557 );
buf ( n170028 , n170027 );
nand ( n2560 , n2553 , n170028 );
buf ( n170030 , n2560 );
buf ( n170031 , n170030 );
xor ( n2563 , n170014 , n170031 );
buf ( n170033 , n169071 );
not ( n2565 , n170033 );
buf ( n2566 , n1321 );
buf ( n170036 , n2566 );
not ( n2568 , n170036 );
or ( n2569 , n2565 , n2568 );
buf ( n170039 , n168806 );
buf ( n170040 , n168779 );
nand ( n2572 , n170039 , n170040 );
buf ( n170042 , n2572 );
buf ( n170043 , n170042 );
nand ( n2575 , n2569 , n170043 );
buf ( n170045 , n2575 );
buf ( n170046 , n170045 );
xor ( n2578 , n2563 , n170046 );
buf ( n170048 , n2578 );
buf ( n170049 , n170048 );
xor ( n2581 , n2532 , n170049 );
buf ( n170051 , n2581 );
xor ( n2583 , n169749 , n2263 );
xor ( n2584 , n2583 , n169770 );
buf ( n170054 , n2584 );
buf ( n170055 , n785 );
buf ( n170056 , n818 );
xor ( n2588 , n170055 , n170056 );
buf ( n170058 , n2588 );
buf ( n170059 , n170058 );
not ( n2591 , n170059 );
buf ( n170061 , n168796 );
not ( n2593 , n170061 );
or ( n2594 , n2591 , n2593 );
buf ( n170064 , n168806 );
buf ( n170065 , n169061 );
nand ( n2597 , n170064 , n170065 );
buf ( n170067 , n2597 );
buf ( n170068 , n170067 );
nand ( n2600 , n2594 , n170068 );
buf ( n170070 , n2600 );
buf ( n170071 , n170070 );
xor ( n2603 , n169202 , n169221 );
buf ( n170073 , n2603 );
xor ( n2605 , n170071 , n170073 );
buf ( n170075 , n168743 );
buf ( n170076 , n799 );
and ( n2608 , n170075 , n170076 );
buf ( n170078 , n2608 );
buf ( n170079 , n170078 );
buf ( n170080 , n776 );
buf ( n170081 , n828 );
xor ( n2613 , n170080 , n170081 );
buf ( n170083 , n2613 );
buf ( n170084 , n170083 );
not ( n2616 , n170084 );
buf ( n170086 , n1742 );
not ( n2618 , n170086 );
or ( n2619 , n2616 , n2618 );
buf ( n170089 , n168559 );
buf ( n170090 , n169207 );
nand ( n2622 , n170089 , n170090 );
buf ( n170092 , n2622 );
buf ( n170093 , n170092 );
nand ( n2625 , n2619 , n170093 );
buf ( n170095 , n2625 );
buf ( n170096 , n170095 );
xor ( n2628 , n170079 , n170096 );
buf ( n170098 , n1679 );
buf ( n2630 , n170098 );
buf ( n170100 , n2630 );
buf ( n170101 , n170100 );
not ( n2633 , n170101 );
buf ( n170103 , n2633 );
buf ( n170104 , n170103 );
buf ( n170105 , n780 );
buf ( n170106 , n824 );
xor ( n2638 , n170105 , n170106 );
buf ( n170108 , n2638 );
buf ( n170109 , n170108 );
not ( n2641 , n170109 );
buf ( n170111 , n2641 );
buf ( n170112 , n170111 );
or ( n2644 , n170104 , n170112 );
buf ( n170114 , n169799 );
buf ( n170115 , n169267 );
not ( n2647 , n170115 );
buf ( n170117 , n2647 );
buf ( n170118 , n170117 );
or ( n2650 , n170114 , n170118 );
nand ( n2651 , n2644 , n2650 );
buf ( n170121 , n2651 );
buf ( n170122 , n170121 );
and ( n2654 , n2628 , n170122 );
and ( n2655 , n170079 , n170096 );
or ( n2656 , n2654 , n2655 );
buf ( n170126 , n2656 );
buf ( n170127 , n170126 );
and ( n2659 , n2605 , n170127 );
and ( n2660 , n170071 , n170073 );
or ( n2661 , n2659 , n2660 );
buf ( n170131 , n2661 );
buf ( n170132 , n170131 );
xor ( n2664 , n170054 , n170132 );
buf ( n170134 , n790 );
buf ( n170135 , n814 );
xor ( n2667 , n170134 , n170135 );
buf ( n170137 , n2667 );
buf ( n170138 , n170137 );
not ( n2670 , n170138 );
buf ( n170140 , n169241 );
not ( n2672 , n170140 );
or ( n2673 , n2670 , n2672 );
buf ( n170143 , n169247 );
buf ( n170144 , n169233 );
nand ( n2676 , n170143 , n170144 );
buf ( n170146 , n2676 );
buf ( n170147 , n170146 );
nand ( n2679 , n2673 , n170147 );
buf ( n170149 , n2679 );
buf ( n170150 , n788 );
buf ( n170151 , n816 );
xor ( n2683 , n170150 , n170151 );
buf ( n170153 , n2683 );
buf ( n170154 , n170153 );
not ( n2686 , n170154 );
buf ( n170156 , n169833 );
not ( n2688 , n170156 );
or ( n2689 , n2686 , n2688 );
buf ( n170159 , n169842 );
buf ( n170160 , n169303 );
nand ( n2692 , n170159 , n170160 );
buf ( n170162 , n2692 );
buf ( n170163 , n170162 );
nand ( n2695 , n2689 , n170163 );
buf ( n170165 , n2695 );
xor ( n2697 , n170149 , n170165 );
buf ( n170167 , n782 );
buf ( n170168 , n822 );
xor ( n2700 , n170167 , n170168 );
buf ( n170170 , n2700 );
buf ( n170171 , n170170 );
not ( n2703 , n170171 );
buf ( n170173 , n169411 );
not ( n2705 , n170173 );
or ( n2706 , n2703 , n2705 );
buf ( n170176 , n169417 );
buf ( n170177 , n169392 );
nand ( n2709 , n170176 , n170177 );
buf ( n170179 , n2709 );
buf ( n170180 , n170179 );
nand ( n2712 , n2706 , n170180 );
buf ( n170182 , n2712 );
and ( n2714 , n2697 , n170182 );
and ( n2715 , n170149 , n170165 );
or ( n2716 , n2714 , n2715 );
not ( n2717 , n2716 );
not ( n2718 , n2048 );
buf ( n170188 , n774 );
buf ( n170189 , n830 );
xor ( n2721 , n170188 , n170189 );
buf ( n170191 , n2721 );
not ( n2723 , n170191 );
or ( n2724 , n2718 , n2723 );
buf ( n170194 , n169522 );
buf ( n170195 , n831 );
nand ( n2727 , n170194 , n170195 );
buf ( n170197 , n2727 );
nand ( n2729 , n2724 , n170197 );
buf ( n170199 , n2729 );
xor ( n2731 , n810 , n794 );
buf ( n170201 , n2731 );
not ( n2733 , n170201 );
not ( n2734 , n810 );
nand ( n2735 , n2734 , n811 );
nand ( n2736 , n168964 , n2735 );
and ( n2737 , n168973 , n2736 );
buf ( n170207 , n2737 );
not ( n2739 , n170207 );
or ( n2740 , n2733 , n2739 );
buf ( n170210 , n168989 );
buf ( n170211 , n169352 );
nand ( n2743 , n170210 , n170211 );
buf ( n170213 , n2743 );
buf ( n170214 , n170213 );
nand ( n2746 , n2740 , n170214 );
buf ( n170216 , n2746 );
buf ( n170217 , n170216 );
xor ( n2749 , n170199 , n170217 );
buf ( n170219 , n792 );
buf ( n170220 , n812 );
xor ( n2752 , n170219 , n170220 );
buf ( n170222 , n2752 );
buf ( n170223 , n170222 );
not ( n2755 , n170223 );
not ( n2756 , n1906 );
not ( n2757 , n2756 );
buf ( n170227 , n2757 );
not ( n2759 , n170227 );
or ( n2760 , n2755 , n2759 );
buf ( n170230 , n1534 );
buf ( n170231 , n169369 );
nand ( n2763 , n170230 , n170231 );
buf ( n170233 , n2763 );
buf ( n170234 , n170233 );
nand ( n2766 , n2760 , n170234 );
buf ( n170236 , n2766 );
buf ( n170237 , n170236 );
and ( n2769 , n2749 , n170237 );
and ( n2770 , n170199 , n170217 );
or ( n2771 , n2769 , n2770 );
buf ( n170241 , n2771 );
not ( n2773 , n170241 );
buf ( n170243 , n796 );
buf ( n170244 , n808 );
xor ( n2776 , n170243 , n170244 );
buf ( n170246 , n2776 );
buf ( n170247 , n170246 );
not ( n2779 , n170247 );
buf ( n170249 , n169545 );
not ( n2781 , n170249 );
or ( n2782 , n2779 , n2781 );
buf ( n170252 , n168619 );
buf ( n170253 , n169536 );
nand ( n2785 , n170252 , n170253 );
buf ( n170255 , n2785 );
buf ( n170256 , n170255 );
nand ( n2788 , n2782 , n170256 );
buf ( n170258 , n2788 );
buf ( n170259 , n170258 );
not ( n2791 , n170259 );
buf ( n170261 , n784 );
buf ( n170262 , n820 );
xor ( n2794 , n170261 , n170262 );
buf ( n170264 , n2794 );
buf ( n170265 , n170264 );
not ( n2797 , n170265 );
buf ( n170267 , n2251 );
not ( n2799 , n170267 );
or ( n2800 , n2797 , n2799 );
buf ( n170270 , n169567 );
buf ( n170271 , n168656 );
nand ( n2803 , n170270 , n170271 );
buf ( n170273 , n2803 );
buf ( n170274 , n170273 );
nand ( n2806 , n2800 , n170274 );
buf ( n170276 , n2806 );
buf ( n170277 , n170276 );
not ( n2809 , n170277 );
or ( n2810 , n2791 , n2809 );
buf ( n170280 , n170276 );
buf ( n170281 , n170258 );
or ( n2813 , n170280 , n170281 );
buf ( n170283 , n798 );
buf ( n170284 , n806 );
xor ( n2816 , n170283 , n170284 );
buf ( n170286 , n2816 );
buf ( n170287 , n170286 );
not ( n2819 , n170287 );
buf ( n170289 , n168713 );
not ( n2821 , n170289 );
or ( n2822 , n2819 , n2821 );
xor ( n2823 , n807 , n808 );
buf ( n170293 , n2823 );
buf ( n170294 , n169626 );
nand ( n2826 , n170293 , n170294 );
buf ( n170296 , n2826 );
buf ( n170297 , n170296 );
nand ( n2829 , n2822 , n170297 );
buf ( n170299 , n2829 );
buf ( n170300 , n170299 );
nand ( n2832 , n2813 , n170300 );
buf ( n170302 , n2832 );
buf ( n170303 , n170302 );
nand ( n2835 , n2810 , n170303 );
buf ( n170305 , n2835 );
not ( n2837 , n170305 );
nand ( n2838 , n2773 , n2837 );
not ( n2839 , n2838 );
or ( n2840 , n2717 , n2839 );
not ( n2841 , n2837 );
nand ( n2842 , n2841 , n170241 );
nand ( n2843 , n2840 , n2842 );
buf ( n170313 , n2843 );
and ( n2845 , n2664 , n170313 );
and ( n2846 , n170054 , n170132 );
or ( n2847 , n2845 , n2846 );
buf ( n170317 , n2847 );
xor ( n2849 , n170051 , n170317 );
xor ( n2850 , n169604 , n169690 );
xor ( n2851 , n2850 , n169713 );
buf ( n170321 , n2851 );
buf ( n170322 , n170321 );
and ( n2854 , n169337 , n169224 );
not ( n2855 , n169337 );
and ( n2856 , n169221 , n169202 );
and ( n2857 , n2855 , n2856 );
nor ( n2858 , n2854 , n2857 );
xor ( n2859 , n169439 , n2858 );
buf ( n170329 , n2859 );
not ( n2861 , n170329 );
buf ( n170331 , n2861 );
buf ( n170332 , n170331 );
or ( n2864 , n170322 , n170332 );
not ( n2865 , n169591 );
xor ( n2866 , n2061 , n2865 );
xnor ( n2867 , n2866 , n2091 );
buf ( n170337 , n2867 );
not ( n2869 , n170337 );
buf ( n170339 , n169663 );
not ( n2871 , n170339 );
buf ( n170341 , n2214 );
not ( n2873 , n170341 );
or ( n2874 , n2871 , n2873 );
buf ( n170344 , n2214 );
buf ( n170345 , n169663 );
or ( n2877 , n170344 , n170345 );
nand ( n2878 , n2874 , n2877 );
buf ( n170348 , n2878 );
buf ( n170349 , n170348 );
buf ( n170350 , n169658 );
and ( n2882 , n170349 , n170350 );
not ( n2883 , n170349 );
buf ( n170353 , n169620 );
and ( n2885 , n2883 , n170353 );
nor ( n2886 , n2882 , n2885 );
buf ( n170356 , n2886 );
buf ( n170357 , n170356 );
not ( n2889 , n170357 );
buf ( n170359 , n2889 );
buf ( n170360 , n170359 );
not ( n2892 , n170360 );
or ( n2893 , n2869 , n2892 );
not ( n2894 , n170356 );
not ( n2895 , n2867 );
not ( n2896 , n2895 );
or ( n2897 , n2894 , n2896 );
buf ( n170367 , n169331 );
buf ( n170368 , n169285 );
and ( n2900 , n170367 , n170368 );
not ( n2901 , n170367 );
buf ( n170371 , n169296 );
and ( n2903 , n2901 , n170371 );
nor ( n2904 , n2900 , n2903 );
buf ( n170374 , n2904 );
buf ( n170375 , n169261 );
buf ( n2907 , n170375 );
buf ( n170377 , n2907 );
not ( n2909 , n170377 );
and ( n2910 , n170374 , n2909 );
not ( n2911 , n170374 );
and ( n2912 , n2911 , n170377 );
nor ( n2913 , n2910 , n2912 );
not ( n2914 , n2913 );
nand ( n2915 , n2897 , n2914 );
buf ( n170385 , n2915 );
nand ( n2917 , n2893 , n170385 );
buf ( n170387 , n2917 );
buf ( n170388 , n170387 );
nand ( n2920 , n2864 , n170388 );
buf ( n170390 , n2920 );
buf ( n170391 , n170390 );
buf ( n170392 , n170331 );
buf ( n170393 , n170321 );
nand ( n2925 , n170392 , n170393 );
buf ( n170395 , n2925 );
buf ( n170396 , n170395 );
nand ( n2928 , n170391 , n170396 );
buf ( n170398 , n2928 );
xor ( n2930 , n2849 , n170398 );
buf ( n170400 , n2930 );
not ( n2932 , n170400 );
or ( n2933 , n2414 , n2932 );
not ( n2934 , n2409 );
nand ( n2935 , n2934 , n169874 );
buf ( n170405 , n2935 );
nand ( n2937 , n2933 , n170405 );
buf ( n170407 , n2937 );
buf ( n170408 , n170407 );
xor ( n2940 , n169871 , n170408 );
buf ( n170410 , n1435 );
buf ( n170411 , n168922 );
and ( n2943 , n170410 , n170411 );
buf ( n170413 , n2943 );
buf ( n170414 , n170413 );
buf ( n170415 , n168875 );
not ( n2947 , n170415 );
buf ( n170417 , n168861 );
buf ( n2949 , n170417 );
buf ( n170419 , n2949 );
buf ( n170420 , n170419 );
not ( n2952 , n170420 );
or ( n2953 , n2947 , n2952 );
buf ( n170423 , n168870 );
xor ( n2955 , n802 , n797 );
buf ( n170425 , n2955 );
nand ( n2957 , n170423 , n170425 );
buf ( n170427 , n2957 );
buf ( n170428 , n170427 );
nand ( n2960 , n2953 , n170428 );
buf ( n170430 , n2960 );
buf ( n170431 , n170430 );
xor ( n2963 , n170414 , n170431 );
xor ( n2964 , n169814 , n169827 );
and ( n2965 , n2964 , n169857 );
and ( n2966 , n169814 , n169827 );
or ( n2967 , n2965 , n2966 );
buf ( n170437 , n2967 );
buf ( n170438 , n170437 );
xor ( n2970 , n2963 , n170438 );
buf ( n170440 , n2970 );
buf ( n170441 , n170440 );
xor ( n2973 , n1994 , n1998 );
and ( n2974 , n2973 , n2044 );
and ( n2975 , n1994 , n1998 );
or ( n2976 , n2974 , n2975 );
buf ( n170446 , n2976 );
xor ( n2978 , n170441 , n170446 );
xor ( n2979 , n169946 , n170000 );
and ( n2980 , n2979 , n170049 );
and ( n2981 , n169946 , n170000 );
or ( n2982 , n2980 , n2981 );
buf ( n170452 , n2982 );
buf ( n170453 , n170452 );
xor ( n2985 , n2978 , n170453 );
buf ( n170455 , n2985 );
buf ( n170456 , n170455 );
xor ( n2988 , n169782 , n169787 );
and ( n2989 , n2988 , n169860 );
and ( n2990 , n169782 , n169787 );
or ( n2991 , n2989 , n2990 );
buf ( n170461 , n2991 );
buf ( n170462 , n170461 );
xor ( n2994 , n169902 , n169916 );
and ( n2995 , n2994 , n169943 );
and ( n2996 , n169902 , n169916 );
or ( n2997 , n2995 , n2996 );
buf ( n170467 , n2997 );
buf ( n170468 , n170467 );
xor ( n3000 , n169966 , n169979 );
and ( n3001 , n3000 , n169997 );
and ( n3002 , n169966 , n169979 );
or ( n3003 , n3001 , n3002 );
buf ( n170473 , n3003 );
buf ( n170474 , n170473 );
xor ( n3006 , n170468 , n170474 );
xor ( n3007 , n170014 , n170031 );
and ( n3008 , n3007 , n170046 );
and ( n3009 , n170014 , n170031 );
or ( n3010 , n3008 , n3009 );
buf ( n170480 , n3010 );
buf ( n170481 , n170480 );
xor ( n3013 , n3006 , n170481 );
buf ( n170483 , n3013 );
buf ( n170484 , n170483 );
xor ( n3016 , n170462 , n170484 );
not ( n3017 , n1457 );
not ( n3018 , n168845 );
or ( n3019 , n3017 , n3018 );
buf ( n170489 , n1457 );
buf ( n170490 , n168845 );
nor ( n3022 , n170489 , n170490 );
buf ( n170492 , n3022 );
or ( n3024 , n170492 , n168887 );
nand ( n3025 , n3019 , n3024 );
buf ( n170495 , n3025 );
buf ( n170496 , n169895 );
not ( n3028 , n170496 );
buf ( n170498 , n1939 );
not ( n3030 , n170498 );
or ( n3031 , n3028 , n3030 );
buf ( n170501 , n169417 );
xor ( n3033 , n822 , n777 );
buf ( n170503 , n3033 );
nand ( n3035 , n170501 , n170503 );
buf ( n170505 , n3035 );
buf ( n170506 , n170505 );
nand ( n3038 , n3031 , n170506 );
buf ( n170508 , n3038 );
buf ( n170509 , n170508 );
not ( n3041 , n170509 );
buf ( n170511 , n2440 );
not ( n3043 , n170511 );
buf ( n170513 , n1907 );
not ( n3045 , n170513 );
or ( n3046 , n3043 , n3045 );
buf ( n170516 , n1534 );
xor ( n3048 , n812 , n787 );
buf ( n170518 , n3048 );
nand ( n3050 , n170516 , n170518 );
buf ( n170520 , n3050 );
buf ( n170521 , n170520 );
nand ( n3053 , n3046 , n170521 );
buf ( n170523 , n3053 );
buf ( n170524 , n170523 );
not ( n3056 , n170524 );
buf ( n170526 , n3056 );
buf ( n170527 , n170526 );
not ( n3059 , n170527 );
or ( n3060 , n3041 , n3059 );
buf ( n170530 , n170526 );
buf ( n170531 , n170508 );
or ( n3063 , n170530 , n170531 );
nand ( n3064 , n3060 , n3063 );
buf ( n170534 , n3064 );
buf ( n170535 , n170534 );
buf ( n170536 , n2490 );
not ( n3068 , n170536 );
buf ( n170538 , n168980 );
not ( n3070 , n170538 );
or ( n3071 , n3068 , n3070 );
buf ( n170541 , n169957 );
xor ( n3073 , n810 , n789 );
buf ( n170543 , n3073 );
nand ( n3075 , n170541 , n170543 );
buf ( n170545 , n3075 );
buf ( n170546 , n170545 );
nand ( n3078 , n3071 , n170546 );
buf ( n170548 , n3078 );
buf ( n170549 , n170548 );
xor ( n3081 , n170535 , n170549 );
buf ( n170551 , n3081 );
buf ( n170552 , n170551 );
xor ( n3084 , n170495 , n170552 );
buf ( n170554 , n169807 );
not ( n3086 , n170554 );
buf ( n170556 , n1806 );
not ( n3088 , n170556 );
or ( n3089 , n3086 , n3088 );
buf ( n170559 , n825 );
buf ( n170560 , n826 );
xnor ( n3092 , n170559 , n170560 );
buf ( n170562 , n3092 );
buf ( n170563 , n170562 );
not ( n3095 , n170563 );
buf ( n170565 , n3095 );
buf ( n170566 , n170565 );
buf ( n170567 , n775 );
buf ( n170568 , n824 );
xor ( n3100 , n170567 , n170568 );
buf ( n170570 , n3100 );
buf ( n170571 , n170570 );
nand ( n3103 , n170566 , n170571 );
buf ( n170573 , n3103 );
buf ( n170574 , n170573 );
nand ( n3106 , n3089 , n170574 );
buf ( n170576 , n3106 );
buf ( n170577 , n169850 );
not ( n3109 , n170577 );
buf ( n170579 , n169836 );
not ( n3111 , n170579 );
or ( n3112 , n3109 , n3111 );
buf ( n170582 , n169320 );
buf ( n170583 , n783 );
buf ( n170584 , n816 );
xor ( n3116 , n170583 , n170584 );
buf ( n170586 , n3116 );
buf ( n170587 , n170586 );
nand ( n3119 , n170582 , n170587 );
buf ( n170589 , n3119 );
buf ( n170590 , n170589 );
nand ( n3122 , n3112 , n170590 );
buf ( n170592 , n3122 );
xor ( n3124 , n170576 , n170592 );
buf ( n170594 , n169936 );
not ( n3126 , n170594 );
buf ( n170596 , n169922 );
not ( n3128 , n170596 );
or ( n3129 , n3126 , n3128 );
buf ( n170599 , n169931 );
buf ( n170600 , n785 );
buf ( n170601 , n814 );
xor ( n3133 , n170600 , n170601 );
buf ( n170603 , n3133 );
buf ( n170604 , n170603 );
nand ( n3136 , n170599 , n170604 );
buf ( n170606 , n3136 );
buf ( n170607 , n170606 );
nand ( n3139 , n3129 , n170607 );
buf ( n170609 , n3139 );
xor ( n3141 , n3124 , n170609 );
buf ( n170611 , n3141 );
xor ( n3143 , n3084 , n170611 );
buf ( n170613 , n3143 );
buf ( n170614 , n170613 );
xor ( n3146 , n3016 , n170614 );
buf ( n170616 , n3146 );
buf ( n170617 , n170616 );
xor ( n3149 , n170456 , n170617 );
xor ( n3150 , n170051 , n170317 );
and ( n3151 , n3150 , n170398 );
and ( n3152 , n170051 , n170317 );
or ( n3153 , n3151 , n3152 );
buf ( n170623 , n3153 );
xor ( n3155 , n3149 , n170623 );
buf ( n170625 , n3155 );
buf ( n170626 , n170625 );
and ( n3158 , n2940 , n170626 );
and ( n3159 , n169871 , n170408 );
or ( n3160 , n3158 , n3159 );
buf ( n170630 , n3160 );
buf ( n170631 , n170630 );
xor ( n3163 , n168524 , n170631 );
buf ( n170633 , n168624 );
not ( n3165 , n170633 );
buf ( n170635 , n169545 );
not ( n3167 , n170635 );
or ( n3168 , n3165 , n3167 );
buf ( n170638 , n790 );
buf ( n170639 , n808 );
xor ( n3171 , n170638 , n170639 );
buf ( n170641 , n3171 );
buf ( n170642 , n170641 );
buf ( n170643 , n168619 );
nand ( n3175 , n170642 , n170643 );
buf ( n170645 , n3175 );
buf ( n170646 , n170645 );
nand ( n3178 , n3168 , n170646 );
buf ( n170648 , n3178 );
buf ( n170649 , n170648 );
buf ( n170650 , n168724 );
not ( n3182 , n170650 );
buf ( n170652 , n168713 );
not ( n3184 , n170652 );
or ( n3185 , n3182 , n3184 );
buf ( n170655 , n169759 );
buf ( n170656 , n792 );
buf ( n170657 , n806 );
xor ( n3189 , n170656 , n170657 );
buf ( n170659 , n3189 );
buf ( n170660 , n170659 );
nand ( n3192 , n170655 , n170660 );
buf ( n170662 , n3192 );
buf ( n170663 , n170662 );
nand ( n3195 , n3185 , n170663 );
buf ( n170665 , n3195 );
buf ( n170666 , n170665 );
xor ( n3198 , n170649 , n170666 );
not ( n3199 , n2513 );
buf ( n170669 , n778 );
buf ( n170670 , n820 );
xor ( n3202 , n170669 , n170670 );
buf ( n170672 , n3202 );
not ( n3204 , n170672 );
or ( n3205 , n3199 , n3204 );
buf ( n170675 , n168654 );
not ( n3207 , n170675 );
buf ( n170677 , n3207 );
or ( n3209 , n169988 , n170677 );
nand ( n3210 , n3205 , n3209 );
buf ( n170680 , n3210 );
xor ( n3212 , n3198 , n170680 );
buf ( n170682 , n3212 );
buf ( n170683 , n170682 );
buf ( n170684 , n3048 );
not ( n3216 , n170684 );
buf ( n170686 , n2757 );
not ( n3218 , n170686 );
or ( n3219 , n3216 , n3218 );
buf ( n3220 , n1534 );
buf ( n170690 , n3220 );
buf ( n170691 , n786 );
buf ( n170692 , n812 );
xor ( n3224 , n170691 , n170692 );
buf ( n170694 , n3224 );
buf ( n170695 , n170694 );
nand ( n3227 , n170690 , n170695 );
buf ( n170697 , n3227 );
buf ( n170698 , n170697 );
nand ( n3230 , n3219 , n170698 );
buf ( n170700 , n3230 );
buf ( n170701 , n3073 );
not ( n3233 , n170701 );
buf ( n170703 , n169951 );
not ( n3235 , n170703 );
or ( n3236 , n3233 , n3235 );
buf ( n170706 , n168986 );
not ( n3238 , n170706 );
buf ( n170708 , n3238 );
buf ( n170709 , n170708 );
buf ( n170710 , n788 );
buf ( n170711 , n810 );
xor ( n3243 , n170710 , n170711 );
buf ( n170713 , n3243 );
buf ( n170714 , n170713 );
nand ( n3246 , n170709 , n170714 );
buf ( n170716 , n3246 );
buf ( n170717 , n170716 );
nand ( n3249 , n3236 , n170717 );
buf ( n170719 , n3249 );
xor ( n3251 , n170700 , n170719 );
buf ( n170721 , n1217 );
not ( n3253 , n170721 );
buf ( n170723 , n1621 );
not ( n3255 , n170723 );
or ( n3256 , n3253 , n3255 );
buf ( n170726 , n169081 );
buf ( n170727 , n772 );
buf ( n170728 , n826 );
xor ( n3260 , n170727 , n170728 );
buf ( n170730 , n3260 );
buf ( n170731 , n170730 );
nand ( n3263 , n170726 , n170731 );
buf ( n170733 , n3263 );
buf ( n170734 , n170733 );
nand ( n3266 , n3256 , n170734 );
buf ( n170736 , n3266 );
xor ( n3268 , n3251 , n170736 );
buf ( n170738 , n3268 );
xor ( n3270 , n170683 , n170738 );
xor ( n3271 , n170468 , n170474 );
and ( n3272 , n3271 , n170481 );
and ( n3273 , n170468 , n170474 );
or ( n3274 , n3272 , n3273 );
buf ( n170744 , n3274 );
buf ( n170745 , n170744 );
xor ( n3277 , n3270 , n170745 );
buf ( n170747 , n3277 );
buf ( n170748 , n170747 );
xor ( n3280 , n170441 , n170446 );
and ( n3281 , n3280 , n170453 );
and ( n3282 , n170441 , n170446 );
or ( n3283 , n3281 , n3282 );
buf ( n170753 , n3283 );
buf ( n170754 , n170753 );
xor ( n3286 , n170748 , n170754 );
xor ( n3287 , n170462 , n170484 );
and ( n3288 , n3287 , n170614 );
and ( n3289 , n170462 , n170484 );
or ( n3290 , n3288 , n3289 );
buf ( n170760 , n3290 );
buf ( n170761 , n170760 );
xor ( n3293 , n3286 , n170761 );
buf ( n170763 , n3293 );
buf ( n170764 , n170763 );
buf ( n170765 , n799 );
buf ( n170766 , n801 );
nand ( n3298 , n170765 , n170766 );
buf ( n170768 , n3298 );
buf ( n170769 , n799 );
buf ( n170770 , n801 );
or ( n3302 , n170769 , n170770 );
buf ( n170772 , n802 );
nand ( n3304 , n3302 , n170772 );
buf ( n170774 , n3304 );
nand ( n3306 , n170768 , n800 , n170774 );
buf ( n170776 , n3306 );
not ( n3308 , n170776 );
buf ( n170778 , n168585 );
not ( n3310 , n170778 );
buf ( n170780 , n1471 );
not ( n3312 , n170780 );
or ( n3313 , n3310 , n3312 );
buf ( n170783 , n768 );
buf ( n170784 , n830 );
xor ( n3316 , n170783 , n170784 );
buf ( n170786 , n3316 );
buf ( n170787 , n170786 );
buf ( n170788 , n831 );
nand ( n3320 , n170787 , n170788 );
buf ( n170790 , n3320 );
buf ( n170791 , n170790 );
nand ( n3323 , n3313 , n170791 );
buf ( n170793 , n3323 );
buf ( n170794 , n170793 );
not ( n3326 , n170794 );
or ( n3327 , n3308 , n3326 );
buf ( n170797 , n170793 );
buf ( n170798 , n3306 );
or ( n3330 , n170797 , n170798 );
nand ( n3331 , n3327 , n3330 );
buf ( n170801 , n3331 );
buf ( n170802 , n170801 );
xor ( n3334 , n168533 , n168571 );
and ( n3335 , n3334 , n168593 );
and ( n3336 , n168533 , n168571 );
or ( n3337 , n3335 , n3336 );
buf ( n170807 , n3337 );
buf ( n170808 , n170807 );
xor ( n3340 , n170802 , n170808 );
not ( n3341 , n170609 );
not ( n3342 , n170576 );
or ( n3343 , n3341 , n3342 );
buf ( n170813 , n170609 );
buf ( n170814 , n170576 );
nor ( n3346 , n170813 , n170814 );
buf ( n170816 , n3346 );
buf ( n170817 , n170592 );
not ( n3349 , n170817 );
buf ( n170819 , n3349 );
or ( n3351 , n170816 , n170819 );
nand ( n3352 , n3343 , n3351 );
buf ( n170822 , n3352 );
xor ( n3354 , n3340 , n170822 );
buf ( n170824 , n3354 );
not ( n3356 , n170508 );
not ( n3357 , n170548 );
or ( n3358 , n3356 , n3357 );
buf ( n170828 , n170508 );
buf ( n170829 , n170548 );
or ( n3361 , n170828 , n170829 );
buf ( n170831 , n170523 );
nand ( n3363 , n3361 , n170831 );
buf ( n170833 , n3363 );
nand ( n3365 , n3358 , n170833 );
not ( n3366 , n3365 );
not ( n3367 , n3366 );
not ( n3368 , n168658 );
not ( n3369 , n168630 );
not ( n3370 , n3369 );
not ( n3371 , n3370 );
or ( n3372 , n3368 , n3371 );
not ( n3373 , n3369 );
not ( n3374 , n168658 );
not ( n3375 , n3374 );
or ( n3376 , n3373 , n3375 );
nand ( n3377 , n3376 , n168692 );
nand ( n3378 , n3372 , n3377 );
not ( n3379 , n3378 );
not ( n3380 , n3379 );
or ( n3381 , n3367 , n3380 );
nand ( n3382 , n3365 , n3378 );
nand ( n3383 , n3381 , n3382 );
not ( n3384 , n168814 );
nand ( n3385 , n1304 , n1262 );
not ( n3386 , n3385 );
or ( n3387 , n3384 , n3386 );
nand ( n3388 , n168770 , n168730 );
nand ( n3389 , n3387 , n3388 );
not ( n3390 , n3389 );
and ( n3391 , n3383 , n3390 );
not ( n3392 , n3383 );
and ( n3393 , n3392 , n3389 );
nor ( n3394 , n3391 , n3393 );
not ( n3395 , n3394 );
xor ( n3396 , n170414 , n170431 );
and ( n3397 , n3396 , n170438 );
and ( n3398 , n170414 , n170431 );
or ( n3399 , n3397 , n3398 );
buf ( n170869 , n3399 );
and ( n3401 , n3395 , n170869 );
not ( n3402 , n3395 );
not ( n3403 , n170869 );
and ( n3404 , n3402 , n3403 );
nor ( n3405 , n3401 , n3404 );
xnor ( n3406 , n170824 , n3405 );
buf ( n170876 , n3406 );
xor ( n3408 , n168596 , n168694 );
and ( n3409 , n3408 , n168820 );
and ( n3410 , n168596 , n168694 );
or ( n3411 , n3409 , n3410 );
buf ( n170881 , n3411 );
buf ( n170882 , n170881 );
xor ( n3414 , n170495 , n170552 );
and ( n3415 , n3414 , n170611 );
and ( n3416 , n170495 , n170552 );
or ( n3417 , n3415 , n3416 );
buf ( n170887 , n3417 );
buf ( n170888 , n170887 );
xor ( n3420 , n170882 , n170888 );
buf ( n170890 , n2955 );
not ( n3422 , n170890 );
buf ( n170892 , n1389 );
not ( n3424 , n170892 );
or ( n3425 , n3422 , n3424 );
buf ( n170895 , n168867 );
buf ( n170896 , n796 );
buf ( n170897 , n802 );
xor ( n3429 , n170896 , n170897 );
buf ( n170899 , n3429 );
buf ( n170900 , n170899 );
nand ( n3432 , n170895 , n170900 );
buf ( n170902 , n3432 );
buf ( n170903 , n170902 );
nand ( n3435 , n3425 , n170903 );
buf ( n170905 , n3435 );
buf ( n170906 , n168764 );
not ( n3438 , n170906 );
buf ( n170908 , n1578 );
not ( n3440 , n170908 );
or ( n3441 , n3438 , n3440 );
buf ( n170911 , n168759 );
buf ( n170912 , n794 );
buf ( n170913 , n804 );
xor ( n3445 , n170912 , n170913 );
buf ( n170915 , n3445 );
buf ( n170916 , n170915 );
nand ( n3448 , n170911 , n170916 );
buf ( n170918 , n3448 );
buf ( n170919 , n170918 );
nand ( n3451 , n3441 , n170919 );
buf ( n170921 , n3451 );
xor ( n3453 , n170905 , n170921 );
buf ( n170923 , n1339 );
not ( n3455 , n170923 );
buf ( n170925 , n1321 );
not ( n3457 , n170925 );
or ( n3458 , n3455 , n3457 );
buf ( n170928 , n168806 );
xor ( n3460 , n818 , n780 );
buf ( n170930 , n3460 );
nand ( n3462 , n170928 , n170930 );
buf ( n170932 , n3462 );
buf ( n170933 , n170932 );
nand ( n3465 , n3458 , n170933 );
buf ( n170935 , n3465 );
xor ( n3467 , n3453 , n170935 );
buf ( n170937 , n3467 );
buf ( n170938 , n170570 );
not ( n3470 , n170938 );
buf ( n170940 , n1806 );
not ( n3472 , n170940 );
or ( n3473 , n3470 , n3472 );
buf ( n170943 , n170565 );
buf ( n170944 , n774 );
buf ( n170945 , n824 );
xor ( n3477 , n170944 , n170945 );
buf ( n170947 , n3477 );
buf ( n170948 , n170947 );
nand ( n3480 , n170943 , n170948 );
buf ( n170950 , n3480 );
buf ( n170951 , n170950 );
nand ( n3483 , n3473 , n170951 );
buf ( n170953 , n3483 );
buf ( n170954 , n170953 );
buf ( n170955 , n799 );
buf ( n170956 , n800 );
xor ( n3488 , n170955 , n170956 );
buf ( n170958 , n3488 );
buf ( n170959 , n170958 );
not ( n3491 , n170959 );
buf ( n170961 , n801 );
buf ( n170962 , n800 );
xnor ( n3494 , n170961 , n170962 );
buf ( n170964 , n3494 );
nor ( n3496 , n170964 , n168528 );
buf ( n3497 , n3496 );
buf ( n170967 , n3497 );
not ( n3499 , n170967 );
or ( n3500 , n3491 , n3499 );
buf ( n170970 , n168528 );
buf ( n3502 , n170970 );
buf ( n170972 , n3502 );
buf ( n170973 , n170972 );
buf ( n170974 , n798 );
buf ( n170975 , n800 );
xor ( n3507 , n170974 , n170975 );
buf ( n170977 , n3507 );
buf ( n170978 , n170977 );
nand ( n3510 , n170973 , n170978 );
buf ( n170980 , n3510 );
buf ( n170981 , n170980 );
nand ( n3513 , n3500 , n170981 );
buf ( n170983 , n3513 );
buf ( n170984 , n170983 );
xor ( n3516 , n170954 , n170984 );
buf ( n170986 , n168564 );
not ( n3518 , n170986 );
buf ( n170988 , n1742 );
buf ( n3520 , n170988 );
buf ( n170990 , n3520 );
buf ( n170991 , n170990 );
not ( n3523 , n170991 );
or ( n3524 , n3518 , n3523 );
buf ( n170994 , n168559 );
buf ( n170995 , n770 );
buf ( n170996 , n828 );
xor ( n3528 , n170995 , n170996 );
buf ( n170998 , n3528 );
buf ( n170999 , n170998 );
nand ( n3531 , n170994 , n170999 );
buf ( n171001 , n3531 );
buf ( n171002 , n171001 );
nand ( n3534 , n3524 , n171002 );
buf ( n171004 , n3534 );
buf ( n171005 , n171004 );
xor ( n3537 , n3516 , n171005 );
buf ( n171007 , n3537 );
buf ( n171008 , n171007 );
xor ( n3540 , n170937 , n171008 );
not ( n3541 , n170603 );
buf ( n171011 , n169241 );
buf ( n3543 , n171011 );
buf ( n171013 , n3543 );
not ( n3545 , n171013 );
or ( n3546 , n3541 , n3545 );
buf ( n171016 , n169931 );
buf ( n171017 , n784 );
buf ( n171018 , n814 );
xor ( n3550 , n171017 , n171018 );
buf ( n171020 , n3550 );
buf ( n171021 , n171020 );
nand ( n3553 , n171016 , n171021 );
buf ( n171023 , n3553 );
nand ( n3555 , n3546 , n171023 );
buf ( n171025 , n170586 );
not ( n3557 , n171025 );
buf ( n171027 , n169314 );
buf ( n3559 , n171027 );
buf ( n171029 , n3559 );
buf ( n171030 , n171029 );
not ( n3562 , n171030 );
or ( n3563 , n3557 , n3562 );
buf ( n171033 , n169845 );
buf ( n171034 , n782 );
buf ( n171035 , n816 );
xor ( n3567 , n171034 , n171035 );
buf ( n171037 , n3567 );
buf ( n171038 , n171037 );
nand ( n3570 , n171033 , n171038 );
buf ( n171040 , n3570 );
buf ( n171041 , n171040 );
nand ( n3573 , n3563 , n171041 );
buf ( n171043 , n3573 );
xor ( n3575 , n3555 , n171043 );
buf ( n171045 , n3033 );
not ( n3577 , n171045 );
buf ( n171047 , n1939 );
buf ( n3579 , n171047 );
buf ( n171049 , n3579 );
buf ( n171050 , n171049 );
not ( n3582 , n171050 );
or ( n3583 , n3577 , n3582 );
buf ( n171053 , n169417 );
buf ( n3585 , n171053 );
buf ( n171055 , n3585 );
buf ( n171056 , n171055 );
buf ( n171057 , n776 );
buf ( n171058 , n822 );
xor ( n3590 , n171057 , n171058 );
buf ( n171060 , n3590 );
buf ( n171061 , n171060 );
nand ( n3593 , n171056 , n171061 );
buf ( n171063 , n3593 );
buf ( n171064 , n171063 );
nand ( n3596 , n3583 , n171064 );
buf ( n171066 , n3596 );
xor ( n3598 , n3575 , n171066 );
buf ( n171068 , n3598 );
xor ( n3600 , n3540 , n171068 );
buf ( n171070 , n3600 );
buf ( n171071 , n171070 );
xor ( n3603 , n3420 , n171071 );
buf ( n171073 , n3603 );
buf ( n171074 , n171073 );
xor ( n3606 , n170876 , n171074 );
xor ( n3607 , n168823 , n169452 );
and ( n3608 , n3607 , n169868 );
and ( n3609 , n168823 , n169452 );
or ( n3610 , n3608 , n3609 );
buf ( n171080 , n3610 );
buf ( n171081 , n171080 );
xor ( n3613 , n3606 , n171081 );
buf ( n171083 , n3613 );
buf ( n171084 , n171083 );
xor ( n3616 , n170764 , n171084 );
xor ( n3617 , n170456 , n170617 );
and ( n3618 , n3617 , n170623 );
and ( n3619 , n170456 , n170617 );
or ( n3620 , n3618 , n3619 );
buf ( n171090 , n3620 );
buf ( n171091 , n171090 );
xor ( n3623 , n3616 , n171091 );
buf ( n171093 , n3623 );
buf ( n171094 , n171093 );
and ( n3626 , n3163 , n171094 );
and ( n3627 , n168524 , n170631 );
or ( n3628 , n3626 , n3627 );
buf ( n171098 , n3628 );
buf ( n171099 , n171098 );
xor ( n3631 , n170764 , n171084 );
and ( n3632 , n3631 , n171091 );
and ( n3633 , n170764 , n171084 );
or ( n3634 , n3632 , n3633 );
buf ( n171104 , n3634 );
buf ( n171105 , n171104 );
not ( n3637 , n171105 );
xor ( n3638 , n170748 , n170754 );
and ( n3639 , n3638 , n170761 );
and ( n3640 , n170748 , n170754 );
or ( n3641 , n3639 , n3640 );
buf ( n171111 , n3641 );
buf ( n171112 , n171111 );
xor ( n3644 , n170876 , n171074 );
and ( n3645 , n3644 , n171081 );
and ( n3646 , n170876 , n171074 );
or ( n3647 , n3645 , n3646 );
buf ( n171117 , n3647 );
buf ( n171118 , n171117 );
xor ( n3650 , n171112 , n171118 );
xor ( n3651 , n170802 , n170808 );
and ( n3652 , n3651 , n170822 );
and ( n3653 , n170802 , n170808 );
or ( n3654 , n3652 , n3653 );
buf ( n171124 , n3654 );
buf ( n171125 , n171124 );
not ( n3657 , n171125 );
buf ( n171127 , n3657 );
buf ( n171128 , n171127 );
buf ( n171129 , n799 );
buf ( n171130 , n800 );
and ( n3662 , n171129 , n171130 );
buf ( n171132 , n3662 );
buf ( n171133 , n171132 );
buf ( n171134 , n170786 );
not ( n3666 , n171134 );
buf ( n171136 , n168471 );
not ( n3668 , n171136 );
or ( n3669 , n3666 , n3668 );
buf ( n171139 , n830 );
buf ( n171140 , n831 );
nand ( n3672 , n171139 , n171140 );
buf ( n171142 , n3672 );
buf ( n171143 , n171142 );
nand ( n3675 , n3669 , n171143 );
buf ( n171145 , n3675 );
buf ( n171146 , n171145 );
xor ( n3678 , n171133 , n171146 );
buf ( n171148 , n170998 );
not ( n3680 , n171148 );
not ( n3681 , n168547 );
xor ( n3682 , n829 , n830 );
nor ( n3683 , n3681 , n3682 );
buf ( n171153 , n3683 );
not ( n3685 , n171153 );
or ( n3686 , n3680 , n3685 );
buf ( n171156 , n168559 );
buf ( n171157 , n769 );
buf ( n171158 , n828 );
xor ( n3690 , n171157 , n171158 );
buf ( n171160 , n3690 );
buf ( n171161 , n171160 );
nand ( n3693 , n171156 , n171161 );
buf ( n171163 , n3693 );
buf ( n171164 , n171163 );
nand ( n3696 , n3686 , n171164 );
buf ( n171166 , n3696 );
buf ( n171167 , n171166 );
xor ( n3699 , n3678 , n171167 );
buf ( n171169 , n3699 );
buf ( n171170 , n171169 );
buf ( n171171 , n170905 );
not ( n3703 , n171171 );
buf ( n171173 , n170921 );
not ( n3705 , n171173 );
or ( n3706 , n3703 , n3705 );
buf ( n171176 , n170921 );
buf ( n171177 , n170905 );
or ( n3709 , n171176 , n171177 );
buf ( n171179 , n170935 );
nand ( n3711 , n3709 , n171179 );
buf ( n171181 , n3711 );
buf ( n171182 , n171181 );
nand ( n3714 , n3706 , n171182 );
buf ( n171184 , n3714 );
buf ( n171185 , n171184 );
xor ( n3717 , n171170 , n171185 );
xor ( n3718 , n170649 , n170666 );
and ( n3719 , n3718 , n170680 );
and ( n3720 , n170649 , n170666 );
or ( n3721 , n3719 , n3720 );
buf ( n171191 , n3721 );
buf ( n171192 , n171191 );
xnor ( n3724 , n3717 , n171192 );
buf ( n171194 , n3724 );
buf ( n171195 , n171194 );
not ( n3727 , n171195 );
buf ( n171197 , n3727 );
buf ( n171198 , n171197 );
xor ( n3730 , n171128 , n171198 );
xor ( n3731 , n170937 , n171008 );
and ( n3732 , n3731 , n171068 );
and ( n3733 , n170937 , n171008 );
or ( n3734 , n3732 , n3733 );
buf ( n171204 , n3734 );
buf ( n171205 , n171204 );
xnor ( n3737 , n3730 , n171205 );
buf ( n171207 , n3737 );
buf ( n171208 , n171207 );
buf ( n171209 , n171060 );
not ( n3741 , n171209 );
buf ( n171211 , n2418 );
not ( n3743 , n171211 );
or ( n3744 , n3741 , n3743 );
buf ( n171214 , n169417 );
buf ( n171215 , n775 );
buf ( n171216 , n822 );
xor ( n3748 , n171215 , n171216 );
buf ( n171218 , n3748 );
buf ( n171219 , n171218 );
nand ( n3751 , n171214 , n171219 );
buf ( n171221 , n3751 );
buf ( n171222 , n171221 );
nand ( n3754 , n3744 , n171222 );
buf ( n171224 , n3754 );
buf ( n171225 , n171224 );
buf ( n171226 , n171020 );
not ( n3758 , n171226 );
not ( n3759 , n814 );
and ( n3760 , n815 , n3759 );
not ( n3761 , n815 );
and ( n3762 , n3761 , n814 );
nor ( n3763 , n3760 , n3762 );
nor ( n3764 , n3763 , n1768 );
buf ( n171234 , n3764 );
not ( n3766 , n171234 );
or ( n3767 , n3758 , n3766 );
buf ( n171237 , n169247 );
buf ( n171238 , n783 );
buf ( n171239 , n814 );
xor ( n3771 , n171238 , n171239 );
buf ( n171241 , n3771 );
buf ( n171242 , n171241 );
nand ( n3774 , n171237 , n171242 );
buf ( n171244 , n3774 );
buf ( n171245 , n171244 );
nand ( n3777 , n3767 , n171245 );
buf ( n171247 , n3777 );
buf ( n171248 , n171247 );
not ( n3780 , n171248 );
buf ( n171250 , n3780 );
buf ( n171251 , n171250 );
and ( n3783 , n171225 , n171251 );
not ( n3784 , n171225 );
buf ( n171254 , n171247 );
and ( n3786 , n3784 , n171254 );
nor ( n3787 , n3783 , n3786 );
buf ( n171257 , n3787 );
buf ( n171258 , n171257 );
buf ( n171259 , n170694 );
not ( n3791 , n171259 );
buf ( n171261 , n2757 );
not ( n3793 , n171261 );
or ( n3794 , n3791 , n3793 );
buf ( n171264 , n1534 );
buf ( n171265 , n785 );
buf ( n171266 , n812 );
xor ( n3798 , n171265 , n171266 );
buf ( n171268 , n3798 );
buf ( n171269 , n171268 );
nand ( n3801 , n171264 , n171269 );
buf ( n171271 , n3801 );
buf ( n171272 , n171271 );
nand ( n3804 , n3794 , n171272 );
buf ( n171274 , n3804 );
buf ( n171275 , n171274 );
and ( n3807 , n171258 , n171275 );
not ( n3808 , n171258 );
buf ( n171278 , n171274 );
not ( n3810 , n171278 );
buf ( n171280 , n3810 );
buf ( n171281 , n171280 );
and ( n3813 , n3808 , n171281 );
nor ( n3814 , n3807 , n3813 );
buf ( n171284 , n3814 );
not ( n3816 , n170672 );
not ( n3817 , n168648 );
or ( n3818 , n3816 , n3817 );
buf ( n171288 , n777 );
buf ( n171289 , n820 );
xor ( n3821 , n171288 , n171289 );
buf ( n171291 , n3821 );
buf ( n171292 , n171291 );
buf ( n171293 , n821 );
buf ( n171294 , n822 );
xor ( n3826 , n171293 , n171294 );
buf ( n171296 , n3826 );
buf ( n171297 , n171296 );
nand ( n3829 , n171292 , n171297 );
buf ( n171299 , n3829 );
nand ( n3831 , n3818 , n171299 );
not ( n3832 , n3831 );
not ( n3833 , n170713 );
not ( n3834 , n2737 );
or ( n3835 , n3833 , n3834 );
buf ( n171305 , n169957 );
buf ( n171306 , n787 );
buf ( n171307 , n810 );
xor ( n3839 , n171306 , n171307 );
buf ( n171309 , n3839 );
buf ( n171310 , n171309 );
nand ( n3842 , n171305 , n171310 );
buf ( n171312 , n3842 );
nand ( n3844 , n3835 , n171312 );
not ( n3845 , n3844 );
or ( n3846 , n3832 , n3845 );
not ( n3847 , n170713 );
not ( n3848 , n2737 );
or ( n3849 , n3847 , n3848 );
nand ( n3850 , n3849 , n171312 );
or ( n3851 , n3850 , n3831 );
nand ( n3852 , n3846 , n3851 );
buf ( n171322 , n169093 );
buf ( n171323 , n170730 );
not ( n3855 , n171323 );
buf ( n171325 , n3855 );
buf ( n171326 , n171325 );
or ( n3858 , n171322 , n171326 );
buf ( n171328 , n169081 );
not ( n3860 , n171328 );
buf ( n171330 , n3860 );
buf ( n171331 , n171330 );
buf ( n171332 , n771 );
buf ( n171333 , n826 );
xor ( n3865 , n171332 , n171333 );
buf ( n171335 , n3865 );
buf ( n171336 , n171335 );
not ( n3868 , n171336 );
buf ( n171338 , n3868 );
buf ( n171339 , n171338 );
or ( n3871 , n171331 , n171339 );
nand ( n3872 , n3858 , n3871 );
buf ( n171342 , n3872 );
and ( n3874 , n3852 , n171342 );
not ( n3875 , n3852 );
buf ( n171345 , n171342 );
not ( n3877 , n171345 );
buf ( n171347 , n3877 );
and ( n3879 , n3875 , n171347 );
nor ( n3880 , n3874 , n3879 );
and ( n3881 , n171284 , n3880 );
not ( n3882 , n171284 );
not ( n3883 , n3880 );
and ( n3884 , n3882 , n3883 );
nor ( n3885 , n3881 , n3884 );
buf ( n171355 , n3885 );
buf ( n171356 , n170641 );
not ( n3888 , n171356 );
buf ( n171358 , n168615 );
not ( n3890 , n171358 );
or ( n3891 , n3888 , n3890 );
buf ( n171361 , n168619 );
buf ( n171362 , n789 );
buf ( n171363 , n808 );
xor ( n3895 , n171362 , n171363 );
buf ( n171365 , n3895 );
buf ( n171366 , n171365 );
nand ( n3898 , n171361 , n171366 );
buf ( n171368 , n3898 );
buf ( n171369 , n171368 );
nand ( n3901 , n3891 , n171369 );
buf ( n171371 , n3901 );
buf ( n171372 , n171371 );
buf ( n171373 , n170659 );
not ( n3905 , n171373 );
buf ( n171375 , n169635 );
not ( n3907 , n171375 );
or ( n3908 , n3905 , n3907 );
buf ( n171378 , n169641 );
buf ( n171379 , n791 );
buf ( n171380 , n806 );
xor ( n3912 , n171379 , n171380 );
buf ( n171382 , n3912 );
buf ( n171383 , n171382 );
nand ( n3915 , n171378 , n171383 );
buf ( n171385 , n3915 );
buf ( n171386 , n171385 );
nand ( n3918 , n3908 , n171386 );
buf ( n171388 , n3918 );
buf ( n171389 , n171388 );
xor ( n3921 , n171372 , n171389 );
buf ( n171391 , n3460 );
not ( n3923 , n171391 );
buf ( n171393 , n1321 );
not ( n3925 , n171393 );
or ( n3926 , n3923 , n3925 );
buf ( n171396 , n168806 );
buf ( n171397 , n779 );
buf ( n171398 , n818 );
xor ( n3930 , n171397 , n171398 );
buf ( n171400 , n3930 );
buf ( n171401 , n171400 );
nand ( n3933 , n171396 , n171401 );
buf ( n171403 , n3933 );
buf ( n171404 , n171403 );
nand ( n3936 , n3926 , n171404 );
buf ( n171406 , n3936 );
buf ( n171407 , n171406 );
xor ( n3939 , n3921 , n171407 );
buf ( n171409 , n3939 );
buf ( n171410 , n171409 );
and ( n3942 , n171355 , n171410 );
not ( n3943 , n171355 );
buf ( n171413 , n171409 );
not ( n3945 , n171413 );
buf ( n171415 , n3945 );
buf ( n171416 , n171415 );
and ( n3948 , n3943 , n171416 );
nor ( n3949 , n3942 , n3948 );
buf ( n171419 , n3949 );
buf ( n171420 , n171419 );
buf ( n171421 , n171066 );
not ( n3953 , n171421 );
buf ( n171423 , n170603 );
not ( n3955 , n171423 );
buf ( n171425 , n171013 );
not ( n3957 , n171425 );
or ( n3958 , n3955 , n3957 );
buf ( n171428 , n171023 );
nand ( n3960 , n3958 , n171428 );
buf ( n171430 , n3960 );
buf ( n171431 , n171430 );
not ( n3963 , n171431 );
or ( n3964 , n3953 , n3963 );
buf ( n171434 , n171066 );
buf ( n171435 , n171430 );
or ( n3967 , n171434 , n171435 );
buf ( n171437 , n171043 );
nand ( n3969 , n3967 , n171437 );
buf ( n171439 , n3969 );
buf ( n171440 , n171439 );
nand ( n3972 , n3964 , n171440 );
buf ( n171442 , n3972 );
buf ( n171443 , n170719 );
not ( n3975 , n171443 );
buf ( n171445 , n170736 );
not ( n3977 , n171445 );
or ( n3978 , n3975 , n3977 );
buf ( n171448 , n170736 );
buf ( n171449 , n170719 );
or ( n3981 , n171448 , n171449 );
buf ( n171451 , n170700 );
nand ( n3983 , n3981 , n171451 );
buf ( n171453 , n3983 );
buf ( n171454 , n171453 );
nand ( n3986 , n3978 , n171454 );
buf ( n171456 , n3986 );
buf ( n171457 , n171456 );
not ( n3989 , n171457 );
buf ( n171459 , n3989 );
xor ( n3991 , n171442 , n171459 );
xor ( n3992 , n170954 , n170984 );
and ( n3993 , n3992 , n171005 );
and ( n3994 , n170954 , n170984 );
or ( n3995 , n3993 , n3994 );
buf ( n171465 , n3995 );
xnor ( n3997 , n3991 , n171465 );
buf ( n171467 , n3997 );
xor ( n3999 , n171420 , n171467 );
xor ( n4000 , n170683 , n170738 );
and ( n4001 , n4000 , n170745 );
and ( n4002 , n170683 , n170738 );
or ( n4003 , n4001 , n4002 );
buf ( n171473 , n4003 );
buf ( n171474 , n171473 );
xor ( n4006 , n3999 , n171474 );
buf ( n171476 , n4006 );
buf ( n171477 , n171476 );
xor ( n4009 , n171208 , n171477 );
buf ( n171479 , n3365 );
not ( n4011 , n171479 );
buf ( n171481 , n3378 );
not ( n4013 , n171481 );
or ( n4014 , n4011 , n4013 );
or ( n4015 , n3365 , n3378 );
nand ( n4016 , n4015 , n3389 );
buf ( n171486 , n4016 );
nand ( n4018 , n4014 , n171486 );
buf ( n171488 , n4018 );
buf ( n171489 , n171488 );
not ( n4021 , n171489 );
buf ( n171491 , n170899 );
not ( n4023 , n171491 );
buf ( n171493 , n1389 );
not ( n4025 , n171493 );
or ( n4026 , n4023 , n4025 );
buf ( n171496 , n168867 );
buf ( n171497 , n795 );
buf ( n171498 , n802 );
xor ( n4030 , n171497 , n171498 );
buf ( n171500 , n4030 );
buf ( n171501 , n171500 );
nand ( n4033 , n171496 , n171501 );
buf ( n171503 , n4033 );
buf ( n171504 , n171503 );
nand ( n4036 , n4026 , n171504 );
buf ( n171506 , n4036 );
buf ( n171507 , n170915 );
not ( n4039 , n171507 );
buf ( n171509 , n168832 );
not ( n4041 , n171509 );
or ( n4042 , n4039 , n4041 );
buf ( n171512 , n168759 );
buf ( n171513 , n793 );
buf ( n171514 , n804 );
xor ( n4046 , n171513 , n171514 );
buf ( n171516 , n4046 );
buf ( n171517 , n171516 );
nand ( n4049 , n171512 , n171517 );
buf ( n171519 , n4049 );
buf ( n171520 , n171519 );
nand ( n4052 , n4042 , n171520 );
buf ( n171522 , n4052 );
xor ( n4054 , n171506 , n171522 );
buf ( n171524 , n3306 );
not ( n4056 , n171524 );
buf ( n171526 , n170793 );
nand ( n4058 , n4056 , n171526 );
buf ( n171528 , n4058 );
and ( n4060 , n4054 , n171528 );
not ( n4061 , n4054 );
buf ( n171531 , n171528 );
not ( n4063 , n171531 );
buf ( n171533 , n4063 );
and ( n4065 , n4061 , n171533 );
nor ( n4066 , n4060 , n4065 );
buf ( n171536 , n4066 );
not ( n4068 , n171536 );
buf ( n171538 , n170977 );
not ( n4070 , n171538 );
buf ( n171540 , n170964 );
buf ( n171541 , n168528 );
nor ( n4073 , n171540 , n171541 );
buf ( n171543 , n4073 );
buf ( n171544 , n171543 );
not ( n4076 , n171544 );
or ( n4077 , n4070 , n4076 );
buf ( n171547 , n168528 );
buf ( n171548 , n797 );
buf ( n171549 , n800 );
xor ( n4081 , n171548 , n171549 );
buf ( n171551 , n4081 );
buf ( n171552 , n171551 );
nand ( n4084 , n171547 , n171552 );
buf ( n171554 , n4084 );
buf ( n171555 , n171554 );
nand ( n4087 , n4077 , n171555 );
buf ( n171557 , n4087 );
buf ( n171558 , n171557 );
buf ( n171559 , n171037 );
not ( n4091 , n171559 );
buf ( n171561 , n169833 );
not ( n4093 , n171561 );
or ( n4094 , n4091 , n4093 );
buf ( n171564 , n169842 );
buf ( n171565 , n781 );
buf ( n171566 , n816 );
xor ( n4098 , n171565 , n171566 );
buf ( n171568 , n4098 );
buf ( n171569 , n171568 );
nand ( n4101 , n171564 , n171569 );
buf ( n171571 , n4101 );
buf ( n171572 , n171571 );
nand ( n4104 , n4094 , n171572 );
buf ( n171574 , n4104 );
buf ( n171575 , n171574 );
xor ( n4107 , n171558 , n171575 );
buf ( n171577 , n170947 );
not ( n4109 , n171577 );
buf ( n171579 , n170100 );
not ( n4111 , n171579 );
or ( n4112 , n4109 , n4111 );
buf ( n171582 , n170565 );
xor ( n4114 , n824 , n773 );
buf ( n171584 , n4114 );
nand ( n4116 , n171582 , n171584 );
buf ( n171586 , n4116 );
buf ( n171587 , n171586 );
nand ( n4119 , n4112 , n171587 );
buf ( n171589 , n4119 );
buf ( n171590 , n171589 );
xor ( n4122 , n4107 , n171590 );
buf ( n171592 , n4122 );
buf ( n171593 , n171592 );
not ( n4125 , n171593 );
and ( n4126 , n4068 , n4125 );
buf ( n171596 , n4066 );
buf ( n171597 , n171592 );
and ( n4129 , n171596 , n171597 );
nor ( n4130 , n4126 , n4129 );
buf ( n171600 , n4130 );
buf ( n171601 , n171600 );
not ( n4133 , n171601 );
or ( n4134 , n4021 , n4133 );
buf ( n171604 , n171600 );
buf ( n171605 , n171488 );
or ( n4137 , n171604 , n171605 );
nand ( n4138 , n4134 , n4137 );
buf ( n171608 , n4138 );
buf ( n171609 , n171608 );
not ( n4141 , n170869 );
not ( n4142 , n170824 );
or ( n4143 , n4141 , n4142 );
buf ( n171613 , n170869 );
buf ( n171614 , n170824 );
or ( n4146 , n171613 , n171614 );
buf ( n171616 , n3394 );
nand ( n4148 , n4146 , n171616 );
buf ( n171618 , n4148 );
nand ( n4150 , n4143 , n171618 );
buf ( n171620 , n4150 );
xor ( n4152 , n171609 , n171620 );
xor ( n4153 , n170882 , n170888 );
and ( n4154 , n4153 , n171071 );
and ( n4155 , n170882 , n170888 );
or ( n4156 , n4154 , n4155 );
buf ( n171626 , n4156 );
buf ( n171627 , n171626 );
xor ( n4159 , n4152 , n171627 );
buf ( n171629 , n4159 );
buf ( n171630 , n171629 );
xor ( n4162 , n4009 , n171630 );
buf ( n171632 , n4162 );
buf ( n171633 , n171632 );
xor ( n4165 , n3650 , n171633 );
buf ( n171635 , n4165 );
buf ( n171636 , n171635 );
not ( n4168 , n171636 );
buf ( n171638 , n4168 );
buf ( n171639 , n171638 );
not ( n4171 , n171639 );
or ( n4172 , n3637 , n4171 );
buf ( n171642 , n171635 );
buf ( n171643 , n171104 );
not ( n4175 , n171643 );
buf ( n171645 , n4175 );
buf ( n171646 , n171645 );
nand ( n4178 , n171642 , n171646 );
buf ( n171648 , n4178 );
buf ( n171649 , n171648 );
nand ( n4181 , n4172 , n171649 );
buf ( n171651 , n4181 );
buf ( n171652 , n171651 );
or ( n4184 , n171099 , n171652 );
buf ( n171654 , n4184 );
buf ( n171655 , n171654 );
buf ( n4187 , n171655 );
buf ( n171657 , n4187 );
buf ( n171658 , n171657 );
nand ( n4190 , n171098 , n171651 );
buf ( n171660 , n4190 );
buf ( n4192 , n171660 );
buf ( n171662 , n4192 );
buf ( n171663 , n171662 );
nand ( n4195 , n171658 , n171663 );
buf ( n171665 , n4195 );
buf ( n171666 , n171665 );
not ( n4198 , n171666 );
xor ( n4199 , n168524 , n170631 );
xor ( n4200 , n4199 , n171094 );
buf ( n171670 , n4200 );
not ( n4202 , n171670 );
buf ( n171672 , n833 );
xor ( n4204 , n169871 , n170408 );
xor ( n4205 , n4204 , n170626 );
buf ( n171675 , n4205 );
buf ( n171676 , n171675 );
xor ( n4208 , n171672 , n171676 );
xor ( n4209 , n169874 , n2409 );
and ( n4210 , n4209 , n2930 );
not ( n4211 , n4209 );
not ( n4212 , n2930 );
and ( n4213 , n4211 , n4212 );
nor ( n4214 , n4210 , n4213 );
not ( n4215 , n4214 );
not ( n4216 , n1631 );
nand ( n4217 , n4216 , n1637 , n1708 );
not ( n4218 , n1708 );
nand ( n4219 , n4218 , n1562 , n1635 );
nand ( n4220 , n1707 , n1631 , n1637 );
nand ( n4221 , n1708 , n1631 , n1562 );
nand ( n4222 , n4217 , n4219 , n4220 , n4221 );
buf ( n171692 , n4222 );
buf ( n171693 , n786 );
buf ( n171694 , n818 );
xor ( n4226 , n171693 , n171694 );
buf ( n171696 , n4226 );
buf ( n171697 , n171696 );
not ( n4229 , n171697 );
buf ( n171699 , n818 );
buf ( n171700 , n819 );
xnor ( n4232 , n171699 , n171700 );
buf ( n171702 , n4232 );
buf ( n171703 , n171702 );
buf ( n171704 , n168788 );
nor ( n4236 , n171703 , n171704 );
buf ( n171706 , n4236 );
buf ( n171707 , n171706 );
not ( n4239 , n171707 );
or ( n4240 , n4229 , n4239 );
buf ( n171710 , n168806 );
buf ( n171711 , n170058 );
nand ( n4243 , n171710 , n171711 );
buf ( n171713 , n4243 );
buf ( n171714 , n171713 );
nand ( n4246 , n4240 , n171714 );
buf ( n171716 , n4246 );
buf ( n171717 , n171716 );
buf ( n171718 , n778 );
buf ( n171719 , n826 );
xor ( n4251 , n171718 , n171719 );
buf ( n171721 , n4251 );
buf ( n171722 , n171721 );
not ( n4254 , n171722 );
buf ( n171724 , n169674 );
not ( n4256 , n171724 );
or ( n4257 , n4254 , n4256 );
buf ( n171727 , n2207 );
buf ( n171728 , n168684 );
nand ( n4260 , n171727 , n171728 );
buf ( n171730 , n4260 );
buf ( n171731 , n171730 );
nand ( n4263 , n4257 , n171731 );
buf ( n171733 , n4263 );
buf ( n171734 , n171733 );
xor ( n4266 , n171717 , n171734 );
not ( n4267 , n170083 );
not ( n4268 , n168559 );
or ( n4269 , n4267 , n4268 );
not ( n4270 , n3682 );
xor ( n4271 , n777 , n828 );
nand ( n4272 , n4270 , n168547 , n4271 );
nand ( n4273 , n4269 , n4272 );
buf ( n171743 , n4273 );
buf ( n171744 , n799 );
buf ( n171745 , n807 );
or ( n4277 , n171744 , n171745 );
buf ( n171747 , n808 );
nand ( n4279 , n4277 , n171747 );
buf ( n171749 , n4279 );
buf ( n171750 , n799 );
buf ( n171751 , n807 );
nand ( n4283 , n171750 , n171751 );
buf ( n171753 , n4283 );
and ( n4285 , n171749 , n171753 , n806 );
buf ( n171755 , n4285 );
and ( n4287 , n171743 , n171755 );
buf ( n171757 , n4287 );
buf ( n171758 , n171757 );
and ( n4290 , n4266 , n171758 );
and ( n4291 , n171717 , n171734 );
or ( n4292 , n4290 , n4291 );
buf ( n171762 , n4292 );
buf ( n171763 , n171762 );
xor ( n4295 , n169365 , n169387 );
xor ( n4296 , n4295 , n169435 );
buf ( n171766 , n4296 );
buf ( n171767 , n171766 );
xor ( n4299 , n171763 , n171767 );
xor ( n4300 , n170071 , n170073 );
xor ( n4301 , n4300 , n170127 );
buf ( n171771 , n4301 );
buf ( n171772 , n171771 );
and ( n4304 , n4299 , n171772 );
and ( n4305 , n171763 , n171767 );
or ( n4306 , n4304 , n4305 );
buf ( n171776 , n4306 );
buf ( n171777 , n171776 );
xor ( n4309 , n171692 , n171777 );
xor ( n4310 , n170199 , n170217 );
xor ( n4311 , n4310 , n170237 );
buf ( n171781 , n4311 );
buf ( n171782 , n171781 );
buf ( n171783 , n799 );
buf ( n171784 , n806 );
xor ( n4316 , n171783 , n171784 );
buf ( n171786 , n4316 );
buf ( n171787 , n171786 );
not ( n4319 , n171787 );
buf ( n171789 , n169635 );
not ( n4321 , n171789 );
or ( n4322 , n4319 , n4321 );
buf ( n171792 , n169641 );
buf ( n171793 , n170286 );
nand ( n4325 , n171792 , n171793 );
buf ( n171795 , n4325 );
buf ( n171796 , n171795 );
nand ( n4328 , n4322 , n171796 );
buf ( n171798 , n4328 );
buf ( n171799 , n171798 );
buf ( n171800 , n779 );
buf ( n171801 , n826 );
xor ( n4333 , n171800 , n171801 );
buf ( n171803 , n4333 );
buf ( n171804 , n171803 );
not ( n4336 , n171804 );
not ( n4337 , n1620 );
buf ( n171807 , n4337 );
not ( n4339 , n171807 );
or ( n4340 , n4336 , n4339 );
buf ( n171810 , n169081 );
buf ( n171811 , n171721 );
nand ( n4343 , n171810 , n171811 );
buf ( n171813 , n4343 );
buf ( n171814 , n171813 );
nand ( n4346 , n4340 , n171814 );
buf ( n171816 , n4346 );
buf ( n171817 , n171816 );
xor ( n4349 , n171799 , n171817 );
buf ( n171819 , n787 );
buf ( n171820 , n818 );
xor ( n4352 , n171819 , n171820 );
buf ( n171822 , n4352 );
buf ( n171823 , n171822 );
not ( n4355 , n171823 );
buf ( n171825 , n1321 );
not ( n4357 , n171825 );
or ( n4358 , n4355 , n4357 );
buf ( n171828 , n168806 );
buf ( n171829 , n171696 );
nand ( n4361 , n171828 , n171829 );
buf ( n171831 , n4361 );
buf ( n171832 , n171831 );
nand ( n4364 , n4358 , n171832 );
buf ( n171834 , n4364 );
buf ( n171835 , n171834 );
and ( n4367 , n4349 , n171835 );
and ( n4368 , n171799 , n171817 );
or ( n4369 , n4367 , n4368 );
buf ( n171839 , n4369 );
buf ( n171840 , n171839 );
xor ( n4372 , n171782 , n171840 );
xor ( n4373 , n170079 , n170096 );
xor ( n4374 , n4373 , n170122 );
buf ( n171844 , n4374 );
buf ( n171845 , n171844 );
and ( n4377 , n4372 , n171845 );
and ( n4378 , n171782 , n171840 );
or ( n4379 , n4377 , n4378 );
buf ( n171849 , n4379 );
buf ( n171850 , n171849 );
not ( n4382 , n2716 );
not ( n4383 , n4382 );
not ( n4384 , n170305 );
not ( n4385 , n170241 );
not ( n4386 , n4385 );
or ( n4387 , n4384 , n4386 );
nand ( n4388 , n2837 , n170241 );
nand ( n4389 , n4387 , n4388 );
not ( n4390 , n4389 );
or ( n4391 , n4383 , n4390 );
or ( n4392 , n4382 , n4389 );
nand ( n4393 , n4391 , n4392 );
buf ( n171863 , n4393 );
or ( n4395 , n171850 , n171863 );
xor ( n4396 , n783 , n822 );
not ( n4397 , n4396 );
not ( n4398 , n1939 );
or ( n4399 , n4397 , n4398 );
buf ( n171869 , n171055 );
buf ( n171870 , n170170 );
nand ( n4402 , n171869 , n171870 );
buf ( n171872 , n4402 );
nand ( n4404 , n4399 , n171872 );
not ( n4405 , n4404 );
xor ( n4406 , n810 , n795 );
buf ( n171876 , n4406 );
not ( n4408 , n171876 );
buf ( n171878 , n168977 );
not ( n4410 , n171878 );
buf ( n171880 , n4410 );
buf ( n171881 , n171880 );
not ( n4413 , n171881 );
or ( n4414 , n4408 , n4413 );
buf ( n171884 , n168989 );
buf ( n171885 , n2731 );
nand ( n4417 , n171884 , n171885 );
buf ( n171887 , n4417 );
buf ( n171888 , n171887 );
nand ( n4420 , n4414 , n171888 );
buf ( n171890 , n4420 );
not ( n4422 , n171890 );
or ( n4423 , n4405 , n4422 );
buf ( n171893 , n171890 );
buf ( n171894 , n4404 );
nor ( n4426 , n171893 , n171894 );
buf ( n171896 , n4426 );
xor ( n4428 , n812 , n793 );
buf ( n171898 , n4428 );
not ( n4430 , n171898 );
buf ( n171900 , n1907 );
not ( n4432 , n171900 );
or ( n4433 , n4430 , n4432 );
buf ( n171903 , n3220 );
buf ( n171904 , n170222 );
nand ( n4436 , n171903 , n171904 );
buf ( n171906 , n4436 );
buf ( n171907 , n171906 );
nand ( n4439 , n4433 , n171907 );
buf ( n171909 , n4439 );
buf ( n171910 , n171909 );
not ( n4442 , n171910 );
buf ( n171912 , n4442 );
or ( n4444 , n171896 , n171912 );
nand ( n4445 , n4423 , n4444 );
buf ( n171915 , n791 );
buf ( n171916 , n814 );
xor ( n4448 , n171915 , n171916 );
buf ( n171918 , n4448 );
buf ( n171919 , n171918 );
not ( n4451 , n171919 );
buf ( n171921 , n169922 );
not ( n4453 , n171921 );
or ( n4454 , n4451 , n4453 );
buf ( n171924 , n169247 );
buf ( n171925 , n170137 );
nand ( n4457 , n171924 , n171925 );
buf ( n171927 , n4457 );
buf ( n171928 , n171927 );
nand ( n4460 , n4454 , n171928 );
buf ( n171930 , n4460 );
buf ( n171931 , n171930 );
not ( n4463 , n171931 );
buf ( n171933 , n781 );
buf ( n171934 , n824 );
xor ( n4466 , n171933 , n171934 );
buf ( n171936 , n4466 );
buf ( n171937 , n171936 );
not ( n4469 , n171937 );
buf ( n171939 , n170100 );
not ( n4471 , n171939 );
or ( n4472 , n4469 , n4471 );
buf ( n171942 , n170565 );
buf ( n171943 , n170108 );
nand ( n4475 , n171942 , n171943 );
buf ( n171945 , n4475 );
buf ( n171946 , n171945 );
nand ( n4478 , n4472 , n171946 );
buf ( n171948 , n4478 );
buf ( n171949 , n171948 );
not ( n4481 , n171949 );
or ( n4482 , n4463 , n4481 );
buf ( n171952 , n171948 );
buf ( n171953 , n171930 );
or ( n4485 , n171952 , n171953 );
buf ( n171955 , n789 );
buf ( n171956 , n816 );
xor ( n4488 , n171955 , n171956 );
buf ( n171958 , n4488 );
buf ( n171959 , n171958 );
not ( n4491 , n171959 );
buf ( n171961 , n169836 );
not ( n4493 , n171961 );
or ( n4494 , n4491 , n4493 );
buf ( n171964 , n169320 );
buf ( n171965 , n170153 );
nand ( n4497 , n171964 , n171965 );
buf ( n171967 , n4497 );
buf ( n171968 , n171967 );
nand ( n4500 , n4494 , n171968 );
buf ( n171970 , n4500 );
buf ( n171971 , n171970 );
nand ( n4503 , n4485 , n171971 );
buf ( n171973 , n4503 );
buf ( n171974 , n171973 );
nand ( n4506 , n4482 , n171974 );
buf ( n171976 , n4506 );
xor ( n4508 , n4445 , n171976 );
buf ( n171978 , n775 );
buf ( n171979 , n830 );
xor ( n4511 , n171978 , n171979 );
buf ( n171981 , n4511 );
buf ( n171982 , n171981 );
not ( n4514 , n171982 );
buf ( n171984 , n1471 );
not ( n4516 , n171984 );
or ( n4517 , n4514 , n4516 );
buf ( n171987 , n170191 );
buf ( n171988 , n831 );
nand ( n4520 , n171987 , n171988 );
buf ( n171990 , n4520 );
buf ( n171991 , n171990 );
nand ( n4523 , n4517 , n171991 );
buf ( n171993 , n4523 );
buf ( n171994 , n171993 );
buf ( n171995 , n797 );
buf ( n171996 , n808 );
xor ( n4528 , n171995 , n171996 );
buf ( n171998 , n4528 );
buf ( n171999 , n171998 );
not ( n4531 , n171999 );
buf ( n172001 , n169545 );
not ( n4533 , n172001 );
or ( n4534 , n4531 , n4533 );
buf ( n172004 , n168619 );
buf ( n172005 , n170246 );
nand ( n4537 , n172004 , n172005 );
buf ( n172007 , n4537 );
buf ( n172008 , n172007 );
nand ( n4540 , n4534 , n172008 );
buf ( n172010 , n4540 );
buf ( n172011 , n172010 );
xor ( n4543 , n171994 , n172011 );
not ( n4544 , n168656 );
not ( n4545 , n170264 );
or ( n4546 , n4544 , n4545 );
buf ( n172016 , n785 );
buf ( n172017 , n820 );
xnor ( n4549 , n172016 , n172017 );
buf ( n172019 , n4549 );
or ( n4551 , n169988 , n172019 );
nand ( n4552 , n4546 , n4551 );
buf ( n172022 , n4552 );
and ( n4554 , n4543 , n172022 );
and ( n4555 , n171994 , n172011 );
or ( n4556 , n4554 , n4555 );
buf ( n172026 , n4556 );
and ( n4558 , n4508 , n172026 );
and ( n4559 , n4445 , n171976 );
or ( n4560 , n4558 , n4559 );
buf ( n172030 , n4560 );
nand ( n4562 , n4395 , n172030 );
buf ( n172032 , n4562 );
buf ( n172033 , n172032 );
buf ( n172034 , n171849 );
buf ( n172035 , n4393 );
nand ( n4567 , n172034 , n172035 );
buf ( n172037 , n4567 );
buf ( n172038 , n172037 );
nand ( n4570 , n172033 , n172038 );
buf ( n172040 , n4570 );
buf ( n172041 , n172040 );
and ( n4573 , n4309 , n172041 );
and ( n4574 , n171692 , n171777 );
or ( n4575 , n4573 , n4574 );
buf ( n172045 , n4575 );
buf ( n172046 , n172045 );
not ( n4578 , n172046 );
buf ( n172048 , n4578 );
not ( n4580 , n172048 );
and ( n4581 , n4215 , n4580 );
buf ( n172051 , n172045 );
not ( n4583 , n172051 );
buf ( n172053 , n4214 );
nand ( n4585 , n4583 , n172053 );
buf ( n172055 , n4585 );
xor ( n4587 , n170054 , n170132 );
xor ( n4588 , n4587 , n170313 );
buf ( n172058 , n4588 );
buf ( n172059 , n172058 );
xor ( n4591 , n171717 , n171734 );
xor ( n4592 , n4591 , n171758 );
buf ( n172062 , n4592 );
not ( n4594 , n172062 );
buf ( n172064 , n4594 );
not ( n4596 , n172064 );
not ( n4597 , n170299 );
not ( n4598 , n4597 );
not ( n4599 , n170276 );
not ( n4600 , n4599 );
or ( n4601 , n4598 , n4600 );
nand ( n4602 , n170299 , n170276 );
nand ( n4603 , n4601 , n4602 );
buf ( n172073 , n170258 );
not ( n4605 , n172073 );
buf ( n172075 , n4605 );
or ( n4607 , n4603 , n172075 );
nand ( n4608 , n4603 , n172075 );
nand ( n4609 , n4607 , n4608 );
buf ( n172079 , n4609 );
not ( n4611 , n172079 );
or ( n4612 , n4596 , n4611 );
xor ( n4613 , n170149 , n170165 );
xor ( n4614 , n4613 , n170182 );
buf ( n4615 , n4614 );
buf ( n172085 , n4615 );
nand ( n4617 , n4612 , n172085 );
buf ( n172087 , n4617 );
buf ( n172088 , n172062 );
not ( n4620 , n4609 );
buf ( n172090 , n4620 );
nand ( n4622 , n172088 , n172090 );
buf ( n172092 , n4622 );
and ( n4624 , n172087 , n172092 );
buf ( n172094 , n4624 );
not ( n4626 , n172094 );
and ( n4627 , n2913 , n2867 );
not ( n4628 , n2913 );
and ( n4629 , n4628 , n2895 );
nor ( n4630 , n4627 , n4629 );
and ( n4631 , n4630 , n170359 );
not ( n4632 , n4630 );
and ( n4633 , n4632 , n170356 );
nor ( n4634 , n4631 , n4633 );
buf ( n172104 , n4634 );
not ( n4636 , n172104 );
or ( n4637 , n4626 , n4636 );
xor ( n4638 , n171763 , n171767 );
xor ( n4639 , n4638 , n171772 );
buf ( n172109 , n4639 );
buf ( n172110 , n172109 );
nand ( n4642 , n4637 , n172110 );
buf ( n172112 , n4642 );
buf ( n172113 , n172112 );
buf ( n172114 , n4634 );
not ( n4646 , n172114 );
buf ( n172116 , n172087 );
buf ( n172117 , n172092 );
nand ( n4649 , n172116 , n172117 );
buf ( n172119 , n4649 );
buf ( n172120 , n172119 );
nand ( n4652 , n4646 , n172120 );
buf ( n172122 , n4652 );
buf ( n172123 , n172122 );
nand ( n4655 , n172113 , n172123 );
buf ( n172125 , n4655 );
buf ( n172126 , n172125 );
xor ( n4658 , n172059 , n172126 );
buf ( n172128 , n170387 );
not ( n4660 , n172128 );
buf ( n172130 , n2859 );
not ( n4662 , n172130 );
or ( n4663 , n4660 , n4662 );
buf ( n172133 , n170387 );
buf ( n172134 , n2859 );
or ( n4666 , n172133 , n172134 );
nand ( n4667 , n4663 , n4666 );
buf ( n172137 , n4667 );
buf ( n172138 , n172137 );
buf ( n172139 , n170321 );
xor ( n4671 , n172138 , n172139 );
buf ( n172141 , n4671 );
buf ( n172142 , n172141 );
and ( n4674 , n4658 , n172142 );
and ( n4675 , n172059 , n172126 );
or ( n4676 , n4674 , n4675 );
buf ( n172146 , n4676 );
buf ( n4678 , n172146 );
and ( n4679 , n172055 , n4678 );
nor ( n4680 , n4581 , n4679 );
buf ( n172150 , n4680 );
not ( n4682 , n172150 );
buf ( n172152 , n4682 );
buf ( n172153 , n172152 );
and ( n4685 , n4208 , n172153 );
and ( n4686 , n171672 , n171676 );
or ( n4687 , n4685 , n4686 );
buf ( n172157 , n4687 );
not ( n4689 , n172157 );
and ( n4690 , n4202 , n4689 );
xor ( n4691 , n171672 , n171676 );
xor ( n4692 , n4691 , n172153 );
buf ( n172162 , n4692 );
buf ( n172163 , n172162 );
buf ( n172164 , n834 );
xor ( n4696 , n171692 , n171777 );
xor ( n4697 , n4696 , n172041 );
buf ( n172167 , n4697 );
buf ( n172168 , n172167 );
xor ( n4700 , n2716 , n4389 );
xnor ( n4701 , n4700 , n4560 );
not ( n4702 , n171849 );
and ( n4703 , n4701 , n4702 );
not ( n4704 , n4701 );
and ( n4705 , n4704 , n171849 );
nor ( n4706 , n4703 , n4705 );
not ( n4707 , n4706 );
xor ( n4708 , n4445 , n171976 );
xor ( n4709 , n4708 , n172026 );
buf ( n172179 , n4709 );
xor ( n4711 , n171782 , n171840 );
xor ( n4712 , n4711 , n171845 );
buf ( n172182 , n4712 );
buf ( n172183 , n172182 );
or ( n4715 , n172179 , n172183 );
and ( n4716 , n4614 , n172062 );
not ( n4717 , n4614 );
and ( n4718 , n4717 , n4594 );
nor ( n4719 , n4716 , n4718 );
buf ( n172189 , n4719 );
buf ( n172190 , n4620 );
and ( n4722 , n172189 , n172190 );
not ( n4723 , n172189 );
not ( n4724 , n4620 );
buf ( n172194 , n4724 );
and ( n4726 , n4723 , n172194 );
nor ( n4727 , n4722 , n4726 );
buf ( n172197 , n4727 );
buf ( n172198 , n172197 );
nand ( n4730 , n4715 , n172198 );
buf ( n172200 , n4730 );
buf ( n172201 , n172182 );
buf ( n172202 , n4709 );
nand ( n4734 , n172201 , n172202 );
buf ( n172204 , n4734 );
nand ( n4736 , n172200 , n172204 );
not ( n4737 , n4736 );
not ( n4738 , n4737 );
not ( n4739 , n4738 );
or ( n4740 , n4707 , n4739 );
or ( n4741 , n4738 , n4706 );
xor ( n4742 , n4404 , n171909 );
xor ( n4743 , n4742 , n171890 );
xor ( n4744 , n171994 , n172011 );
xor ( n4745 , n4744 , n172022 );
buf ( n172215 , n4745 );
xor ( n4747 , n4743 , n172215 );
xnor ( n4748 , n171948 , n171970 );
xnor ( n4749 , n171930 , n4748 );
and ( n4750 , n4747 , n4749 );
and ( n4751 , n4743 , n172215 );
or ( n4752 , n4750 , n4751 );
not ( n4753 , n4752 );
buf ( n172223 , n792 );
buf ( n172224 , n814 );
xor ( n4756 , n172223 , n172224 );
buf ( n172226 , n4756 );
buf ( n172227 , n172226 );
not ( n4759 , n172227 );
buf ( n172229 , n171013 );
not ( n4761 , n172229 );
or ( n4762 , n4759 , n4761 );
buf ( n172232 , n169250 );
buf ( n172233 , n171918 );
nand ( n4765 , n172232 , n172233 );
buf ( n172235 , n4765 );
buf ( n172236 , n172235 );
nand ( n4768 , n4762 , n172236 );
buf ( n172238 , n4768 );
buf ( n172239 , n172238 );
buf ( n172240 , n790 );
buf ( n172241 , n816 );
xor ( n4773 , n172240 , n172241 );
buf ( n172243 , n4773 );
buf ( n172244 , n172243 );
not ( n4776 , n172244 );
buf ( n172246 , n171029 );
not ( n4778 , n172246 );
or ( n4779 , n4776 , n4778 );
buf ( n172249 , n169845 );
buf ( n172250 , n171958 );
nand ( n4782 , n172249 , n172250 );
buf ( n172252 , n4782 );
buf ( n172253 , n172252 );
nand ( n4785 , n4779 , n172253 );
buf ( n172255 , n4785 );
buf ( n172256 , n172255 );
xor ( n4788 , n172239 , n172256 );
xor ( n4789 , n822 , n784 );
buf ( n172259 , n4789 );
not ( n4791 , n172259 );
buf ( n172261 , n169411 );
not ( n4793 , n172261 );
or ( n4794 , n4791 , n4793 );
nand ( n4795 , n169423 , n4396 );
buf ( n172265 , n4795 );
nand ( n4797 , n4794 , n172265 );
buf ( n172267 , n4797 );
buf ( n172268 , n172267 );
and ( n4800 , n4788 , n172268 );
and ( n4801 , n172239 , n172256 );
or ( n4802 , n4800 , n4801 );
buf ( n172272 , n4802 );
buf ( n172273 , n172272 );
not ( n4805 , n172273 );
buf ( n172275 , n4805 );
buf ( n172276 , n172275 );
xor ( n4808 , n830 , n776 );
buf ( n172278 , n4808 );
not ( n4810 , n172278 );
buf ( n172280 , n168471 );
not ( n4812 , n172280 );
or ( n4813 , n4810 , n4812 );
buf ( n172283 , n171981 );
buf ( n172284 , n831 );
nand ( n4816 , n172283 , n172284 );
buf ( n172286 , n4816 );
buf ( n172287 , n172286 );
nand ( n4819 , n4813 , n172287 );
buf ( n172289 , n4819 );
buf ( n172290 , n172289 );
xor ( n4822 , n810 , n796 );
buf ( n172292 , n4822 );
not ( n4824 , n172292 );
buf ( n172294 , n168980 );
not ( n4826 , n172294 );
or ( n4827 , n4824 , n4826 );
buf ( n172297 , n169957 );
buf ( n172298 , n4406 );
nand ( n4830 , n172297 , n172298 );
buf ( n172300 , n4830 );
buf ( n172301 , n172300 );
nand ( n4833 , n4827 , n172301 );
buf ( n172303 , n4833 );
buf ( n172304 , n172303 );
xor ( n4836 , n172290 , n172304 );
buf ( n172306 , n794 );
buf ( n172307 , n812 );
xor ( n4839 , n172306 , n172307 );
buf ( n172309 , n4839 );
buf ( n172310 , n172309 );
not ( n4842 , n172310 );
buf ( n172312 , n1907 );
not ( n4844 , n172312 );
or ( n4845 , n4842 , n4844 );
buf ( n172315 , n1534 );
buf ( n172316 , n4428 );
nand ( n4848 , n172315 , n172316 );
buf ( n172318 , n4848 );
buf ( n172319 , n172318 );
nand ( n4851 , n4845 , n172319 );
buf ( n172321 , n4851 );
buf ( n172322 , n172321 );
and ( n4854 , n4836 , n172322 );
and ( n4855 , n172290 , n172304 );
or ( n4856 , n4854 , n4855 );
buf ( n172326 , n4856 );
xor ( n4858 , n4285 , n4273 );
nor ( n4859 , n172326 , n4858 );
buf ( n172329 , n4859 );
or ( n4861 , n172276 , n172329 );
nand ( n4862 , n172326 , n4858 );
buf ( n172332 , n4862 );
nand ( n4864 , n4861 , n172332 );
buf ( n172334 , n4864 );
not ( n4866 , n172334 );
buf ( n172336 , n168719 );
buf ( n172337 , n799 );
and ( n4869 , n172336 , n172337 );
buf ( n172339 , n4869 );
buf ( n172340 , n172339 );
buf ( n172341 , n778 );
buf ( n172342 , n828 );
xor ( n4874 , n172341 , n172342 );
buf ( n172344 , n4874 );
buf ( n172345 , n172344 );
not ( n4877 , n172345 );
buf ( n172347 , n168549 );
not ( n4879 , n172347 );
or ( n4880 , n4877 , n4879 );
buf ( n172350 , n168559 );
buf ( n172351 , n4271 );
nand ( n4883 , n172350 , n172351 );
buf ( n172353 , n4883 );
buf ( n172354 , n172353 );
nand ( n4886 , n4880 , n172354 );
buf ( n172356 , n4886 );
buf ( n172357 , n172356 );
xor ( n4889 , n172340 , n172357 );
xor ( n4890 , n824 , n782 );
buf ( n172360 , n4890 );
not ( n4892 , n172360 );
buf ( n172362 , n1806 );
not ( n4894 , n172362 );
or ( n4895 , n4892 , n4894 );
buf ( n172365 , n170565 );
buf ( n172366 , n171936 );
nand ( n4898 , n172365 , n172366 );
buf ( n172368 , n4898 );
buf ( n172369 , n172368 );
nand ( n4901 , n4895 , n172369 );
buf ( n172371 , n4901 );
buf ( n172372 , n172371 );
and ( n4904 , n4889 , n172372 );
and ( n4905 , n172340 , n172357 );
or ( n4906 , n4904 , n4905 );
buf ( n172376 , n4906 );
buf ( n172377 , n172376 );
buf ( n172378 , n798 );
buf ( n172379 , n808 );
xor ( n4911 , n172378 , n172379 );
buf ( n172381 , n4911 );
buf ( n172382 , n172381 );
not ( n4914 , n172382 );
buf ( n172384 , n168615 );
not ( n4916 , n172384 );
or ( n4917 , n4914 , n4916 );
buf ( n172387 , n168619 );
buf ( n172388 , n171998 );
nand ( n4920 , n172387 , n172388 );
buf ( n172390 , n4920 );
buf ( n172391 , n172390 );
nand ( n4923 , n4917 , n172391 );
buf ( n172393 , n4923 );
buf ( n172394 , n172393 );
buf ( n172395 , n786 );
buf ( n172396 , n820 );
xor ( n4928 , n172395 , n172396 );
buf ( n172398 , n4928 );
not ( n4930 , n172398 );
not ( n4931 , n168648 );
or ( n4932 , n4930 , n4931 );
not ( n4933 , n172019 );
nand ( n4934 , n4933 , n171296 );
nand ( n4935 , n4932 , n4934 );
buf ( n172405 , n4935 );
xor ( n4937 , n172394 , n172405 );
not ( n4938 , n171803 );
or ( n4939 , n4938 , n169681 );
and ( n4940 , n826 , n780 );
not ( n4941 , n826 );
and ( n4942 , n4941 , n168631 );
nor ( n4943 , n4940 , n4942 );
nand ( n4944 , n4943 , n168666 );
nand ( n4945 , n4939 , n4944 );
buf ( n172415 , n4945 );
and ( n4947 , n4937 , n172415 );
and ( n4948 , n172394 , n172405 );
or ( n4949 , n4947 , n4948 );
buf ( n172419 , n4949 );
buf ( n172420 , n172419 );
xor ( n4952 , n172377 , n172420 );
xor ( n4953 , n171799 , n171817 );
xor ( n4954 , n4953 , n171835 );
buf ( n172424 , n4954 );
buf ( n172425 , n172424 );
and ( n4957 , n4952 , n172425 );
and ( n4958 , n172377 , n172420 );
or ( n4959 , n4957 , n4958 );
buf ( n172429 , n4959 );
not ( n4961 , n172429 );
nand ( n4962 , n4866 , n4961 );
not ( n4963 , n4962 );
or ( n4964 , n4753 , n4963 );
not ( n4965 , n4866 );
nand ( n4966 , n4965 , n172429 );
nand ( n4967 , n4964 , n4966 );
buf ( n4968 , n4967 );
nand ( n4969 , n4741 , n4968 );
nand ( n4970 , n4740 , n4969 );
buf ( n172440 , n4970 );
xor ( n4972 , n172168 , n172440 );
xor ( n4973 , n172059 , n172126 );
xor ( n4974 , n4973 , n172142 );
buf ( n172444 , n4974 );
buf ( n172445 , n172444 );
and ( n4977 , n4972 , n172445 );
and ( n4978 , n172168 , n172440 );
or ( n4979 , n4977 , n4978 );
buf ( n172449 , n4979 );
buf ( n172450 , n172449 );
xor ( n4982 , n172164 , n172450 );
not ( n4983 , n4214 );
buf ( n172453 , n4983 );
not ( n4985 , n172453 );
buf ( n172455 , n172146 );
not ( n4987 , n172455 );
buf ( n172457 , n172048 );
not ( n4989 , n172457 );
and ( n4990 , n4987 , n4989 );
buf ( n172460 , n172146 );
buf ( n172461 , n172048 );
and ( n4993 , n172460 , n172461 );
nor ( n4994 , n4990 , n4993 );
buf ( n172464 , n4994 );
buf ( n172465 , n172464 );
not ( n4997 , n172465 );
or ( n4998 , n4985 , n4997 );
buf ( n172468 , n172464 );
not ( n5000 , n172468 );
buf ( n172470 , n5000 );
buf ( n172471 , n172470 );
not ( n5003 , n4983 );
buf ( n172473 , n5003 );
nand ( n5005 , n172471 , n172473 );
buf ( n172475 , n5005 );
buf ( n172476 , n172475 );
nand ( n5008 , n4998 , n172476 );
buf ( n172478 , n5008 );
buf ( n172479 , n172478 );
and ( n5011 , n4982 , n172479 );
and ( n5012 , n172164 , n172450 );
or ( n5013 , n5011 , n5012 );
buf ( n172483 , n5013 );
buf ( n172484 , n172483 );
nor ( n5016 , n172163 , n172484 );
buf ( n172486 , n5016 );
nor ( n5018 , n4690 , n172486 );
buf ( n172488 , n5018 );
xor ( n5020 , n172164 , n172450 );
xor ( n5021 , n5020 , n172479 );
buf ( n172491 , n5021 );
buf ( n172492 , n172491 );
not ( n5024 , n172492 );
buf ( n172494 , n5024 );
buf ( n172495 , n172494 );
buf ( n172496 , n835 );
buf ( n172497 , n4634 );
not ( n5029 , n172497 );
buf ( n172499 , n5029 );
xor ( n5031 , n4624 , n172499 );
xnor ( n5032 , n5031 , n172109 );
buf ( n172502 , n5032 );
buf ( n172503 , n788 );
buf ( n172504 , n818 );
xor ( n5036 , n172503 , n172504 );
buf ( n172506 , n5036 );
buf ( n172507 , n172506 );
not ( n5039 , n172507 );
buf ( n172509 , n1321 );
not ( n5041 , n172509 );
or ( n5042 , n5039 , n5041 );
buf ( n172512 , n168806 );
buf ( n172513 , n171822 );
nand ( n5045 , n172512 , n172513 );
buf ( n172515 , n5045 );
buf ( n172516 , n172515 );
nand ( n5048 , n5042 , n172516 );
buf ( n172518 , n5048 );
buf ( n172519 , n172518 );
buf ( n172520 , n799 );
buf ( n172521 , n809 );
or ( n5053 , n172520 , n172521 );
buf ( n172523 , n810 );
nand ( n5055 , n5053 , n172523 );
buf ( n172525 , n5055 );
buf ( n172526 , n172525 );
buf ( n172527 , n799 );
buf ( n172528 , n809 );
nand ( n5060 , n172527 , n172528 );
buf ( n172530 , n5060 );
buf ( n172531 , n172530 );
buf ( n172532 , n808 );
and ( n5064 , n172526 , n172531 , n172532 );
buf ( n172534 , n5064 );
buf ( n172535 , n172534 );
buf ( n172536 , n779 );
buf ( n172537 , n828 );
xor ( n5069 , n172536 , n172537 );
buf ( n172539 , n5069 );
buf ( n172540 , n172539 );
not ( n5072 , n172540 );
buf ( n172542 , n168549 );
not ( n5074 , n172542 );
or ( n5075 , n5072 , n5074 );
buf ( n172545 , n168559 );
buf ( n172546 , n172344 );
nand ( n5078 , n172545 , n172546 );
buf ( n172548 , n5078 );
buf ( n172549 , n172548 );
nand ( n5081 , n5075 , n172549 );
buf ( n172551 , n5081 );
buf ( n172552 , n172551 );
and ( n5084 , n172535 , n172552 );
buf ( n172554 , n5084 );
buf ( n172555 , n172554 );
xor ( n5087 , n172519 , n172555 );
buf ( n172557 , n795 );
buf ( n172558 , n812 );
xor ( n5090 , n172557 , n172558 );
buf ( n172560 , n5090 );
buf ( n172561 , n172560 );
not ( n5093 , n172561 );
buf ( n172563 , n1553 );
not ( n5095 , n172563 );
or ( n5096 , n5093 , n5095 );
buf ( n172566 , n1534 );
buf ( n172567 , n172309 );
nand ( n5099 , n172566 , n172567 );
buf ( n172569 , n5099 );
buf ( n172570 , n172569 );
nand ( n5102 , n5096 , n172570 );
buf ( n172572 , n5102 );
buf ( n172573 , n172572 );
xor ( n5105 , n810 , n797 );
buf ( n172575 , n5105 );
not ( n5107 , n172575 );
buf ( n172577 , n169951 );
not ( n5109 , n172577 );
or ( n5110 , n5107 , n5109 );
buf ( n172580 , n168986 );
not ( n5112 , n172580 );
buf ( n172582 , n5112 );
buf ( n172583 , n172582 );
buf ( n172584 , n4822 );
nand ( n5116 , n172583 , n172584 );
buf ( n172586 , n5116 );
buf ( n172587 , n172586 );
nand ( n5119 , n5110 , n172587 );
buf ( n172589 , n5119 );
buf ( n172590 , n172589 );
xor ( n5122 , n172573 , n172590 );
xor ( n5123 , n822 , n785 );
buf ( n172593 , n5123 );
not ( n5125 , n172593 );
buf ( n172595 , n171049 );
not ( n5127 , n172595 );
or ( n5128 , n5125 , n5127 );
buf ( n172598 , n169423 );
buf ( n172599 , n4789 );
nand ( n5131 , n172598 , n172599 );
buf ( n172601 , n5131 );
buf ( n172602 , n172601 );
nand ( n5134 , n5128 , n172602 );
buf ( n172604 , n5134 );
buf ( n172605 , n172604 );
and ( n5137 , n5122 , n172605 );
and ( n5138 , n172573 , n172590 );
or ( n5139 , n5137 , n5138 );
buf ( n172609 , n5139 );
buf ( n172610 , n172609 );
and ( n5142 , n5087 , n172610 );
and ( n5143 , n172519 , n172555 );
or ( n5144 , n5142 , n5143 );
buf ( n172614 , n5144 );
buf ( n172615 , n172614 );
xor ( n5147 , n172377 , n172420 );
xor ( n5148 , n5147 , n172425 );
buf ( n172618 , n5148 );
buf ( n172619 , n172618 );
xor ( n5151 , n172615 , n172619 );
xor ( n5152 , n172340 , n172357 );
xor ( n5153 , n5152 , n172372 );
buf ( n172623 , n5153 );
buf ( n172624 , n172623 );
xor ( n5156 , n172290 , n172304 );
xor ( n5157 , n5156 , n172322 );
buf ( n172627 , n5157 );
buf ( n172628 , n172627 );
xor ( n5160 , n172624 , n172628 );
xor ( n5161 , n172239 , n172256 );
xor ( n5162 , n5161 , n172268 );
buf ( n172632 , n5162 );
buf ( n172633 , n172632 );
and ( n5165 , n5160 , n172633 );
and ( n5166 , n172624 , n172628 );
or ( n5167 , n5165 , n5166 );
buf ( n172637 , n5167 );
buf ( n172638 , n172637 );
and ( n5170 , n5151 , n172638 );
and ( n5171 , n172615 , n172619 );
or ( n5172 , n5170 , n5171 );
buf ( n172642 , n5172 );
buf ( n172643 , n172642 );
not ( n5175 , n831 );
not ( n5176 , n4808 );
or ( n5177 , n5175 , n5176 );
xor ( n5178 , n830 , n777 );
nand ( n5179 , n2048 , n5178 );
nand ( n5180 , n5177 , n5179 );
buf ( n172650 , n799 );
buf ( n172651 , n808 );
xor ( n5183 , n172650 , n172651 );
buf ( n172653 , n5183 );
buf ( n172654 , n172653 );
not ( n5186 , n172654 );
buf ( n172656 , n169545 );
not ( n5188 , n172656 );
or ( n5189 , n5186 , n5188 );
buf ( n172659 , n168619 );
buf ( n172660 , n172381 );
nand ( n5192 , n172659 , n172660 );
buf ( n172662 , n5192 );
buf ( n172663 , n172662 );
nand ( n5195 , n5189 , n172663 );
buf ( n172665 , n5195 );
xor ( n5197 , n5180 , n172665 );
buf ( n172667 , n781 );
buf ( n172668 , n826 );
xor ( n5200 , n172667 , n172668 );
buf ( n172670 , n5200 );
buf ( n172671 , n172670 );
not ( n5203 , n172671 );
buf ( n172673 , n4337 );
not ( n5205 , n172673 );
or ( n5206 , n5203 , n5205 );
buf ( n172676 , n168684 );
buf ( n172677 , n4943 );
nand ( n5209 , n172676 , n172677 );
buf ( n172679 , n5209 );
buf ( n172680 , n172679 );
nand ( n5212 , n5206 , n172680 );
buf ( n172682 , n5212 );
and ( n5214 , n5197 , n172682 );
and ( n5215 , n5180 , n172665 );
or ( n5216 , n5214 , n5215 );
buf ( n172686 , n793 );
buf ( n172687 , n814 );
xor ( n5219 , n172686 , n172687 );
buf ( n172689 , n5219 );
buf ( n172690 , n172689 );
not ( n5222 , n172690 );
buf ( n172692 , n3764 );
not ( n5224 , n172692 );
or ( n5225 , n5222 , n5224 );
buf ( n172695 , n169247 );
buf ( n172696 , n172226 );
nand ( n5228 , n172695 , n172696 );
buf ( n172698 , n5228 );
buf ( n172699 , n172698 );
nand ( n5231 , n5225 , n172699 );
buf ( n172701 , n5231 );
buf ( n172702 , n172701 );
xor ( n5234 , n824 , n783 );
buf ( n172704 , n5234 );
not ( n5236 , n172704 );
buf ( n172706 , n170100 );
not ( n5238 , n172706 );
or ( n5239 , n5236 , n5238 );
buf ( n172709 , n169802 );
buf ( n172710 , n4890 );
nand ( n5242 , n172709 , n172710 );
buf ( n172712 , n5242 );
buf ( n172713 , n172712 );
nand ( n5245 , n5239 , n172713 );
buf ( n172715 , n5245 );
buf ( n172716 , n172715 );
xor ( n5248 , n172702 , n172716 );
buf ( n172718 , n791 );
buf ( n172719 , n816 );
xor ( n5251 , n172718 , n172719 );
buf ( n172721 , n5251 );
buf ( n172722 , n172721 );
not ( n5254 , n172722 );
buf ( n172724 , n171029 );
not ( n5256 , n172724 );
or ( n5257 , n5254 , n5256 );
buf ( n172727 , n169320 );
buf ( n172728 , n172243 );
nand ( n5260 , n172727 , n172728 );
buf ( n172730 , n5260 );
buf ( n172731 , n172730 );
nand ( n5263 , n5257 , n172731 );
buf ( n172733 , n5263 );
buf ( n172734 , n172733 );
and ( n5266 , n5248 , n172734 );
and ( n5267 , n172702 , n172716 );
or ( n5268 , n5266 , n5267 );
buf ( n172738 , n5268 );
xor ( n5270 , n5216 , n172738 );
xor ( n5271 , n172394 , n172405 );
xor ( n5272 , n5271 , n172415 );
buf ( n172742 , n5272 );
and ( n5274 , n5270 , n172742 );
and ( n5275 , n5216 , n172738 );
or ( n5276 , n5274 , n5275 );
not ( n5277 , n5276 );
not ( n5278 , n172272 );
not ( n5279 , n4858 );
and ( n5280 , n5279 , n172326 );
not ( n5281 , n5279 );
not ( n5282 , n172326 );
and ( n5283 , n5281 , n5282 );
nor ( n5284 , n5280 , n5283 );
not ( n5285 , n5284 );
not ( n5286 , n5285 );
or ( n5287 , n5278 , n5286 );
nand ( n5288 , n172275 , n5284 );
nand ( n5289 , n5287 , n5288 );
not ( n5290 , n5289 );
not ( n5291 , n5290 );
or ( n5292 , n5277 , n5291 );
not ( n5293 , n5276 );
not ( n5294 , n5293 );
not ( n5295 , n5289 );
or ( n5296 , n5294 , n5295 );
xor ( n5297 , n4743 , n172215 );
xor ( n5298 , n5297 , n4749 );
nand ( n5299 , n5296 , n5298 );
nand ( n5300 , n5292 , n5299 );
buf ( n172770 , n5300 );
xor ( n5302 , n172643 , n172770 );
not ( n5303 , n172334 );
xor ( n5304 , n172429 , n5303 );
xnor ( n5305 , n5304 , n4752 );
buf ( n172775 , n5305 );
and ( n5307 , n5302 , n172775 );
and ( n5308 , n172643 , n172770 );
or ( n5309 , n5307 , n5308 );
buf ( n172779 , n5309 );
buf ( n172780 , n172779 );
xor ( n5312 , n172502 , n172780 );
not ( n5313 , n4736 );
not ( n5314 , n5313 );
not ( n5315 , n4967 );
or ( n5316 , n5314 , n5315 );
or ( n5317 , n4737 , n4967 );
nand ( n5318 , n5316 , n5317 );
and ( n5319 , n5318 , n4706 );
not ( n5320 , n5318 );
not ( n5321 , n4706 );
and ( n5322 , n5320 , n5321 );
nor ( n5323 , n5319 , n5322 );
buf ( n172793 , n5323 );
and ( n5325 , n5312 , n172793 );
and ( n5326 , n172502 , n172780 );
or ( n5327 , n5325 , n5326 );
buf ( n172797 , n5327 );
buf ( n172798 , n172797 );
xor ( n5330 , n172496 , n172798 );
xor ( n5331 , n172168 , n172440 );
xor ( n5332 , n5331 , n172445 );
buf ( n172802 , n5332 );
buf ( n172803 , n172802 );
and ( n5335 , n5330 , n172803 );
and ( n5336 , n172496 , n172798 );
or ( n5337 , n5335 , n5336 );
buf ( n172807 , n5337 );
buf ( n172808 , n172807 );
not ( n5340 , n172808 );
buf ( n172810 , n5340 );
buf ( n172811 , n172810 );
nand ( n5343 , n172495 , n172811 );
buf ( n172813 , n5343 );
buf ( n172814 , n172813 );
buf ( n172815 , n836 );
buf ( n172816 , n172197 );
buf ( n172817 , n4709 );
not ( n5349 , n172817 );
buf ( n172819 , n5349 );
buf ( n172820 , n172819 );
and ( n5352 , n172816 , n172820 );
not ( n5353 , n172816 );
buf ( n172823 , n4709 );
and ( n5355 , n5353 , n172823 );
nor ( n5356 , n5352 , n5355 );
buf ( n172826 , n5356 );
buf ( n172827 , n172826 );
buf ( n172828 , n172182 );
buf ( n5360 , n172828 );
buf ( n172830 , n5360 );
buf ( n172831 , n172830 );
not ( n5363 , n172831 );
buf ( n172833 , n5363 );
buf ( n172834 , n172833 );
and ( n5366 , n172827 , n172834 );
not ( n5367 , n172827 );
buf ( n172837 , n172830 );
and ( n5369 , n5367 , n172837 );
nor ( n5370 , n5366 , n5369 );
buf ( n172840 , n5370 );
buf ( n172841 , n172840 );
buf ( n172842 , n789 );
buf ( n172843 , n818 );
xor ( n5375 , n172842 , n172843 );
buf ( n172845 , n5375 );
buf ( n172846 , n172845 );
not ( n5378 , n172846 );
buf ( n172848 , n1321 );
not ( n5380 , n172848 );
or ( n5381 , n5378 , n5380 );
buf ( n172851 , n168806 );
buf ( n172852 , n172506 );
nand ( n5384 , n172851 , n172852 );
buf ( n172854 , n5384 );
buf ( n172855 , n172854 );
nand ( n5387 , n5381 , n172855 );
buf ( n172857 , n5387 );
buf ( n172858 , n172857 );
buf ( n172859 , n787 );
buf ( n172860 , n820 );
xor ( n5392 , n172859 , n172860 );
buf ( n172862 , n5392 );
buf ( n172863 , n172862 );
not ( n5395 , n172863 );
buf ( n172865 , n2108 );
not ( n5397 , n172865 );
or ( n5398 , n5395 , n5397 );
buf ( n172868 , n168656 );
buf ( n172869 , n172398 );
nand ( n5401 , n172868 , n172869 );
buf ( n172871 , n5401 );
buf ( n172872 , n172871 );
nand ( n5404 , n5398 , n172872 );
buf ( n172874 , n5404 );
buf ( n172875 , n172874 );
xor ( n5407 , n172858 , n172875 );
xor ( n5408 , n172535 , n172552 );
buf ( n172878 , n5408 );
buf ( n172879 , n172878 );
and ( n5411 , n5407 , n172879 );
and ( n5412 , n172858 , n172875 );
or ( n5413 , n5411 , n5412 );
buf ( n172883 , n5413 );
buf ( n172884 , n172883 );
xor ( n5416 , n824 , n784 );
buf ( n172886 , n5416 );
not ( n5418 , n172886 );
buf ( n172888 , n1806 );
not ( n5420 , n172888 );
or ( n5421 , n5418 , n5420 );
buf ( n172891 , n170565 );
buf ( n172892 , n5234 );
nand ( n5424 , n172891 , n172892 );
buf ( n172894 , n5424 );
buf ( n172895 , n172894 );
nand ( n5427 , n5421 , n172895 );
buf ( n172897 , n5427 );
buf ( n172898 , n172897 );
buf ( n172899 , n168619 );
not ( n5431 , n172899 );
buf ( n172901 , n168466 );
nor ( n5433 , n5431 , n172901 );
buf ( n172903 , n5433 );
buf ( n172904 , n172903 );
or ( n5436 , n172898 , n172904 );
not ( n5437 , n172539 );
not ( n5438 , n168559 );
or ( n5439 , n5437 , n5438 );
buf ( n172909 , n780 );
buf ( n172910 , n828 );
xor ( n5442 , n172909 , n172910 );
buf ( n172912 , n5442 );
nand ( n5444 , n172912 , n3683 );
nand ( n5445 , n5439 , n5444 );
buf ( n172915 , n5445 );
nand ( n5447 , n5436 , n172915 );
buf ( n172917 , n5447 );
buf ( n172918 , n172917 );
buf ( n172919 , n172897 );
buf ( n172920 , n168619 );
buf ( n172921 , n799 );
and ( n5453 , n172920 , n172921 );
buf ( n172923 , n5453 );
buf ( n172924 , n172923 );
nand ( n5456 , n172919 , n172924 );
buf ( n172926 , n5456 );
buf ( n172927 , n172926 );
nand ( n5459 , n172918 , n172927 );
buf ( n172929 , n5459 );
buf ( n172930 , n172929 );
not ( n5462 , n2048 );
buf ( n172932 , n778 );
buf ( n172933 , n830 );
xor ( n5465 , n172932 , n172933 );
buf ( n172935 , n5465 );
not ( n5467 , n172935 );
or ( n5468 , n5462 , n5467 );
nand ( n5469 , n5178 , n831 );
nand ( n5470 , n5468 , n5469 );
buf ( n172940 , n5470 );
buf ( n172941 , n796 );
buf ( n172942 , n812 );
xor ( n5474 , n172941 , n172942 );
buf ( n172944 , n5474 );
buf ( n172945 , n172944 );
not ( n5477 , n172945 );
buf ( n172947 , n1553 );
not ( n5479 , n172947 );
or ( n5480 , n5477 , n5479 );
buf ( n172950 , n1534 );
buf ( n172951 , n172560 );
nand ( n5483 , n172950 , n172951 );
buf ( n172953 , n5483 );
buf ( n172954 , n172953 );
nand ( n5486 , n5480 , n172954 );
buf ( n172956 , n5486 );
buf ( n172957 , n172956 );
xor ( n5489 , n172940 , n172957 );
xor ( n5490 , n810 , n798 );
buf ( n172960 , n5490 );
not ( n5492 , n172960 );
buf ( n172962 , n169951 );
not ( n5494 , n172962 );
or ( n5495 , n5492 , n5494 );
buf ( n172965 , n168989 );
buf ( n172966 , n5105 );
nand ( n5498 , n172965 , n172966 );
buf ( n172968 , n5498 );
buf ( n172969 , n172968 );
nand ( n5501 , n5495 , n172969 );
buf ( n172971 , n5501 );
buf ( n172972 , n172971 );
and ( n5504 , n5489 , n172972 );
and ( n5505 , n172940 , n172957 );
or ( n5506 , n5504 , n5505 );
buf ( n172976 , n5506 );
buf ( n172977 , n172976 );
xor ( n5509 , n172930 , n172977 );
buf ( n172979 , n782 );
buf ( n172980 , n826 );
xor ( n5512 , n172979 , n172980 );
buf ( n172982 , n5512 );
buf ( n172983 , n172982 );
not ( n5515 , n172983 );
buf ( n172985 , n169674 );
not ( n5517 , n172985 );
or ( n5518 , n5515 , n5517 );
buf ( n172988 , n168684 );
buf ( n172989 , n172670 );
nand ( n5521 , n172988 , n172989 );
buf ( n172991 , n5521 );
buf ( n172992 , n172991 );
nand ( n5524 , n5518 , n172992 );
buf ( n172994 , n5524 );
not ( n5526 , n172994 );
buf ( n172996 , n5526 );
not ( n5528 , n172996 );
buf ( n172998 , n788 );
buf ( n172999 , n820 );
xor ( n5531 , n172998 , n172999 );
buf ( n173001 , n5531 );
not ( n5533 , n173001 );
not ( n5534 , n168648 );
or ( n5535 , n5533 , n5534 );
buf ( n173005 , n172862 );
buf ( n173006 , n171296 );
nand ( n5538 , n173005 , n173006 );
buf ( n173008 , n5538 );
nand ( n5540 , n5535 , n173008 );
not ( n5541 , n5540 );
buf ( n173011 , n5541 );
not ( n5543 , n173011 );
or ( n5544 , n5528 , n5543 );
buf ( n173014 , n790 );
buf ( n173015 , n818 );
xor ( n5547 , n173014 , n173015 );
buf ( n173017 , n5547 );
buf ( n173018 , n173017 );
not ( n5550 , n173018 );
buf ( n173020 , n1321 );
not ( n5552 , n173020 );
or ( n5553 , n5550 , n5552 );
buf ( n173023 , n168806 );
buf ( n173024 , n172845 );
nand ( n5556 , n173023 , n173024 );
buf ( n173026 , n5556 );
buf ( n173027 , n173026 );
nand ( n5559 , n5553 , n173027 );
buf ( n173029 , n5559 );
buf ( n173030 , n173029 );
nand ( n5562 , n5544 , n173030 );
buf ( n173032 , n5562 );
buf ( n173033 , n173032 );
buf ( n173034 , n5540 );
buf ( n173035 , n172994 );
nand ( n5567 , n173034 , n173035 );
buf ( n173037 , n5567 );
buf ( n173038 , n173037 );
nand ( n5570 , n173033 , n173038 );
buf ( n173040 , n5570 );
buf ( n173041 , n173040 );
and ( n5573 , n5509 , n173041 );
and ( n5574 , n172930 , n172977 );
or ( n5575 , n5573 , n5574 );
buf ( n173045 , n5575 );
buf ( n173046 , n173045 );
xor ( n5578 , n172884 , n173046 );
xor ( n5579 , n172519 , n172555 );
xor ( n5580 , n5579 , n172610 );
buf ( n173050 , n5580 );
buf ( n173051 , n173050 );
and ( n5583 , n5578 , n173051 );
and ( n5584 , n172884 , n173046 );
or ( n5585 , n5583 , n5584 );
buf ( n173055 , n5585 );
buf ( n173056 , n173055 );
xor ( n5588 , n172615 , n172619 );
xor ( n5589 , n5588 , n172638 );
buf ( n173059 , n5589 );
buf ( n173060 , n173059 );
xor ( n5592 , n173056 , n173060 );
xor ( n5593 , n172624 , n172628 );
xor ( n5594 , n5593 , n172633 );
buf ( n173064 , n5594 );
not ( n5596 , n173064 );
not ( n5597 , n5596 );
not ( n5598 , n5597 );
xor ( n5599 , n5180 , n172665 );
xor ( n5600 , n5599 , n172682 );
buf ( n173070 , n5600 );
buf ( n173071 , n792 );
buf ( n173072 , n816 );
xor ( n5604 , n173071 , n173072 );
buf ( n173074 , n5604 );
buf ( n173075 , n173074 );
not ( n5607 , n173075 );
buf ( n173077 , n169314 );
not ( n5609 , n173077 );
or ( n5610 , n5607 , n5609 );
buf ( n173080 , n169845 );
buf ( n173081 , n172721 );
nand ( n5613 , n173080 , n173081 );
buf ( n173083 , n5613 );
buf ( n173084 , n173083 );
nand ( n5616 , n5610 , n173084 );
buf ( n173086 , n5616 );
buf ( n173087 , n173086 );
not ( n5619 , n173087 );
buf ( n173089 , n5619 );
buf ( n173090 , n173089 );
buf ( n5622 , n173090 );
buf ( n173092 , n5622 );
buf ( n173093 , n173092 );
buf ( n173094 , n794 );
buf ( n173095 , n814 );
xor ( n5627 , n173094 , n173095 );
buf ( n173097 , n5627 );
buf ( n173098 , n173097 );
not ( n5630 , n173098 );
buf ( n173100 , n169241 );
not ( n5632 , n173100 );
or ( n5633 , n5630 , n5632 );
buf ( n173103 , n169247 );
buf ( n173104 , n172689 );
nand ( n5636 , n173103 , n173104 );
buf ( n173106 , n5636 );
buf ( n173107 , n173106 );
nand ( n5639 , n5633 , n173107 );
buf ( n173109 , n5639 );
buf ( n173110 , n173109 );
xor ( n5642 , n822 , n786 );
buf ( n173112 , n5642 );
not ( n5644 , n173112 );
buf ( n173114 , n1939 );
not ( n5646 , n173114 );
or ( n5647 , n5644 , n5646 );
buf ( n173117 , n169423 );
buf ( n173118 , n5123 );
nand ( n5650 , n173117 , n173118 );
buf ( n173120 , n5650 );
buf ( n173121 , n173120 );
nand ( n5653 , n5647 , n173121 );
buf ( n173123 , n5653 );
buf ( n173124 , n173123 );
nor ( n5656 , n173110 , n173124 );
buf ( n173126 , n5656 );
buf ( n173127 , n173126 );
or ( n5659 , n173093 , n173127 );
buf ( n173129 , n173109 );
buf ( n173130 , n173123 );
nand ( n5662 , n173129 , n173130 );
buf ( n173132 , n5662 );
buf ( n173133 , n173132 );
nand ( n5665 , n5659 , n173133 );
buf ( n173135 , n5665 );
buf ( n173136 , n173135 );
xor ( n5668 , n173070 , n173136 );
xor ( n5669 , n172573 , n172590 );
xor ( n5670 , n5669 , n172605 );
buf ( n173140 , n5670 );
buf ( n173141 , n173140 );
and ( n5673 , n5668 , n173141 );
and ( n5674 , n173070 , n173136 );
or ( n5675 , n5673 , n5674 );
buf ( n173145 , n5675 );
not ( n5677 , n173145 );
or ( n5678 , n5598 , n5677 );
not ( n5679 , n173145 );
not ( n5680 , n5679 );
not ( n5681 , n5596 );
or ( n5682 , n5680 , n5681 );
xor ( n5683 , n5216 , n172738 );
xor ( n5684 , n5683 , n172742 );
nand ( n5685 , n5682 , n5684 );
nand ( n5686 , n5678 , n5685 );
buf ( n173156 , n5686 );
and ( n5688 , n5592 , n173156 );
and ( n5689 , n173056 , n173060 );
or ( n5690 , n5688 , n5689 );
buf ( n173160 , n5690 );
buf ( n173161 , n173160 );
xor ( n5693 , n172841 , n173161 );
xor ( n5694 , n172643 , n172770 );
xor ( n5695 , n5694 , n172775 );
buf ( n173165 , n5695 );
buf ( n173166 , n173165 );
and ( n5698 , n5693 , n173166 );
and ( n5699 , n172841 , n173161 );
or ( n5700 , n5698 , n5699 );
buf ( n173170 , n5700 );
buf ( n173171 , n173170 );
xor ( n5703 , n172815 , n173171 );
xor ( n5704 , n172502 , n172780 );
xor ( n5705 , n5704 , n172793 );
buf ( n173175 , n5705 );
buf ( n173176 , n173175 );
and ( n5708 , n5703 , n173176 );
and ( n5709 , n172815 , n173171 );
or ( n5710 , n5708 , n5709 );
buf ( n173180 , n5710 );
not ( n5712 , n173180 );
xor ( n5713 , n172496 , n172798 );
xor ( n5714 , n5713 , n172803 );
buf ( n173184 , n5714 );
buf ( n173185 , n173184 );
not ( n5717 , n173185 );
buf ( n173187 , n5717 );
nand ( n5719 , n5712 , n173187 );
buf ( n173189 , n5719 );
nand ( n5721 , n172814 , n173189 );
buf ( n173191 , n5721 );
buf ( n173192 , n173191 );
not ( n5724 , n173192 );
buf ( n173194 , n5724 );
buf ( n173195 , n173194 );
nand ( n5727 , n172488 , n173195 );
buf ( n173197 , n5727 );
buf ( n173198 , n173197 );
not ( n5730 , n173198 );
buf ( n173200 , n837 );
buf ( n173201 , n5298 );
not ( n5733 , n173201 );
buf ( n173203 , n5733 );
not ( n5735 , n5293 );
not ( n5736 , n5290 );
or ( n5737 , n5735 , n5736 );
nand ( n5738 , n5289 , n5276 );
nand ( n5739 , n5737 , n5738 );
or ( n5740 , n173203 , n5739 );
nand ( n5741 , n5739 , n173203 );
nand ( n5742 , n5740 , n5741 );
buf ( n173212 , n5742 );
xor ( n5744 , n172702 , n172716 );
xor ( n5745 , n5744 , n172734 );
buf ( n173215 , n5745 );
buf ( n173216 , n173215 );
xor ( n5748 , n172858 , n172875 );
xor ( n5749 , n5748 , n172879 );
buf ( n173219 , n5749 );
buf ( n173220 , n173219 );
xor ( n5752 , n173216 , n173220 );
buf ( n173222 , n799 );
buf ( n173223 , n811 );
or ( n5755 , n173222 , n173223 );
buf ( n173225 , n812 );
nand ( n5757 , n5755 , n173225 );
buf ( n173227 , n5757 );
buf ( n173228 , n173227 );
buf ( n173229 , n799 );
buf ( n173230 , n811 );
nand ( n5762 , n173229 , n173230 );
buf ( n173232 , n5762 );
buf ( n173233 , n173232 );
buf ( n173234 , n810 );
and ( n5766 , n173228 , n173233 , n173234 );
buf ( n173236 , n5766 );
buf ( n173237 , n173236 );
xor ( n5769 , n828 , n781 );
buf ( n173239 , n5769 );
not ( n5771 , n173239 );
buf ( n173241 , n168549 );
not ( n5773 , n173241 );
or ( n5774 , n5771 , n5773 );
buf ( n173244 , n168559 );
buf ( n173245 , n172912 );
nand ( n5777 , n173244 , n173245 );
buf ( n173247 , n5777 );
buf ( n173248 , n173247 );
nand ( n5780 , n5774 , n173248 );
buf ( n173250 , n5780 );
buf ( n173251 , n173250 );
and ( n5783 , n173237 , n173251 );
buf ( n173253 , n5783 );
xor ( n5785 , n822 , n787 );
buf ( n173255 , n5785 );
not ( n5787 , n173255 );
buf ( n173257 , n1939 );
not ( n5789 , n173257 );
or ( n5790 , n5787 , n5789 );
buf ( n173260 , n169417 );
buf ( n173261 , n5642 );
nand ( n5793 , n173260 , n173261 );
buf ( n173263 , n5793 );
buf ( n173264 , n173263 );
nand ( n5796 , n5790 , n173264 );
buf ( n173266 , n5796 );
xor ( n5798 , n812 , n797 );
buf ( n173268 , n5798 );
not ( n5800 , n173268 );
buf ( n173270 , n1553 );
not ( n5802 , n173270 );
or ( n5803 , n5800 , n5802 );
buf ( n173273 , n1534 );
buf ( n173274 , n172944 );
nand ( n5806 , n173273 , n173274 );
buf ( n173276 , n5806 );
buf ( n173277 , n173276 );
nand ( n5809 , n5803 , n173277 );
buf ( n173279 , n5809 );
or ( n5811 , n173266 , n173279 );
not ( n5812 , n5811 );
buf ( n173282 , n810 );
not ( n5814 , n173282 );
buf ( n173284 , n799 );
nand ( n5816 , n5814 , n173284 );
buf ( n173286 , n5816 );
buf ( n173287 , n173286 );
not ( n5819 , n173287 );
buf ( n173289 , n799 );
not ( n5821 , n173289 );
buf ( n173291 , n810 );
nand ( n5823 , n5821 , n173291 );
buf ( n173293 , n5823 );
buf ( n173294 , n173293 );
not ( n5826 , n173294 );
or ( n5827 , n5819 , n5826 );
buf ( n173297 , n169951 );
nand ( n5829 , n5827 , n173297 );
buf ( n173299 , n5829 );
buf ( n173300 , n173299 );
buf ( n173301 , n172582 );
buf ( n173302 , n5490 );
nand ( n5834 , n173301 , n173302 );
buf ( n173304 , n5834 );
buf ( n173305 , n173304 );
nand ( n5837 , n173300 , n173305 );
buf ( n173307 , n5837 );
not ( n5839 , n173307 );
or ( n5840 , n5812 , n5839 );
nand ( n5841 , n173279 , n173266 );
nand ( n5842 , n5840 , n5841 );
nand ( n5843 , n173253 , n5842 );
buf ( n173313 , n779 );
buf ( n173314 , n830 );
xor ( n5846 , n173313 , n173314 );
buf ( n173316 , n5846 );
buf ( n173317 , n173316 );
not ( n5849 , n173317 );
buf ( n173319 , n168471 );
not ( n5851 , n173319 );
or ( n5852 , n5849 , n5851 );
buf ( n173322 , n172935 );
buf ( n173323 , n831 );
nand ( n5855 , n173322 , n173323 );
buf ( n173325 , n5855 );
buf ( n173326 , n173325 );
nand ( n5858 , n5852 , n173326 );
buf ( n173328 , n5858 );
buf ( n173329 , n173328 );
buf ( n173330 , n783 );
buf ( n173331 , n826 );
xor ( n5863 , n173330 , n173331 );
buf ( n173333 , n5863 );
buf ( n173334 , n173333 );
not ( n5866 , n173334 );
buf ( n173336 , n4337 );
not ( n5868 , n173336 );
or ( n5869 , n5866 , n5868 );
buf ( n173339 , n168684 );
buf ( n173340 , n172982 );
nand ( n5872 , n173339 , n173340 );
buf ( n173342 , n5872 );
buf ( n173343 , n173342 );
nand ( n5875 , n5869 , n173343 );
buf ( n173345 , n5875 );
buf ( n173346 , n173345 );
xor ( n5878 , n173329 , n173346 );
not ( n5879 , n168656 );
not ( n5880 , n173001 );
or ( n5881 , n5879 , n5880 );
buf ( n173351 , n789 );
buf ( n173352 , n820 );
xor ( n5884 , n173351 , n173352 );
buf ( n173354 , n5884 );
buf ( n173355 , n173354 );
not ( n5887 , n173355 );
buf ( n173357 , n5887 );
or ( n5889 , n169988 , n173357 );
nand ( n5890 , n5881 , n5889 );
buf ( n173360 , n5890 );
and ( n5892 , n5878 , n173360 );
and ( n5893 , n173329 , n173346 );
or ( n5894 , n5892 , n5893 );
buf ( n173364 , n5894 );
nand ( n5896 , n173253 , n173364 );
nand ( n5897 , n5842 , n173364 );
nand ( n5898 , n5843 , n5896 , n5897 );
buf ( n173368 , n5898 );
and ( n5900 , n5752 , n173368 );
and ( n5901 , n173216 , n173220 );
or ( n5902 , n5900 , n5901 );
buf ( n173372 , n5902 );
buf ( n173373 , n173372 );
xor ( n5905 , n172884 , n173046 );
xor ( n5906 , n5905 , n173051 );
buf ( n173376 , n5906 );
buf ( n173377 , n173376 );
xor ( n5909 , n173373 , n173377 );
xor ( n5910 , n172930 , n172977 );
xor ( n5911 , n5910 , n173041 );
buf ( n173381 , n5911 );
buf ( n173382 , n173381 );
buf ( n173383 , n173109 );
buf ( n173384 , n173089 );
and ( n5916 , n173383 , n173384 );
not ( n5917 , n173383 );
buf ( n173387 , n173086 );
and ( n5919 , n5917 , n173387 );
nor ( n5920 , n5916 , n5919 );
buf ( n173390 , n5920 );
not ( n5922 , n173390 );
and ( n5923 , n5922 , n173123 );
not ( n5924 , n5922 );
not ( n5925 , n173123 );
and ( n5926 , n5924 , n5925 );
nor ( n5927 , n5923 , n5926 );
not ( n5928 , n5927 );
buf ( n173398 , n173097 );
not ( n5930 , n173398 );
buf ( n173400 , n169250 );
not ( n5932 , n173400 );
or ( n5933 , n5930 , n5932 );
buf ( n173403 , n171013 );
xor ( n5935 , n814 , n795 );
buf ( n173405 , n5935 );
nand ( n5937 , n173403 , n173405 );
buf ( n173407 , n5937 );
buf ( n173408 , n173407 );
nand ( n5940 , n5933 , n173408 );
buf ( n173410 , n5940 );
not ( n5942 , n173410 );
xor ( n5943 , n824 , n785 );
buf ( n173413 , n5943 );
not ( n5945 , n173413 );
buf ( n173415 , n169793 );
not ( n5947 , n173415 );
or ( n5948 , n5945 , n5947 );
buf ( n173418 , n169169 );
buf ( n173419 , n5416 );
nand ( n5951 , n173418 , n173419 );
buf ( n173421 , n5951 );
buf ( n173422 , n173421 );
nand ( n5954 , n5948 , n173422 );
buf ( n173424 , n5954 );
not ( n5956 , n173424 );
buf ( n173426 , n793 );
buf ( n173427 , n816 );
xor ( n5959 , n173426 , n173427 );
buf ( n173429 , n5959 );
buf ( n173430 , n173429 );
not ( n5962 , n173430 );
xnor ( n5963 , n817 , n816 );
nor ( n5964 , n5963 , n169310 );
buf ( n173434 , n5964 );
not ( n5966 , n173434 );
or ( n5967 , n5962 , n5966 );
buf ( n173437 , n169842 );
buf ( n173438 , n173074 );
nand ( n5970 , n173437 , n173438 );
buf ( n173440 , n5970 );
buf ( n173441 , n173440 );
nand ( n5973 , n5967 , n173441 );
buf ( n173443 , n5973 );
not ( n5975 , n173443 );
nand ( n5976 , n5956 , n5975 );
not ( n5977 , n5976 );
or ( n5978 , n5942 , n5977 );
not ( n5979 , n5975 );
nand ( n5980 , n5979 , n173424 );
nand ( n5981 , n5978 , n5980 );
not ( n5982 , n5981 );
or ( n5983 , n5928 , n5982 );
not ( n5984 , n5981 );
not ( n5985 , n5984 );
not ( n5986 , n5925 );
not ( n5987 , n173390 );
or ( n5988 , n5986 , n5987 );
not ( n5989 , n5922 );
or ( n5990 , n5925 , n5989 );
nand ( n5991 , n5988 , n5990 );
not ( n5992 , n5991 );
or ( n5993 , n5985 , n5992 );
and ( n5994 , n5541 , n5526 );
not ( n5995 , n5541 );
and ( n5996 , n5995 , n172994 );
nor ( n5997 , n5994 , n5996 );
not ( n5998 , n173029 );
xor ( n5999 , n5997 , n5998 );
buf ( n173469 , n5999 );
not ( n6001 , n173469 );
buf ( n173471 , n6001 );
nand ( n6003 , n5993 , n173471 );
nand ( n6004 , n5983 , n6003 );
buf ( n173474 , n6004 );
xor ( n6006 , n173382 , n173474 );
xor ( n6007 , n173070 , n173136 );
xor ( n6008 , n6007 , n173141 );
buf ( n173478 , n6008 );
buf ( n173479 , n173478 );
and ( n6011 , n6006 , n173479 );
and ( n6012 , n173382 , n173474 );
or ( n6013 , n6011 , n6012 );
buf ( n173483 , n6013 );
buf ( n173484 , n173483 );
and ( n6016 , n5909 , n173484 );
and ( n6017 , n173373 , n173377 );
or ( n6018 , n6016 , n6017 );
buf ( n173488 , n6018 );
buf ( n173489 , n173488 );
xor ( n6021 , n173212 , n173489 );
xor ( n6022 , n173056 , n173060 );
xor ( n6023 , n6022 , n173156 );
buf ( n173493 , n6023 );
buf ( n173494 , n173493 );
and ( n6026 , n6021 , n173494 );
and ( n6027 , n173212 , n173489 );
or ( n6028 , n6026 , n6027 );
buf ( n173498 , n6028 );
buf ( n173499 , n173498 );
xor ( n6031 , n173200 , n173499 );
xor ( n6032 , n172841 , n173161 );
xor ( n6033 , n6032 , n173166 );
buf ( n173503 , n6033 );
buf ( n173504 , n173503 );
xor ( n6036 , n6031 , n173504 );
buf ( n173506 , n6036 );
buf ( n173507 , n173506 );
buf ( n173508 , n838 );
xor ( n6040 , n5684 , n173145 );
xor ( n6041 , n6040 , n5597 );
buf ( n173511 , n6041 );
xor ( n6043 , n5445 , n172923 );
xor ( n6044 , n6043 , n172897 );
buf ( n173514 , n6044 );
xor ( n6046 , n172940 , n172957 );
xor ( n6047 , n6046 , n172972 );
buf ( n173517 , n6047 );
buf ( n173518 , n173517 );
xor ( n6050 , n173514 , n173518 );
buf ( n173520 , n791 );
buf ( n173521 , n818 );
xor ( n6053 , n173520 , n173521 );
buf ( n173523 , n6053 );
buf ( n173524 , n173523 );
not ( n6056 , n173524 );
buf ( n173526 , n1321 );
not ( n6058 , n173526 );
or ( n6059 , n6056 , n6058 );
buf ( n173529 , n168806 );
buf ( n173530 , n173017 );
nand ( n6062 , n173529 , n173530 );
buf ( n173532 , n6062 );
buf ( n173533 , n173532 );
nand ( n6065 , n6059 , n173533 );
buf ( n173535 , n6065 );
buf ( n173536 , n173535 );
xor ( n6068 , n173237 , n173251 );
buf ( n173538 , n6068 );
buf ( n173539 , n173538 );
xor ( n6071 , n173536 , n173539 );
xor ( n6072 , n794 , n816 );
not ( n6073 , n6072 );
not ( n6074 , n5964 );
or ( n6075 , n6073 , n6074 );
buf ( n173545 , n169842 );
buf ( n173546 , n173429 );
nand ( n6078 , n173545 , n173546 );
buf ( n173548 , n6078 );
nand ( n6080 , n6075 , n173548 );
buf ( n173550 , n6080 );
buf ( n173551 , n796 );
buf ( n173552 , n814 );
xor ( n6084 , n173551 , n173552 );
buf ( n173554 , n6084 );
buf ( n173555 , n173554 );
not ( n6087 , n173555 );
buf ( n173557 , n3764 );
not ( n6089 , n173557 );
or ( n6090 , n6087 , n6089 );
buf ( n173560 , n169247 );
buf ( n173561 , n5935 );
nand ( n6093 , n173560 , n173561 );
buf ( n173563 , n6093 );
buf ( n173564 , n173563 );
nand ( n6096 , n6090 , n173564 );
buf ( n173566 , n6096 );
buf ( n173567 , n173566 );
xor ( n6099 , n173550 , n173567 );
buf ( n173569 , n782 );
buf ( n173570 , n828 );
xor ( n6102 , n173569 , n173570 );
buf ( n173572 , n6102 );
buf ( n173573 , n173572 );
not ( n6105 , n173573 );
buf ( n173575 , n1742 );
not ( n6107 , n173575 );
or ( n6108 , n6105 , n6107 );
buf ( n173578 , n168559 );
buf ( n173579 , n5769 );
nand ( n6111 , n173578 , n173579 );
buf ( n173581 , n6111 );
buf ( n173582 , n173581 );
nand ( n6114 , n6108 , n173582 );
buf ( n173584 , n6114 );
buf ( n173585 , n173584 );
and ( n6117 , n6099 , n173585 );
and ( n6118 , n173550 , n173567 );
or ( n6119 , n6117 , n6118 );
buf ( n173589 , n6119 );
buf ( n173590 , n173589 );
and ( n6122 , n6071 , n173590 );
and ( n6123 , n173536 , n173539 );
or ( n6124 , n6122 , n6123 );
buf ( n173594 , n6124 );
buf ( n173595 , n173594 );
and ( n6127 , n6050 , n173595 );
and ( n6128 , n173514 , n173518 );
or ( n6129 , n6127 , n6128 );
buf ( n173599 , n6129 );
buf ( n173600 , n173599 );
xor ( n6132 , n173216 , n173220 );
xor ( n6133 , n6132 , n173368 );
buf ( n173603 , n6133 );
buf ( n173604 , n173603 );
xor ( n6136 , n173600 , n173604 );
xor ( n6137 , n173382 , n173474 );
xor ( n6138 , n6137 , n173479 );
buf ( n173608 , n6138 );
buf ( n173609 , n173608 );
and ( n6141 , n6136 , n173609 );
and ( n6142 , n173600 , n173604 );
or ( n6143 , n6141 , n6142 );
buf ( n173613 , n6143 );
buf ( n173614 , n173613 );
xor ( n6146 , n173511 , n173614 );
xor ( n6147 , n173373 , n173377 );
xor ( n6148 , n6147 , n173484 );
buf ( n173618 , n6148 );
buf ( n173619 , n173618 );
and ( n6151 , n6146 , n173619 );
and ( n6152 , n173511 , n173614 );
or ( n6153 , n6151 , n6152 );
buf ( n173623 , n6153 );
buf ( n173624 , n173623 );
xor ( n6156 , n173508 , n173624 );
xor ( n6157 , n173212 , n173489 );
xor ( n6158 , n6157 , n173494 );
buf ( n173628 , n6158 );
buf ( n173629 , n173628 );
and ( n6161 , n6156 , n173629 );
and ( n6162 , n173508 , n173624 );
or ( n6163 , n6161 , n6162 );
buf ( n173633 , n6163 );
buf ( n173634 , n173633 );
nand ( n6166 , n173507 , n173634 );
buf ( n173636 , n6166 );
buf ( n173637 , n173636 );
not ( n6169 , n173637 );
buf ( n173639 , n6169 );
not ( n6171 , n173639 );
xor ( n6172 , n172815 , n173171 );
xor ( n6173 , n6172 , n173176 );
buf ( n173643 , n6173 );
xor ( n6175 , n173200 , n173499 );
and ( n6176 , n6175 , n173504 );
and ( n6177 , n173200 , n173499 );
or ( n6178 , n6176 , n6177 );
buf ( n173648 , n6178 );
nor ( n6180 , n173643 , n173648 );
not ( n6181 , n6180 );
not ( n6182 , n6181 );
or ( n6183 , n6171 , n6182 );
buf ( n173653 , n173643 );
buf ( n6185 , n173653 );
buf ( n173655 , n6185 );
buf ( n173656 , n173655 );
buf ( n173657 , n173648 );
buf ( n6189 , n173657 );
buf ( n173659 , n6189 );
buf ( n173660 , n173659 );
nand ( n6192 , n173656 , n173660 );
buf ( n173662 , n6192 );
nand ( n6194 , n6183 , n173662 );
not ( n6195 , n6194 );
xor ( n6196 , n173508 , n173624 );
xor ( n6197 , n6196 , n173629 );
buf ( n173667 , n6197 );
buf ( n173668 , n173667 );
buf ( n173669 , n839 );
xor ( n6201 , n173253 , n5842 );
xor ( n6202 , n6201 , n173364 );
buf ( n173672 , n6202 );
buf ( n173673 , n168989 );
buf ( n173674 , n799 );
nand ( n6206 , n173673 , n173674 );
buf ( n173676 , n6206 );
buf ( n173677 , n173676 );
not ( n6209 , n173677 );
not ( n6210 , n831 );
not ( n6211 , n173316 );
or ( n6212 , n6210 , n6211 );
nand ( n6213 , n168469 , n830 );
not ( n6214 , n6213 );
and ( n6215 , n830 , n780 );
not ( n6216 , n830 );
and ( n6217 , n6216 , n168631 );
nor ( n6218 , n6215 , n6217 );
nand ( n6219 , n6214 , n6218 );
nand ( n6220 , n6212 , n6219 );
buf ( n173690 , n6220 );
not ( n6222 , n173690 );
buf ( n173692 , n6222 );
buf ( n173693 , n173692 );
not ( n6225 , n173693 );
or ( n6226 , n6209 , n6225 );
buf ( n173696 , n786 );
buf ( n173697 , n824 );
xor ( n6229 , n173696 , n173697 );
buf ( n173699 , n6229 );
buf ( n173700 , n173699 );
not ( n6232 , n173700 );
buf ( n173702 , n1806 );
not ( n6234 , n173702 );
or ( n6235 , n6232 , n6234 );
buf ( n173705 , n170565 );
buf ( n173706 , n5943 );
nand ( n6238 , n173705 , n173706 );
buf ( n173708 , n6238 );
buf ( n173709 , n173708 );
nand ( n6241 , n6235 , n173709 );
buf ( n173711 , n6241 );
buf ( n173712 , n173711 );
nand ( n6244 , n6226 , n173712 );
buf ( n173714 , n6244 );
buf ( n173715 , n173714 );
buf ( n173716 , n173676 );
not ( n6248 , n173716 );
buf ( n173718 , n6220 );
nand ( n6250 , n6248 , n173718 );
buf ( n173720 , n6250 );
buf ( n173721 , n173720 );
nand ( n6253 , n173715 , n173721 );
buf ( n173723 , n6253 );
buf ( n173724 , n173723 );
xor ( n6256 , n173329 , n173346 );
xor ( n6257 , n6256 , n173360 );
buf ( n173727 , n6257 );
buf ( n173728 , n173727 );
xor ( n6260 , n173724 , n173728 );
buf ( n173730 , n788 );
buf ( n173731 , n822 );
xor ( n6263 , n173730 , n173731 );
buf ( n173733 , n6263 );
buf ( n173734 , n173733 );
not ( n6266 , n173734 );
buf ( n173736 , n1939 );
not ( n6268 , n173736 );
or ( n6269 , n6266 , n6268 );
buf ( n173739 , n169417 );
buf ( n173740 , n5785 );
nand ( n6272 , n173739 , n173740 );
buf ( n173742 , n6272 );
buf ( n173743 , n173742 );
nand ( n6275 , n6269 , n173743 );
buf ( n173745 , n6275 );
buf ( n173746 , n173745 );
buf ( n173747 , n798 );
buf ( n173748 , n812 );
xor ( n6280 , n173747 , n173748 );
buf ( n173750 , n6280 );
buf ( n173751 , n173750 );
not ( n6283 , n173751 );
buf ( n173753 , n2757 );
not ( n6285 , n173753 );
or ( n6286 , n6283 , n6285 );
buf ( n6287 , n1534 );
buf ( n173757 , n6287 );
buf ( n173758 , n5798 );
nand ( n6290 , n173757 , n173758 );
buf ( n173760 , n6290 );
buf ( n173761 , n173760 );
nand ( n6293 , n6286 , n173761 );
buf ( n173763 , n6293 );
buf ( n173764 , n173763 );
xor ( n6296 , n173746 , n173764 );
buf ( n173766 , n173333 );
not ( n6298 , n173766 );
buf ( n173768 , n169081 );
not ( n6300 , n173768 );
or ( n6301 , n6298 , n6300 );
buf ( n173771 , n4337 );
not ( n6303 , n173771 );
buf ( n173773 , n6303 );
buf ( n173774 , n173773 );
xor ( n6306 , n826 , n784 );
buf ( n173776 , n6306 );
not ( n6308 , n173776 );
buf ( n173778 , n6308 );
buf ( n173779 , n173778 );
or ( n6311 , n173774 , n173779 );
nand ( n6312 , n6301 , n6311 );
buf ( n173782 , n6312 );
buf ( n173783 , n173782 );
and ( n6315 , n6296 , n173783 );
and ( n6316 , n173746 , n173764 );
or ( n6317 , n6315 , n6316 );
buf ( n173787 , n6317 );
buf ( n173788 , n173787 );
and ( n6320 , n6260 , n173788 );
and ( n6321 , n173724 , n173728 );
or ( n6322 , n6320 , n6321 );
buf ( n173792 , n6322 );
buf ( n173793 , n173792 );
xor ( n6325 , n173672 , n173793 );
xor ( n6326 , n5975 , n173424 );
xor ( n6327 , n6326 , n173410 );
not ( n6328 , n6327 );
not ( n6329 , n6328 );
buf ( n6330 , n173266 );
xor ( n6331 , n173279 , n6330 );
xnor ( n6332 , n6331 , n173307 );
not ( n6333 , n6332 );
not ( n6334 , n6333 );
or ( n6335 , n6329 , n6334 );
not ( n6336 , n6332 );
not ( n6337 , n6327 );
or ( n6338 , n6336 , n6337 );
xor ( n6339 , n820 , n790 );
buf ( n173809 , n6339 );
not ( n6341 , n173809 );
buf ( n173811 , n2251 );
not ( n6343 , n173811 );
or ( n6344 , n6341 , n6343 );
buf ( n173814 , n168656 );
buf ( n173815 , n173354 );
nand ( n6347 , n173814 , n173815 );
buf ( n173817 , n6347 );
buf ( n173818 , n173817 );
nand ( n6350 , n6344 , n173818 );
buf ( n173820 , n6350 );
not ( n6352 , n173820 );
buf ( n173822 , n792 );
buf ( n173823 , n818 );
xor ( n6355 , n173822 , n173823 );
buf ( n173825 , n6355 );
buf ( n173826 , n173825 );
not ( n6358 , n173826 );
buf ( n173828 , n1321 );
not ( n6360 , n173828 );
or ( n6361 , n6358 , n6360 );
buf ( n173831 , n168806 );
buf ( n173832 , n173523 );
nand ( n6364 , n173831 , n173832 );
buf ( n173834 , n6364 );
buf ( n173835 , n173834 );
nand ( n6367 , n6361 , n173835 );
buf ( n173837 , n6367 );
not ( n6369 , n173837 );
or ( n6370 , n6352 , n6369 );
or ( n6371 , n173837 , n173820 );
buf ( n173841 , n799 );
buf ( n173842 , n813 );
or ( n6374 , n173841 , n173842 );
buf ( n173844 , n814 );
nand ( n6376 , n6374 , n173844 );
buf ( n173846 , n6376 );
buf ( n173847 , n799 );
buf ( n173848 , n813 );
nand ( n6380 , n173847 , n173848 );
buf ( n173850 , n6380 );
and ( n6382 , n173846 , n173850 , n812 );
not ( n6383 , n1471 );
buf ( n173853 , n781 );
buf ( n173854 , n830 );
xor ( n6386 , n173853 , n173854 );
buf ( n173856 , n6386 );
not ( n6388 , n173856 );
or ( n6389 , n6383 , n6388 );
buf ( n173859 , n6218 );
buf ( n173860 , n831 );
nand ( n6392 , n173859 , n173860 );
buf ( n173862 , n6392 );
nand ( n6394 , n6389 , n173862 );
and ( n6395 , n6382 , n6394 );
nand ( n6396 , n6371 , n6395 );
nand ( n6397 , n6370 , n6396 );
nand ( n6398 , n6338 , n6397 );
nand ( n6399 , n6335 , n6398 );
buf ( n173869 , n6399 );
and ( n6401 , n6325 , n173869 );
and ( n6402 , n173672 , n173793 );
or ( n6403 , n6401 , n6402 );
buf ( n173873 , n6403 );
buf ( n173874 , n173873 );
and ( n6406 , n5999 , n5984 );
not ( n6407 , n5999 );
and ( n6408 , n6407 , n5981 );
nor ( n6409 , n6406 , n6408 );
buf ( n173879 , n6409 );
buf ( n173880 , n5927 );
and ( n6412 , n173879 , n173880 );
not ( n6413 , n173879 );
buf ( n6414 , n5991 );
buf ( n173884 , n6414 );
and ( n6416 , n6413 , n173884 );
nor ( n6417 , n6412 , n6416 );
buf ( n173887 , n6417 );
buf ( n173888 , n173887 );
xor ( n6420 , n173514 , n173518 );
xor ( n6421 , n6420 , n173595 );
buf ( n173891 , n6421 );
buf ( n173892 , n173891 );
xor ( n6424 , n173888 , n173892 );
xor ( n6425 , n173536 , n173539 );
xor ( n6426 , n6425 , n173590 );
buf ( n173896 , n6426 );
buf ( n173897 , n173896 );
buf ( n173898 , n787 );
buf ( n173899 , n824 );
xor ( n6431 , n173898 , n173899 );
buf ( n173901 , n6431 );
not ( n6433 , n173901 );
not ( n6434 , n1679 );
or ( n6435 , n6433 , n6434 );
not ( n6436 , n170562 );
nand ( n6437 , n6436 , n173699 );
nand ( n6438 , n6435 , n6437 );
buf ( n173908 , n6438 );
not ( n6440 , n173908 );
xor ( n6441 , n814 , n797 );
buf ( n173911 , n6441 );
not ( n6443 , n173911 );
buf ( n173913 , n169241 );
not ( n6445 , n173913 );
or ( n6446 , n6443 , n6445 );
buf ( n173916 , n169247 );
buf ( n173917 , n173554 );
nand ( n6449 , n173916 , n173917 );
buf ( n173919 , n6449 );
buf ( n173920 , n173919 );
nand ( n6452 , n6446 , n173920 );
buf ( n173922 , n6452 );
buf ( n173923 , n173922 );
not ( n6455 , n173923 );
or ( n6456 , n6440 , n6455 );
buf ( n173926 , n6438 );
buf ( n173927 , n173922 );
or ( n6459 , n173926 , n173927 );
xor ( n6460 , n795 , n816 );
not ( n6461 , n6460 );
not ( n6462 , n5964 );
or ( n6463 , n6461 , n6462 );
nand ( n6464 , n169842 , n6072 );
nand ( n6465 , n6463 , n6464 );
buf ( n173935 , n6465 );
nand ( n6467 , n6459 , n173935 );
buf ( n173937 , n6467 );
buf ( n173938 , n173937 );
nand ( n6470 , n6456 , n173938 );
buf ( n173940 , n6470 );
buf ( n173941 , n173940 );
buf ( n173942 , n789 );
buf ( n173943 , n822 );
xor ( n6475 , n173942 , n173943 );
buf ( n173945 , n6475 );
buf ( n173946 , n173945 );
not ( n6478 , n173946 );
buf ( n173948 , n1939 );
not ( n6480 , n173948 );
or ( n6481 , n6478 , n6480 );
buf ( n173951 , n169417 );
buf ( n173952 , n173733 );
nand ( n6484 , n173951 , n173952 );
buf ( n173954 , n6484 );
buf ( n173955 , n173954 );
nand ( n6487 , n6481 , n173955 );
buf ( n173957 , n6487 );
not ( n6489 , n173957 );
buf ( n173959 , n783 );
buf ( n173960 , n828 );
xor ( n6492 , n173959 , n173960 );
buf ( n173962 , n6492 );
buf ( n173963 , n173962 );
not ( n6495 , n173963 );
buf ( n173965 , n168549 );
not ( n6497 , n173965 );
or ( n6498 , n6495 , n6497 );
buf ( n173968 , n168559 );
buf ( n173969 , n173572 );
nand ( n6501 , n173968 , n173969 );
buf ( n173971 , n6501 );
buf ( n173972 , n173971 );
nand ( n6504 , n6498 , n173972 );
buf ( n173974 , n6504 );
not ( n6506 , n173974 );
or ( n6507 , n6489 , n6506 );
buf ( n173977 , n173974 );
buf ( n173978 , n173957 );
nor ( n6510 , n173977 , n173978 );
buf ( n173980 , n6510 );
buf ( n173981 , n799 );
buf ( n173982 , n812 );
xor ( n6514 , n173981 , n173982 );
buf ( n173984 , n6514 );
buf ( n173985 , n173984 );
not ( n6517 , n173985 );
buf ( n173987 , n2757 );
not ( n6519 , n173987 );
or ( n6520 , n6517 , n6519 );
buf ( n173990 , n1534 );
buf ( n173991 , n173750 );
nand ( n6523 , n173990 , n173991 );
buf ( n173993 , n6523 );
buf ( n173994 , n173993 );
nand ( n6526 , n6520 , n173994 );
buf ( n173996 , n6526 );
buf ( n173997 , n173996 );
not ( n6529 , n173997 );
buf ( n173999 , n6529 );
or ( n6531 , n173980 , n173999 );
nand ( n6532 , n6507 , n6531 );
buf ( n174002 , n6532 );
xor ( n6534 , n173941 , n174002 );
xor ( n6535 , n820 , n791 );
not ( n6536 , n6535 );
not ( n6537 , n2251 );
or ( n6538 , n6536 , n6537 );
buf ( n174008 , n2513 );
buf ( n174009 , n6339 );
nand ( n6541 , n174008 , n174009 );
buf ( n174011 , n6541 );
nand ( n6543 , n6538 , n174011 );
not ( n6544 , n6543 );
xor ( n6545 , n818 , n793 );
not ( n6546 , n6545 );
not ( n6547 , n1321 );
or ( n6548 , n6546 , n6547 );
buf ( n174018 , n168806 );
buf ( n174019 , n173825 );
nand ( n6551 , n174018 , n174019 );
buf ( n174021 , n6551 );
nand ( n6553 , n6548 , n174021 );
not ( n6554 , n6553 );
or ( n6555 , n6544 , n6554 );
nor ( n6556 , n6543 , n6553 );
xor ( n6557 , n826 , n785 );
not ( n6558 , n6557 );
not ( n6559 , n169674 );
or ( n6560 , n6558 , n6559 );
buf ( n174030 , n169081 );
buf ( n174031 , n6306 );
nand ( n6563 , n174030 , n174031 );
buf ( n174033 , n6563 );
nand ( n6565 , n6560 , n174033 );
not ( n6566 , n6565 );
or ( n6567 , n6556 , n6566 );
nand ( n6568 , n6555 , n6567 );
buf ( n174038 , n6568 );
and ( n6570 , n6534 , n174038 );
and ( n6571 , n173941 , n174002 );
or ( n6572 , n6570 , n6571 );
buf ( n174042 , n6572 );
buf ( n174043 , n174042 );
xor ( n6575 , n173897 , n174043 );
xor ( n6576 , n173724 , n173728 );
xor ( n6577 , n6576 , n173788 );
buf ( n174047 , n6577 );
buf ( n174048 , n174047 );
and ( n6580 , n6575 , n174048 );
and ( n6581 , n173897 , n174043 );
or ( n6582 , n6580 , n6581 );
buf ( n174052 , n6582 );
buf ( n174053 , n174052 );
and ( n6585 , n6424 , n174053 );
and ( n6586 , n173888 , n173892 );
or ( n6587 , n6585 , n6586 );
buf ( n174057 , n6587 );
buf ( n174058 , n174057 );
xor ( n6590 , n173874 , n174058 );
xor ( n6591 , n173600 , n173604 );
xor ( n6592 , n6591 , n173609 );
buf ( n174062 , n6592 );
buf ( n174063 , n174062 );
and ( n6595 , n6590 , n174063 );
and ( n6596 , n173874 , n174058 );
or ( n6597 , n6595 , n6596 );
buf ( n174067 , n6597 );
buf ( n174068 , n174067 );
xor ( n6600 , n173669 , n174068 );
xor ( n6601 , n173511 , n173614 );
xor ( n6602 , n6601 , n173619 );
buf ( n174072 , n6602 );
buf ( n174073 , n174072 );
and ( n6605 , n6600 , n174073 );
and ( n6606 , n173669 , n174068 );
or ( n6607 , n6605 , n6606 );
buf ( n174077 , n6607 );
buf ( n174078 , n174077 );
nor ( n6610 , n173668 , n174078 );
buf ( n174080 , n6610 );
buf ( n174081 , n174080 );
xor ( n6613 , n173669 , n174068 );
xor ( n6614 , n6613 , n174073 );
buf ( n174084 , n6614 );
buf ( n174085 , n174084 );
buf ( n174086 , n840 );
xor ( n6618 , n173672 , n173793 );
xor ( n6619 , n6618 , n173869 );
buf ( n174089 , n6619 );
buf ( n174090 , n174089 );
xor ( n6622 , n173888 , n173892 );
xor ( n6623 , n6622 , n174053 );
buf ( n174093 , n6623 );
buf ( n174094 , n174093 );
xor ( n6626 , n174090 , n174094 );
buf ( n174096 , n173711 );
not ( n6628 , n174096 );
buf ( n174098 , n6220 );
not ( n6630 , n174098 );
buf ( n174100 , n173676 );
not ( n6632 , n174100 );
and ( n6633 , n6630 , n6632 );
buf ( n174103 , n6220 );
buf ( n174104 , n173676 );
and ( n6636 , n174103 , n174104 );
nor ( n6637 , n6633 , n6636 );
buf ( n174107 , n6637 );
buf ( n174108 , n174107 );
not ( n6640 , n174108 );
or ( n6641 , n6628 , n6640 );
buf ( n174111 , n174107 );
buf ( n174112 , n173711 );
or ( n6644 , n174111 , n174112 );
nand ( n6645 , n6641 , n6644 );
buf ( n174115 , n6645 );
buf ( n174116 , n174115 );
xor ( n6648 , n173550 , n173567 );
xor ( n6649 , n6648 , n173585 );
buf ( n174119 , n6649 );
buf ( n174120 , n174119 );
xor ( n6652 , n174116 , n174120 );
xor ( n6653 , n173746 , n173764 );
xor ( n6654 , n6653 , n173783 );
buf ( n174124 , n6654 );
buf ( n174125 , n174124 );
and ( n6657 , n6652 , n174125 );
and ( n6658 , n174116 , n174120 );
or ( n6659 , n6657 , n6658 );
buf ( n174129 , n6659 );
buf ( n174130 , n174129 );
nand ( n6662 , n6328 , n6397 , n6333 );
not ( n6663 , n6397 );
nand ( n6664 , n6327 , n6663 , n6333 );
nand ( n6665 , n6328 , n6663 , n6332 );
nand ( n6666 , n6332 , n6397 , n6327 );
nand ( n6667 , n6662 , n6664 , n6665 , n6666 );
buf ( n174137 , n6667 );
xor ( n6669 , n174130 , n174137 );
xor ( n6670 , n173897 , n174043 );
xor ( n6671 , n6670 , n174048 );
buf ( n174141 , n6671 );
buf ( n174142 , n174141 );
and ( n6674 , n6669 , n174142 );
and ( n6675 , n174130 , n174137 );
or ( n6676 , n6674 , n6675 );
buf ( n174146 , n6676 );
buf ( n174147 , n174146 );
and ( n6679 , n6626 , n174147 );
and ( n6680 , n174090 , n174094 );
or ( n6681 , n6679 , n6680 );
buf ( n174151 , n6681 );
buf ( n174152 , n174151 );
xor ( n6684 , n174086 , n174152 );
xor ( n6685 , n173874 , n174058 );
xor ( n6686 , n6685 , n174063 );
buf ( n174156 , n6686 );
buf ( n174157 , n174156 );
and ( n6689 , n6684 , n174157 );
and ( n6690 , n174086 , n174152 );
or ( n6691 , n6689 , n6690 );
buf ( n174161 , n6691 );
buf ( n174162 , n174161 );
nor ( n6694 , n174085 , n174162 );
buf ( n174164 , n6694 );
buf ( n174165 , n174164 );
nor ( n6697 , n174081 , n174165 );
buf ( n174167 , n6697 );
buf ( n174168 , n174167 );
buf ( n6700 , n174168 );
buf ( n174170 , n6700 );
buf ( n174171 , n174170 );
not ( n6703 , n174171 );
buf ( n174173 , n6703 );
buf ( n174174 , n174084 );
buf ( n174175 , n174161 );
nand ( n6707 , n174174 , n174175 );
buf ( n174177 , n6707 );
buf ( n174178 , n174177 );
not ( n6710 , n174178 );
buf ( n174180 , n6710 );
not ( n6712 , n174180 );
buf ( n174182 , n174080 );
not ( n6714 , n174182 );
buf ( n174184 , n6714 );
not ( n6716 , n174184 );
or ( n6717 , n6712 , n6716 );
buf ( n174187 , n173667 );
buf ( n6719 , n174187 );
buf ( n174189 , n6719 );
buf ( n174190 , n174189 );
buf ( n174191 , n174077 );
nand ( n6723 , n174190 , n174191 );
buf ( n174193 , n6723 );
nand ( n6725 , n6717 , n174193 );
not ( n6726 , n6725 );
nand ( n6727 , n6195 , n174173 , n6726 );
buf ( n174197 , n6727 );
xor ( n6729 , n174086 , n174152 );
xor ( n6730 , n6729 , n174157 );
buf ( n174200 , n6730 );
buf ( n174201 , n174200 );
buf ( n174202 , n841 );
xor ( n6734 , n173837 , n173820 );
xor ( n6735 , n6734 , n6395 );
buf ( n174205 , n788 );
buf ( n174206 , n824 );
xor ( n6738 , n174205 , n174206 );
buf ( n174208 , n6738 );
not ( n6740 , n174208 );
not ( n6741 , n170100 );
or ( n6742 , n6740 , n6741 );
buf ( n174212 , n170565 );
buf ( n174213 , n173901 );
nand ( n6745 , n174212 , n174213 );
buf ( n174215 , n6745 );
nand ( n6747 , n6742 , n174215 );
not ( n6748 , n6747 );
buf ( n174218 , n1534 );
buf ( n174219 , n799 );
and ( n6751 , n174218 , n174219 );
buf ( n174221 , n6751 );
not ( n6753 , n174221 );
buf ( n174223 , n782 );
buf ( n174224 , n830 );
xor ( n6756 , n174223 , n174224 );
buf ( n174226 , n6756 );
buf ( n174227 , n174226 );
not ( n6759 , n174227 );
buf ( n174229 , n168471 );
not ( n6761 , n174229 );
or ( n6762 , n6759 , n6761 );
buf ( n174232 , n173856 );
buf ( n174233 , n831 );
nand ( n6765 , n174232 , n174233 );
buf ( n174235 , n6765 );
buf ( n174236 , n174235 );
nand ( n6768 , n6762 , n174236 );
buf ( n174238 , n6768 );
not ( n6770 , n174238 );
nand ( n6771 , n6753 , n6770 );
not ( n6772 , n6771 );
or ( n6773 , n6748 , n6772 );
nand ( n6774 , n174238 , n174221 );
nand ( n6775 , n6773 , n6774 );
not ( n6776 , n6775 );
xor ( n6777 , n6382 , n6394 );
not ( n6778 , n6777 );
nand ( n6779 , n6776 , n6778 );
not ( n6780 , n6779 );
buf ( n174250 , n796 );
buf ( n174251 , n816 );
xor ( n6783 , n174250 , n174251 );
buf ( n174253 , n6783 );
buf ( n174254 , n174253 );
not ( n6786 , n174254 );
buf ( n174256 , n169836 );
not ( n6788 , n174256 );
or ( n6789 , n6786 , n6788 );
nand ( n6790 , n6460 , n169320 );
buf ( n174260 , n6790 );
nand ( n6792 , n6789 , n174260 );
buf ( n174262 , n6792 );
buf ( n174263 , n174262 );
not ( n6795 , n174263 );
buf ( n174265 , n6795 );
buf ( n174266 , n174265 );
not ( n6798 , n174266 );
buf ( n174268 , n798 );
buf ( n174269 , n814 );
xor ( n6801 , n174268 , n174269 );
buf ( n174271 , n6801 );
buf ( n174272 , n174271 );
not ( n174273 , n174272 );
buf ( n174274 , n171013 );
not ( n174275 , n174274 );
or ( n6807 , n174273 , n174275 );
buf ( n174277 , n169250 );
buf ( n174278 , n6441 );
nand ( n174279 , n174277 , n174278 );
buf ( n174280 , n174279 );
buf ( n174281 , n174280 );
nand ( n6813 , n6807 , n174281 );
buf ( n174283 , n6813 );
buf ( n174284 , n174283 );
not ( n174285 , n174284 );
buf ( n174286 , n174285 );
buf ( n174287 , n174286 );
not ( n6819 , n174287 );
or ( n174289 , n6798 , n6819 );
buf ( n174290 , n784 );
buf ( n174291 , n828 );
xor ( n6823 , n174290 , n174291 );
buf ( n174293 , n6823 );
buf ( n174294 , n174293 );
not ( n174295 , n174294 );
buf ( n174296 , n170990 );
not ( n174297 , n174296 );
or ( n6829 , n174295 , n174297 );
buf ( n174299 , n168559 );
buf ( n174300 , n173962 );
nand ( n174301 , n174299 , n174300 );
buf ( n174302 , n174301 );
buf ( n174303 , n174302 );
nand ( n6835 , n6829 , n174303 );
buf ( n174305 , n6835 );
buf ( n174306 , n174305 );
nand ( n174307 , n174289 , n174306 );
buf ( n174308 , n174307 );
buf ( n174309 , n174271 );
not ( n6841 , n174309 );
buf ( n174311 , n171013 );
not ( n6843 , n174311 );
or ( n174313 , n6841 , n6843 );
buf ( n174314 , n174280 );
nand ( n174315 , n174313 , n174314 );
buf ( n174316 , n174315 );
buf ( n174317 , n174316 );
buf ( n174318 , n174262 );
nand ( n174319 , n174317 , n174318 );
buf ( n174320 , n174319 );
nand ( n174321 , n174308 , n174320 );
not ( n6853 , n174321 );
or ( n174323 , n6780 , n6853 );
nand ( n6855 , n6777 , n6775 );
nand ( n174325 , n174323 , n6855 );
xor ( n6857 , n6735 , n174325 );
buf ( n174327 , n6438 );
not ( n6859 , n174327 );
buf ( n174329 , n6465 );
not ( n6861 , n174329 );
buf ( n174331 , n6861 );
buf ( n174332 , n174331 );
not ( n174333 , n174332 );
or ( n6865 , n6859 , n174333 );
buf ( n174335 , n174331 );
buf ( n174336 , n6438 );
or ( n174337 , n174335 , n174336 );
nand ( n6869 , n6865 , n174337 );
buf ( n174339 , n6869 );
buf ( n174340 , n174339 );
buf ( n174341 , n173922 );
and ( n6873 , n174340 , n174341 );
not ( n174343 , n174340 );
buf ( n174344 , n173922 );
not ( n174345 , n174344 );
buf ( n174346 , n174345 );
buf ( n174347 , n174346 );
and ( n6879 , n174343 , n174347 );
nor ( n174349 , n6873 , n6879 );
buf ( n174350 , n174349 );
buf ( n174351 , n174350 );
buf ( n174352 , n790 );
buf ( n174353 , n822 );
xor ( n6885 , n174352 , n174353 );
buf ( n174355 , n6885 );
buf ( n174356 , n174355 );
not ( n174357 , n174356 );
buf ( n174358 , n1939 );
not ( n174359 , n174358 );
or ( n6891 , n174357 , n174359 );
buf ( n174361 , n169417 );
buf ( n174362 , n173945 );
nand ( n174363 , n174361 , n174362 );
buf ( n174364 , n174363 );
buf ( n174365 , n174364 );
nand ( n6897 , n6891 , n174365 );
buf ( n174367 , n6897 );
buf ( n174368 , n174367 );
xor ( n174369 , n820 , n792 );
not ( n6901 , n174369 );
not ( n174371 , n2251 );
or ( n6903 , n6901 , n174371 );
nand ( n174373 , n6535 , n168655 );
nand ( n6905 , n6903 , n174373 );
buf ( n174375 , n6905 );
xor ( n6907 , n174368 , n174375 );
buf ( n174377 , n6557 );
not ( n6909 , n174377 );
buf ( n174379 , n169081 );
not ( n6911 , n174379 );
or ( n174381 , n6909 , n6911 );
buf ( n174382 , n169093 );
buf ( n174383 , n786 );
buf ( n174384 , n826 );
xor ( n174385 , n174383 , n174384 );
buf ( n174386 , n174385 );
buf ( n174387 , n174386 );
not ( n6919 , n174387 );
buf ( n174389 , n6919 );
buf ( n174390 , n174389 );
or ( n174391 , n174382 , n174390 );
nand ( n6923 , n174381 , n174391 );
buf ( n174393 , n6923 );
buf ( n174394 , n174393 );
and ( n174395 , n6907 , n174394 );
and ( n6927 , n174368 , n174375 );
or ( n174397 , n174395 , n6927 );
buf ( n174398 , n174397 );
buf ( n174399 , n174398 );
xor ( n174400 , n174351 , n174399 );
xor ( n6932 , n6565 , n6553 );
xor ( n174402 , n6932 , n6543 );
buf ( n174403 , n174402 );
and ( n6935 , n174400 , n174403 );
and ( n174405 , n174351 , n174399 );
or ( n6937 , n6935 , n174405 );
buf ( n174407 , n6937 );
and ( n174408 , n6857 , n174407 );
and ( n174409 , n6735 , n174325 );
or ( n6941 , n174408 , n174409 );
buf ( n174411 , n6941 );
xor ( n6943 , n173941 , n174002 );
xor ( n6944 , n6943 , n174038 );
buf ( n174414 , n6944 );
not ( n6946 , n174414 );
xor ( n6947 , n174116 , n174120 );
xor ( n174417 , n6947 , n174125 );
buf ( n174418 , n174417 );
not ( n174419 , n174418 );
nand ( n6954 , n6946 , n174419 );
not ( n6955 , n6954 );
xor ( n6956 , n6735 , n174325 );
xor ( n6957 , n6956 , n174407 );
not ( n6958 , n6957 );
or ( n174425 , n6955 , n6958 );
not ( n6960 , n174419 );
nand ( n6961 , n6960 , n174414 );
nand ( n6962 , n174425 , n6961 );
buf ( n174429 , n6962 );
xor ( n6964 , n174411 , n174429 );
xor ( n6965 , n174130 , n174137 );
xor ( n174432 , n6965 , n174142 );
buf ( n174433 , n174432 );
buf ( n174434 , n174433 );
and ( n6969 , n6964 , n174434 );
and ( n6970 , n174411 , n174429 );
or ( n6971 , n6969 , n6970 );
buf ( n174438 , n6971 );
buf ( n174439 , n174438 );
xor ( n6974 , n174202 , n174439 );
xor ( n6975 , n174090 , n174094 );
xor ( n6976 , n6975 , n174147 );
buf ( n174443 , n6976 );
buf ( n174444 , n174443 );
and ( n174445 , n6974 , n174444 );
and ( n6980 , n174202 , n174439 );
or ( n6981 , n174445 , n6980 );
buf ( n174448 , n6981 );
buf ( n174449 , n174448 );
nor ( n6984 , n174201 , n174449 );
buf ( n174451 , n6984 );
xor ( n174452 , n174202 , n174439 );
xor ( n6987 , n174452 , n174444 );
buf ( n174454 , n6987 );
buf ( n174455 , n174454 );
buf ( n174456 , n842 );
xor ( n6991 , n173996 , n173974 );
xor ( n174458 , n6991 , n173957 );
buf ( n174459 , n174458 );
xor ( n6997 , n6778 , n6775 );
xnor ( n174461 , n6997 , n174321 );
buf ( n174462 , n174461 );
xor ( n7000 , n174459 , n174462 );
buf ( n174464 , n6545 );
not ( n7002 , n174464 );
buf ( n174466 , n168806 );
not ( n7004 , n174466 );
or ( n7005 , n7002 , n7004 );
buf ( n174469 , n1321 );
buf ( n174470 , n794 );
buf ( n174471 , n818 );
xor ( n7009 , n174470 , n174471 );
buf ( n174473 , n7009 );
buf ( n174474 , n174473 );
nand ( n7012 , n174469 , n174474 );
buf ( n174476 , n7012 );
buf ( n174477 , n174476 );
nand ( n7015 , n7005 , n174477 );
buf ( n174479 , n7015 );
not ( n174480 , n174479 );
buf ( n174481 , n783 );
buf ( n174482 , n830 );
xor ( n7020 , n174481 , n174482 );
buf ( n174484 , n7020 );
buf ( n174485 , n174484 );
not ( n7023 , n174485 );
buf ( n174487 , n1471 );
not ( n7025 , n174487 );
or ( n7026 , n7023 , n7025 );
buf ( n174490 , n174226 );
buf ( n174491 , n831 );
nand ( n174492 , n174490 , n174491 );
buf ( n174493 , n174492 );
buf ( n174494 , n174493 );
nand ( n7032 , n7026 , n174494 );
buf ( n174496 , n7032 );
buf ( n174497 , n799 );
buf ( n174498 , n815 );
or ( n7036 , n174497 , n174498 );
buf ( n174500 , n816 );
nand ( n174501 , n7036 , n174500 );
buf ( n174502 , n174501 );
buf ( n174503 , n174502 );
buf ( n174504 , n799 );
buf ( n174505 , n815 );
nand ( n7046 , n174504 , n174505 );
buf ( n174507 , n7046 );
buf ( n174508 , n174507 );
buf ( n174509 , n814 );
nand ( n7050 , n174503 , n174508 , n174509 );
buf ( n174511 , n7050 );
not ( n7052 , n174511 );
and ( n7053 , n174496 , n7052 );
not ( n174514 , n7053 );
nand ( n7055 , n174480 , n174514 );
buf ( n174516 , n7055 );
not ( n7057 , n174516 );
buf ( n174518 , n170565 );
buf ( n174519 , n174208 );
nand ( n7060 , n174518 , n174519 );
buf ( n174521 , n7060 );
buf ( n174522 , n789 );
buf ( n174523 , n824 );
xor ( n7064 , n174522 , n174523 );
buf ( n174525 , n7064 );
nand ( n7066 , n170100 , n174525 );
and ( n7067 , n174521 , n7066 );
not ( n174528 , n7067 );
buf ( n174529 , n799 );
buf ( n174530 , n814 );
xor ( n7071 , n174529 , n174530 );
buf ( n174532 , n7071 );
not ( n7073 , n174532 );
not ( n7074 , n169922 );
or ( n7075 , n7073 , n7074 );
buf ( n174536 , n169250 );
buf ( n174537 , n174271 );
nand ( n7078 , n174536 , n174537 );
buf ( n174539 , n7078 );
nand ( n7080 , n7075 , n174539 );
or ( n7081 , n174528 , n7080 );
buf ( n174542 , n797 );
buf ( n174543 , n816 );
xor ( n7084 , n174542 , n174543 );
buf ( n174545 , n7084 );
not ( n7086 , n174545 );
not ( n7087 , n169836 );
or ( n7088 , n7086 , n7087 );
buf ( n174549 , n169320 );
buf ( n174550 , n174253 );
nand ( n7091 , n174549 , n174550 );
buf ( n174552 , n7091 );
nand ( n7093 , n7088 , n174552 );
nand ( n7094 , n7081 , n7093 );
nand ( n7095 , n174528 , n7080 );
nand ( n7096 , n7094 , n7095 );
buf ( n174557 , n7096 );
not ( n7098 , n174557 );
or ( n7099 , n7057 , n7098 );
nand ( n7100 , n174479 , n7053 );
buf ( n174561 , n7100 );
nand ( n7102 , n7099 , n174561 );
buf ( n174563 , n7102 );
buf ( n174564 , n174563 );
and ( n7105 , n7000 , n174564 );
and ( n7106 , n174459 , n174462 );
or ( n7107 , n7105 , n7106 );
buf ( n174568 , n7107 );
xor ( n7109 , n174351 , n174399 );
xor ( n7110 , n7109 , n174403 );
buf ( n174571 , n7110 );
xor ( n174572 , n174221 , n6770 );
xnor ( n7116 , n174572 , n6747 );
buf ( n174574 , n791 );
buf ( n174575 , n822 );
xor ( n7119 , n174574 , n174575 );
buf ( n174577 , n7119 );
buf ( n174578 , n174577 );
not ( n7122 , n174578 );
buf ( n174580 , n169411 );
not ( n174581 , n174580 );
or ( n7125 , n7122 , n174581 );
buf ( n174583 , n169417 );
buf ( n174584 , n174355 );
nand ( n7128 , n174583 , n174584 );
buf ( n174586 , n7128 );
buf ( n174587 , n174586 );
nand ( n7131 , n7125 , n174587 );
buf ( n174589 , n7131 );
not ( n7133 , n174589 );
not ( n174591 , n168663 );
not ( n7135 , n168661 );
or ( n7136 , n174591 , n7135 );
nand ( n7137 , n7136 , n168665 );
buf ( n174595 , n7137 );
not ( n7139 , n174595 );
buf ( n174597 , n787 );
buf ( n174598 , n826 );
xnor ( n7142 , n174597 , n174598 );
buf ( n174600 , n7142 );
buf ( n174601 , n174600 );
not ( n7145 , n174601 );
and ( n7146 , n7139 , n7145 );
buf ( n174604 , n169081 );
buf ( n174605 , n174386 );
and ( n7149 , n174604 , n174605 );
nor ( n7150 , n7146 , n7149 );
buf ( n174608 , n7150 );
not ( n174609 , n174608 );
not ( n7153 , n174609 );
or ( n7154 , n7133 , n7153 );
not ( n174612 , n174608 );
buf ( n174613 , n174577 );
not ( n7157 , n174613 );
buf ( n174615 , n169411 );
not ( n7159 , n174615 );
or ( n7160 , n7157 , n7159 );
buf ( n174618 , n174586 );
nand ( n7162 , n7160 , n174618 );
buf ( n174620 , n7162 );
buf ( n174621 , n174620 );
not ( n174622 , n174621 );
buf ( n174623 , n174622 );
not ( n7167 , n174623 );
or ( n7168 , n174612 , n7167 );
buf ( n174626 , n785 );
buf ( n174627 , n828 );
xor ( n7171 , n174626 , n174627 );
buf ( n174629 , n7171 );
buf ( n174630 , n174629 );
not ( n7174 , n174630 );
buf ( n174632 , n170990 );
not ( n7176 , n174632 );
or ( n7177 , n7174 , n7176 );
buf ( n174635 , n168559 );
buf ( n174636 , n174293 );
nand ( n7183 , n174635 , n174636 );
buf ( n174638 , n7183 );
buf ( n174639 , n174638 );
nand ( n7186 , n7177 , n174639 );
buf ( n174641 , n7186 );
nand ( n7188 , n7168 , n174641 );
nand ( n7189 , n7154 , n7188 );
xor ( n7190 , n7116 , n7189 );
xor ( n174645 , n174368 , n174375 );
xor ( n7192 , n174645 , n174394 );
buf ( n174647 , n7192 );
and ( n7194 , n7190 , n174647 );
and ( n174649 , n7116 , n7189 );
or ( n7196 , n7194 , n174649 );
xor ( n7197 , n174571 , n7196 );
buf ( n174652 , n174286 );
not ( n7199 , n174652 );
buf ( n174654 , n174262 );
not ( n174655 , n174654 );
and ( n7202 , n7199 , n174655 );
buf ( n174657 , n174262 );
buf ( n174658 , n174286 );
and ( n7205 , n174657 , n174658 );
nor ( n7206 , n7202 , n7205 );
buf ( n174661 , n7206 );
buf ( n174662 , n174661 );
buf ( n174663 , n174305 );
not ( n7210 , n174663 );
buf ( n174665 , n7210 );
buf ( n174666 , n174665 );
and ( n7213 , n174662 , n174666 );
not ( n7214 , n174662 );
buf ( n174669 , n174305 );
and ( n7216 , n7214 , n174669 );
nor ( n7217 , n7213 , n7216 );
buf ( n174672 , n7217 );
not ( n7219 , n174672 );
xor ( n7220 , n820 , n793 );
buf ( n174675 , n7220 );
not ( n7222 , n174675 );
buf ( n174677 , n2251 );
not ( n7224 , n174677 );
or ( n7225 , n7222 , n7224 );
buf ( n174680 , n2513 );
buf ( n174681 , n174369 );
nand ( n7228 , n174680 , n174681 );
buf ( n174683 , n7228 );
buf ( n174684 , n174683 );
nand ( n7231 , n7225 , n174684 );
buf ( n174686 , n7231 );
buf ( n174687 , n174686 );
not ( n7234 , n174687 );
buf ( n174689 , n174511 );
not ( n174690 , n174689 );
buf ( n174691 , n174496 );
not ( n7238 , n174691 );
or ( n7239 , n174690 , n7238 );
buf ( n174694 , n174496 );
buf ( n174695 , n174511 );
or ( n7242 , n174694 , n174695 );
nand ( n7243 , n7239 , n7242 );
buf ( n174698 , n7243 );
buf ( n174699 , n174698 );
not ( n174700 , n174699 );
or ( n7247 , n7234 , n174700 );
buf ( n174702 , n174698 );
buf ( n174703 , n174686 );
or ( n7250 , n174702 , n174703 );
buf ( n174705 , n795 );
buf ( n174706 , n818 );
xor ( n7253 , n174705 , n174706 );
buf ( n174708 , n7253 );
buf ( n174709 , n174708 );
not ( n7256 , n174709 );
buf ( n174711 , n1321 );
not ( n7258 , n174711 );
or ( n7259 , n7256 , n7258 );
buf ( n174714 , n168806 );
buf ( n174715 , n174473 );
nand ( n7262 , n174714 , n174715 );
buf ( n174717 , n7262 );
buf ( n174718 , n174717 );
nand ( n7265 , n7259 , n174718 );
buf ( n174720 , n7265 );
buf ( n174721 , n174720 );
nand ( n7268 , n7250 , n174721 );
buf ( n174723 , n7268 );
buf ( n174724 , n174723 );
nand ( n7271 , n7247 , n174724 );
buf ( n174726 , n7271 );
not ( n7276 , n174726 );
or ( n7277 , n7219 , n7276 );
buf ( n174729 , n174672 );
buf ( n174730 , n174726 );
nor ( n7280 , n174729 , n174730 );
buf ( n174732 , n7280 );
and ( n7282 , n174514 , n174479 );
not ( n7283 , n174514 );
and ( n7284 , n7283 , n174480 );
nor ( n7285 , n7282 , n7284 );
xor ( n7286 , n7096 , n7285 );
or ( n7287 , n174732 , n7286 );
nand ( n7288 , n7277 , n7287 );
and ( n7289 , n7197 , n7288 );
and ( n7290 , n174571 , n7196 );
or ( n174742 , n7289 , n7290 );
xor ( n7292 , n174568 , n174742 );
not ( n7293 , n174418 );
and ( n7294 , n174414 , n7293 );
not ( n7295 , n174414 );
and ( n7296 , n7295 , n174418 );
nor ( n7297 , n7294 , n7296 );
not ( n7298 , n6957 );
and ( n7299 , n7297 , n7298 );
not ( n7300 , n7297 );
and ( n174752 , n7300 , n6957 );
nor ( n7302 , n7299 , n174752 );
and ( n7303 , n7292 , n7302 );
and ( n7304 , n174568 , n174742 );
or ( n7305 , n7303 , n7304 );
buf ( n174757 , n7305 );
xor ( n7307 , n174456 , n174757 );
xor ( n7308 , n174411 , n174429 );
xor ( n7309 , n7308 , n174434 );
buf ( n174761 , n7309 );
buf ( n174762 , n174761 );
and ( n7312 , n7307 , n174762 );
and ( n7313 , n174456 , n174757 );
or ( n7314 , n7312 , n7313 );
buf ( n174766 , n7314 );
buf ( n174767 , n174766 );
nor ( n174768 , n174455 , n174767 );
buf ( n174769 , n174768 );
nor ( n7319 , n174451 , n174769 );
xor ( n7320 , n174456 , n174757 );
xor ( n7321 , n7320 , n174762 );
buf ( n174773 , n7321 );
buf ( n174774 , n174773 );
buf ( n174775 , n843 );
xor ( n7325 , n174459 , n174462 );
xor ( n7326 , n7325 , n174564 );
buf ( n174778 , n7326 );
buf ( n174779 , n169247 );
buf ( n174780 , n799 );
nand ( n7330 , n174779 , n174780 );
buf ( n174782 , n7330 );
buf ( n174783 , n174782 );
not ( n7333 , n174783 );
not ( n7334 , n831 );
not ( n7335 , n174484 );
or ( n7336 , n7334 , n7335 );
not ( n7337 , n1470 );
buf ( n174789 , n784 );
buf ( n174790 , n830 );
xor ( n7340 , n174789 , n174790 );
buf ( n174792 , n7340 );
nand ( n174793 , n7337 , n174792 );
nand ( n7343 , n7336 , n174793 );
buf ( n174795 , n7343 );
not ( n7345 , n174795 );
buf ( n174797 , n7345 );
buf ( n174798 , n174797 );
not ( n7348 , n174798 );
or ( n7349 , n7333 , n7348 );
buf ( n174801 , n786 );
buf ( n174802 , n828 );
xor ( n7352 , n174801 , n174802 );
buf ( n174804 , n7352 );
buf ( n174805 , n174804 );
not ( n7355 , n174805 );
buf ( n174807 , n168549 );
not ( n7357 , n174807 );
or ( n174809 , n7355 , n7357 );
buf ( n174810 , n168559 );
buf ( n174811 , n174629 );
nand ( n7364 , n174810 , n174811 );
buf ( n174813 , n7364 );
buf ( n174814 , n174813 );
nand ( n174815 , n174809 , n174814 );
buf ( n174816 , n174815 );
buf ( n174817 , n174816 );
nand ( n7370 , n7349 , n174817 );
buf ( n174819 , n7370 );
buf ( n174820 , n174819 );
buf ( n174821 , n174782 );
not ( n7374 , n174821 );
buf ( n174823 , n7343 );
nand ( n7376 , n7374 , n174823 );
buf ( n174825 , n7376 );
buf ( n174826 , n174825 );
nand ( n7379 , n174820 , n174826 );
buf ( n174828 , n7379 );
buf ( n174829 , n174828 );
not ( n7382 , n174829 );
buf ( n174831 , n7382 );
buf ( n174832 , n174831 );
not ( n7385 , n174832 );
buf ( n174834 , n788 );
buf ( n174835 , n826 );
xor ( n7388 , n174834 , n174835 );
buf ( n174837 , n7388 );
buf ( n174838 , n174837 );
not ( n7391 , n174838 );
buf ( n174840 , n7391 );
or ( n7393 , n174840 , n168667 );
or ( n7394 , n171330 , n174600 );
nand ( n7395 , n7393 , n7394 );
buf ( n174844 , n7395 );
not ( n7397 , n174844 );
xor ( n7398 , n820 , n794 );
buf ( n174847 , n7398 );
not ( n7400 , n174847 );
buf ( n174849 , n2251 );
not ( n7402 , n174849 );
or ( n7403 , n7400 , n7402 );
buf ( n174852 , n2513 );
buf ( n174853 , n7220 );
nand ( n7406 , n174852 , n174853 );
buf ( n174855 , n7406 );
buf ( n174856 , n174855 );
nand ( n7409 , n7403 , n174856 );
buf ( n174858 , n7409 );
buf ( n174859 , n174858 );
not ( n7412 , n174859 );
or ( n7413 , n7397 , n7412 );
buf ( n174862 , n7395 );
buf ( n174863 , n174858 );
or ( n7416 , n174862 , n174863 );
buf ( n174865 , n796 );
buf ( n174866 , n818 );
xor ( n7419 , n174865 , n174866 );
buf ( n174868 , n7419 );
buf ( n174869 , n174868 );
not ( n174870 , n174869 );
buf ( n174871 , n1321 );
not ( n7424 , n174871 );
or ( n7425 , n174870 , n7424 );
buf ( n174874 , n168806 );
buf ( n174875 , n174708 );
nand ( n7428 , n174874 , n174875 );
buf ( n174877 , n7428 );
buf ( n174878 , n174877 );
nand ( n7431 , n7425 , n174878 );
buf ( n174880 , n7431 );
buf ( n174881 , n174880 );
nand ( n7434 , n7416 , n174881 );
buf ( n174883 , n7434 );
buf ( n174884 , n174883 );
nand ( n7437 , n7413 , n174884 );
buf ( n174886 , n7437 );
not ( n7439 , n174886 );
buf ( n174888 , n7439 );
not ( n7441 , n174888 );
or ( n7442 , n7385 , n7441 );
buf ( n174891 , n790 );
buf ( n174892 , n824 );
xor ( n7445 , n174891 , n174892 );
buf ( n174894 , n7445 );
buf ( n174895 , n174894 );
not ( n7448 , n174895 );
buf ( n174897 , n170100 );
not ( n7450 , n174897 );
or ( n7451 , n7448 , n7450 );
buf ( n174900 , n169802 );
buf ( n174901 , n174525 );
nand ( n7454 , n174900 , n174901 );
buf ( n174903 , n7454 );
buf ( n174904 , n174903 );
nand ( n7457 , n7451 , n174904 );
buf ( n174906 , n7457 );
not ( n7459 , n174906 );
buf ( n174908 , n171049 );
xor ( n7461 , n822 , n792 );
buf ( n174910 , n7461 );
and ( n7463 , n174908 , n174910 );
buf ( n174912 , n171055 );
buf ( n174913 , n174577 );
and ( n7466 , n174912 , n174913 );
nor ( n7467 , n7463 , n7466 );
buf ( n174916 , n7467 );
buf ( n174917 , n174916 );
not ( n7470 , n174917 );
buf ( n174919 , n7470 );
not ( n174920 , n174919 );
or ( n7476 , n7459 , n174920 );
buf ( n174922 , n174916 );
not ( n7478 , n174922 );
buf ( n174924 , n174906 );
not ( n7480 , n174924 );
buf ( n174926 , n7480 );
buf ( n174927 , n174926 );
not ( n7483 , n174927 );
or ( n7484 , n7478 , n7483 );
buf ( n174930 , n798 );
buf ( n174931 , n816 );
xor ( n7487 , n174930 , n174931 );
buf ( n174933 , n7487 );
buf ( n174934 , n174933 );
not ( n7490 , n174934 );
buf ( n174936 , n169836 );
buf ( n7492 , n174936 );
buf ( n174938 , n7492 );
buf ( n174939 , n174938 );
not ( n7495 , n174939 );
or ( n7496 , n7490 , n7495 );
buf ( n174942 , n169320 );
buf ( n174943 , n174545 );
nand ( n7499 , n174942 , n174943 );
buf ( n174945 , n7499 );
buf ( n174946 , n174945 );
nand ( n7502 , n7496 , n174946 );
buf ( n174948 , n7502 );
buf ( n174949 , n174948 );
nand ( n7505 , n7484 , n174949 );
buf ( n174951 , n7505 );
nand ( n7507 , n7476 , n174951 );
buf ( n174953 , n7507 );
nand ( n7509 , n7442 , n174953 );
buf ( n174955 , n7509 );
buf ( n174956 , n174955 );
buf ( n174957 , n174886 );
buf ( n174958 , n174828 );
nand ( n7514 , n174957 , n174958 );
buf ( n174960 , n7514 );
buf ( n174961 , n174960 );
nand ( n7517 , n174956 , n174961 );
buf ( n174963 , n7517 );
not ( n7519 , n174963 );
xor ( n7520 , n7116 , n7189 );
xor ( n7521 , n7520 , n174647 );
not ( n7522 , n7521 );
or ( n7523 , n7519 , n7522 );
or ( n7524 , n7521 , n174963 );
not ( n7525 , n7093 );
not ( n7526 , n7067 );
or ( n174972 , n7525 , n7526 );
or ( n7528 , n7067 , n7093 );
nand ( n7529 , n174972 , n7528 );
buf ( n174975 , n7529 );
buf ( n174976 , n7080 );
xnor ( n7532 , n174975 , n174976 );
buf ( n174978 , n7532 );
buf ( n174979 , n174978 );
not ( n7535 , n174979 );
buf ( n174981 , n7535 );
buf ( n174982 , n174981 );
not ( n7538 , n174982 );
xor ( n7539 , n174720 , n174686 );
buf ( n174985 , n7539 );
buf ( n174986 , n174698 );
xnor ( n7542 , n174985 , n174986 );
buf ( n174988 , n7542 );
not ( n174989 , n174988 );
buf ( n174990 , n174989 );
not ( n7546 , n174990 );
or ( n7547 , n7538 , n7546 );
buf ( n174993 , n174988 );
not ( n7549 , n174993 );
buf ( n174995 , n174978 );
not ( n7551 , n174995 );
or ( n7552 , n7549 , n7551 );
xor ( n7553 , n174623 , n174641 );
buf ( n174999 , n7553 );
buf ( n7555 , n174608 );
buf ( n175001 , n7555 );
and ( n7557 , n174999 , n175001 );
not ( n7558 , n174999 );
not ( n7559 , n7555 );
buf ( n175005 , n7559 );
and ( n7561 , n7558 , n175005 );
nor ( n7562 , n7557 , n7561 );
buf ( n175008 , n7562 );
buf ( n175009 , n175008 );
nand ( n7565 , n7552 , n175009 );
buf ( n175011 , n7565 );
buf ( n175012 , n175011 );
nand ( n7568 , n7547 , n175012 );
buf ( n175014 , n7568 );
nand ( n7570 , n7524 , n175014 );
nand ( n7571 , n7523 , n7570 );
xor ( n7572 , n174778 , n7571 );
xor ( n7573 , n174571 , n7196 );
xor ( n7574 , n7573 , n7288 );
and ( n7575 , n7572 , n7574 );
and ( n7576 , n174778 , n7571 );
or ( n7577 , n7575 , n7576 );
buf ( n175023 , n7577 );
xor ( n7582 , n174775 , n175023 );
xor ( n7583 , n174568 , n174742 );
xor ( n7584 , n7583 , n7302 );
buf ( n175027 , n7584 );
and ( n7586 , n7582 , n175027 );
and ( n175029 , n174775 , n175023 );
or ( n7588 , n7586 , n175029 );
buf ( n175031 , n7588 );
buf ( n175032 , n175031 );
nor ( n7591 , n174774 , n175032 );
buf ( n175034 , n7591 );
xor ( n7593 , n174775 , n175023 );
xor ( n7594 , n7593 , n175027 );
buf ( n175037 , n7594 );
buf ( n175038 , n844 );
buf ( n175039 , n7286 );
not ( n7598 , n175039 );
xor ( n7599 , n174726 , n174672 );
buf ( n175042 , n7599 );
not ( n7601 , n175042 );
or ( n7602 , n7598 , n7601 );
buf ( n175045 , n7599 );
buf ( n175046 , n7286 );
or ( n175047 , n175045 , n175046 );
nand ( n7606 , n7602 , n175047 );
buf ( n175049 , n7606 );
buf ( n7608 , n175049 );
not ( n7609 , n7608 );
buf ( n175052 , n799 );
buf ( n175053 , n817 );
or ( n7612 , n175052 , n175053 );
buf ( n175055 , n818 );
nand ( n7614 , n7612 , n175055 );
buf ( n175057 , n7614 );
buf ( n175058 , n175057 );
buf ( n175059 , n799 );
buf ( n175060 , n817 );
nand ( n7619 , n175059 , n175060 );
buf ( n175062 , n7619 );
buf ( n175063 , n175062 );
buf ( n175064 , n816 );
and ( n7623 , n175058 , n175063 , n175064 );
buf ( n175066 , n7623 );
buf ( n175067 , n175066 );
buf ( n175068 , n785 );
buf ( n175069 , n830 );
xor ( n7628 , n175068 , n175069 );
buf ( n175071 , n7628 );
buf ( n175072 , n175071 );
not ( n7631 , n175072 );
buf ( n175074 , n168471 );
not ( n7633 , n175074 );
or ( n7634 , n7631 , n7633 );
buf ( n175077 , n174792 );
buf ( n175078 , n831 );
nand ( n7637 , n175077 , n175078 );
buf ( n175080 , n7637 );
buf ( n175081 , n175080 );
nand ( n7640 , n7634 , n175081 );
buf ( n175083 , n7640 );
buf ( n175084 , n175083 );
and ( n7643 , n175067 , n175084 );
buf ( n175086 , n7643 );
buf ( n175087 , n791 );
buf ( n175088 , n824 );
xor ( n175089 , n175087 , n175088 );
buf ( n175090 , n175089 );
buf ( n175091 , n175090 );
not ( n7650 , n175091 );
buf ( n175093 , n170100 );
not ( n175094 , n175093 );
or ( n7653 , n7650 , n175094 );
buf ( n175096 , n169802 );
buf ( n175097 , n174894 );
nand ( n7656 , n175096 , n175097 );
buf ( n175099 , n7656 );
buf ( n175100 , n175099 );
nand ( n7659 , n7653 , n175100 );
buf ( n175102 , n7659 );
not ( n7661 , n175102 );
not ( n7662 , n169320 );
not ( n7663 , n174933 );
or ( n7664 , n7662 , n7663 );
not ( n7665 , n169836 );
buf ( n175108 , n799 );
buf ( n175109 , n816 );
xor ( n7668 , n175108 , n175109 );
buf ( n175111 , n7668 );
not ( n175112 , n175111 );
or ( n7671 , n7665 , n175112 );
nand ( n7672 , n7664 , n7671 );
not ( n7673 , n7672 );
or ( n7674 , n7661 , n7673 );
or ( n7675 , n7672 , n175102 );
buf ( n175118 , n787 );
buf ( n175119 , n828 );
xor ( n7678 , n175118 , n175119 );
buf ( n175121 , n7678 );
buf ( n175122 , n175121 );
not ( n7681 , n175122 );
buf ( n175124 , n168549 );
not ( n7683 , n175124 );
or ( n7684 , n7681 , n7683 );
buf ( n175127 , n168559 );
buf ( n175128 , n174804 );
nand ( n7687 , n175127 , n175128 );
buf ( n175130 , n7687 );
buf ( n175131 , n175130 );
nand ( n7690 , n7684 , n175131 );
buf ( n175133 , n7690 );
nand ( n7692 , n7675 , n175133 );
nand ( n7693 , n7674 , n7692 );
xor ( n7694 , n175086 , n7693 );
buf ( n175137 , n795 );
buf ( n175138 , n820 );
xor ( n7697 , n175137 , n175138 );
buf ( n175140 , n7697 );
buf ( n175141 , n175140 );
not ( n7700 , n175141 );
buf ( n175143 , n2251 );
not ( n7702 , n175143 );
or ( n7703 , n7700 , n7702 );
buf ( n175146 , n7398 );
buf ( n175147 , n168656 );
nand ( n7706 , n175146 , n175147 );
buf ( n175149 , n7706 );
buf ( n175150 , n175149 );
nand ( n7709 , n7703 , n175150 );
buf ( n175152 , n7709 );
buf ( n175153 , n175152 );
not ( n175154 , n169411 );
xor ( n7716 , n822 , n793 );
not ( n7717 , n7716 );
or ( n7718 , n175154 , n7717 );
buf ( n175158 , n169423 );
buf ( n175159 , n7461 );
nand ( n175160 , n175158 , n175159 );
buf ( n175161 , n175160 );
nand ( n7723 , n7718 , n175161 );
buf ( n175163 , n7723 );
or ( n7725 , n175153 , n175163 );
buf ( n175165 , n789 );
buf ( n175166 , n826 );
xor ( n7728 , n175165 , n175166 );
buf ( n175168 , n7728 );
buf ( n175169 , n175168 );
not ( n7731 , n175169 );
buf ( n175171 , n1621 );
not ( n7733 , n175171 );
or ( n7734 , n7731 , n7733 );
buf ( n175174 , n169081 );
buf ( n175175 , n174837 );
nand ( n7737 , n175174 , n175175 );
buf ( n175177 , n7737 );
buf ( n175178 , n175177 );
nand ( n7740 , n7734 , n175178 );
buf ( n175180 , n7740 );
buf ( n175181 , n175180 );
nand ( n7743 , n7725 , n175181 );
buf ( n175183 , n7743 );
buf ( n175184 , n175183 );
buf ( n175185 , n175152 );
buf ( n175186 , n7723 );
nand ( n7748 , n175185 , n175186 );
buf ( n175188 , n7748 );
buf ( n175189 , n175188 );
nand ( n7751 , n175184 , n175189 );
buf ( n175191 , n7751 );
and ( n7753 , n7694 , n175191 );
and ( n7754 , n175086 , n7693 );
or ( n7755 , n7753 , n7754 );
buf ( n175195 , n7755 );
not ( n7757 , n175195 );
not ( n7758 , n174886 );
not ( n7759 , n174828 );
or ( n175199 , n7758 , n7759 );
nand ( n7761 , n174831 , n7439 );
nand ( n7762 , n175199 , n7761 );
xor ( n7763 , n7762 , n7507 );
not ( n7764 , n7763 );
buf ( n175204 , n7764 );
not ( n7766 , n175204 );
or ( n7767 , n7757 , n7766 );
buf ( n175207 , n7763 );
not ( n7769 , n175207 );
buf ( n175209 , n7755 );
not ( n7771 , n175209 );
buf ( n175211 , n7771 );
buf ( n175212 , n175211 );
not ( n7774 , n175212 );
or ( n7775 , n7769 , n7774 );
not ( n7776 , n174782 );
not ( n175216 , n7776 );
not ( n7778 , n7343 );
or ( n7779 , n175216 , n7778 );
or ( n7780 , n7776 , n7343 );
nand ( n7781 , n7779 , n7780 );
xnor ( n175221 , n174816 , n7781 );
buf ( n175222 , n175221 );
not ( n7784 , n7395 );
not ( n7785 , n7784 );
not ( n7786 , n174858 );
not ( n7787 , n174880 );
not ( n7788 , n7787 );
or ( n7789 , n7786 , n7788 );
not ( n175229 , n174858 );
nand ( n7791 , n175229 , n174880 );
nand ( n7792 , n7789 , n7791 );
not ( n7793 , n7792 );
or ( n7794 , n7785 , n7793 );
or ( n7795 , n7792 , n7784 );
nand ( n7796 , n7794 , n7795 );
buf ( n175236 , n7796 );
xor ( n7798 , n175222 , n175236 );
xor ( n7799 , n174926 , n174948 );
xnor ( n7800 , n7799 , n174919 );
buf ( n175240 , n7800 );
and ( n7802 , n7798 , n175240 );
and ( n7803 , n175222 , n175236 );
or ( n7804 , n7802 , n7803 );
buf ( n175244 , n7804 );
buf ( n175245 , n175244 );
nand ( n7807 , n7775 , n175245 );
buf ( n175247 , n7807 );
buf ( n175248 , n175247 );
nand ( n7810 , n7767 , n175248 );
buf ( n175250 , n7810 );
not ( n7812 , n175250 );
or ( n7813 , n7609 , n7812 );
or ( n7814 , n175250 , n7608 );
xor ( n7815 , n174963 , n7521 );
xor ( n7816 , n7815 , n175014 );
nand ( n7817 , n7814 , n7816 );
nand ( n7818 , n7813 , n7817 );
buf ( n175258 , n7818 );
xor ( n7820 , n175038 , n175258 );
xor ( n175260 , n174778 , n7571 );
xor ( n7822 , n175260 , n7574 );
buf ( n175262 , n7822 );
and ( n7824 , n7820 , n175262 );
and ( n7825 , n175038 , n175258 );
or ( n7826 , n7824 , n7825 );
buf ( n175266 , n7826 );
nor ( n7828 , n175037 , n175266 );
nor ( n7829 , n175034 , n7828 );
nand ( n7830 , n7319 , n7829 );
not ( n7831 , n7830 );
buf ( n175271 , n845 );
buf ( n175272 , n174978 );
not ( n7834 , n175272 );
buf ( n175274 , n175008 );
not ( n7836 , n175274 );
and ( n7837 , n7834 , n7836 );
buf ( n175277 , n174978 );
buf ( n175278 , n175008 );
and ( n7843 , n175277 , n175278 );
nor ( n7844 , n7837 , n7843 );
buf ( n175281 , n7844 );
buf ( n175282 , n175281 );
not ( n175283 , n174989 );
buf ( n175284 , n175283 );
and ( n7849 , n175282 , n175284 );
not ( n7850 , n175282 );
buf ( n175287 , n174989 );
and ( n7852 , n7850 , n175287 );
nor ( n7853 , n7849 , n7852 );
buf ( n175290 , n7853 );
buf ( n175291 , n175290 );
buf ( n175292 , n797 );
buf ( n175293 , n818 );
xor ( n7858 , n175292 , n175293 );
buf ( n175295 , n7858 );
buf ( n175296 , n175295 );
not ( n7861 , n175296 );
buf ( n175298 , n2566 );
not ( n7863 , n175298 );
or ( n7864 , n7861 , n7863 );
buf ( n175301 , n168806 );
buf ( n175302 , n174868 );
nand ( n7867 , n175301 , n175302 );
buf ( n175304 , n7867 );
buf ( n175305 , n175304 );
nand ( n7870 , n7864 , n175305 );
buf ( n175307 , n7870 );
buf ( n175308 , n175307 );
xor ( n7873 , n175067 , n175084 );
buf ( n175310 , n7873 );
buf ( n175311 , n175310 );
xor ( n7876 , n175308 , n175311 );
buf ( n175313 , n169320 );
buf ( n175314 , n799 );
and ( n7879 , n175313 , n175314 );
buf ( n175316 , n7879 );
buf ( n175317 , n175316 );
buf ( n175318 , n786 );
buf ( n175319 , n830 );
xor ( n7884 , n175318 , n175319 );
buf ( n175321 , n7884 );
buf ( n175322 , n175321 );
not ( n7887 , n175322 );
buf ( n175324 , n1471 );
not ( n7889 , n175324 );
or ( n175326 , n7887 , n7889 );
buf ( n175327 , n175071 );
buf ( n175328 , n831 );
nand ( n7893 , n175327 , n175328 );
buf ( n175330 , n7893 );
buf ( n175331 , n175330 );
nand ( n7896 , n175326 , n175331 );
buf ( n175333 , n7896 );
buf ( n175334 , n175333 );
xor ( n7899 , n175317 , n175334 );
buf ( n175336 , n788 );
buf ( n175337 , n828 );
xor ( n7902 , n175336 , n175337 );
buf ( n175339 , n7902 );
buf ( n175340 , n175339 );
not ( n7905 , n175340 );
buf ( n175342 , n1742 );
not ( n7907 , n175342 );
or ( n7908 , n7905 , n7907 );
buf ( n175345 , n168559 );
buf ( n175346 , n175121 );
nand ( n7911 , n175345 , n175346 );
buf ( n175348 , n7911 );
buf ( n175349 , n175348 );
nand ( n7914 , n7908 , n175349 );
buf ( n175351 , n7914 );
buf ( n175352 , n175351 );
and ( n175353 , n7899 , n175352 );
and ( n7918 , n175317 , n175334 );
or ( n7919 , n175353 , n7918 );
buf ( n175356 , n7919 );
buf ( n175357 , n175356 );
and ( n175358 , n7876 , n175357 );
and ( n7923 , n175308 , n175311 );
or ( n7924 , n175358 , n7923 );
buf ( n175361 , n7924 );
buf ( n175362 , n175361 );
xor ( n7927 , n175086 , n7693 );
xor ( n7928 , n7927 , n175191 );
buf ( n175365 , n7928 );
xor ( n7930 , n175362 , n175365 );
buf ( n175367 , n794 );
buf ( n175368 , n822 );
xor ( n7933 , n175367 , n175368 );
buf ( n175370 , n7933 );
not ( n7935 , n175370 );
not ( n7936 , n171049 );
or ( n7937 , n7935 , n7936 );
buf ( n175374 , n169423 );
buf ( n175375 , n7716 );
nand ( n7940 , n175374 , n175375 );
buf ( n175377 , n7940 );
nand ( n7942 , n7937 , n175377 );
not ( n7943 , n7942 );
buf ( n175380 , n792 );
buf ( n175381 , n824 );
xor ( n7946 , n175380 , n175381 );
buf ( n175383 , n7946 );
not ( n7948 , n175383 );
not ( n7949 , n170100 );
or ( n7950 , n7948 , n7949 );
buf ( n175387 , n169802 );
buf ( n175388 , n175090 );
nand ( n7953 , n175387 , n175388 );
buf ( n175390 , n7953 );
nand ( n7955 , n7950 , n175390 );
not ( n7956 , n7955 );
or ( n7957 , n7943 , n7956 );
or ( n7958 , n7955 , n7942 );
xor ( n7959 , n826 , n790 );
buf ( n175396 , n7959 );
not ( n7961 , n175396 );
buf ( n175398 , n173773 );
not ( n7963 , n175398 );
buf ( n175400 , n7963 );
buf ( n175401 , n175400 );
not ( n7966 , n175401 );
or ( n7967 , n7961 , n7966 );
buf ( n175404 , n169081 );
buf ( n175405 , n175168 );
nand ( n7970 , n175404 , n175405 );
buf ( n175407 , n7970 );
buf ( n175408 , n175407 );
nand ( n7973 , n7967 , n175408 );
buf ( n175410 , n7973 );
nand ( n7975 , n7958 , n175410 );
nand ( n7976 , n7957 , n7975 );
buf ( n175413 , n7976 );
xor ( n7978 , n175102 , n175133 );
xor ( n7979 , n7978 , n7672 );
buf ( n175416 , n7979 );
xor ( n7981 , n175413 , n175416 );
buf ( n175418 , n7723 );
not ( n7983 , n175418 );
not ( n7984 , n175180 );
xor ( n7985 , n175152 , n7984 );
buf ( n175422 , n7985 );
not ( n7987 , n175422 );
or ( n7988 , n7983 , n7987 );
buf ( n175425 , n7985 );
buf ( n175426 , n7723 );
or ( n7991 , n175425 , n175426 );
nand ( n175428 , n7988 , n7991 );
buf ( n175429 , n175428 );
buf ( n175430 , n175429 );
and ( n7998 , n7981 , n175430 );
and ( n7999 , n175413 , n175416 );
or ( n8000 , n7998 , n7999 );
buf ( n175434 , n8000 );
buf ( n175435 , n175434 );
and ( n8003 , n7930 , n175435 );
and ( n8004 , n175362 , n175365 );
or ( n175438 , n8003 , n8004 );
buf ( n175439 , n175438 );
buf ( n175440 , n175439 );
xor ( n8008 , n175291 , n175440 );
buf ( n175442 , n7764 );
not ( n8010 , n175442 );
buf ( n175444 , n175211 );
not ( n8012 , n175444 );
or ( n8013 , n8010 , n8012 );
buf ( n175447 , n7763 );
buf ( n175448 , n7755 );
nand ( n8016 , n175447 , n175448 );
buf ( n175450 , n8016 );
buf ( n175451 , n175450 );
nand ( n8019 , n8013 , n175451 );
buf ( n175453 , n8019 );
buf ( n175454 , n175453 );
buf ( n175455 , n175244 );
and ( n8023 , n175454 , n175455 );
not ( n8024 , n175454 );
buf ( n175458 , n175244 );
not ( n8026 , n175458 );
buf ( n175460 , n8026 );
buf ( n175461 , n175460 );
and ( n8029 , n8024 , n175461 );
nor ( n8030 , n8023 , n8029 );
buf ( n175464 , n8030 );
buf ( n175465 , n175464 );
and ( n8033 , n8008 , n175465 );
and ( n8034 , n175291 , n175440 );
or ( n8035 , n8033 , n8034 );
buf ( n175469 , n8035 );
buf ( n175470 , n175469 );
xor ( n8038 , n175271 , n175470 );
xor ( n8039 , n175049 , n175250 );
xor ( n8040 , n8039 , n7816 );
buf ( n175474 , n8040 );
xor ( n8042 , n8038 , n175474 );
buf ( n175476 , n8042 );
buf ( n175477 , n175476 );
buf ( n175478 , n846 );
xor ( n8046 , n175222 , n175236 );
xor ( n8047 , n8046 , n175240 );
buf ( n175481 , n8047 );
buf ( n175482 , n175481 );
buf ( n175483 , n787 );
buf ( n175484 , n830 );
xor ( n8052 , n175483 , n175484 );
buf ( n175486 , n8052 );
buf ( n175487 , n175486 );
not ( n8055 , n175487 );
buf ( n175489 , n168471 );
not ( n8057 , n175489 );
or ( n8058 , n8055 , n8057 );
buf ( n175492 , n175321 );
buf ( n175493 , n831 );
nand ( n8061 , n175492 , n175493 );
buf ( n175495 , n8061 );
buf ( n175496 , n175495 );
nand ( n8064 , n8058 , n175496 );
buf ( n175498 , n8064 );
buf ( n175499 , n175498 );
buf ( n175500 , n799 );
buf ( n175501 , n819 );
or ( n8069 , n175500 , n175501 );
buf ( n175503 , n820 );
nand ( n8071 , n8069 , n175503 );
buf ( n175505 , n8071 );
buf ( n175506 , n175505 );
buf ( n175507 , n799 );
buf ( n175508 , n819 );
nand ( n175509 , n175507 , n175508 );
buf ( n175510 , n175509 );
buf ( n175511 , n175510 );
buf ( n175512 , n818 );
nand ( n8080 , n175506 , n175511 , n175512 );
buf ( n175514 , n8080 );
buf ( n175515 , n175514 );
not ( n8083 , n175515 );
buf ( n175517 , n8083 );
buf ( n175518 , n175517 );
and ( n8086 , n175499 , n175518 );
buf ( n175520 , n8086 );
buf ( n175521 , n175520 );
xor ( n8089 , n820 , n796 );
buf ( n175523 , n8089 );
not ( n8091 , n175523 );
buf ( n175525 , n2108 );
not ( n8093 , n175525 );
or ( n8094 , n8091 , n8093 );
buf ( n175528 , n2513 );
buf ( n175529 , n175140 );
nand ( n8097 , n175528 , n175529 );
buf ( n175531 , n8097 );
buf ( n175532 , n175531 );
nand ( n8100 , n8094 , n175532 );
buf ( n175534 , n8100 );
buf ( n175535 , n175534 );
nor ( n8103 , n175521 , n175535 );
buf ( n175537 , n8103 );
buf ( n175538 , n175537 );
buf ( n175539 , n798 );
buf ( n175540 , n818 );
xor ( n175541 , n175539 , n175540 );
buf ( n175542 , n175541 );
buf ( n175543 , n175542 );
not ( n8111 , n175543 );
buf ( n175545 , n1321 );
not ( n8113 , n175545 );
or ( n8114 , n8111 , n8113 );
buf ( n175548 , n168806 );
buf ( n175549 , n175295 );
nand ( n8117 , n175548 , n175549 );
buf ( n175551 , n8117 );
buf ( n175552 , n175551 );
nand ( n8120 , n8114 , n175552 );
buf ( n175554 , n8120 );
buf ( n175555 , n175554 );
not ( n8123 , n175555 );
buf ( n175557 , n8123 );
buf ( n175558 , n175557 );
or ( n8126 , n175538 , n175558 );
buf ( n175560 , n175534 );
buf ( n175561 , n175520 );
nand ( n8129 , n175560 , n175561 );
buf ( n175563 , n8129 );
buf ( n175564 , n175563 );
nand ( n8132 , n8126 , n175564 );
buf ( n175566 , n8132 );
buf ( n175567 , n175566 );
xor ( n8135 , n175308 , n175311 );
xor ( n8136 , n8135 , n175357 );
buf ( n175570 , n8136 );
buf ( n175571 , n175570 );
xor ( n8142 , n175567 , n175571 );
xor ( n8143 , n175317 , n175334 );
xor ( n8144 , n8143 , n175352 );
buf ( n175575 , n8144 );
xor ( n8146 , n826 , n791 );
buf ( n175577 , n8146 );
not ( n8148 , n175577 );
buf ( n175579 , n4337 );
not ( n8150 , n175579 );
or ( n8151 , n8148 , n8150 );
buf ( n175582 , n169081 );
buf ( n175583 , n7959 );
nand ( n8154 , n175582 , n175583 );
buf ( n175585 , n8154 );
buf ( n175586 , n175585 );
nand ( n8157 , n8151 , n175586 );
buf ( n175588 , n8157 );
buf ( n175589 , n175588 );
not ( n8160 , n175589 );
xor ( n175591 , n820 , n797 );
buf ( n175592 , n175591 );
not ( n8163 , n175592 );
buf ( n175594 , n2251 );
not ( n8165 , n175594 );
or ( n8166 , n8163 , n8165 );
buf ( n175597 , n168656 );
buf ( n175598 , n8089 );
nand ( n8169 , n175597 , n175598 );
buf ( n175600 , n8169 );
buf ( n175601 , n175600 );
nand ( n8172 , n8166 , n175601 );
buf ( n175603 , n8172 );
buf ( n175604 , n175603 );
not ( n8175 , n175604 );
or ( n8176 , n8160 , n8175 );
buf ( n175607 , n175603 );
buf ( n175608 , n175588 );
or ( n8179 , n175607 , n175608 );
buf ( n175610 , n799 );
buf ( n175611 , n818 );
xor ( n8182 , n175610 , n175611 );
buf ( n175613 , n8182 );
buf ( n175614 , n175613 );
not ( n8185 , n175614 );
buf ( n175616 , n1321 );
not ( n8187 , n175616 );
or ( n8188 , n8185 , n8187 );
buf ( n175619 , n168806 );
buf ( n175620 , n175542 );
nand ( n8191 , n175619 , n175620 );
buf ( n175622 , n8191 );
buf ( n175623 , n175622 );
nand ( n8194 , n8188 , n175623 );
buf ( n175625 , n8194 );
buf ( n175626 , n175625 );
nand ( n8197 , n8179 , n175626 );
buf ( n175628 , n8197 );
buf ( n175629 , n175628 );
nand ( n8200 , n8176 , n175629 );
buf ( n175631 , n8200 );
and ( n8202 , n175575 , n175631 );
not ( n8203 , n8202 );
not ( n8204 , n175575 );
not ( n8205 , n8204 );
not ( n8206 , n175631 );
not ( n8207 , n8206 );
or ( n8208 , n8205 , n8207 );
xor ( n8209 , n828 , n789 );
buf ( n175640 , n8209 );
not ( n8211 , n175640 );
buf ( n175642 , n170990 );
not ( n8213 , n175642 );
or ( n8214 , n8211 , n8213 );
buf ( n175645 , n168559 );
buf ( n175646 , n175339 );
nand ( n8217 , n175645 , n175646 );
buf ( n175648 , n8217 );
buf ( n175649 , n175648 );
nand ( n8220 , n8214 , n175649 );
buf ( n175651 , n8220 );
not ( n8222 , n175651 );
buf ( n175653 , n793 );
buf ( n175654 , n824 );
xor ( n8225 , n175653 , n175654 );
buf ( n175656 , n8225 );
buf ( n175657 , n175656 );
not ( n8228 , n175657 );
buf ( n175659 , n170100 );
not ( n8230 , n175659 );
or ( n8231 , n8228 , n8230 );
buf ( n175662 , n169799 );
not ( n8233 , n175662 );
buf ( n175664 , n8233 );
buf ( n175665 , n175664 );
buf ( n175666 , n175383 );
nand ( n8237 , n175665 , n175666 );
buf ( n175668 , n8237 );
buf ( n175669 , n175668 );
nand ( n175670 , n8231 , n175669 );
buf ( n175671 , n175670 );
not ( n8242 , n175671 );
nand ( n8243 , n8222 , n8242 );
not ( n8244 , n8243 );
buf ( n175675 , n795 );
buf ( n175676 , n822 );
xor ( n8247 , n175675 , n175676 );
buf ( n175678 , n8247 );
buf ( n175679 , n175678 );
not ( n8250 , n175679 );
buf ( n175681 , n171049 );
not ( n8252 , n175681 );
or ( n8253 , n8250 , n8252 );
buf ( n175684 , n171055 );
buf ( n175685 , n175370 );
nand ( n8256 , n175684 , n175685 );
buf ( n175687 , n8256 );
buf ( n175688 , n175687 );
nand ( n8259 , n8253 , n175688 );
buf ( n175690 , n8259 );
not ( n8261 , n175690 );
or ( n8262 , n8244 , n8261 );
nand ( n8263 , n175671 , n175651 );
nand ( n8264 , n8262 , n8263 );
nand ( n8265 , n8208 , n8264 );
nand ( n8266 , n8203 , n8265 );
buf ( n175697 , n8266 );
and ( n8268 , n8142 , n175697 );
and ( n8269 , n175567 , n175571 );
or ( n8270 , n8268 , n8269 );
buf ( n175701 , n8270 );
buf ( n175702 , n175701 );
xor ( n8273 , n175482 , n175702 );
xor ( n8274 , n175362 , n175365 );
xor ( n8275 , n8274 , n175435 );
buf ( n175706 , n8275 );
buf ( n175707 , n175706 );
and ( n8278 , n8273 , n175707 );
and ( n8279 , n175482 , n175702 );
or ( n8280 , n8278 , n8279 );
buf ( n175711 , n8280 );
buf ( n175712 , n175711 );
xor ( n8283 , n175478 , n175712 );
xor ( n8284 , n175291 , n175440 );
xor ( n8285 , n8284 , n175465 );
buf ( n175716 , n8285 );
buf ( n175717 , n175716 );
and ( n8288 , n8283 , n175717 );
and ( n8289 , n175478 , n175712 );
or ( n8290 , n8288 , n8289 );
buf ( n175721 , n8290 );
buf ( n175722 , n175721 );
nor ( n8293 , n175477 , n175722 );
buf ( n175724 , n8293 );
xor ( n8295 , n175271 , n175470 );
and ( n8296 , n8295 , n175474 );
and ( n8297 , n175271 , n175470 );
or ( n8298 , n8296 , n8297 );
buf ( n175729 , n8298 );
buf ( n175730 , n175729 );
xor ( n8301 , n175038 , n175258 );
xor ( n8302 , n8301 , n175262 );
buf ( n175733 , n8302 );
buf ( n175734 , n175733 );
nor ( n8305 , n175730 , n175734 );
buf ( n175736 , n8305 );
nor ( n8307 , n175724 , n175736 );
not ( n8308 , n8307 );
buf ( n175739 , n848 );
not ( n8310 , n8264 );
not ( n8311 , n8204 );
not ( n175742 , n175631 );
or ( n8316 , n8311 , n175742 );
nand ( n8317 , n8206 , n175575 );
nand ( n8318 , n8316 , n8317 );
nand ( n8319 , n8310 , n8318 );
nand ( n8320 , n8202 , n8264 );
nand ( n175748 , n8264 , n8204 , n8206 );
nand ( n8322 , n8319 , n8320 , n175748 );
buf ( n175750 , n8322 );
xor ( n8324 , n175651 , n8242 );
not ( n8325 , n175690 );
xor ( n8326 , n8324 , n8325 );
xor ( n8327 , n175625 , n175588 );
xor ( n8328 , n8327 , n175603 );
xor ( n8329 , n8326 , n8328 );
buf ( n175757 , n826 );
buf ( n175758 , n792 );
xor ( n8332 , n175757 , n175758 );
buf ( n175760 , n8332 );
buf ( n175761 , n175760 );
not ( n8335 , n175761 );
buf ( n175763 , n1621 );
not ( n8337 , n175763 );
or ( n175765 , n8335 , n8337 );
buf ( n175766 , n169081 );
buf ( n175767 , n8146 );
nand ( n8341 , n175766 , n175767 );
buf ( n175769 , n8341 );
buf ( n175770 , n175769 );
nand ( n8344 , n175765 , n175770 );
buf ( n175772 , n8344 );
buf ( n175773 , n175772 );
buf ( n175774 , n791 );
buf ( n175775 , n828 );
xor ( n8349 , n175774 , n175775 );
buf ( n175777 , n8349 );
buf ( n175778 , n175777 );
not ( n8352 , n175778 );
buf ( n175780 , n170990 );
not ( n8354 , n175780 );
or ( n8355 , n8352 , n8354 );
buf ( n175783 , n168559 );
xor ( n8357 , n828 , n790 );
buf ( n175785 , n8357 );
nand ( n8359 , n175783 , n175785 );
buf ( n175787 , n8359 );
buf ( n175788 , n175787 );
nand ( n8362 , n8355 , n175788 );
buf ( n175790 , n8362 );
buf ( n175791 , n175790 );
not ( n8365 , n175791 );
buf ( n175793 , n799 );
buf ( n175794 , n821 );
or ( n8368 , n175793 , n175794 );
buf ( n175796 , n822 );
nand ( n8370 , n8368 , n175796 );
buf ( n175798 , n8370 );
buf ( n175799 , n175798 );
buf ( n175800 , n799 );
buf ( n175801 , n821 );
nand ( n8375 , n175800 , n175801 );
buf ( n175803 , n8375 );
buf ( n175804 , n175803 );
buf ( n175805 , n820 );
nand ( n8379 , n175799 , n175804 , n175805 );
buf ( n175807 , n8379 );
buf ( n175808 , n175807 );
nor ( n8382 , n8365 , n175808 );
buf ( n175810 , n8382 );
buf ( n175811 , n175810 );
xor ( n8385 , n175773 , n175811 );
buf ( n175813 , n789 );
buf ( n175814 , n830 );
xor ( n8388 , n175813 , n175814 );
buf ( n175816 , n8388 );
buf ( n175817 , n175816 );
not ( n8391 , n175817 );
buf ( n175819 , n168471 );
not ( n8393 , n175819 );
or ( n8394 , n8391 , n8393 );
buf ( n175822 , n788 );
buf ( n175823 , n830 );
xor ( n175824 , n175822 , n175823 );
buf ( n175825 , n175824 );
buf ( n175826 , n175825 );
buf ( n175827 , n831 );
nand ( n8401 , n175826 , n175827 );
buf ( n175829 , n8401 );
buf ( n175830 , n175829 );
nand ( n8404 , n8394 , n175830 );
buf ( n175832 , n8404 );
buf ( n175833 , n175832 );
buf ( n175834 , n795 );
buf ( n175835 , n824 );
xor ( n8409 , n175834 , n175835 );
buf ( n175837 , n8409 );
buf ( n175838 , n175837 );
not ( n8412 , n175838 );
buf ( n175840 , n170100 );
not ( n8414 , n175840 );
or ( n8415 , n8412 , n8414 );
buf ( n175843 , n175664 );
buf ( n175844 , n794 );
buf ( n175845 , n824 );
xor ( n175846 , n175844 , n175845 );
buf ( n175847 , n175846 );
buf ( n175848 , n175847 );
nand ( n8422 , n175843 , n175848 );
buf ( n175850 , n8422 );
buf ( n175851 , n175850 );
nand ( n8425 , n8415 , n175851 );
buf ( n175853 , n8425 );
buf ( n175854 , n175853 );
xor ( n8428 , n175833 , n175854 );
buf ( n175856 , n797 );
buf ( n175857 , n822 );
xor ( n8431 , n175856 , n175857 );
buf ( n175859 , n8431 );
buf ( n175860 , n175859 );
not ( n8434 , n175860 );
buf ( n175862 , n169411 );
not ( n8436 , n175862 );
or ( n8437 , n8434 , n8436 );
buf ( n175865 , n171055 );
buf ( n175866 , n796 );
buf ( n175867 , n822 );
xor ( n8441 , n175866 , n175867 );
buf ( n175869 , n8441 );
buf ( n175870 , n175869 );
nand ( n8444 , n175865 , n175870 );
buf ( n175872 , n8444 );
buf ( n175873 , n175872 );
nand ( n8447 , n8437 , n175873 );
buf ( n175875 , n8447 );
buf ( n175876 , n175875 );
and ( n8450 , n8428 , n175876 );
and ( n8451 , n175833 , n175854 );
or ( n8452 , n8450 , n8451 );
buf ( n175880 , n8452 );
buf ( n175881 , n175880 );
and ( n8455 , n8385 , n175881 );
and ( n8456 , n175773 , n175811 );
or ( n8457 , n8455 , n8456 );
buf ( n175885 , n8457 );
and ( n8459 , n8329 , n175885 );
and ( n8460 , n8326 , n8328 );
or ( n8461 , n8459 , n8460 );
buf ( n175889 , n8461 );
xor ( n8463 , n175750 , n175889 );
xor ( n8464 , n7955 , n7942 );
xor ( n8465 , n8464 , n175410 );
buf ( n175893 , n8465 );
buf ( n175894 , n175537 );
not ( n8468 , n175894 );
buf ( n175896 , n175563 );
nand ( n8470 , n8468 , n175896 );
buf ( n175898 , n8470 );
buf ( n175899 , n175898 );
buf ( n175900 , n175557 );
and ( n8474 , n175899 , n175900 );
not ( n8475 , n175899 );
buf ( n175903 , n175554 );
and ( n8477 , n8475 , n175903 );
nor ( n175905 , n8474 , n8477 );
buf ( n175906 , n175905 );
buf ( n175907 , n175906 );
xor ( n8484 , n175893 , n175907 );
buf ( n175909 , n175498 );
buf ( n175910 , n175517 );
and ( n175911 , n175909 , n175910 );
not ( n8488 , n175909 );
buf ( n175913 , n175514 );
and ( n8490 , n8488 , n175913 );
nor ( n8491 , n175911 , n8490 );
buf ( n175916 , n8491 );
buf ( n175917 , n175916 );
buf ( n175918 , n168806 );
buf ( n175919 , n799 );
and ( n8496 , n175918 , n175919 );
buf ( n175921 , n8496 );
buf ( n175922 , n175921 );
buf ( n175923 , n175847 );
not ( n8500 , n175923 );
buf ( n175925 , n170100 );
not ( n8502 , n175925 );
or ( n8503 , n8500 , n8502 );
buf ( n175928 , n169802 );
buf ( n175929 , n175656 );
nand ( n8506 , n175928 , n175929 );
buf ( n175931 , n8506 );
buf ( n175932 , n175931 );
nand ( n8509 , n8503 , n175932 );
buf ( n175934 , n8509 );
buf ( n175935 , n175934 );
xor ( n8512 , n175922 , n175935 );
buf ( n175937 , n8357 );
not ( n8514 , n175937 );
buf ( n175939 , n170990 );
not ( n8516 , n175939 );
or ( n8517 , n8514 , n8516 );
buf ( n175942 , n168559 );
buf ( n175943 , n8209 );
nand ( n8520 , n175942 , n175943 );
buf ( n175945 , n8520 );
buf ( n175946 , n175945 );
nand ( n8523 , n8517 , n175946 );
buf ( n175948 , n8523 );
buf ( n175949 , n175948 );
and ( n8526 , n8512 , n175949 );
and ( n8527 , n175922 , n175935 );
or ( n8528 , n8526 , n8527 );
buf ( n175953 , n8528 );
buf ( n175954 , n175953 );
xor ( n8531 , n175917 , n175954 );
buf ( n175956 , n175825 );
not ( n8533 , n175956 );
buf ( n175958 , n168471 );
not ( n8535 , n175958 );
or ( n8536 , n8533 , n8535 );
buf ( n175961 , n175486 );
buf ( n175962 , n831 );
nand ( n8539 , n175961 , n175962 );
buf ( n175964 , n8539 );
buf ( n175965 , n175964 );
nand ( n8542 , n8536 , n175965 );
buf ( n175967 , n8542 );
buf ( n175968 , n175967 );
buf ( n175969 , n798 );
buf ( n175970 , n820 );
xor ( n175971 , n175969 , n175970 );
buf ( n175972 , n175971 );
buf ( n175973 , n175972 );
not ( n8550 , n175973 );
buf ( n175975 , n2251 );
not ( n8552 , n175975 );
or ( n8553 , n8550 , n8552 );
buf ( n175978 , n2513 );
buf ( n175979 , n175591 );
nand ( n8556 , n175978 , n175979 );
buf ( n175981 , n8556 );
buf ( n175982 , n175981 );
nand ( n8559 , n8553 , n175982 );
buf ( n175984 , n8559 );
buf ( n175985 , n175984 );
xor ( n8562 , n175968 , n175985 );
buf ( n175987 , n175869 );
not ( n8564 , n175987 );
buf ( n175989 , n171049 );
not ( n8566 , n175989 );
or ( n8567 , n8564 , n8566 );
buf ( n175992 , n171055 );
buf ( n175993 , n175678 );
nand ( n8570 , n175992 , n175993 );
buf ( n175995 , n8570 );
buf ( n175996 , n175995 );
nand ( n8573 , n8567 , n175996 );
buf ( n175998 , n8573 );
buf ( n175999 , n175998 );
and ( n8576 , n8562 , n175999 );
and ( n176001 , n175968 , n175985 );
or ( n8578 , n8576 , n176001 );
buf ( n176003 , n8578 );
buf ( n176004 , n176003 );
and ( n8581 , n8531 , n176004 );
and ( n176006 , n175917 , n175954 );
or ( n8583 , n8581 , n176006 );
buf ( n176008 , n8583 );
buf ( n176009 , n176008 );
xor ( n8586 , n8484 , n176009 );
buf ( n176011 , n8586 );
buf ( n176012 , n176011 );
and ( n8589 , n8463 , n176012 );
and ( n8590 , n175750 , n175889 );
or ( n8591 , n8589 , n8590 );
buf ( n176016 , n8591 );
buf ( n176017 , n176016 );
xor ( n8594 , n175739 , n176017 );
xor ( n8595 , n175413 , n175416 );
xor ( n8596 , n8595 , n175430 );
buf ( n176021 , n8596 );
buf ( n176022 , n176021 );
xor ( n8599 , n175567 , n175571 );
xor ( n8600 , n8599 , n175697 );
buf ( n176025 , n8600 );
buf ( n176026 , n176025 );
xor ( n8603 , n176022 , n176026 );
xor ( n8604 , n175893 , n175907 );
and ( n8605 , n8604 , n176009 );
and ( n8606 , n175893 , n175907 );
or ( n8607 , n8605 , n8606 );
buf ( n176032 , n8607 );
buf ( n176033 , n176032 );
xor ( n8610 , n8603 , n176033 );
buf ( n176035 , n8610 );
buf ( n176036 , n176035 );
and ( n8613 , n8594 , n176036 );
and ( n8614 , n175739 , n176017 );
or ( n8615 , n8613 , n8614 );
buf ( n176040 , n8615 );
buf ( n176041 , n176040 );
buf ( n176042 , n847 );
xor ( n8619 , n176022 , n176026 );
and ( n8620 , n8619 , n176033 );
and ( n8621 , n176022 , n176026 );
or ( n8622 , n8620 , n8621 );
buf ( n176047 , n8622 );
buf ( n176048 , n176047 );
xor ( n8625 , n176042 , n176048 );
xor ( n8626 , n175482 , n175702 );
xor ( n8627 , n8626 , n175707 );
buf ( n176052 , n8627 );
buf ( n176053 , n176052 );
xor ( n8630 , n8625 , n176053 );
buf ( n176055 , n8630 );
buf ( n176056 , n176055 );
nand ( n8633 , n176041 , n176056 );
buf ( n176058 , n8633 );
buf ( n176059 , n176058 );
not ( n8636 , n176059 );
xor ( n8637 , n175478 , n175712 );
xor ( n8638 , n8637 , n175717 );
buf ( n176063 , n8638 );
buf ( n176064 , n176063 );
xor ( n8641 , n176042 , n176048 );
and ( n176066 , n8641 , n176053 );
and ( n8643 , n176042 , n176048 );
or ( n8644 , n176066 , n8643 );
buf ( n176069 , n8644 );
buf ( n176070 , n176069 );
nand ( n8647 , n176064 , n176070 );
buf ( n176072 , n8647 );
buf ( n176073 , n176072 );
not ( n8650 , n176073 );
or ( n8651 , n8636 , n8650 );
or ( n8652 , n176063 , n176069 );
buf ( n176077 , n8652 );
nand ( n8654 , n8651 , n176077 );
buf ( n176079 , n8654 );
buf ( n176080 , n176079 );
not ( n8657 , n176080 );
buf ( n176082 , n8657 );
not ( n8659 , n176082 );
or ( n8660 , n8308 , n8659 );
buf ( n176085 , n175736 );
not ( n8662 , n176085 );
buf ( n176087 , n8662 );
buf ( n176088 , n176087 );
buf ( n176089 , n175476 );
not ( n8666 , n176089 );
buf ( n176091 , n8666 );
buf ( n176092 , n176091 );
buf ( n176093 , n175721 );
not ( n8670 , n176093 );
buf ( n176095 , n8670 );
buf ( n176096 , n176095 );
nor ( n8676 , n176092 , n176096 );
buf ( n176098 , n8676 );
buf ( n176099 , n176098 );
and ( n8679 , n176088 , n176099 );
buf ( n176101 , n175733 );
buf ( n176102 , n175729 );
and ( n8682 , n176101 , n176102 );
buf ( n176104 , n8682 );
buf ( n176105 , n176104 );
nor ( n8685 , n8679 , n176105 );
buf ( n176107 , n8685 );
nand ( n8687 , n8660 , n176107 );
nand ( n8688 , n7831 , n8687 );
not ( n176110 , n174200 );
not ( n8690 , n174448 );
and ( n8691 , n176110 , n8690 );
buf ( n176113 , n174766 );
buf ( n176114 , n174454 );
nor ( n8694 , n176113 , n176114 );
buf ( n176116 , n8694 );
nor ( n8696 , n8691 , n176116 );
buf ( n176118 , n8696 );
not ( n8698 , n176118 );
buf ( n176120 , n175037 );
buf ( n176121 , n175266 );
and ( n8701 , n176120 , n176121 );
buf ( n176123 , n8701 );
buf ( n176124 , n176123 );
not ( n8704 , n176124 );
not ( n8705 , n175031 );
buf ( n176127 , n174773 );
not ( n8707 , n176127 );
buf ( n176129 , n8707 );
nand ( n8709 , n8705 , n176129 );
buf ( n176131 , n8709 );
not ( n8711 , n176131 );
or ( n8712 , n8704 , n8711 );
not ( n8713 , n176129 );
nand ( n8714 , n8713 , n175031 );
buf ( n176136 , n8714 );
nand ( n8716 , n8712 , n176136 );
buf ( n176138 , n8716 );
buf ( n176139 , n176138 );
not ( n8719 , n176139 );
or ( n8720 , n8698 , n8719 );
buf ( n176142 , n174451 );
not ( n8722 , n176142 );
buf ( n176144 , n8722 );
buf ( n176145 , n176144 );
buf ( n176146 , n174454 );
buf ( n176147 , n174766 );
nand ( n8727 , n176146 , n176147 );
buf ( n176149 , n8727 );
buf ( n176150 , n176149 );
not ( n8730 , n176150 );
buf ( n176152 , n8730 );
buf ( n176153 , n176152 );
and ( n8733 , n176145 , n176153 );
buf ( n176155 , n174448 );
buf ( n176156 , n174200 );
and ( n8736 , n176155 , n176156 );
buf ( n176158 , n8736 );
buf ( n176159 , n176158 );
nor ( n8739 , n8733 , n176159 );
buf ( n176161 , n8739 );
buf ( n176162 , n176161 );
nand ( n8742 , n8720 , n176162 );
buf ( n176164 , n8742 );
nor ( n8744 , n6725 , n176164 );
nand ( n8745 , n6195 , n8688 , n8744 );
buf ( n176167 , n8745 );
buf ( n176168 , n173506 );
buf ( n176169 , n173633 );
nor ( n8749 , n176168 , n176169 );
buf ( n176171 , n8749 );
nor ( n8751 , n6180 , n176171 );
buf ( n176173 , n8751 );
buf ( n8753 , n176173 );
buf ( n176175 , n8753 );
not ( n8755 , n176175 );
nand ( n8756 , n8755 , n6195 );
buf ( n176178 , n8756 );
nand ( n8758 , n5730 , n174197 , n176167 , n176178 );
buf ( n176180 , n8758 );
buf ( n176181 , n176180 );
buf ( n176182 , n176091 );
buf ( n176183 , n176095 );
nand ( n8763 , n176182 , n176183 );
buf ( n176185 , n8763 );
buf ( n176186 , n176185 );
not ( n8766 , n176063 );
not ( n176188 , n176069 );
and ( n8768 , n8766 , n176188 );
buf ( n176190 , n176040 );
buf ( n176191 , n176055 );
nor ( n8771 , n176190 , n176191 );
buf ( n176193 , n8771 );
nor ( n8773 , n8768 , n176193 );
buf ( n176195 , n8773 );
buf ( n176196 , n176087 );
and ( n8776 , n176186 , n176195 , n176196 );
buf ( n176198 , n8776 );
buf ( n176199 , n176198 );
not ( n8779 , n176199 );
buf ( n176201 , n8779 );
buf ( n176202 , n176201 );
not ( n8782 , n176202 );
buf ( n176204 , n8782 );
not ( n8784 , n7830 );
and ( n8785 , n173194 , n176204 , n174170 , n8784 );
buf ( n176207 , n8785 );
buf ( n176208 , n5018 );
buf ( n176209 , n176175 );
xor ( n8789 , n175739 , n176017 );
xor ( n176211 , n8789 , n176036 );
buf ( n176212 , n176211 );
buf ( n176213 , n176212 );
buf ( n176214 , n849 );
xor ( n8794 , n175917 , n175954 );
xor ( n8795 , n8794 , n176004 );
buf ( n176217 , n8795 );
buf ( n176218 , n176217 );
xor ( n8798 , n175922 , n175935 );
xor ( n8799 , n8798 , n175949 );
buf ( n176221 , n8799 );
buf ( n176222 , n176221 );
xor ( n8802 , n175968 , n175985 );
xor ( n8803 , n8802 , n175999 );
buf ( n176225 , n8803 );
buf ( n176226 , n176225 );
xor ( n8806 , n176222 , n176226 );
buf ( n176228 , n799 );
buf ( n176229 , n820 );
xor ( n8809 , n176228 , n176229 );
buf ( n176231 , n8809 );
buf ( n176232 , n176231 );
not ( n8812 , n176232 );
buf ( n176234 , n2251 );
not ( n8814 , n176234 );
or ( n8815 , n8812 , n8814 );
buf ( n176237 , n2513 );
buf ( n176238 , n175972 );
nand ( n8818 , n176237 , n176238 );
buf ( n176240 , n8818 );
buf ( n176241 , n176240 );
nand ( n8821 , n8815 , n176241 );
buf ( n176243 , n8821 );
buf ( n176244 , n176243 );
xor ( n8824 , n826 , n793 );
buf ( n176246 , n8824 );
not ( n8826 , n176246 );
buf ( n176248 , n175400 );
not ( n8828 , n176248 );
or ( n8829 , n8826 , n8828 );
buf ( n176251 , n169081 );
buf ( n176252 , n175760 );
nand ( n8832 , n176251 , n176252 );
buf ( n176254 , n8832 );
buf ( n176255 , n176254 );
nand ( n8835 , n8829 , n176255 );
buf ( n176257 , n8835 );
buf ( n176258 , n176257 );
xor ( n8838 , n176244 , n176258 );
buf ( n176260 , n175807 );
not ( n8840 , n176260 );
buf ( n176262 , n175790 );
not ( n8842 , n176262 );
or ( n8843 , n8840 , n8842 );
buf ( n176265 , n175790 );
buf ( n176266 , n175807 );
or ( n8846 , n176265 , n176266 );
nand ( n8847 , n8843 , n8846 );
buf ( n176269 , n8847 );
buf ( n176270 , n176269 );
and ( n8850 , n8838 , n176270 );
and ( n8851 , n176244 , n176258 );
or ( n8852 , n8850 , n8851 );
buf ( n176274 , n8852 );
buf ( n176275 , n176274 );
and ( n8855 , n8806 , n176275 );
and ( n8856 , n176222 , n176226 );
or ( n8857 , n8855 , n8856 );
buf ( n176279 , n8857 );
buf ( n176280 , n176279 );
xor ( n8863 , n176218 , n176280 );
xor ( n8864 , n8326 , n8328 );
xor ( n8865 , n8864 , n175885 );
buf ( n176284 , n8865 );
and ( n176285 , n8863 , n176284 );
and ( n8868 , n176218 , n176280 );
or ( n8869 , n176285 , n8868 );
buf ( n176288 , n8869 );
buf ( n176289 , n176288 );
xor ( n8872 , n176214 , n176289 );
xor ( n8873 , n175750 , n175889 );
xor ( n8874 , n8873 , n176012 );
buf ( n176293 , n8874 );
buf ( n176294 , n176293 );
and ( n8877 , n8872 , n176294 );
and ( n8878 , n176214 , n176289 );
or ( n8879 , n8877 , n8878 );
buf ( n176298 , n8879 );
buf ( n176299 , n176298 );
nor ( n8882 , n176213 , n176299 );
buf ( n176301 , n8882 );
buf ( n176302 , n176301 );
xor ( n8885 , n176214 , n176289 );
xor ( n8886 , n8885 , n176294 );
buf ( n176305 , n8886 );
buf ( n176306 , n176305 );
buf ( n176307 , n850 );
xor ( n8890 , n175773 , n175811 );
xor ( n8891 , n8890 , n175881 );
buf ( n176310 , n8891 );
buf ( n176311 , n176310 );
buf ( n176312 , n168656 );
buf ( n176313 , n799 );
and ( n8896 , n176312 , n176313 );
buf ( n176315 , n8896 );
buf ( n176316 , n176315 );
buf ( n176317 , n792 );
buf ( n176318 , n828 );
xor ( n8901 , n176317 , n176318 );
buf ( n176320 , n8901 );
buf ( n176321 , n176320 );
not ( n8904 , n176321 );
buf ( n176323 , n170990 );
not ( n8906 , n176323 );
or ( n8907 , n8904 , n8906 );
buf ( n176326 , n168559 );
buf ( n176327 , n175777 );
nand ( n8910 , n176326 , n176327 );
buf ( n176329 , n8910 );
buf ( n176330 , n176329 );
nand ( n8913 , n8907 , n176330 );
buf ( n176332 , n8913 );
buf ( n176333 , n176332 );
xor ( n8916 , n176316 , n176333 );
buf ( n176335 , n796 );
buf ( n176336 , n824 );
xor ( n8919 , n176335 , n176336 );
buf ( n176338 , n8919 );
buf ( n176339 , n176338 );
not ( n8922 , n176339 );
buf ( n176341 , n170100 );
not ( n8924 , n176341 );
or ( n8925 , n8922 , n8924 );
buf ( n176344 , n175664 );
buf ( n176345 , n175837 );
nand ( n8928 , n176344 , n176345 );
buf ( n176347 , n8928 );
buf ( n176348 , n176347 );
nand ( n8931 , n8925 , n176348 );
buf ( n176350 , n8931 );
buf ( n176351 , n176350 );
and ( n8934 , n8916 , n176351 );
and ( n8935 , n176316 , n176333 );
or ( n8936 , n8934 , n8935 );
buf ( n176355 , n8936 );
buf ( n176356 , n176355 );
buf ( n176357 , n790 );
buf ( n176358 , n830 );
xor ( n8941 , n176357 , n176358 );
buf ( n176360 , n8941 );
buf ( n176361 , n176360 );
not ( n8944 , n176361 );
buf ( n176363 , n168471 );
not ( n8946 , n176363 );
or ( n8947 , n8944 , n8946 );
buf ( n176366 , n175816 );
buf ( n176367 , n831 );
nand ( n8950 , n176366 , n176367 );
buf ( n176369 , n8950 );
buf ( n176370 , n176369 );
nand ( n8953 , n8947 , n176370 );
buf ( n176372 , n8953 );
buf ( n176373 , n176372 );
buf ( n176374 , n798 );
buf ( n176375 , n822 );
xor ( n8958 , n176374 , n176375 );
buf ( n176377 , n8958 );
buf ( n176378 , n176377 );
not ( n8961 , n176378 );
buf ( n176380 , n171049 );
not ( n8963 , n176380 );
or ( n8964 , n8961 , n8963 );
buf ( n176383 , n171055 );
buf ( n176384 , n175859 );
nand ( n176385 , n176383 , n176384 );
buf ( n176386 , n176385 );
buf ( n176387 , n176386 );
nand ( n8970 , n8964 , n176387 );
buf ( n176389 , n8970 );
buf ( n176390 , n176389 );
xor ( n8973 , n176373 , n176390 );
buf ( n176392 , n8824 );
not ( n8975 , n176392 );
buf ( n176394 , n169081 );
not ( n8977 , n176394 );
or ( n8978 , n8975 , n8977 );
buf ( n176397 , n169093 );
buf ( n176398 , n794 );
buf ( n176399 , n826 );
xor ( n8982 , n176398 , n176399 );
buf ( n176401 , n8982 );
buf ( n176402 , n176401 );
not ( n8985 , n176402 );
buf ( n176404 , n8985 );
buf ( n176405 , n176404 );
or ( n176406 , n176397 , n176405 );
nand ( n8989 , n8978 , n176406 );
buf ( n176408 , n8989 );
buf ( n176409 , n176408 );
and ( n8992 , n8973 , n176409 );
and ( n8993 , n176373 , n176390 );
or ( n8994 , n8992 , n8993 );
buf ( n176413 , n8994 );
buf ( n176414 , n176413 );
xor ( n8997 , n176356 , n176414 );
xor ( n8998 , n175833 , n175854 );
xor ( n8999 , n8998 , n175876 );
buf ( n176418 , n8999 );
buf ( n176419 , n176418 );
and ( n9002 , n8997 , n176419 );
and ( n9003 , n176356 , n176414 );
or ( n9004 , n9002 , n9003 );
buf ( n176423 , n9004 );
buf ( n176424 , n176423 );
xor ( n9007 , n176311 , n176424 );
xor ( n9008 , n176222 , n176226 );
xor ( n9009 , n9008 , n176275 );
buf ( n176428 , n9009 );
buf ( n176429 , n176428 );
and ( n9012 , n9007 , n176429 );
and ( n9013 , n176311 , n176424 );
or ( n9014 , n9012 , n9013 );
buf ( n176433 , n9014 );
buf ( n176434 , n176433 );
xor ( n176435 , n176307 , n176434 );
xor ( n9018 , n176218 , n176280 );
xor ( n9019 , n9018 , n176284 );
buf ( n176438 , n9019 );
buf ( n176439 , n176438 );
and ( n9022 , n176435 , n176439 );
and ( n9023 , n176307 , n176434 );
or ( n9024 , n9022 , n9023 );
buf ( n176443 , n9024 );
buf ( n176444 , n176443 );
nor ( n9027 , n176306 , n176444 );
buf ( n176446 , n9027 );
buf ( n176447 , n176446 );
nor ( n9030 , n176302 , n176447 );
buf ( n176449 , n9030 );
buf ( n176450 , n176449 );
xor ( n9033 , n176307 , n176434 );
xor ( n9034 , n9033 , n176439 );
buf ( n176453 , n9034 );
not ( n9036 , n176453 );
buf ( n176455 , n851 );
xor ( n9038 , n176244 , n176258 );
xor ( n9039 , n9038 , n176270 );
buf ( n176458 , n9039 );
buf ( n176459 , n176458 );
buf ( n176460 , n793 );
buf ( n176461 , n828 );
xor ( n9044 , n176460 , n176461 );
buf ( n176463 , n9044 );
buf ( n176464 , n176463 );
not ( n9047 , n176464 );
buf ( n176466 , n170990 );
not ( n9049 , n176466 );
or ( n9050 , n9047 , n9049 );
buf ( n176469 , n168559 );
buf ( n176470 , n176320 );
nand ( n9053 , n176469 , n176470 );
buf ( n176472 , n9053 );
buf ( n176473 , n176472 );
nand ( n9056 , n9050 , n176473 );
buf ( n176475 , n9056 );
buf ( n176476 , n176475 );
not ( n9059 , n176476 );
buf ( n176478 , n799 );
buf ( n176479 , n823 );
or ( n9062 , n176478 , n176479 );
buf ( n176481 , n824 );
nand ( n9064 , n9062 , n176481 );
buf ( n176483 , n9064 );
buf ( n176484 , n176483 );
buf ( n176485 , n799 );
buf ( n176486 , n823 );
nand ( n9069 , n176485 , n176486 );
buf ( n176488 , n9069 );
buf ( n176489 , n176488 );
buf ( n176490 , n822 );
nand ( n9076 , n176484 , n176489 , n176490 );
buf ( n176492 , n9076 );
buf ( n176493 , n176492 );
nor ( n9079 , n9059 , n176493 );
buf ( n176495 , n9079 );
buf ( n176496 , n176495 );
xor ( n9082 , n176316 , n176333 );
xor ( n9083 , n9082 , n176351 );
buf ( n176499 , n9083 );
buf ( n176500 , n176499 );
xor ( n9086 , n176496 , n176500 );
buf ( n176502 , n791 );
buf ( n176503 , n830 );
xor ( n9089 , n176502 , n176503 );
buf ( n176505 , n9089 );
buf ( n176506 , n176505 );
not ( n9092 , n176506 );
buf ( n176508 , n168471 );
not ( n9094 , n176508 );
or ( n9095 , n9092 , n9094 );
buf ( n176511 , n176360 );
buf ( n176512 , n831 );
nand ( n9098 , n176511 , n176512 );
buf ( n176514 , n9098 );
buf ( n176515 , n176514 );
nand ( n9101 , n9095 , n176515 );
buf ( n176517 , n9101 );
xor ( n9103 , n824 , n797 );
buf ( n176519 , n9103 );
not ( n9105 , n176519 );
buf ( n176521 , n170100 );
not ( n9107 , n176521 );
or ( n9108 , n9105 , n9107 );
buf ( n176524 , n169169 );
buf ( n176525 , n176338 );
nand ( n9111 , n176524 , n176525 );
buf ( n176527 , n9111 );
buf ( n176528 , n176527 );
nand ( n9114 , n9108 , n176528 );
buf ( n176530 , n9114 );
xor ( n9116 , n176517 , n176530 );
xor ( n9117 , n822 , n799 );
not ( n9118 , n9117 );
not ( n9119 , n171049 );
or ( n9120 , n9118 , n9119 );
buf ( n176536 , n171055 );
buf ( n176537 , n176377 );
nand ( n9123 , n176536 , n176537 );
buf ( n176539 , n9123 );
nand ( n9125 , n9120 , n176539 );
and ( n9126 , n9116 , n9125 );
and ( n9127 , n176517 , n176530 );
or ( n9128 , n9126 , n9127 );
buf ( n176544 , n9128 );
and ( n9130 , n9086 , n176544 );
and ( n9131 , n176496 , n176500 );
or ( n9132 , n9130 , n9131 );
buf ( n176548 , n9132 );
buf ( n176549 , n176548 );
xor ( n9135 , n176459 , n176549 );
xor ( n9136 , n176356 , n176414 );
xor ( n9137 , n9136 , n176419 );
buf ( n176553 , n9137 );
buf ( n176554 , n176553 );
and ( n9140 , n9135 , n176554 );
and ( n9141 , n176459 , n176549 );
or ( n9142 , n9140 , n9141 );
buf ( n176558 , n9142 );
buf ( n176559 , n176558 );
xor ( n9145 , n176455 , n176559 );
xor ( n9146 , n176311 , n176424 );
xor ( n9147 , n9146 , n176429 );
buf ( n176563 , n9147 );
buf ( n176564 , n176563 );
and ( n9150 , n9145 , n176564 );
and ( n9151 , n176455 , n176559 );
or ( n9152 , n9150 , n9151 );
buf ( n176568 , n9152 );
not ( n9154 , n176568 );
and ( n9155 , n9036 , n9154 );
xor ( n9156 , n176455 , n176559 );
xor ( n9157 , n9156 , n176564 );
buf ( n176573 , n9157 );
buf ( n176574 , n176573 );
buf ( n176575 , n852 );
xor ( n9161 , n176373 , n176390 );
xor ( n9162 , n9161 , n176409 );
buf ( n176578 , n9162 );
buf ( n176579 , n176578 );
buf ( n176580 , n795 );
buf ( n176581 , n826 );
xor ( n9167 , n176580 , n176581 );
buf ( n176583 , n9167 );
buf ( n176584 , n176583 );
not ( n9170 , n176584 );
buf ( n176586 , n175400 );
not ( n9172 , n176586 );
or ( n9173 , n9170 , n9172 );
buf ( n176589 , n169081 );
buf ( n176590 , n176401 );
nand ( n9176 , n176589 , n176590 );
buf ( n176592 , n9176 );
buf ( n176593 , n176592 );
nand ( n9179 , n9173 , n176593 );
buf ( n176595 , n9179 );
buf ( n176596 , n176595 );
buf ( n176597 , n169417 );
buf ( n176598 , n799 );
and ( n9184 , n176597 , n176598 );
buf ( n176600 , n9184 );
buf ( n176601 , n176600 );
buf ( n176602 , n792 );
buf ( n176603 , n830 );
xor ( n9189 , n176602 , n176603 );
buf ( n176605 , n9189 );
buf ( n176606 , n176605 );
not ( n9192 , n176606 );
buf ( n176608 , n168471 );
not ( n9194 , n176608 );
or ( n9195 , n9192 , n9194 );
buf ( n176611 , n176505 );
buf ( n176612 , n831 );
nand ( n9198 , n176611 , n176612 );
buf ( n176614 , n9198 );
buf ( n176615 , n176614 );
nand ( n9201 , n9195 , n176615 );
buf ( n176617 , n9201 );
buf ( n176618 , n176617 );
xor ( n9204 , n176601 , n176618 );
xor ( n9205 , n824 , n798 );
buf ( n176621 , n9205 );
not ( n9207 , n176621 );
buf ( n176623 , n170100 );
not ( n9209 , n176623 );
or ( n9210 , n9207 , n9209 );
buf ( n176626 , n175664 );
buf ( n176627 , n9103 );
nand ( n9213 , n176626 , n176627 );
buf ( n176629 , n9213 );
buf ( n176630 , n176629 );
nand ( n9216 , n9210 , n176630 );
buf ( n176632 , n9216 );
buf ( n176633 , n176632 );
and ( n9219 , n9204 , n176633 );
and ( n9220 , n176601 , n176618 );
or ( n9221 , n9219 , n9220 );
buf ( n176637 , n9221 );
buf ( n176638 , n176637 );
xor ( n9224 , n176596 , n176638 );
buf ( n176640 , n176492 );
not ( n9226 , n176640 );
buf ( n176642 , n176475 );
not ( n9228 , n176642 );
or ( n9229 , n9226 , n9228 );
buf ( n176645 , n176475 );
buf ( n176646 , n176492 );
or ( n9232 , n176645 , n176646 );
nand ( n9233 , n9229 , n9232 );
buf ( n176649 , n9233 );
buf ( n176650 , n176649 );
and ( n9236 , n9224 , n176650 );
and ( n9237 , n176596 , n176638 );
or ( n9238 , n9236 , n9237 );
buf ( n176654 , n9238 );
buf ( n176655 , n176654 );
xor ( n9241 , n176579 , n176655 );
xor ( n9242 , n176496 , n176500 );
xor ( n9243 , n9242 , n176544 );
buf ( n176659 , n9243 );
buf ( n176660 , n176659 );
and ( n9246 , n9241 , n176660 );
and ( n9247 , n176579 , n176655 );
or ( n9248 , n9246 , n9247 );
buf ( n176664 , n9248 );
buf ( n176665 , n176664 );
xor ( n9251 , n176575 , n176665 );
xor ( n9252 , n176459 , n176549 );
xor ( n9253 , n9252 , n176554 );
buf ( n176669 , n9253 );
buf ( n176670 , n176669 );
and ( n9256 , n9251 , n176670 );
and ( n9257 , n176575 , n176665 );
or ( n9258 , n9256 , n9257 );
buf ( n176674 , n9258 );
buf ( n176675 , n176674 );
nor ( n9261 , n176574 , n176675 );
buf ( n176677 , n9261 );
nor ( n9263 , n9155 , n176677 );
buf ( n176679 , n9263 );
and ( n9265 , n176450 , n176679 );
buf ( n176681 , n9265 );
buf ( n176682 , n176681 );
not ( n9268 , n176682 );
xor ( n9269 , n176575 , n176665 );
xor ( n9270 , n9269 , n176670 );
buf ( n176686 , n9270 );
buf ( n176687 , n176686 );
not ( n9273 , n176687 );
buf ( n176689 , n9273 );
buf ( n176690 , n176689 );
buf ( n176691 , n793 );
buf ( n176692 , n830 );
xor ( n176693 , n176691 , n176692 );
buf ( n176694 , n176693 );
buf ( n176695 , n176694 );
not ( n9284 , n176695 );
buf ( n176697 , n168471 );
not ( n9286 , n176697 );
or ( n176699 , n9284 , n9286 );
buf ( n176700 , n176605 );
buf ( n176701 , n831 );
nand ( n9290 , n176700 , n176701 );
buf ( n176703 , n9290 );
buf ( n176704 , n176703 );
nand ( n9293 , n176699 , n176704 );
buf ( n176706 , n9293 );
buf ( n176707 , n176706 );
buf ( n176708 , n799 );
buf ( n176709 , n825 );
or ( n9298 , n176708 , n176709 );
buf ( n176711 , n826 );
nand ( n9300 , n9298 , n176711 );
buf ( n176713 , n9300 );
buf ( n176714 , n176713 );
buf ( n176715 , n799 );
buf ( n176716 , n825 );
nand ( n9305 , n176715 , n176716 );
buf ( n176718 , n9305 );
buf ( n176719 , n176718 );
buf ( n176720 , n824 );
nand ( n9309 , n176714 , n176719 , n176720 );
buf ( n176722 , n9309 );
buf ( n176723 , n176722 );
not ( n9312 , n176723 );
buf ( n176725 , n9312 );
buf ( n176726 , n176725 );
nand ( n9315 , n176707 , n176726 );
buf ( n176728 , n9315 );
buf ( n176729 , n176728 );
not ( n9318 , n176729 );
buf ( n176731 , n796 );
buf ( n176732 , n826 );
xor ( n9321 , n176731 , n176732 );
buf ( n176734 , n9321 );
buf ( n176735 , n176734 );
not ( n9324 , n176735 );
buf ( n176737 , n1621 );
not ( n9326 , n176737 );
or ( n9327 , n9324 , n9326 );
buf ( n176740 , n169081 );
buf ( n176741 , n176583 );
nand ( n9330 , n176740 , n176741 );
buf ( n176743 , n9330 );
buf ( n176744 , n176743 );
nand ( n9333 , n9327 , n176744 );
buf ( n176746 , n9333 );
buf ( n176747 , n176746 );
not ( n9336 , n176747 );
buf ( n176749 , n9336 );
buf ( n176750 , n176749 );
not ( n9339 , n176750 );
or ( n9340 , n9318 , n9339 );
buf ( n176753 , n794 );
buf ( n176754 , n828 );
xor ( n9343 , n176753 , n176754 );
buf ( n176756 , n9343 );
buf ( n176757 , n176756 );
not ( n9346 , n176757 );
buf ( n176759 , n170990 );
not ( n9348 , n176759 );
or ( n9349 , n9346 , n9348 );
buf ( n176762 , n168559 );
not ( n9351 , n176762 );
buf ( n176764 , n9351 );
buf ( n176765 , n176764 );
not ( n9354 , n176765 );
buf ( n176767 , n9354 );
buf ( n176768 , n176767 );
buf ( n176769 , n176463 );
nand ( n9358 , n176768 , n176769 );
buf ( n176771 , n9358 );
buf ( n176772 , n176771 );
nand ( n9361 , n9349 , n176772 );
buf ( n176774 , n9361 );
buf ( n176775 , n176774 );
nand ( n9364 , n9340 , n176775 );
buf ( n176777 , n9364 );
buf ( n176778 , n176777 );
buf ( n176779 , n176728 );
not ( n9368 , n176779 );
buf ( n176781 , n176746 );
nand ( n9370 , n9368 , n176781 );
buf ( n176783 , n9370 );
buf ( n176784 , n176783 );
nand ( n9373 , n176778 , n176784 );
buf ( n176786 , n9373 );
buf ( n176787 , n176786 );
xor ( n9376 , n176517 , n176530 );
xor ( n9377 , n9376 , n9125 );
buf ( n176790 , n9377 );
xor ( n9379 , n176787 , n176790 );
xor ( n9380 , n176596 , n176638 );
xor ( n9381 , n9380 , n176650 );
buf ( n176794 , n9381 );
buf ( n176795 , n176794 );
and ( n9384 , n9379 , n176795 );
and ( n9385 , n176787 , n176790 );
or ( n9386 , n9384 , n9385 );
buf ( n176799 , n9386 );
buf ( n176800 , n176799 );
buf ( n9389 , n176800 );
buf ( n176802 , n9389 );
buf ( n176803 , n176802 );
not ( n9392 , n176803 );
xor ( n9393 , n176579 , n176655 );
xor ( n9394 , n9393 , n176660 );
buf ( n176807 , n9394 );
buf ( n9396 , n176807 );
buf ( n176809 , n9396 );
not ( n9398 , n176809 );
or ( n9399 , n9392 , n9398 );
buf ( n176812 , n9396 );
buf ( n176813 , n176802 );
or ( n176814 , n176812 , n176813 );
buf ( n176815 , n853 );
nand ( n9404 , n176814 , n176815 );
buf ( n176817 , n9404 );
buf ( n176818 , n176817 );
nand ( n9407 , n9399 , n176818 );
buf ( n176820 , n9407 );
buf ( n176821 , n176820 );
not ( n9410 , n176821 );
buf ( n176823 , n9410 );
buf ( n176824 , n176823 );
nand ( n9413 , n176690 , n176824 );
buf ( n176826 , n9413 );
buf ( n176827 , n176799 );
not ( n9416 , n176827 );
buf ( n176829 , n9416 );
and ( n9418 , n853 , n176829 );
not ( n9419 , n853 );
and ( n9420 , n9419 , n176799 );
or ( n9421 , n9418 , n9420 );
buf ( n176834 , n9421 );
buf ( n176835 , n9396 );
and ( n9424 , n176834 , n176835 );
not ( n9425 , n176834 );
buf ( n176838 , n9396 );
not ( n9427 , n176838 );
buf ( n176840 , n9427 );
buf ( n176841 , n176840 );
and ( n9430 , n9425 , n176841 );
nor ( n9431 , n9424 , n9430 );
buf ( n176844 , n9431 );
buf ( n176845 , n176844 );
not ( n9434 , n176845 );
buf ( n176847 , n9434 );
buf ( n176848 , n176847 );
buf ( n176849 , n854 );
xor ( n9438 , n176601 , n176618 );
xor ( n9439 , n9438 , n176633 );
buf ( n176852 , n9439 );
buf ( n176853 , n176852 );
buf ( n176854 , n797 );
buf ( n176855 , n826 );
xor ( n9444 , n176854 , n176855 );
buf ( n176857 , n9444 );
buf ( n176858 , n176857 );
not ( n9447 , n176858 );
buf ( n176860 , n1621 );
not ( n9449 , n176860 );
or ( n9450 , n9447 , n9449 );
buf ( n176863 , n169081 );
buf ( n176864 , n176734 );
nand ( n9453 , n176863 , n176864 );
buf ( n176866 , n9453 );
buf ( n176867 , n176866 );
nand ( n9456 , n9450 , n176867 );
buf ( n176869 , n9456 );
buf ( n176870 , n176869 );
xor ( n9459 , n824 , n799 );
buf ( n176872 , n9459 );
not ( n9461 , n176872 );
buf ( n176874 , n170100 );
not ( n9463 , n176874 );
or ( n9464 , n9461 , n9463 );
buf ( n176877 , n169802 );
buf ( n176878 , n9205 );
nand ( n9467 , n176877 , n176878 );
buf ( n176880 , n9467 );
buf ( n176881 , n176880 );
nand ( n9470 , n9464 , n176881 );
buf ( n176883 , n9470 );
buf ( n176884 , n176883 );
or ( n9473 , n176870 , n176884 );
buf ( n176886 , n795 );
buf ( n176887 , n828 );
xor ( n9476 , n176886 , n176887 );
buf ( n176889 , n9476 );
buf ( n176890 , n176889 );
not ( n9479 , n176890 );
buf ( n176892 , n170990 );
not ( n9481 , n176892 );
or ( n9482 , n9479 , n9481 );
buf ( n176895 , n176767 );
buf ( n176896 , n176756 );
nand ( n9485 , n176895 , n176896 );
buf ( n176898 , n9485 );
buf ( n176899 , n176898 );
nand ( n9488 , n9482 , n176899 );
buf ( n176901 , n9488 );
buf ( n176902 , n176901 );
nand ( n9491 , n9473 , n176902 );
buf ( n176904 , n9491 );
buf ( n176905 , n176904 );
buf ( n176906 , n176869 );
buf ( n176907 , n176883 );
nand ( n9496 , n176906 , n176907 );
buf ( n176909 , n9496 );
buf ( n176910 , n176909 );
nand ( n9499 , n176905 , n176910 );
buf ( n176912 , n9499 );
buf ( n176913 , n176912 );
xor ( n9502 , n176853 , n176913 );
xor ( n9503 , n176728 , n176746 );
buf ( n176916 , n9503 );
buf ( n176917 , n176774 );
xnor ( n9506 , n176916 , n176917 );
buf ( n176919 , n9506 );
buf ( n176920 , n176919 );
and ( n9509 , n9502 , n176920 );
and ( n9510 , n176853 , n176913 );
or ( n9511 , n9509 , n9510 );
buf ( n176924 , n9511 );
buf ( n176925 , n176924 );
xor ( n9517 , n176849 , n176925 );
xor ( n9518 , n176787 , n176790 );
xor ( n9519 , n9518 , n176795 );
buf ( n176929 , n9519 );
buf ( n176930 , n176929 );
and ( n9522 , n9517 , n176930 );
and ( n9523 , n176849 , n176925 );
or ( n9524 , n9522 , n9523 );
buf ( n176934 , n9524 );
buf ( n176935 , n176934 );
not ( n9527 , n176935 );
buf ( n176937 , n9527 );
buf ( n176938 , n176937 );
nand ( n9530 , n176848 , n176938 );
buf ( n176940 , n9530 );
buf ( n176941 , n855 );
buf ( n176942 , n176706 );
buf ( n176943 , n176725 );
and ( n9535 , n176942 , n176943 );
not ( n9536 , n176942 );
buf ( n176946 , n176722 );
and ( n9538 , n9536 , n176946 );
nor ( n9539 , n9535 , n9538 );
buf ( n176949 , n9539 );
buf ( n176950 , n176949 );
not ( n9542 , n176950 );
buf ( n176952 , n9542 );
buf ( n176953 , n175664 );
buf ( n176954 , n799 );
nand ( n9546 , n176953 , n176954 );
buf ( n176956 , n9546 );
buf ( n176957 , n176956 );
not ( n9549 , n176957 );
buf ( n176959 , n9549 );
buf ( n176960 , n176959 );
not ( n9552 , n176960 );
buf ( n176962 , n794 );
buf ( n176963 , n830 );
xor ( n9555 , n176962 , n176963 );
buf ( n176965 , n9555 );
buf ( n176966 , n176965 );
not ( n176967 , n176966 );
buf ( n176968 , n168471 );
not ( n9560 , n176968 );
or ( n9561 , n176967 , n9560 );
buf ( n176971 , n176694 );
buf ( n176972 , n831 );
nand ( n9564 , n176971 , n176972 );
buf ( n176974 , n9564 );
buf ( n176975 , n176974 );
nand ( n9567 , n9561 , n176975 );
buf ( n176977 , n9567 );
buf ( n176978 , n176977 );
not ( n9570 , n176978 );
or ( n9571 , n9552 , n9570 );
buf ( n176981 , n176956 );
not ( n9573 , n176981 );
buf ( n176983 , n176977 );
not ( n9575 , n176983 );
buf ( n176985 , n9575 );
buf ( n176986 , n176985 );
not ( n9578 , n176986 );
or ( n9579 , n9573 , n9578 );
buf ( n176989 , n796 );
buf ( n176990 , n828 );
xor ( n9582 , n176989 , n176990 );
buf ( n176992 , n9582 );
buf ( n176993 , n176992 );
not ( n9585 , n176993 );
buf ( n176995 , n170990 );
not ( n9587 , n176995 );
or ( n9588 , n9585 , n9587 );
buf ( n176998 , n176889 );
buf ( n176999 , n168559 );
nand ( n9591 , n176998 , n176999 );
buf ( n177001 , n9591 );
buf ( n177002 , n177001 );
nand ( n9594 , n9588 , n177002 );
buf ( n177004 , n9594 );
buf ( n177005 , n177004 );
nand ( n9597 , n9579 , n177005 );
buf ( n177007 , n9597 );
buf ( n177008 , n177007 );
nand ( n9600 , n9571 , n177008 );
buf ( n177010 , n9600 );
not ( n9602 , n177010 );
and ( n9603 , n176952 , n9602 );
not ( n9604 , n9603 );
buf ( n177014 , n9604 );
not ( n9606 , n177014 );
xor ( n9607 , n176869 , n176883 );
xnor ( n9608 , n9607 , n176901 );
buf ( n177018 , n9608 );
not ( n9610 , n177018 );
buf ( n177020 , n9610 );
buf ( n177021 , n177020 );
not ( n9613 , n177021 );
or ( n9614 , n9606 , n9613 );
buf ( n177024 , n177010 );
buf ( n177025 , n176949 );
nand ( n9617 , n177024 , n177025 );
buf ( n177027 , n9617 );
buf ( n177028 , n177027 );
nand ( n9620 , n9614 , n177028 );
buf ( n177030 , n9620 );
buf ( n177031 , n177030 );
xor ( n9623 , n176941 , n177031 );
xor ( n9624 , n176853 , n176913 );
xor ( n9625 , n9624 , n176920 );
buf ( n177035 , n9625 );
buf ( n177036 , n177035 );
and ( n9628 , n9623 , n177036 );
and ( n9629 , n176941 , n177031 );
or ( n9630 , n9628 , n9629 );
buf ( n177040 , n9630 );
buf ( n177041 , n177040 );
xor ( n9633 , n176849 , n176925 );
xor ( n9634 , n9633 , n176930 );
buf ( n177044 , n9634 );
buf ( n177045 , n177044 );
nor ( n9637 , n177041 , n177045 );
buf ( n177047 , n9637 );
buf ( n177048 , n177047 );
xor ( n9640 , n176941 , n177031 );
xor ( n9641 , n9640 , n177036 );
buf ( n177051 , n9641 );
buf ( n177052 , n177051 );
buf ( n177053 , n799 );
buf ( n177054 , n827 );
or ( n9646 , n177053 , n177054 );
buf ( n177056 , n828 );
nand ( n9648 , n9646 , n177056 );
buf ( n177058 , n9648 );
buf ( n177059 , n177058 );
buf ( n177060 , n799 );
buf ( n177061 , n827 );
nand ( n9653 , n177060 , n177061 );
buf ( n177063 , n9653 );
buf ( n177064 , n177063 );
buf ( n177065 , n826 );
and ( n9657 , n177059 , n177064 , n177065 );
buf ( n177067 , n9657 );
buf ( n177068 , n177067 );
buf ( n177069 , n795 );
buf ( n177070 , n830 );
xor ( n9662 , n177069 , n177070 );
buf ( n177072 , n9662 );
buf ( n177073 , n177072 );
not ( n9665 , n177073 );
buf ( n177075 , n168471 );
not ( n9667 , n177075 );
or ( n9668 , n9665 , n9667 );
buf ( n177078 , n176965 );
buf ( n177079 , n831 );
nand ( n9671 , n177078 , n177079 );
buf ( n177081 , n9671 );
buf ( n177082 , n177081 );
nand ( n9674 , n9668 , n177082 );
buf ( n177084 , n9674 );
buf ( n177085 , n177084 );
and ( n9677 , n177068 , n177085 );
buf ( n177087 , n9677 );
buf ( n177088 , n798 );
buf ( n177089 , n826 );
xor ( n9681 , n177088 , n177089 );
buf ( n177091 , n9681 );
buf ( n177092 , n177091 );
not ( n9684 , n177092 );
buf ( n177094 , n175400 );
not ( n9686 , n177094 );
or ( n9687 , n9684 , n9686 );
buf ( n177097 , n169081 );
buf ( n177098 , n176857 );
nand ( n9690 , n177097 , n177098 );
buf ( n177100 , n9690 );
buf ( n177101 , n177100 );
nand ( n9693 , n9687 , n177101 );
buf ( n177103 , n9693 );
xor ( n9695 , n177087 , n177103 );
xor ( n9696 , n176956 , n176977 );
xnor ( n9697 , n9696 , n177004 );
and ( n9698 , n9695 , n9697 );
and ( n9699 , n177087 , n177103 );
or ( n9700 , n9698 , n9699 );
buf ( n177110 , n9700 );
buf ( n9702 , n177110 );
buf ( n177112 , n9702 );
buf ( n177113 , n177112 );
not ( n9705 , n177113 );
not ( n9706 , n177010 );
xor ( n9707 , n176952 , n9706 );
buf ( n177117 , n9707 );
not ( n9709 , n177117 );
buf ( n177119 , n9709 );
buf ( n177120 , n177119 );
not ( n9712 , n177120 );
buf ( n177122 , n177020 );
not ( n9714 , n177122 );
or ( n9715 , n9712 , n9714 );
buf ( n177125 , n9707 );
buf ( n177126 , n9608 );
nand ( n9718 , n177125 , n177126 );
buf ( n177128 , n9718 );
buf ( n177129 , n177128 );
nand ( n9721 , n9715 , n177129 );
buf ( n177131 , n9721 );
buf ( n9723 , n177131 );
buf ( n177133 , n9723 );
buf ( n9725 , n177133 );
buf ( n177135 , n9725 );
buf ( n177136 , n177135 );
not ( n9728 , n177136 );
or ( n9729 , n9705 , n9728 );
buf ( n177139 , n177135 );
buf ( n177140 , n177112 );
or ( n9732 , n177139 , n177140 );
buf ( n177142 , n856 );
nand ( n9734 , n9732 , n177142 );
buf ( n177144 , n9734 );
buf ( n177145 , n177144 );
nand ( n9737 , n9729 , n177145 );
buf ( n177147 , n9737 );
buf ( n177148 , n177147 );
nor ( n9743 , n177052 , n177148 );
buf ( n177150 , n9743 );
buf ( n177151 , n177150 );
nor ( n9746 , n177048 , n177151 );
buf ( n177153 , n9746 );
and ( n9748 , n176826 , n176940 , n177153 );
buf ( n177155 , n856 );
not ( n9750 , n177155 );
buf ( n177157 , n9700 );
not ( n9752 , n177157 );
buf ( n177159 , n9752 );
buf ( n177160 , n177159 );
not ( n9755 , n177160 );
or ( n9756 , n9750 , n9755 );
not ( n9757 , n856 );
nand ( n9758 , n9757 , n9700 );
buf ( n177165 , n9758 );
nand ( n9760 , n9756 , n177165 );
buf ( n177167 , n9760 );
buf ( n177168 , n177167 );
buf ( n177169 , n9723 );
and ( n9764 , n177168 , n177169 );
not ( n9765 , n177168 );
buf ( n177172 , n9723 );
not ( n9767 , n177172 );
buf ( n177174 , n9767 );
buf ( n177175 , n177174 );
and ( n9770 , n9765 , n177175 );
nor ( n9771 , n9764 , n9770 );
buf ( n177178 , n9771 );
buf ( n177179 , n177178 );
buf ( n177180 , n857 );
buf ( n177181 , n797 );
buf ( n177182 , n828 );
xor ( n9777 , n177181 , n177182 );
buf ( n177184 , n9777 );
buf ( n177185 , n177184 );
not ( n9780 , n177185 );
buf ( n177187 , n170990 );
not ( n9782 , n177187 );
or ( n9783 , n9780 , n9782 );
buf ( n177190 , n168559 );
buf ( n177191 , n176992 );
nand ( n9786 , n177190 , n177191 );
buf ( n177193 , n9786 );
buf ( n177194 , n177193 );
nand ( n9789 , n9783 , n177194 );
buf ( n177196 , n9789 );
buf ( n177197 , n177196 );
xor ( n9792 , n177068 , n177085 );
buf ( n177199 , n9792 );
buf ( n177200 , n177199 );
xor ( n9795 , n177197 , n177200 );
buf ( n177202 , n826 );
buf ( n177203 , n799 );
xor ( n9798 , n177202 , n177203 );
buf ( n177205 , n9798 );
buf ( n177206 , n177205 );
not ( n9801 , n177206 );
buf ( n177208 , n175400 );
not ( n9803 , n177208 );
or ( n9804 , n9801 , n9803 );
buf ( n177211 , n169081 );
buf ( n177212 , n177091 );
nand ( n9807 , n177211 , n177212 );
buf ( n177214 , n9807 );
buf ( n177215 , n177214 );
nand ( n9810 , n9804 , n177215 );
buf ( n177217 , n9810 );
buf ( n177218 , n177217 );
and ( n9813 , n9795 , n177218 );
and ( n9814 , n177197 , n177200 );
or ( n9815 , n9813 , n9814 );
buf ( n177222 , n9815 );
buf ( n177223 , n177222 );
xor ( n9818 , n177180 , n177223 );
xor ( n9819 , n177087 , n177103 );
xor ( n9820 , n9819 , n9697 );
buf ( n177227 , n9820 );
and ( n9822 , n9818 , n177227 );
and ( n9823 , n177180 , n177223 );
or ( n9824 , n9822 , n9823 );
buf ( n177231 , n9824 );
buf ( n177232 , n177231 );
or ( n9827 , n177179 , n177232 );
buf ( n177234 , n9827 );
buf ( n177235 , n177234 );
xor ( n9830 , n177180 , n177223 );
xor ( n9831 , n9830 , n177227 );
buf ( n177238 , n9831 );
buf ( n177239 , n177238 );
buf ( n177240 , n858 );
buf ( n177241 , n796 );
buf ( n177242 , n830 );
xor ( n9837 , n177241 , n177242 );
buf ( n177244 , n9837 );
buf ( n177245 , n177244 );
not ( n9840 , n177245 );
buf ( n177247 , n168471 );
not ( n9842 , n177247 );
or ( n9843 , n9840 , n9842 );
buf ( n177250 , n177072 );
buf ( n177251 , n831 );
nand ( n9846 , n177250 , n177251 );
buf ( n177253 , n9846 );
buf ( n177254 , n177253 );
nand ( n9849 , n9843 , n177254 );
buf ( n177256 , n9849 );
not ( n9851 , n177256 );
buf ( n177258 , n799 );
buf ( n177259 , n169081 );
nand ( n9854 , n177258 , n177259 );
buf ( n177261 , n9854 );
buf ( n177262 , n177261 );
not ( n9857 , n177262 );
buf ( n177264 , n9857 );
not ( n9859 , n177264 );
or ( n9860 , n9851 , n9859 );
buf ( n177267 , n177261 );
not ( n9862 , n177267 );
buf ( n177269 , n177256 );
not ( n9864 , n177269 );
buf ( n177271 , n9864 );
buf ( n177272 , n177271 );
not ( n177273 , n177272 );
or ( n9868 , n9862 , n177273 );
buf ( n177275 , n798 );
buf ( n177276 , n828 );
xor ( n9871 , n177275 , n177276 );
buf ( n177278 , n9871 );
buf ( n177279 , n177278 );
not ( n9874 , n177279 );
buf ( n177281 , n170990 );
not ( n9876 , n177281 );
or ( n9877 , n9874 , n9876 );
buf ( n177284 , n168559 );
buf ( n177285 , n177184 );
nand ( n9880 , n177284 , n177285 );
buf ( n177287 , n9880 );
buf ( n177288 , n177287 );
nand ( n9883 , n9877 , n177288 );
buf ( n177290 , n9883 );
buf ( n177291 , n177290 );
nand ( n9886 , n9868 , n177291 );
buf ( n177293 , n9886 );
nand ( n9888 , n9860 , n177293 );
buf ( n177295 , n9888 );
xor ( n9890 , n177240 , n177295 );
xor ( n9891 , n177197 , n177200 );
xor ( n9892 , n9891 , n177218 );
buf ( n177299 , n9892 );
buf ( n177300 , n177299 );
and ( n9895 , n9890 , n177300 );
and ( n9896 , n177240 , n177295 );
or ( n9897 , n9895 , n9896 );
buf ( n177304 , n9897 );
buf ( n177305 , n177304 );
nand ( n9900 , n177239 , n177305 );
buf ( n177307 , n9900 );
buf ( n177308 , n177307 );
not ( n9903 , n177308 );
buf ( n177310 , n9903 );
buf ( n177311 , n177310 );
and ( n9906 , n177235 , n177311 );
buf ( n177313 , n177178 );
buf ( n177314 , n177231 );
and ( n9909 , n177313 , n177314 );
buf ( n177316 , n9909 );
buf ( n177317 , n177316 );
nor ( n9912 , n9906 , n177317 );
buf ( n177319 , n9912 );
buf ( n177320 , n177319 );
buf ( n177321 , n177234 );
buf ( n177322 , n859 );
buf ( n177323 , n168471 );
not ( n9918 , n177323 );
buf ( n177325 , n797 );
buf ( n177326 , n830 );
xor ( n9921 , n177325 , n177326 );
buf ( n177328 , n9921 );
buf ( n177329 , n177328 );
not ( n9924 , n177329 );
or ( n9925 , n9918 , n9924 );
buf ( n177332 , n177244 );
buf ( n177333 , n831 );
nand ( n9928 , n177332 , n177333 );
buf ( n177335 , n9928 );
buf ( n177336 , n177335 );
nand ( n9931 , n9925 , n177336 );
buf ( n177338 , n9931 );
buf ( n177339 , n177338 );
buf ( n177340 , n799 );
buf ( n177341 , n829 );
or ( n9936 , n177340 , n177341 );
buf ( n177343 , n830 );
nand ( n9938 , n9936 , n177343 );
buf ( n177345 , n9938 );
buf ( n177346 , n177345 );
buf ( n177347 , n799 );
buf ( n177348 , n829 );
nand ( n9943 , n177347 , n177348 );
buf ( n177350 , n9943 );
buf ( n177351 , n177350 );
buf ( n177352 , n828 );
nand ( n9947 , n177346 , n177351 , n177352 );
buf ( n177354 , n9947 );
buf ( n177355 , n177354 );
not ( n9950 , n177355 );
buf ( n177357 , n9950 );
buf ( n177358 , n177357 );
and ( n9953 , n177339 , n177358 );
buf ( n177360 , n9953 );
buf ( n177361 , n177360 );
xor ( n9956 , n177322 , n177361 );
xor ( n9957 , n177264 , n177271 );
xnor ( n9958 , n9957 , n177290 );
buf ( n177365 , n9958 );
and ( n9960 , n9956 , n177365 );
and ( n9961 , n177322 , n177361 );
or ( n9962 , n9960 , n9961 );
buf ( n177369 , n9962 );
buf ( n177370 , n177369 );
xor ( n9965 , n177240 , n177295 );
xor ( n9966 , n9965 , n177300 );
buf ( n177373 , n9966 );
buf ( n177374 , n177373 );
nor ( n9969 , n177370 , n177374 );
buf ( n177376 , n9969 );
buf ( n177377 , n177376 );
xor ( n9972 , n177322 , n177361 );
xor ( n9973 , n9972 , n177365 );
buf ( n177380 , n9973 );
buf ( n177381 , n177380 );
buf ( n177382 , n860 );
buf ( n177383 , n799 );
buf ( n177384 , n828 );
xor ( n9979 , n177383 , n177384 );
buf ( n177386 , n9979 );
buf ( n177387 , n177386 );
not ( n9982 , n177387 );
buf ( n177389 , n170990 );
not ( n9984 , n177389 );
or ( n9985 , n9982 , n9984 );
buf ( n177392 , n168559 );
buf ( n177393 , n177278 );
nand ( n9988 , n177392 , n177393 );
buf ( n177395 , n9988 );
buf ( n177396 , n177395 );
nand ( n9991 , n9985 , n177396 );
buf ( n177398 , n9991 );
buf ( n177399 , n177398 );
xor ( n9997 , n177382 , n177399 );
buf ( n177401 , n177354 );
not ( n9999 , n177401 );
buf ( n177403 , n177338 );
not ( n177404 , n177403 );
or ( n10002 , n9999 , n177404 );
buf ( n10003 , n6213 );
buf ( n177407 , n10003 );
buf ( n177408 , n177328 );
not ( n10006 , n177408 );
buf ( n177410 , n10006 );
buf ( n177411 , n177410 );
or ( n10009 , n177407 , n177411 );
not ( n10010 , n831 );
buf ( n177414 , n10010 );
buf ( n177415 , n177244 );
not ( n10013 , n177415 );
buf ( n177417 , n10013 );
buf ( n177418 , n177417 );
or ( n10016 , n177414 , n177418 );
buf ( n177420 , n177357 );
nand ( n10018 , n10009 , n10016 , n177420 );
buf ( n177422 , n10018 );
buf ( n177423 , n177422 );
nand ( n10021 , n10002 , n177423 );
buf ( n177425 , n10021 );
buf ( n177426 , n177425 );
and ( n10024 , n9997 , n177426 );
and ( n10025 , n177382 , n177399 );
or ( n10026 , n10024 , n10025 );
buf ( n177430 , n10026 );
buf ( n177431 , n177430 );
nand ( n10029 , n177381 , n177431 );
buf ( n177433 , n10029 );
buf ( n177434 , n177433 );
or ( n10032 , n177377 , n177434 );
buf ( n177436 , n177373 );
buf ( n10034 , n177436 );
buf ( n177438 , n10034 );
buf ( n177439 , n177438 );
buf ( n177440 , n177369 );
nand ( n10038 , n177439 , n177440 );
buf ( n177442 , n10038 );
buf ( n177443 , n177442 );
nand ( n10041 , n10032 , n177443 );
buf ( n177445 , n10041 );
buf ( n177446 , n177445 );
buf ( n177447 , n177238 );
buf ( n177448 , n177304 );
nor ( n10046 , n177447 , n177448 );
buf ( n177450 , n10046 );
buf ( n177451 , n177450 );
not ( n10049 , n177451 );
buf ( n177453 , n10049 );
buf ( n177454 , n177453 );
nand ( n10052 , n177321 , n177446 , n177454 );
buf ( n177456 , n10052 );
buf ( n177457 , n177456 );
buf ( n177458 , n177234 );
buf ( n177459 , n177373 );
buf ( n177460 , n177369 );
nor ( n10058 , n177459 , n177460 );
buf ( n177462 , n10058 );
buf ( n177463 , n177462 );
buf ( n177464 , n177380 );
buf ( n177465 , n177430 );
nor ( n10063 , n177464 , n177465 );
buf ( n177467 , n10063 );
buf ( n177468 , n177467 );
nor ( n10066 , n177463 , n177468 );
buf ( n177470 , n10066 );
buf ( n177471 , n177470 );
buf ( n177472 , n861 );
buf ( n177473 , n168478 );
not ( n10071 , n177473 );
buf ( n177475 , n168471 );
not ( n10073 , n177475 );
or ( n10074 , n10071 , n10073 );
buf ( n177478 , n831 );
buf ( n177479 , n177328 );
nand ( n10077 , n177478 , n177479 );
buf ( n177481 , n10077 );
buf ( n177482 , n177481 );
nand ( n10080 , n10074 , n177482 );
buf ( n177484 , n10080 );
buf ( n177485 , n177484 );
xor ( n10083 , n177472 , n177485 );
buf ( n177487 , n176767 );
buf ( n177488 , n799 );
and ( n10086 , n177487 , n177488 );
buf ( n177490 , n10086 );
buf ( n177491 , n177490 );
xor ( n177492 , n10083 , n177491 );
buf ( n177493 , n177492 );
buf ( n177494 , n177493 );
and ( n10092 , n168512 , n168513 );
buf ( n177496 , n10092 );
buf ( n177497 , n177496 );
nor ( n10095 , n177494 , n177497 );
buf ( n177499 , n10095 );
buf ( n177500 , n177499 );
buf ( n177501 , n168485 );
not ( n10099 , n177501 );
buf ( n177503 , n168518 );
nand ( n10101 , n10099 , n177503 );
buf ( n177505 , n10101 );
buf ( n177506 , n168511 );
not ( n10104 , n177506 );
buf ( n177508 , n10104 );
and ( n10106 , n177505 , n177508 );
and ( n10107 , n168485 , n168515 );
nor ( n10108 , n10106 , n10107 );
buf ( n177512 , n10108 );
nor ( n10110 , n177500 , n177512 );
buf ( n177514 , n10110 );
buf ( n177515 , n177514 );
not ( n10113 , n177515 );
buf ( n177517 , n177493 );
buf ( n177518 , n177496 );
nand ( n10116 , n177517 , n177518 );
buf ( n177520 , n10116 );
buf ( n177521 , n177520 );
nand ( n10119 , n10113 , n177521 );
buf ( n177523 , n10119 );
not ( n10121 , n177523 );
xor ( n177525 , n177382 , n177399 );
xor ( n10123 , n177525 , n177426 );
buf ( n177527 , n10123 );
buf ( n177528 , n177527 );
xor ( n10126 , n177472 , n177485 );
and ( n10127 , n10126 , n177491 );
and ( n10128 , n177472 , n177485 );
or ( n10129 , n10127 , n10128 );
buf ( n177533 , n10129 );
buf ( n177534 , n177533 );
nor ( n10132 , n177528 , n177534 );
buf ( n177536 , n10132 );
buf ( n177537 , n177536 );
not ( n10135 , n177537 );
buf ( n177539 , n10135 );
not ( n10137 , n177539 );
or ( n10138 , n10121 , n10137 );
buf ( n177542 , n177527 );
buf ( n10140 , n177542 );
buf ( n177544 , n10140 );
buf ( n177545 , n177544 );
buf ( n177546 , n177533 );
nand ( n10144 , n177545 , n177546 );
buf ( n177548 , n10144 );
nand ( n10146 , n10138 , n177548 );
buf ( n177550 , n10146 );
and ( n10148 , n177471 , n177550 );
buf ( n177552 , n10148 );
buf ( n177553 , n177552 );
buf ( n177554 , n177453 );
nand ( n10152 , n177458 , n177553 , n177554 );
buf ( n177556 , n10152 );
buf ( n177557 , n177556 );
nand ( n10155 , n177320 , n177457 , n177557 );
buf ( n177559 , n10155 );
buf ( n177560 , n177559 );
not ( n10158 , n177560 );
buf ( n177562 , n10158 );
buf ( n177563 , n177562 );
not ( n10161 , n177563 );
buf ( n177565 , n10161 );
nand ( n10163 , n9748 , n177565 );
buf ( n177567 , n177047 );
buf ( n177568 , n177051 );
buf ( n177569 , n177147 );
nand ( n10167 , n177568 , n177569 );
buf ( n177571 , n10167 );
buf ( n177572 , n177571 );
or ( n10170 , n177567 , n177572 );
buf ( n177574 , n177044 );
buf ( n177575 , n177040 );
nand ( n10173 , n177574 , n177575 );
buf ( n177577 , n10173 );
buf ( n177578 , n177577 );
nand ( n10176 , n10170 , n177578 );
buf ( n177580 , n10176 );
buf ( n177581 , n177580 );
not ( n10179 , n177581 );
not ( n10180 , n176686 );
not ( n10181 , n176820 );
and ( n10182 , n10180 , n10181 );
buf ( n177586 , n176844 );
buf ( n177587 , n176934 );
nor ( n10185 , n177586 , n177587 );
buf ( n177589 , n10185 );
nor ( n10187 , n10182 , n177589 );
buf ( n177591 , n10187 );
not ( n10189 , n177591 );
or ( n10190 , n10179 , n10189 );
buf ( n177594 , n176826 );
buf ( n177595 , n176844 );
buf ( n177596 , n176934 );
nand ( n10194 , n177595 , n177596 );
buf ( n177598 , n10194 );
buf ( n177599 , n177598 );
not ( n10197 , n177599 );
buf ( n177601 , n10197 );
buf ( n177602 , n177601 );
and ( n10200 , n177594 , n177602 );
buf ( n177604 , n176689 );
buf ( n177605 , n176823 );
nor ( n177606 , n177604 , n177605 );
buf ( n177607 , n177606 );
buf ( n177608 , n177607 );
nor ( n10206 , n10200 , n177608 );
buf ( n177610 , n10206 );
buf ( n177611 , n177610 );
nand ( n10209 , n10190 , n177611 );
buf ( n177613 , n10209 );
buf ( n177614 , n177613 );
not ( n10212 , n177614 );
buf ( n177616 , n10212 );
nand ( n10214 , n10163 , n177616 );
buf ( n177618 , n10214 );
not ( n10216 , n177618 );
or ( n10217 , n9268 , n10216 );
buf ( n177621 , n176453 );
buf ( n177622 , n176568 );
nor ( n10220 , n177621 , n177622 );
buf ( n177624 , n10220 );
buf ( n177625 , n177624 );
buf ( n177626 , n176573 );
buf ( n177627 , n176674 );
nand ( n10225 , n177626 , n177627 );
buf ( n177629 , n10225 );
buf ( n177630 , n177629 );
or ( n10228 , n177625 , n177630 );
buf ( n177632 , n176453 );
buf ( n177633 , n176568 );
nand ( n10231 , n177632 , n177633 );
buf ( n177635 , n10231 );
buf ( n177636 , n177635 );
nand ( n10234 , n10228 , n177636 );
buf ( n177638 , n10234 );
not ( n10236 , n177638 );
not ( n10237 , n176449 );
or ( n177641 , n10236 , n10237 );
buf ( n177642 , n176305 );
buf ( n177643 , n176443 );
and ( n10244 , n177642 , n177643 );
buf ( n177645 , n10244 );
buf ( n177646 , n177645 );
buf ( n177647 , n176298 );
not ( n10248 , n177647 );
buf ( n177649 , n176212 );
not ( n10250 , n177649 );
buf ( n177651 , n10250 );
buf ( n177652 , n177651 );
nand ( n10253 , n10248 , n177652 );
buf ( n177654 , n10253 );
buf ( n177655 , n177654 );
and ( n10256 , n177646 , n177655 );
buf ( n177657 , n176298 );
not ( n10258 , n177657 );
buf ( n177659 , n177651 );
nor ( n10260 , n10258 , n177659 );
buf ( n177661 , n10260 );
buf ( n177662 , n177661 );
nor ( n10263 , n10256 , n177662 );
buf ( n177664 , n10263 );
nand ( n10265 , n177641 , n177664 );
not ( n10266 , n10265 );
buf ( n177667 , n10266 );
nand ( n10268 , n10217 , n177667 );
buf ( n177669 , n10268 );
buf ( n177670 , n177669 );
and ( n10271 , n176208 , n176209 , n177670 );
buf ( n177672 , n10271 );
buf ( n177673 , n177672 );
and ( n10274 , n176207 , n177673 );
buf ( n177675 , n173180 );
not ( n10276 , n177675 );
buf ( n177677 , n173187 );
nor ( n10278 , n10276 , n177677 );
buf ( n177679 , n10278 );
buf ( n177680 , n177679 );
not ( n10281 , n177680 );
buf ( n177682 , n172813 );
not ( n10283 , n177682 );
or ( n10284 , n10281 , n10283 );
buf ( n177685 , n172807 );
buf ( n177686 , n172491 );
nand ( n177687 , n177685 , n177686 );
buf ( n177688 , n177687 );
buf ( n177689 , n177688 );
nand ( n10290 , n10284 , n177689 );
buf ( n177691 , n10290 );
buf ( n177692 , n177691 );
not ( n10293 , n177692 );
buf ( n177694 , n5018 );
not ( n10295 , n177694 );
or ( n10296 , n10293 , n10295 );
not ( n10297 , n172157 );
not ( n10298 , n171670 );
nand ( n10299 , n10297 , n10298 );
buf ( n177700 , n172162 );
buf ( n177701 , n172483 );
nand ( n10302 , n177700 , n177701 );
buf ( n177703 , n10302 );
buf ( n177704 , n177703 );
not ( n10305 , n177704 );
buf ( n177706 , n10305 );
and ( n10307 , n10299 , n177706 );
buf ( n177708 , n171670 );
buf ( n177709 , n172157 );
nand ( n10310 , n177708 , n177709 );
buf ( n177711 , n10310 );
buf ( n177712 , n177711 );
not ( n10313 , n177712 );
buf ( n177714 , n10313 );
nor ( n10315 , n10307 , n177714 );
buf ( n177716 , n10315 );
nand ( n10317 , n10296 , n177716 );
buf ( n177718 , n10317 );
buf ( n177719 , n177718 );
nor ( n10320 , n10274 , n177719 );
buf ( n177721 , n10320 );
buf ( n177722 , n177721 );
nand ( n10323 , n176181 , n177722 );
buf ( n177724 , n10323 );
buf ( n177725 , n177724 );
buf ( n10326 , n177725 );
buf ( n177727 , n10326 );
buf ( n177728 , n177727 );
not ( n10329 , n177728 );
or ( n177730 , n4198 , n10329 );
buf ( n177731 , n176180 );
buf ( n177732 , n177721 );
nand ( n10333 , n177731 , n177732 );
buf ( n177734 , n10333 );
buf ( n177735 , n177734 );
buf ( n10336 , n177735 );
buf ( n177737 , n10336 );
buf ( n177738 , n177737 );
buf ( n10339 , n177738 );
buf ( n177740 , n10339 );
buf ( n177741 , n177740 );
buf ( n177742 , n171665 );
or ( n10343 , n177741 , n177742 );
nand ( n10344 , n177730 , n10343 );
buf ( n177745 , n10344 );
buf ( n10346 , n177745 );
buf ( n177747 , n795 );
buf ( n177748 , n800 );
and ( n10349 , n177747 , n177748 );
buf ( n177750 , n10349 );
buf ( n177751 , n177750 );
buf ( n177752 , n794 );
buf ( n177753 , n800 );
xor ( n10354 , n177752 , n177753 );
buf ( n177755 , n10354 );
buf ( n177756 , n177755 );
not ( n10357 , n177756 );
buf ( n177758 , n3497 );
not ( n10359 , n177758 );
or ( n10360 , n10357 , n10359 );
buf ( n177761 , n170972 );
xor ( n10362 , n800 , n793 );
buf ( n177763 , n10362 );
nand ( n10364 , n177761 , n177763 );
buf ( n177765 , n10364 );
buf ( n177766 , n177765 );
nand ( n10367 , n10360 , n177766 );
buf ( n177768 , n10367 );
buf ( n177769 , n177768 );
xor ( n10370 , n177751 , n177769 );
buf ( n177771 , n768 );
buf ( n177772 , n826 );
xor ( n10373 , n177771 , n177772 );
buf ( n177774 , n10373 );
buf ( n177775 , n177774 );
not ( n10376 , n177775 );
buf ( n177777 , n4337 );
not ( n10378 , n177777 );
or ( n10379 , n10376 , n10378 );
buf ( n177780 , n169081 );
buf ( n177781 , n826 );
nand ( n177782 , n177780 , n177781 );
buf ( n177783 , n177782 );
buf ( n177784 , n177783 );
nand ( n10385 , n10379 , n177784 );
buf ( n177786 , n10385 );
buf ( n177787 , n177786 );
not ( n10388 , n177787 );
buf ( n177789 , n10388 );
buf ( n177790 , n177789 );
xor ( n10391 , n10370 , n177790 );
buf ( n177792 , n10391 );
buf ( n177793 , n177792 );
buf ( n177794 , n768 );
buf ( n177795 , n828 );
xor ( n10396 , n177794 , n177795 );
buf ( n177797 , n10396 );
buf ( n177798 , n177797 );
not ( n10399 , n177798 );
buf ( n177800 , n170990 );
not ( n10401 , n177800 );
or ( n10402 , n10399 , n10401 );
buf ( n177803 , n828 );
buf ( n177804 , n168559 );
nand ( n10405 , n177803 , n177804 );
buf ( n177806 , n10405 );
buf ( n177807 , n177806 );
nand ( n10408 , n10402 , n177807 );
buf ( n177809 , n10408 );
buf ( n177810 , n177809 );
buf ( n177811 , n795 );
buf ( n177812 , n800 );
xor ( n10413 , n177811 , n177812 );
buf ( n177814 , n10413 );
buf ( n177815 , n177814 );
not ( n10416 , n177815 );
buf ( n177817 , n3497 );
buf ( n10418 , n177817 );
buf ( n177819 , n10418 );
buf ( n177820 , n177819 );
not ( n10421 , n177820 );
or ( n177822 , n10416 , n10421 );
buf ( n177823 , n170972 );
buf ( n177824 , n177755 );
nand ( n10425 , n177823 , n177824 );
buf ( n177826 , n10425 );
buf ( n177827 , n177826 );
nand ( n10428 , n177822 , n177827 );
buf ( n177829 , n10428 );
buf ( n177830 , n177829 );
xor ( n10431 , n177810 , n177830 );
buf ( n177832 , n797 );
buf ( n177833 , n800 );
and ( n10434 , n177832 , n177833 );
buf ( n177835 , n10434 );
buf ( n177836 , n177835 );
buf ( n177837 , n774 );
buf ( n177838 , n822 );
xor ( n10439 , n177837 , n177838 );
buf ( n177840 , n10439 );
buf ( n177841 , n177840 );
not ( n10442 , n177841 );
buf ( n177843 , n2418 );
not ( n10444 , n177843 );
or ( n10445 , n10442 , n10444 );
buf ( n177846 , n169417 );
buf ( n177847 , n773 );
buf ( n177848 , n822 );
xor ( n10449 , n177847 , n177848 );
buf ( n177850 , n10449 );
buf ( n177851 , n177850 );
nand ( n10452 , n177846 , n177851 );
buf ( n177853 , n10452 );
buf ( n177854 , n177853 );
nand ( n10455 , n10445 , n177854 );
buf ( n177856 , n10455 );
buf ( n177857 , n177856 );
xor ( n10458 , n177836 , n177857 );
buf ( n177859 , n770 );
buf ( n177860 , n826 );
xor ( n10461 , n177859 , n177860 );
buf ( n177862 , n10461 );
buf ( n177863 , n177862 );
not ( n10464 , n177863 );
buf ( n177865 , n1621 );
not ( n10466 , n177865 );
or ( n10467 , n10464 , n10466 );
buf ( n177868 , n168684 );
buf ( n177869 , n769 );
buf ( n177870 , n826 );
xor ( n10471 , n177869 , n177870 );
buf ( n177872 , n10471 );
buf ( n177873 , n177872 );
nand ( n10474 , n177868 , n177873 );
buf ( n177875 , n10474 );
buf ( n177876 , n177875 );
nand ( n10477 , n10467 , n177876 );
buf ( n177878 , n10477 );
buf ( n177879 , n177878 );
and ( n10480 , n10458 , n177879 );
and ( n10481 , n177836 , n177857 );
or ( n10482 , n10480 , n10481 );
buf ( n177883 , n10482 );
buf ( n177884 , n177883 );
and ( n10485 , n10431 , n177884 );
and ( n10486 , n177810 , n177830 );
or ( n10487 , n10485 , n10486 );
buf ( n177888 , n10487 );
buf ( n177889 , n177888 );
xor ( n10490 , n177793 , n177889 );
buf ( n177891 , n782 );
buf ( n177892 , n814 );
xor ( n10493 , n177891 , n177892 );
buf ( n177894 , n10493 );
buf ( n177895 , n177894 );
not ( n10496 , n177895 );
buf ( n177897 , n169241 );
not ( n10498 , n177897 );
or ( n10499 , n10496 , n10498 );
buf ( n177900 , n169931 );
buf ( n177901 , n781 );
buf ( n177902 , n814 );
xor ( n10503 , n177901 , n177902 );
buf ( n177904 , n10503 );
buf ( n177905 , n177904 );
nand ( n10506 , n177900 , n177905 );
buf ( n177907 , n10506 );
buf ( n177908 , n177907 );
nand ( n10509 , n10499 , n177908 );
buf ( n177910 , n10509 );
buf ( n177911 , n177910 );
not ( n177912 , n177911 );
not ( n10516 , n168656 );
xor ( n10517 , n820 , n775 );
not ( n10518 , n10517 );
or ( n10519 , n10516 , n10518 );
buf ( n177917 , n776 );
buf ( n177918 , n820 );
xnor ( n10522 , n177917 , n177918 );
buf ( n177920 , n10522 );
or ( n10524 , n169988 , n177920 );
nand ( n10525 , n10519 , n10524 );
buf ( n177923 , n10525 );
not ( n10527 , n177923 );
or ( n10528 , n177912 , n10527 );
buf ( n177926 , n177910 );
buf ( n177927 , n10525 );
or ( n10531 , n177926 , n177927 );
buf ( n177929 , n784 );
buf ( n177930 , n812 );
xor ( n10534 , n177929 , n177930 );
buf ( n177932 , n10534 );
buf ( n177933 , n177932 );
not ( n10537 , n177933 );
buf ( n177935 , n1553 );
not ( n10539 , n177935 );
or ( n10540 , n10537 , n10539 );
buf ( n177938 , n1534 );
buf ( n177939 , n783 );
buf ( n177940 , n812 );
xor ( n10544 , n177939 , n177940 );
buf ( n177942 , n10544 );
buf ( n177943 , n177942 );
nand ( n177944 , n177938 , n177943 );
buf ( n177945 , n177944 );
buf ( n177946 , n177945 );
nand ( n10550 , n10540 , n177946 );
buf ( n177948 , n10550 );
buf ( n177949 , n177948 );
nand ( n10553 , n10531 , n177949 );
buf ( n177951 , n10553 );
buf ( n177952 , n177951 );
nand ( n10556 , n10528 , n177952 );
buf ( n177954 , n10556 );
buf ( n177955 , n177954 );
buf ( n177956 , n772 );
buf ( n177957 , n824 );
xor ( n10561 , n177956 , n177957 );
buf ( n177959 , n10561 );
buf ( n177960 , n177959 );
not ( n10564 , n177960 );
buf ( n177962 , n169154 );
not ( n10566 , n177962 );
or ( n10567 , n10564 , n10566 );
buf ( n177965 , n170565 );
buf ( n177966 , n771 );
buf ( n177967 , n824 );
xor ( n10571 , n177966 , n177967 );
buf ( n177969 , n10571 );
buf ( n177970 , n177969 );
nand ( n10574 , n177965 , n177970 );
buf ( n177972 , n10574 );
buf ( n177973 , n177972 );
nand ( n10577 , n10567 , n177973 );
buf ( n177975 , n10577 );
buf ( n177976 , n788 );
buf ( n177977 , n808 );
xor ( n10581 , n177976 , n177977 );
buf ( n177979 , n10581 );
buf ( n177980 , n177979 );
not ( n10584 , n177980 );
buf ( n177982 , n169542 );
not ( n10586 , n177982 );
buf ( n177984 , n10586 );
buf ( n177985 , n177984 );
not ( n10589 , n177985 );
or ( n10590 , n10584 , n10589 );
buf ( n177988 , n168619 );
buf ( n177989 , n787 );
buf ( n177990 , n808 );
xor ( n10594 , n177989 , n177990 );
buf ( n177992 , n10594 );
buf ( n177993 , n177992 );
nand ( n10597 , n177988 , n177993 );
buf ( n177995 , n10597 );
buf ( n177996 , n177995 );
nand ( n10600 , n10590 , n177996 );
buf ( n177998 , n10600 );
or ( n10602 , n177975 , n177998 );
buf ( n178000 , n786 );
buf ( n178001 , n810 );
xor ( n10605 , n178000 , n178001 );
buf ( n178003 , n10605 );
buf ( n178004 , n178003 );
not ( n10608 , n178004 );
buf ( n178006 , n2737 );
not ( n10610 , n178006 );
or ( n10611 , n10608 , n10610 );
buf ( n178009 , n169957 );
buf ( n178010 , n785 );
buf ( n178011 , n810 );
xor ( n10615 , n178010 , n178011 );
buf ( n178013 , n10615 );
buf ( n178014 , n178013 );
nand ( n10618 , n178009 , n178014 );
buf ( n178016 , n10618 );
buf ( n178017 , n178016 );
nand ( n10621 , n10611 , n178017 );
buf ( n178019 , n10621 );
nand ( n10623 , n10602 , n178019 );
buf ( n178021 , n177975 );
buf ( n178022 , n177998 );
nand ( n10626 , n178021 , n178022 );
buf ( n178024 , n10626 );
nand ( n10628 , n10623 , n178024 );
buf ( n178026 , n10628 );
or ( n10630 , n177955 , n178026 );
buf ( n178028 , n790 );
buf ( n178029 , n806 );
xor ( n10633 , n178028 , n178029 );
buf ( n178031 , n10633 );
buf ( n178032 , n178031 );
not ( n10636 , n178032 );
buf ( n178034 , n169635 );
not ( n10638 , n178034 );
or ( n10639 , n10636 , n10638 );
buf ( n178037 , n169641 );
buf ( n178038 , n789 );
buf ( n178039 , n806 );
xor ( n10643 , n178038 , n178039 );
buf ( n178041 , n10643 );
buf ( n178042 , n178041 );
nand ( n10646 , n178037 , n178042 );
buf ( n178044 , n10646 );
buf ( n178045 , n178044 );
nand ( n10649 , n10639 , n178045 );
buf ( n178047 , n10649 );
buf ( n178048 , n178047 );
buf ( n178049 , n792 );
buf ( n178050 , n804 );
xor ( n10654 , n178049 , n178050 );
buf ( n178052 , n10654 );
buf ( n178053 , n178052 );
not ( n10657 , n178053 );
buf ( n178055 , n168832 );
not ( n10659 , n178055 );
or ( n10660 , n10657 , n10659 );
buf ( n178058 , n168759 );
buf ( n178059 , n791 );
buf ( n178060 , n804 );
xor ( n10664 , n178059 , n178060 );
buf ( n178062 , n10664 );
buf ( n178063 , n178062 );
nand ( n10667 , n178058 , n178063 );
buf ( n178065 , n10667 );
buf ( n178066 , n178065 );
nand ( n10670 , n10660 , n178066 );
buf ( n178068 , n10670 );
buf ( n178069 , n178068 );
xor ( n10673 , n178048 , n178069 );
buf ( n178071 , n778 );
buf ( n178072 , n818 );
xor ( n10676 , n178071 , n178072 );
buf ( n178074 , n10676 );
buf ( n178075 , n178074 );
not ( n10679 , n178075 );
buf ( n178077 , n1321 );
not ( n10681 , n178077 );
or ( n10682 , n10679 , n10681 );
buf ( n178080 , n168806 );
xor ( n10684 , n777 , n818 );
buf ( n178082 , n10684 );
nand ( n10686 , n178080 , n178082 );
buf ( n178084 , n10686 );
buf ( n178085 , n178084 );
nand ( n10689 , n10682 , n178085 );
buf ( n178087 , n10689 );
buf ( n178088 , n178087 );
and ( n10692 , n10673 , n178088 );
and ( n10693 , n178048 , n178069 );
or ( n10694 , n10692 , n10693 );
buf ( n178092 , n10694 );
buf ( n178093 , n178092 );
nand ( n10697 , n10630 , n178093 );
buf ( n178095 , n10697 );
buf ( n178096 , n178095 );
buf ( n178097 , n177954 );
buf ( n178098 , n10628 );
nand ( n10702 , n178097 , n178098 );
buf ( n178100 , n10702 );
buf ( n178101 , n178100 );
nand ( n10705 , n178096 , n178101 );
buf ( n178103 , n10705 );
buf ( n178104 , n178103 );
and ( n10708 , n10490 , n178104 );
and ( n10709 , n177793 , n177889 );
or ( n10710 , n10708 , n10709 );
buf ( n178108 , n10710 );
buf ( n178109 , n178108 );
buf ( n178110 , n796 );
buf ( n178111 , n800 );
and ( n10715 , n178110 , n178111 );
buf ( n178113 , n10715 );
buf ( n178114 , n178113 );
buf ( n178115 , n177942 );
not ( n10719 , n178115 );
buf ( n178117 , n1553 );
not ( n10721 , n178117 );
or ( n10722 , n10719 , n10721 );
buf ( n178120 , n1534 );
buf ( n178121 , n782 );
buf ( n178122 , n812 );
xor ( n10726 , n178121 , n178122 );
buf ( n178124 , n10726 );
buf ( n178125 , n178124 );
nand ( n10729 , n178120 , n178125 );
buf ( n178127 , n10729 );
buf ( n178128 , n178127 );
nand ( n10732 , n10722 , n178128 );
buf ( n178130 , n10732 );
buf ( n178131 , n178130 );
xor ( n10735 , n178114 , n178131 );
buf ( n178133 , n177904 );
not ( n10737 , n178133 );
buf ( n178135 , n169241 );
not ( n10739 , n178135 );
or ( n10740 , n10737 , n10739 );
buf ( n178138 , n169247 );
buf ( n178139 , n780 );
buf ( n178140 , n814 );
xor ( n10744 , n178139 , n178140 );
buf ( n178142 , n10744 );
buf ( n178143 , n178142 );
nand ( n10747 , n178138 , n178143 );
buf ( n178145 , n10747 );
buf ( n178146 , n178145 );
nand ( n10750 , n10740 , n178146 );
buf ( n178148 , n10750 );
buf ( n178149 , n178148 );
xnor ( n10753 , n10735 , n178149 );
buf ( n178151 , n10753 );
buf ( n178152 , n178151 );
not ( n10756 , n178152 );
buf ( n178154 , n829 );
buf ( n178155 , n830 );
xnor ( n10759 , n178154 , n178155 );
buf ( n178157 , n10759 );
buf ( n178158 , n178157 );
buf ( n178159 , n168547 );
nand ( n10763 , n178158 , n178159 );
buf ( n178161 , n10763 );
buf ( n178162 , n178161 );
not ( n10766 , n178162 );
buf ( n178164 , n176764 );
not ( n10768 , n178164 );
or ( n10769 , n10766 , n10768 );
buf ( n178167 , n828 );
nand ( n10771 , n10769 , n178167 );
buf ( n178169 , n10771 );
buf ( n178170 , n178169 );
not ( n10774 , n178170 );
buf ( n178172 , n10774 );
buf ( n178173 , n177872 );
not ( n10777 , n178173 );
buf ( n178175 , n169674 );
not ( n10782 , n178175 );
or ( n10783 , n10777 , n10782 );
buf ( n178178 , n177774 );
buf ( n178179 , n169081 );
nand ( n10786 , n178178 , n178179 );
buf ( n178181 , n10786 );
buf ( n178182 , n178181 );
nand ( n10789 , n10783 , n178182 );
buf ( n178184 , n10789 );
xor ( n10791 , n178172 , n178184 );
buf ( n178186 , n177850 );
not ( n10793 , n178186 );
buf ( n178188 , n1939 );
not ( n10795 , n178188 );
or ( n10796 , n10793 , n10795 );
buf ( n178191 , n169417 );
buf ( n178192 , n772 );
buf ( n178193 , n822 );
xor ( n10800 , n178192 , n178193 );
buf ( n178195 , n10800 );
buf ( n178196 , n178195 );
nand ( n178197 , n178191 , n178196 );
buf ( n178198 , n178197 );
buf ( n178199 , n178198 );
nand ( n10806 , n10796 , n178199 );
buf ( n178201 , n10806 );
and ( n10808 , n10791 , n178201 );
not ( n10809 , n10791 );
buf ( n178204 , n178201 );
not ( n10811 , n178204 );
buf ( n178206 , n10811 );
and ( n10813 , n10809 , n178206 );
nor ( n10814 , n10808 , n10813 );
buf ( n178209 , n10814 );
not ( n10816 , n178209 );
or ( n10817 , n10756 , n10816 );
buf ( n178212 , n794 );
buf ( n178213 , n802 );
xor ( n10820 , n178212 , n178213 );
buf ( n178215 , n10820 );
buf ( n178216 , n178215 );
not ( n10823 , n178216 );
buf ( n178218 , n802 );
not ( n10825 , n178218 );
buf ( n178220 , n803 );
not ( n10827 , n178220 );
and ( n10828 , n10825 , n10827 );
buf ( n178223 , n802 );
buf ( n178224 , n803 );
and ( n10831 , n178223 , n178224 );
nor ( n10832 , n10828 , n10831 );
buf ( n178227 , n10832 );
buf ( n178228 , n178227 );
not ( n10835 , n178228 );
buf ( n178230 , n168857 );
nor ( n10837 , n10835 , n178230 );
buf ( n178232 , n10837 );
buf ( n178233 , n178232 );
not ( n10840 , n178233 );
or ( n10841 , n10823 , n10840 );
buf ( n178236 , n168867 );
buf ( n178237 , n793 );
buf ( n178238 , n802 );
xor ( n10845 , n178237 , n178238 );
buf ( n178240 , n10845 );
buf ( n178241 , n178240 );
nand ( n10848 , n178236 , n178241 );
buf ( n178243 , n10848 );
buf ( n178244 , n178243 );
nand ( n10851 , n10841 , n178244 );
buf ( n178246 , n10851 );
buf ( n178247 , n178246 );
buf ( n178248 , n796 );
buf ( n178249 , n800 );
xor ( n10856 , n178248 , n178249 );
buf ( n178251 , n10856 );
buf ( n178252 , n178251 );
not ( n10859 , n178252 );
buf ( n178254 , n3497 );
not ( n10861 , n178254 );
or ( n10862 , n10859 , n10861 );
buf ( n178257 , n170972 );
buf ( n178258 , n177814 );
nand ( n10865 , n178257 , n178258 );
buf ( n178260 , n10865 );
buf ( n178261 , n178260 );
nand ( n10868 , n10862 , n178261 );
buf ( n178263 , n10868 );
buf ( n178264 , n178263 );
xor ( n10871 , n178247 , n178264 );
buf ( n178266 , n780 );
buf ( n178267 , n816 );
xor ( n10874 , n178266 , n178267 );
buf ( n178269 , n10874 );
buf ( n178270 , n178269 );
not ( n10877 , n178270 );
buf ( n178272 , n169836 );
not ( n10879 , n178272 );
or ( n10880 , n10877 , n10879 );
buf ( n178275 , n779 );
buf ( n178276 , n816 );
xor ( n10883 , n178275 , n178276 );
buf ( n178278 , n10883 );
buf ( n178279 , n178278 );
buf ( n178280 , n169320 );
nand ( n10887 , n178279 , n178280 );
buf ( n178282 , n10887 );
buf ( n178283 , n178282 );
nand ( n10890 , n10880 , n178283 );
buf ( n178285 , n10890 );
buf ( n178286 , n178285 );
and ( n10893 , n10871 , n178286 );
and ( n10894 , n178247 , n178264 );
or ( n10895 , n10893 , n10894 );
buf ( n178290 , n10895 );
buf ( n178291 , n178290 );
nand ( n10898 , n10817 , n178291 );
buf ( n178293 , n10898 );
buf ( n178294 , n178293 );
buf ( n178295 , n178113 );
buf ( n178296 , n178130 );
xor ( n10903 , n178295 , n178296 );
buf ( n178298 , n178148 );
xnor ( n10905 , n10903 , n178298 );
buf ( n178300 , n10905 );
buf ( n178301 , n178300 );
not ( n10908 , n178301 );
buf ( n178303 , n10814 );
not ( n10910 , n178303 );
buf ( n178305 , n10910 );
buf ( n178306 , n178305 );
nand ( n10913 , n10908 , n178306 );
buf ( n178308 , n10913 );
buf ( n178309 , n178308 );
nand ( n10916 , n178294 , n178309 );
buf ( n178311 , n10916 );
buf ( n178312 , n178311 );
not ( n10919 , n178148 );
not ( n10920 , n178113 );
or ( n10921 , n10919 , n10920 );
buf ( n178316 , n178148 );
buf ( n178317 , n178113 );
nor ( n10924 , n178316 , n178317 );
buf ( n178319 , n10924 );
buf ( n178320 , n178130 );
not ( n178321 , n178320 );
buf ( n178322 , n178321 );
or ( n10929 , n178319 , n178322 );
nand ( n10930 , n10921 , n10929 );
buf ( n178325 , n10930 );
buf ( n178326 , n178184 );
buf ( n178327 , n178201 );
nor ( n10934 , n178326 , n178327 );
buf ( n178329 , n10934 );
buf ( n178330 , n178329 );
buf ( n178331 , n178172 );
or ( n10938 , n178330 , n178331 );
buf ( n178333 , n178184 );
buf ( n178334 , n178201 );
nand ( n10941 , n178333 , n178334 );
buf ( n178336 , n10941 );
buf ( n178337 , n178336 );
nand ( n10944 , n10938 , n178337 );
buf ( n178339 , n10944 );
buf ( n178340 , n178339 );
xor ( n10947 , n178325 , n178340 );
buf ( n178342 , n177992 );
not ( n10949 , n178342 );
buf ( n178344 , n177984 );
not ( n10951 , n178344 );
or ( n10952 , n10949 , n10951 );
buf ( n178347 , n168619 );
xor ( n10954 , n808 , n786 );
buf ( n178349 , n10954 );
nand ( n10956 , n178347 , n178349 );
buf ( n178351 , n10956 );
buf ( n178352 , n178351 );
nand ( n10959 , n10952 , n178352 );
buf ( n178354 , n10959 );
buf ( n178355 , n178354 );
buf ( n178356 , n178013 );
not ( n10963 , n178356 );
buf ( n178358 , n168977 );
not ( n10965 , n178358 );
buf ( n178360 , n10965 );
buf ( n178361 , n178360 );
not ( n10968 , n178361 );
or ( n10969 , n10963 , n10968 );
buf ( n178364 , n170708 );
xor ( n10971 , n810 , n784 );
buf ( n178366 , n10971 );
nand ( n10973 , n178364 , n178366 );
buf ( n178368 , n10973 );
buf ( n178369 , n178368 );
nand ( n10976 , n10969 , n178369 );
buf ( n178371 , n10976 );
buf ( n178372 , n178371 );
xor ( n10979 , n178355 , n178372 );
not ( n10980 , n2513 );
xor ( n178375 , n820 , n774 );
not ( n10982 , n178375 );
or ( n10983 , n10980 , n10982 );
buf ( n178378 , n10517 );
not ( n10985 , n178378 );
buf ( n178380 , n10985 );
or ( n10987 , n169991 , n178380 );
nand ( n10988 , n10983 , n10987 );
buf ( n178383 , n10988 );
and ( n10990 , n10979 , n178383 );
and ( n10991 , n178355 , n178372 );
or ( n10992 , n10990 , n10991 );
buf ( n178387 , n10992 );
buf ( n178388 , n178387 );
xor ( n10995 , n10947 , n178388 );
buf ( n178390 , n10995 );
buf ( n178391 , n178390 );
xor ( n10998 , n178312 , n178391 );
buf ( n178393 , n177969 );
not ( n11000 , n178393 );
buf ( n178395 , n1806 );
not ( n11002 , n178395 );
or ( n11003 , n11000 , n11002 );
buf ( n178398 , n170565 );
buf ( n178399 , n770 );
buf ( n178400 , n824 );
xor ( n11007 , n178399 , n178400 );
buf ( n178402 , n11007 );
buf ( n178403 , n178402 );
nand ( n11010 , n178398 , n178403 );
buf ( n178405 , n11010 );
buf ( n178406 , n178405 );
nand ( n11013 , n11003 , n178406 );
buf ( n178408 , n11013 );
buf ( n178409 , n178408 );
not ( n11016 , n168806 );
xor ( n11017 , n818 , n776 );
not ( n11018 , n11017 );
or ( n11019 , n11016 , n11018 );
not ( n11020 , n1315 );
not ( n11021 , n168788 );
nand ( n11022 , n11020 , n11021 , n10684 );
nand ( n11023 , n11019 , n11022 );
buf ( n178418 , n11023 );
xor ( n11025 , n178409 , n178418 );
buf ( n178420 , n178041 );
not ( n11027 , n178420 );
buf ( n178422 , n168713 );
not ( n11029 , n178422 );
or ( n11030 , n11027 , n11029 );
buf ( n178425 , n169641 );
buf ( n178426 , n788 );
buf ( n178427 , n806 );
xor ( n11034 , n178426 , n178427 );
buf ( n178429 , n11034 );
buf ( n178430 , n178429 );
nand ( n11037 , n178425 , n178430 );
buf ( n178432 , n11037 );
buf ( n178433 , n178432 );
nand ( n11040 , n11030 , n178433 );
buf ( n178435 , n11040 );
buf ( n178436 , n178435 );
and ( n11043 , n11025 , n178436 );
and ( n11044 , n178409 , n178418 );
or ( n11045 , n11043 , n11044 );
buf ( n178440 , n11045 );
buf ( n178441 , n178440 );
not ( n11048 , n178062 );
not ( n11049 , n168750 );
or ( n11050 , n11048 , n11049 );
buf ( n178445 , n168759 );
buf ( n11052 , n178445 );
buf ( n178447 , n11052 );
buf ( n178448 , n178447 );
xor ( n11055 , n804 , n790 );
buf ( n178450 , n11055 );
nand ( n11057 , n178448 , n178450 );
buf ( n178452 , n11057 );
nand ( n11059 , n11050 , n178452 );
buf ( n178454 , n178240 );
not ( n11061 , n178454 );
buf ( n178456 , n168861 );
not ( n11063 , n178456 );
or ( n11064 , n11061 , n11063 );
buf ( n178459 , n168870 );
buf ( n178460 , n792 );
buf ( n178461 , n802 );
xor ( n11068 , n178460 , n178461 );
buf ( n178463 , n11068 );
buf ( n178464 , n178463 );
nand ( n11071 , n178459 , n178464 );
buf ( n178466 , n11071 );
buf ( n178467 , n178466 );
nand ( n11077 , n11064 , n178467 );
buf ( n178469 , n11077 );
or ( n11079 , n11059 , n178469 );
not ( n11080 , n178278 );
not ( n178472 , n169836 );
or ( n11082 , n11080 , n178472 );
buf ( n178474 , n169845 );
buf ( n178475 , n778 );
buf ( n178476 , n816 );
xor ( n11086 , n178475 , n178476 );
buf ( n178478 , n11086 );
buf ( n178479 , n178478 );
nand ( n11089 , n178474 , n178479 );
buf ( n178481 , n11089 );
nand ( n11091 , n11082 , n178481 );
nand ( n11092 , n11079 , n11091 );
buf ( n178484 , n11092 );
buf ( n178485 , n11059 );
buf ( n178486 , n178469 );
nand ( n11096 , n178485 , n178486 );
buf ( n178488 , n11096 );
buf ( n178489 , n178488 );
nand ( n11099 , n178484 , n178489 );
buf ( n178491 , n11099 );
buf ( n178492 , n178491 );
xor ( n11102 , n178441 , n178492 );
buf ( n178494 , n178402 );
not ( n11104 , n178494 );
buf ( n178496 , n169793 );
not ( n11106 , n178496 );
or ( n11107 , n11104 , n11106 );
buf ( n178499 , n175664 );
buf ( n178500 , n769 );
not ( n11110 , n178500 );
buf ( n178502 , n11110 );
and ( n11112 , n824 , n178502 );
not ( n11113 , n824 );
and ( n11114 , n11113 , n769 );
or ( n11115 , n11112 , n11114 );
buf ( n178507 , n11115 );
nand ( n11117 , n178499 , n178507 );
buf ( n178509 , n11117 );
buf ( n178510 , n178509 );
nand ( n11120 , n11107 , n178510 );
buf ( n178512 , n11120 );
buf ( n178513 , n178512 );
buf ( n178514 , n178124 );
not ( n11124 , n178514 );
buf ( n178516 , n1907 );
not ( n11126 , n178516 );
or ( n11127 , n11124 , n11126 );
buf ( n178519 , n3220 );
xor ( n11129 , n812 , n781 );
buf ( n178521 , n11129 );
nand ( n11131 , n178519 , n178521 );
buf ( n178523 , n11131 );
buf ( n178524 , n178523 );
nand ( n11134 , n11127 , n178524 );
buf ( n178526 , n11134 );
buf ( n178527 , n178526 );
xor ( n11137 , n178513 , n178527 );
buf ( n178529 , n178375 );
not ( n11139 , n178529 );
buf ( n178531 , n2251 );
not ( n11141 , n178531 );
or ( n11142 , n11139 , n11141 );
buf ( n178534 , n2513 );
buf ( n178535 , n773 );
buf ( n178536 , n820 );
xor ( n11146 , n178535 , n178536 );
buf ( n178538 , n11146 );
buf ( n178539 , n178538 );
nand ( n11149 , n178534 , n178539 );
buf ( n178541 , n11149 );
buf ( n178542 , n178541 );
nand ( n11152 , n11142 , n178542 );
buf ( n178544 , n11152 );
buf ( n178545 , n178544 );
xor ( n11155 , n11137 , n178545 );
buf ( n178547 , n11155 );
buf ( n178548 , n178547 );
xor ( n11158 , n11102 , n178548 );
buf ( n178550 , n11158 );
buf ( n178551 , n178550 );
and ( n11161 , n10998 , n178551 );
and ( n11162 , n178312 , n178391 );
or ( n11163 , n11161 , n11162 );
buf ( n178555 , n11163 );
buf ( n178556 , n178555 );
xor ( n11166 , n178109 , n178556 );
buf ( n178558 , n177786 );
buf ( n178559 , n11017 );
not ( n11169 , n178559 );
buf ( n178561 , n171706 );
not ( n11171 , n178561 );
or ( n11172 , n11169 , n11171 );
buf ( n178564 , n168803 );
buf ( n178565 , n775 );
buf ( n178566 , n818 );
xor ( n11176 , n178565 , n178566 );
buf ( n178568 , n11176 );
buf ( n178569 , n178568 );
nand ( n11179 , n178564 , n178569 );
buf ( n178571 , n11179 );
buf ( n178572 , n178571 );
nand ( n11182 , n11172 , n178572 );
buf ( n178574 , n11182 );
buf ( n178575 , n178574 );
not ( n11185 , n168615 );
not ( n11186 , n10954 );
or ( n11187 , n11185 , n11186 );
buf ( n178579 , n168619 );
xor ( n11189 , n808 , n785 );
buf ( n178581 , n11189 );
nand ( n11191 , n178579 , n178581 );
buf ( n178583 , n11191 );
nand ( n11193 , n11187 , n178583 );
buf ( n178585 , n11193 );
xor ( n11195 , n178575 , n178585 );
buf ( n178587 , n10971 );
not ( n11197 , n178587 );
buf ( n178589 , n171880 );
not ( n11199 , n178589 );
or ( n11200 , n11197 , n11199 );
buf ( n178592 , n172582 );
xor ( n11202 , n810 , n783 );
buf ( n178594 , n11202 );
nand ( n11204 , n178592 , n178594 );
buf ( n178596 , n11204 );
buf ( n178597 , n178596 );
nand ( n11207 , n11200 , n178597 );
buf ( n178599 , n11207 );
buf ( n178600 , n178599 );
and ( n11210 , n11195 , n178600 );
and ( n11211 , n178575 , n178585 );
or ( n11212 , n11210 , n11211 );
buf ( n178604 , n11212 );
buf ( n178605 , n178604 );
xor ( n11215 , n178558 , n178605 );
xor ( n11216 , n178513 , n178527 );
and ( n178608 , n11216 , n178545 );
and ( n11218 , n178513 , n178527 );
or ( n11219 , n178608 , n11218 );
buf ( n178611 , n11219 );
buf ( n178612 , n178611 );
xor ( n178613 , n11215 , n178612 );
buf ( n178614 , n178613 );
xor ( n11224 , n178441 , n178492 );
and ( n11225 , n11224 , n178548 );
and ( n11226 , n178441 , n178492 );
or ( n11227 , n11225 , n11226 );
buf ( n178619 , n11227 );
xor ( n11229 , n178614 , n178619 );
buf ( n178621 , n11055 );
not ( n11231 , n178621 );
buf ( n178623 , n1578 );
not ( n11233 , n178623 );
or ( n11234 , n11231 , n11233 );
buf ( n178626 , n168743 );
buf ( n178627 , n789 );
buf ( n178628 , n804 );
xor ( n11238 , n178627 , n178628 );
buf ( n178630 , n11238 );
buf ( n178631 , n178630 );
nand ( n11241 , n178626 , n178631 );
buf ( n178633 , n11241 );
buf ( n178634 , n178633 );
nand ( n11244 , n11234 , n178634 );
buf ( n178636 , n11244 );
not ( n11246 , n178636 );
buf ( n178638 , n178142 );
not ( n11248 , n178638 );
buf ( n178640 , n169241 );
not ( n11250 , n178640 );
or ( n11251 , n11248 , n11250 );
buf ( n178643 , n169931 );
buf ( n178644 , n779 );
buf ( n178645 , n814 );
xor ( n11255 , n178644 , n178645 );
buf ( n178647 , n11255 );
buf ( n178648 , n178647 );
nand ( n11258 , n178643 , n178648 );
buf ( n178650 , n11258 );
buf ( n178651 , n178650 );
nand ( n11261 , n11251 , n178651 );
buf ( n178653 , n11261 );
not ( n11263 , n178653 );
or ( n11264 , n11246 , n11263 );
or ( n11265 , n178636 , n178653 );
not ( n11266 , n178463 );
not ( n11267 , n178232 );
or ( n11268 , n11266 , n11267 );
buf ( n178660 , n168867 );
buf ( n178661 , n791 );
buf ( n178662 , n802 );
xor ( n11272 , n178661 , n178662 );
buf ( n178664 , n11272 );
buf ( n178665 , n178664 );
nand ( n11275 , n178660 , n178665 );
buf ( n178667 , n11275 );
nand ( n11277 , n11268 , n178667 );
nand ( n11278 , n11265 , n11277 );
nand ( n11279 , n11264 , n11278 );
buf ( n178671 , n11279 );
buf ( n178672 , n178429 );
not ( n11282 , n178672 );
buf ( n178674 , n168713 );
not ( n11284 , n178674 );
or ( n11285 , n11282 , n11284 );
buf ( n178677 , n169641 );
buf ( n178678 , n787 );
buf ( n178679 , n806 );
xor ( n11289 , n178678 , n178679 );
buf ( n178681 , n11289 );
buf ( n178682 , n178681 );
nand ( n11292 , n178677 , n178682 );
buf ( n178684 , n11292 );
buf ( n178685 , n178684 );
nand ( n11295 , n11285 , n178685 );
buf ( n178687 , n11295 );
buf ( n178688 , n178687 );
not ( n178689 , n178688 );
buf ( n178690 , n178195 );
not ( n11300 , n178690 );
buf ( n178692 , n169411 );
not ( n11302 , n178692 );
or ( n11303 , n11300 , n11302 );
buf ( n178695 , n169417 );
xor ( n11305 , n822 , n771 );
buf ( n178697 , n11305 );
nand ( n11307 , n178695 , n178697 );
buf ( n178699 , n11307 );
buf ( n178700 , n178699 );
nand ( n11310 , n11303 , n178700 );
buf ( n178702 , n11310 );
buf ( n178703 , n178702 );
not ( n11313 , n178703 );
or ( n11314 , n178689 , n11313 );
buf ( n178706 , n178702 );
buf ( n178707 , n178687 );
or ( n11317 , n178706 , n178707 );
buf ( n178709 , n178478 );
not ( n11319 , n178709 );
buf ( n178711 , n169836 );
not ( n11321 , n178711 );
or ( n11322 , n11319 , n11321 );
buf ( n178714 , n169320 );
buf ( n178715 , n777 );
buf ( n178716 , n816 );
xor ( n11326 , n178715 , n178716 );
buf ( n178718 , n11326 );
buf ( n178719 , n178718 );
nand ( n11329 , n178714 , n178719 );
buf ( n178721 , n11329 );
buf ( n178722 , n178721 );
nand ( n11332 , n11322 , n178722 );
buf ( n178724 , n11332 );
buf ( n178725 , n178724 );
nand ( n11335 , n11317 , n178725 );
buf ( n178727 , n11335 );
buf ( n178728 , n178727 );
nand ( n11338 , n11314 , n178728 );
buf ( n178730 , n11338 );
buf ( n178731 , n178730 );
xor ( n11341 , n178671 , n178731 );
buf ( n178733 , n178568 );
not ( n11343 , n178733 );
buf ( n178735 , n1321 );
not ( n11345 , n178735 );
or ( n11346 , n11343 , n11345 );
buf ( n178738 , n168806 );
buf ( n178739 , n774 );
buf ( n178740 , n818 );
xor ( n11350 , n178739 , n178740 );
buf ( n178742 , n11350 );
buf ( n178743 , n178742 );
nand ( n11353 , n178738 , n178743 );
buf ( n178745 , n11353 );
buf ( n178746 , n178745 );
nand ( n11356 , n11346 , n178746 );
buf ( n178748 , n11356 );
buf ( n178749 , n178748 );
buf ( n178750 , n11202 );
not ( n11363 , n178750 );
buf ( n178752 , n171880 );
not ( n11365 , n178752 );
or ( n11366 , n11363 , n11365 );
buf ( n178755 , n170708 );
buf ( n178756 , n782 );
buf ( n178757 , n810 );
xor ( n11370 , n178756 , n178757 );
buf ( n178759 , n11370 );
buf ( n178760 , n178759 );
nand ( n11373 , n178755 , n178760 );
buf ( n178762 , n11373 );
buf ( n178763 , n178762 );
nand ( n11376 , n11366 , n178763 );
buf ( n178765 , n11376 );
buf ( n178766 , n178765 );
xor ( n11379 , n178749 , n178766 );
buf ( n178768 , n11129 );
not ( n11381 , n178768 );
buf ( n178770 , n1907 );
not ( n178771 , n178770 );
or ( n11384 , n11381 , n178771 );
buf ( n178773 , n1535 );
buf ( n178774 , n780 );
buf ( n178775 , n812 );
xor ( n11388 , n178774 , n178775 );
buf ( n178777 , n11388 );
buf ( n178778 , n178777 );
nand ( n11391 , n178773 , n178778 );
buf ( n178780 , n11391 );
buf ( n178781 , n178780 );
nand ( n11394 , n11384 , n178781 );
buf ( n178783 , n11394 );
buf ( n178784 , n178783 );
xor ( n11397 , n11379 , n178784 );
buf ( n178786 , n11397 );
buf ( n178787 , n178786 );
xor ( n11400 , n11341 , n178787 );
buf ( n178789 , n11400 );
xor ( n11402 , n11229 , n178789 );
buf ( n178791 , n11402 );
xor ( n11404 , n11166 , n178791 );
buf ( n178793 , n11404 );
buf ( n178794 , n178793 );
xor ( n178795 , n178409 , n178418 );
xor ( n11408 , n178795 , n178436 );
buf ( n178797 , n11408 );
buf ( n178798 , n178797 );
xor ( n11411 , n178355 , n178372 );
xor ( n11412 , n11411 , n178383 );
buf ( n178801 , n11412 );
buf ( n178802 , n178801 );
xor ( n11415 , n178798 , n178802 );
not ( n11416 , n178469 );
not ( n11417 , n11091 );
not ( n11418 , n11059 );
or ( n11419 , n11417 , n11418 );
or ( n11420 , n11059 , n11091 );
nand ( n11421 , n11419 , n11420 );
not ( n11422 , n11421 );
or ( n11423 , n11416 , n11422 );
or ( n11424 , n11421 , n178469 );
nand ( n11425 , n11423 , n11424 );
buf ( n178814 , n11425 );
and ( n11427 , n11415 , n178814 );
and ( n11428 , n178798 , n178802 );
or ( n11429 , n11427 , n11428 );
buf ( n178818 , n11429 );
buf ( n178819 , n178818 );
xor ( n11432 , n11277 , n178636 );
buf ( n178821 , n11432 );
buf ( n178822 , n178653 );
buf ( n11435 , n178822 );
buf ( n178824 , n11435 );
buf ( n178825 , n178824 );
xnor ( n11438 , n178821 , n178825 );
buf ( n178827 , n11438 );
not ( n11440 , n178827 );
xor ( n11441 , n178575 , n178585 );
xor ( n11442 , n11441 , n178600 );
buf ( n178831 , n11442 );
not ( n11444 , n178831 );
and ( n11445 , n11440 , n11444 );
and ( n11446 , n178827 , n178831 );
nor ( n11447 , n11445 , n11446 );
xor ( n11448 , n178724 , n178702 );
buf ( n178837 , n11448 );
buf ( n178838 , n178687 );
and ( n11451 , n178837 , n178838 );
not ( n11452 , n178837 );
buf ( n178841 , n178687 );
not ( n11454 , n178841 );
buf ( n178843 , n11454 );
buf ( n178844 , n178843 );
and ( n11457 , n11452 , n178844 );
nor ( n11458 , n11451 , n11457 );
buf ( n178847 , n11458 );
and ( n11460 , n11447 , n178847 );
not ( n11461 , n11447 );
buf ( n178850 , n178847 );
not ( n11463 , n178850 );
buf ( n178852 , n11463 );
and ( n11465 , n11461 , n178852 );
nor ( n11466 , n11460 , n11465 );
buf ( n178855 , n11466 );
not ( n11468 , n178855 );
buf ( n178857 , n11468 );
buf ( n178858 , n178857 );
or ( n11471 , n178819 , n178858 );
buf ( n178860 , n177809 );
buf ( n178861 , n830 );
nand ( n11474 , n178860 , n178861 );
buf ( n178863 , n11474 );
buf ( n178864 , n178863 );
not ( n11477 , n178864 );
buf ( n178866 , n798 );
buf ( n178867 , n800 );
and ( n11480 , n178866 , n178867 );
buf ( n178869 , n11480 );
buf ( n178870 , n178869 );
buf ( n178871 , n171551 );
not ( n11484 , n178871 );
buf ( n178873 , n3497 );
not ( n11486 , n178873 );
or ( n11487 , n11484 , n11486 );
buf ( n178876 , n170972 );
buf ( n178877 , n178251 );
nand ( n11490 , n178876 , n178877 );
buf ( n178879 , n11490 );
buf ( n178880 , n178879 );
nand ( n11493 , n11487 , n178880 );
buf ( n178882 , n11493 );
buf ( n178883 , n178882 );
xor ( n11496 , n178870 , n178883 );
buf ( n178885 , n171568 );
not ( n11498 , n178885 );
buf ( n178887 , n169836 );
not ( n11500 , n178887 );
or ( n11501 , n11498 , n11500 );
buf ( n178890 , n169320 );
buf ( n178891 , n178269 );
nand ( n11504 , n178890 , n178891 );
buf ( n178893 , n11504 );
buf ( n178894 , n178893 );
nand ( n11507 , n11501 , n178894 );
buf ( n178896 , n11507 );
buf ( n178897 , n178896 );
and ( n11510 , n11496 , n178897 );
and ( n11511 , n178870 , n178883 );
or ( n11512 , n11510 , n11511 );
buf ( n178901 , n11512 );
buf ( n178902 , n178901 );
not ( n11515 , n178902 );
or ( n11516 , n11477 , n11515 );
buf ( n178905 , n177809 );
not ( n11518 , n178905 );
buf ( n178907 , n830 );
not ( n11520 , n178907 );
buf ( n178909 , n11520 );
buf ( n178910 , n178909 );
nand ( n11523 , n11518 , n178910 );
buf ( n178912 , n11523 );
buf ( n178913 , n178912 );
nand ( n178914 , n11516 , n178913 );
buf ( n178915 , n178914 );
buf ( n178916 , n178915 );
xor ( n11529 , n177810 , n177830 );
xor ( n11530 , n11529 , n177884 );
buf ( n178919 , n11530 );
buf ( n178920 , n178919 );
xor ( n11533 , n178916 , n178920 );
buf ( n178922 , n171309 );
not ( n11535 , n178922 );
buf ( n178924 , n171880 );
not ( n11537 , n178924 );
or ( n178926 , n11535 , n11537 );
buf ( n178927 , n169957 );
buf ( n178928 , n178003 );
nand ( n11541 , n178927 , n178928 );
buf ( n178930 , n11541 );
buf ( n178931 , n178930 );
nand ( n11544 , n178926 , n178931 );
buf ( n178933 , n11544 );
buf ( n178934 , n178933 );
buf ( n178935 , n171218 );
not ( n11548 , n178935 );
buf ( n178937 , n1939 );
not ( n11550 , n178937 );
or ( n11551 , n11548 , n11550 );
buf ( n178940 , n169417 );
buf ( n178941 , n177840 );
nand ( n11554 , n178940 , n178941 );
buf ( n178943 , n11554 );
buf ( n178944 , n178943 );
nand ( n11557 , n11551 , n178944 );
buf ( n178946 , n11557 );
buf ( n178947 , n178946 );
or ( n11560 , n178934 , n178947 );
buf ( n178949 , n171268 );
not ( n178950 , n178949 );
buf ( n178951 , n1907 );
not ( n11564 , n178951 );
or ( n11565 , n178950 , n11564 );
buf ( n178954 , n1534 );
buf ( n178955 , n177932 );
nand ( n11568 , n178954 , n178955 );
buf ( n178957 , n11568 );
buf ( n178958 , n178957 );
nand ( n11571 , n11565 , n178958 );
buf ( n178960 , n11571 );
buf ( n178961 , n178960 );
nand ( n11574 , n11560 , n178961 );
buf ( n178963 , n11574 );
buf ( n178964 , n178946 );
buf ( n178965 , n178933 );
nand ( n11578 , n178964 , n178965 );
buf ( n178967 , n11578 );
nand ( n11580 , n178963 , n178967 );
buf ( n178969 , n11580 );
buf ( n178970 , n171241 );
not ( n11583 , n178970 );
buf ( n178972 , n3764 );
not ( n11585 , n178972 );
or ( n11586 , n11583 , n11585 );
buf ( n178975 , n169247 );
buf ( n178976 , n177894 );
nand ( n11589 , n178975 , n178976 );
buf ( n178978 , n11589 );
buf ( n178979 , n178978 );
nand ( n11592 , n11586 , n178979 );
buf ( n178981 , n11592 );
not ( n11594 , n178981 );
buf ( n178983 , n4114 );
not ( n11596 , n178983 );
buf ( n178985 , n170100 );
not ( n11598 , n178985 );
or ( n11599 , n11596 , n11598 );
buf ( n178988 , n169802 );
buf ( n178989 , n177959 );
nand ( n11602 , n178988 , n178989 );
buf ( n178991 , n11602 );
buf ( n178992 , n178991 );
nand ( n11605 , n11599 , n178992 );
buf ( n178994 , n11605 );
not ( n11607 , n178994 );
or ( n11608 , n11594 , n11607 );
or ( n11609 , n178981 , n178994 );
buf ( n178998 , n171160 );
not ( n11611 , n178998 );
buf ( n179000 , n3683 );
not ( n11613 , n179000 );
or ( n11614 , n11611 , n11613 );
buf ( n179003 , n168559 );
buf ( n179004 , n177797 );
nand ( n11617 , n179003 , n179004 );
buf ( n179006 , n11617 );
buf ( n179007 , n179006 );
nand ( n11620 , n11614 , n179007 );
buf ( n179009 , n11620 );
nand ( n11622 , n11609 , n179009 );
nand ( n11623 , n11608 , n11622 );
buf ( n179012 , n11623 );
or ( n11625 , n178969 , n179012 );
buf ( n179014 , n171291 );
not ( n11627 , n179014 );
buf ( n179016 , n168648 );
not ( n11629 , n179016 );
or ( n11630 , n11627 , n11629 );
buf ( n179019 , n177920 );
not ( n11632 , n179019 );
buf ( n179021 , n171296 );
nand ( n11634 , n11632 , n179021 );
buf ( n179023 , n11634 );
buf ( n179024 , n179023 );
nand ( n11637 , n11630 , n179024 );
buf ( n179026 , n11637 );
buf ( n179027 , n179026 );
buf ( n179028 , n171365 );
not ( n11641 , n179028 );
buf ( n179030 , n169545 );
not ( n11643 , n179030 );
or ( n11644 , n11641 , n11643 );
buf ( n179033 , n168619 );
buf ( n179034 , n177979 );
nand ( n11647 , n179033 , n179034 );
buf ( n179036 , n11647 );
buf ( n179037 , n179036 );
nand ( n11650 , n11644 , n179037 );
buf ( n179039 , n11650 );
buf ( n179040 , n179039 );
xor ( n11653 , n179027 , n179040 );
buf ( n179042 , n171335 );
not ( n11655 , n179042 );
buf ( n179044 , n4337 );
not ( n11657 , n179044 );
or ( n11658 , n11655 , n11657 );
buf ( n179047 , n168684 );
buf ( n179048 , n177862 );
nand ( n11661 , n179047 , n179048 );
buf ( n179050 , n11661 );
buf ( n179051 , n179050 );
nand ( n11664 , n11658 , n179051 );
buf ( n179053 , n11664 );
buf ( n179054 , n179053 );
and ( n11667 , n11653 , n179054 );
and ( n11668 , n179027 , n179040 );
or ( n11669 , n11667 , n11668 );
buf ( n179058 , n11669 );
buf ( n179059 , n179058 );
nand ( n179060 , n11625 , n179059 );
buf ( n179061 , n179060 );
buf ( n179062 , n179061 );
buf ( n179063 , n11580 );
buf ( n179064 , n11623 );
nand ( n11680 , n179063 , n179064 );
buf ( n179066 , n11680 );
buf ( n179067 , n179066 );
nand ( n11683 , n179062 , n179067 );
buf ( n179069 , n11683 );
buf ( n179070 , n179069 );
and ( n11686 , n11533 , n179070 );
and ( n11687 , n178916 , n178920 );
or ( n11688 , n11686 , n11687 );
buf ( n179074 , n11688 );
buf ( n179075 , n179074 );
nand ( n11691 , n11471 , n179075 );
buf ( n179077 , n11691 );
buf ( n179078 , n179077 );
buf ( n179079 , n178857 );
buf ( n179080 , n178818 );
nand ( n11696 , n179079 , n179080 );
buf ( n179082 , n11696 );
buf ( n179083 , n179082 );
nand ( n11699 , n179078 , n179083 );
buf ( n179085 , n11699 );
buf ( n179086 , n179085 );
not ( n11702 , n178831 );
nand ( n11703 , n11702 , n178827 );
not ( n11704 , n11703 );
not ( n11705 , n178847 );
or ( n11706 , n11704 , n11705 );
buf ( n179092 , n178827 );
not ( n11708 , n179092 );
buf ( n179094 , n178831 );
nand ( n11710 , n11708 , n179094 );
buf ( n179096 , n11710 );
nand ( n11712 , n11706 , n179096 );
buf ( n179098 , n11712 );
not ( n11714 , n178664 );
not ( n11715 , n178232 );
or ( n11716 , n11714 , n11715 );
buf ( n179102 , n168867 );
buf ( n179103 , n790 );
buf ( n179104 , n802 );
xor ( n11720 , n179103 , n179104 );
buf ( n179106 , n11720 );
buf ( n179107 , n179106 );
nand ( n11723 , n179102 , n179107 );
buf ( n179109 , n11723 );
nand ( n11725 , n11716 , n179109 );
buf ( n179111 , n1578 );
not ( n11727 , n179111 );
buf ( n179113 , n11727 );
buf ( n179114 , n179113 );
not ( n11730 , n179114 );
buf ( n179116 , n178630 );
not ( n11732 , n179116 );
buf ( n179118 , n11732 );
buf ( n179119 , n179118 );
not ( n11735 , n179119 );
and ( n11736 , n11730 , n11735 );
buf ( n179122 , n168743 );
xor ( n11738 , n804 , n788 );
buf ( n179124 , n11738 );
and ( n11740 , n179122 , n179124 );
buf ( n179126 , n11740 );
buf ( n179127 , n179126 );
nor ( n11743 , n11736 , n179127 );
buf ( n179129 , n11743 );
not ( n11745 , n179129 );
xor ( n11746 , n11725 , n11745 );
buf ( n179132 , n178718 );
not ( n11748 , n179132 );
buf ( n179134 , n169836 );
not ( n11750 , n179134 );
or ( n11751 , n11748 , n11750 );
buf ( n179137 , n169320 );
buf ( n179138 , n776 );
buf ( n179139 , n816 );
xor ( n11755 , n179138 , n179139 );
buf ( n179141 , n11755 );
buf ( n179142 , n179141 );
nand ( n11758 , n179137 , n179142 );
buf ( n179144 , n11758 );
buf ( n179145 , n179144 );
nand ( n11761 , n11751 , n179145 );
buf ( n179147 , n11761 );
xnor ( n11763 , n11746 , n179147 );
not ( n11764 , n10362 );
not ( n11765 , n3497 );
or ( n11766 , n11764 , n11765 );
buf ( n179152 , n170972 );
xor ( n11768 , n800 , n792 );
buf ( n179154 , n11768 );
nand ( n11770 , n179152 , n179154 );
buf ( n179156 , n11770 );
nand ( n11772 , n11766 , n179156 );
buf ( n179158 , n794 );
buf ( n179159 , n800 );
and ( n11775 , n179158 , n179159 );
buf ( n179161 , n11775 );
or ( n11777 , n11772 , n179161 );
buf ( n179163 , n11772 );
buf ( n179164 , n179161 );
nand ( n11780 , n179163 , n179164 );
buf ( n179166 , n11780 );
nand ( n11782 , n11777 , n179166 );
buf ( n179168 , n178647 );
not ( n11784 , n179168 );
buf ( n179170 , n171013 );
not ( n11786 , n179170 );
or ( n11787 , n11784 , n11786 );
buf ( n179173 , n169250 );
buf ( n179174 , n778 );
buf ( n179175 , n814 );
xor ( n11791 , n179174 , n179175 );
buf ( n179177 , n11791 );
buf ( n179178 , n179177 );
nand ( n11794 , n179173 , n179178 );
buf ( n179180 , n11794 );
buf ( n179181 , n179180 );
nand ( n11797 , n11787 , n179181 );
buf ( n179183 , n11797 );
xor ( n11799 , n11782 , n179183 );
xor ( n11800 , n11763 , n11799 );
buf ( n179186 , n2202 );
not ( n11802 , n179186 );
buf ( n179188 , n169681 );
not ( n11804 , n179188 );
or ( n11805 , n11802 , n11804 );
buf ( n179191 , n826 );
nand ( n11807 , n11805 , n179191 );
buf ( n179193 , n11807 );
buf ( n179194 , n178538 );
not ( n11810 , n179194 );
buf ( n179196 , n2108 );
not ( n11812 , n179196 );
or ( n11813 , n11810 , n11812 );
buf ( n179199 , n168656 );
buf ( n179200 , n772 );
buf ( n179201 , n820 );
xor ( n11817 , n179200 , n179201 );
buf ( n179203 , n11817 );
buf ( n179204 , n179203 );
nand ( n11820 , n179199 , n179204 );
buf ( n179206 , n11820 );
buf ( n179207 , n179206 );
nand ( n11823 , n11813 , n179207 );
buf ( n179209 , n11823 );
xnor ( n11825 , n179193 , n179209 );
buf ( n179211 , n11825 );
buf ( n179212 , n11115 );
not ( n11828 , n179212 );
buf ( n179214 , n170100 );
not ( n11830 , n179214 );
or ( n11831 , n11828 , n11830 );
buf ( n179217 , n175664 );
buf ( n179218 , n768 );
buf ( n179219 , n824 );
xor ( n11835 , n179218 , n179219 );
buf ( n179221 , n11835 );
buf ( n179222 , n179221 );
nand ( n11838 , n179217 , n179222 );
buf ( n179224 , n11838 );
buf ( n179225 , n179224 );
nand ( n11841 , n11831 , n179225 );
buf ( n179227 , n11841 );
buf ( n179228 , n179227 );
and ( n11844 , n179211 , n179228 );
not ( n11845 , n179211 );
buf ( n179231 , n179227 );
not ( n11847 , n179231 );
buf ( n179233 , n11847 );
buf ( n179234 , n179233 );
and ( n11850 , n11845 , n179234 );
or ( n11851 , n11844 , n11850 );
buf ( n179237 , n11851 );
xor ( n11853 , n11800 , n179237 );
buf ( n179239 , n11853 );
xor ( n11855 , n179098 , n179239 );
xor ( n11856 , n177751 , n177769 );
and ( n11857 , n11856 , n177790 );
and ( n11858 , n177751 , n177769 );
or ( n11859 , n11857 , n11858 );
buf ( n179245 , n11859 );
buf ( n179246 , n179245 );
buf ( n179247 , n11189 );
not ( n11863 , n179247 );
buf ( n179249 , n169545 );
not ( n11865 , n179249 );
or ( n11866 , n11863 , n11865 );
buf ( n179252 , n168619 );
buf ( n179253 , n784 );
buf ( n179254 , n808 );
xor ( n11870 , n179253 , n179254 );
buf ( n179256 , n11870 );
buf ( n179257 , n179256 );
nand ( n11873 , n179252 , n179257 );
buf ( n179259 , n11873 );
buf ( n179260 , n179259 );
nand ( n11876 , n11866 , n179260 );
buf ( n179262 , n11876 );
buf ( n179263 , n11305 );
not ( n11879 , n179263 );
buf ( n179265 , n1939 );
not ( n11881 , n179265 );
or ( n11882 , n11879 , n11881 );
buf ( n179268 , n169417 );
xor ( n11884 , n822 , n770 );
buf ( n179270 , n11884 );
nand ( n11886 , n179268 , n179270 );
buf ( n179272 , n11886 );
buf ( n179273 , n179272 );
nand ( n11889 , n11882 , n179273 );
buf ( n179275 , n11889 );
xor ( n11891 , n179262 , n179275 );
buf ( n179277 , n178681 );
not ( n11893 , n179277 );
buf ( n179279 , n168713 );
not ( n11895 , n179279 );
or ( n11896 , n11893 , n11895 );
buf ( n179282 , n169641 );
xor ( n11898 , n806 , n786 );
buf ( n179284 , n11898 );
nand ( n11900 , n179282 , n179284 );
buf ( n179286 , n11900 );
buf ( n179287 , n179286 );
nand ( n11903 , n11896 , n179287 );
buf ( n179289 , n11903 );
xor ( n11905 , n11891 , n179289 );
buf ( n179291 , n11905 );
xor ( n11907 , n179246 , n179291 );
xor ( n11908 , n178325 , n178340 );
and ( n11909 , n11908 , n178388 );
and ( n11910 , n178325 , n178340 );
or ( n11911 , n11909 , n11910 );
buf ( n179297 , n11911 );
buf ( n179298 , n179297 );
xor ( n11914 , n11907 , n179298 );
buf ( n179300 , n11914 );
buf ( n179301 , n179300 );
xor ( n11917 , n11855 , n179301 );
buf ( n179303 , n11917 );
buf ( n179304 , n179303 );
xor ( n11920 , n179086 , n179304 );
xor ( n11921 , n177793 , n177889 );
xor ( n11922 , n11921 , n178104 );
buf ( n179308 , n11922 );
buf ( n179309 , n179308 );
xor ( n11925 , n178312 , n178391 );
xor ( n11926 , n11925 , n178551 );
buf ( n179312 , n11926 );
buf ( n179313 , n179312 );
or ( n11929 , n179309 , n179313 );
buf ( n179315 , n171382 );
not ( n11931 , n179315 );
buf ( n179317 , n169635 );
not ( n11933 , n179317 );
or ( n11934 , n11931 , n11933 );
buf ( n179320 , n2823 );
buf ( n179321 , n178031 );
nand ( n11937 , n179320 , n179321 );
buf ( n179323 , n11937 );
buf ( n179324 , n179323 );
nand ( n11940 , n11934 , n179324 );
buf ( n179326 , n11940 );
buf ( n179327 , n179326 );
buf ( n179328 , n171400 );
not ( n11944 , n179328 );
buf ( n179330 , n1321 );
not ( n11946 , n179330 );
or ( n11947 , n11944 , n11946 );
buf ( n179333 , n168806 );
buf ( n179334 , n178074 );
nand ( n11950 , n179333 , n179334 );
buf ( n179336 , n11950 );
buf ( n179337 , n179336 );
nand ( n11953 , n11947 , n179337 );
buf ( n179339 , n11953 );
buf ( n179340 , n179339 );
xor ( n11956 , n179327 , n179340 );
buf ( n179342 , n171516 );
not ( n11958 , n179342 );
buf ( n179344 , n168750 );
not ( n11960 , n179344 );
or ( n11961 , n11958 , n11960 );
buf ( n179347 , n168838 );
buf ( n179348 , n178052 );
nand ( n11964 , n179347 , n179348 );
buf ( n179350 , n11964 );
buf ( n179351 , n179350 );
nand ( n11967 , n11961 , n179351 );
buf ( n179353 , n11967 );
buf ( n179354 , n179353 );
and ( n11970 , n11956 , n179354 );
and ( n11971 , n179327 , n179340 );
or ( n11972 , n11970 , n11971 );
buf ( n179358 , n11972 );
buf ( n179359 , n179358 );
xor ( n11975 , n178247 , n178264 );
xor ( n11976 , n11975 , n178286 );
buf ( n179362 , n11976 );
buf ( n179363 , n179362 );
xor ( n11982 , n179359 , n179363 );
xor ( n11983 , n10525 , n177910 );
xor ( n11984 , n11983 , n177948 );
buf ( n179367 , n11984 );
and ( n11986 , n11982 , n179367 );
and ( n179369 , n179359 , n179363 );
or ( n11988 , n11986 , n179369 );
buf ( n179371 , n11988 );
not ( n11990 , n179371 );
buf ( n179373 , n11990 );
not ( n11992 , n179373 );
buf ( n179375 , n177954 );
buf ( n179376 , n10628 );
and ( n11995 , n179375 , n179376 );
not ( n11996 , n179375 );
buf ( n179379 , n10628 );
not ( n11998 , n179379 );
buf ( n179381 , n11998 );
buf ( n179382 , n179381 );
and ( n12001 , n11996 , n179382 );
nor ( n12002 , n11995 , n12001 );
buf ( n179385 , n12002 );
buf ( n179386 , n179385 );
buf ( n179387 , n178092 );
not ( n12006 , n179387 );
buf ( n179389 , n12006 );
buf ( n179390 , n179389 );
and ( n179391 , n179386 , n179390 );
not ( n12010 , n179386 );
buf ( n179393 , n178092 );
and ( n12012 , n12010 , n179393 );
nor ( n12013 , n179391 , n12012 );
buf ( n179396 , n12013 );
buf ( n179397 , n179396 );
not ( n12016 , n179397 );
or ( n12017 , n11992 , n12016 );
xor ( n12018 , n177836 , n177857 );
xor ( n12019 , n12018 , n177879 );
buf ( n179402 , n12019 );
buf ( n179403 , n179402 );
xor ( n12022 , n178048 , n178069 );
xor ( n12023 , n12022 , n178088 );
buf ( n179406 , n12023 );
buf ( n179407 , n179406 );
xor ( n12026 , n179403 , n179407 );
buf ( n179409 , n178019 );
not ( n12028 , n179409 );
buf ( n179411 , n12028 );
xor ( n12030 , n177998 , n179411 );
xnor ( n12031 , n12030 , n177975 );
buf ( n179414 , n12031 );
and ( n12033 , n12026 , n179414 );
and ( n12034 , n179403 , n179407 );
or ( n12035 , n12033 , n12034 );
buf ( n179418 , n12035 );
buf ( n179419 , n179418 );
nand ( n12038 , n12017 , n179419 );
buf ( n179421 , n12038 );
buf ( n179422 , n179421 );
buf ( n179423 , n179396 );
not ( n12042 , n179423 );
buf ( n179425 , n179371 );
nand ( n12044 , n12042 , n179425 );
buf ( n179427 , n12044 );
buf ( n179428 , n179427 );
nand ( n12047 , n179422 , n179428 );
buf ( n179430 , n12047 );
buf ( n179431 , n179430 );
nand ( n12050 , n11929 , n179431 );
buf ( n179433 , n12050 );
buf ( n179434 , n179433 );
buf ( n179435 , n179312 );
buf ( n179436 , n179308 );
nand ( n12055 , n179435 , n179436 );
buf ( n179438 , n12055 );
buf ( n179439 , n179438 );
nand ( n12058 , n179434 , n179439 );
buf ( n179441 , n12058 );
buf ( n179442 , n179441 );
xor ( n12061 , n11920 , n179442 );
buf ( n179444 , n12061 );
buf ( n179445 , n179444 );
xor ( n12064 , n178794 , n179445 );
buf ( n179447 , n178290 );
not ( n12066 , n179447 );
buf ( n179449 , n178151 );
not ( n12068 , n179449 );
and ( n12069 , n12066 , n12068 );
buf ( n179452 , n178290 );
buf ( n179453 , n178300 );
and ( n12072 , n179452 , n179453 );
nor ( n12073 , n12069 , n12072 );
buf ( n179456 , n12073 );
buf ( n179457 , n179456 );
buf ( n179458 , n178305 );
buf ( n12077 , n179458 );
buf ( n179460 , n12077 );
buf ( n179461 , n179460 );
xnor ( n12080 , n179457 , n179461 );
buf ( n179463 , n12080 );
buf ( n179464 , n179463 );
xor ( n12083 , n178798 , n178802 );
xor ( n12084 , n12083 , n178814 );
buf ( n179467 , n12084 );
buf ( n179468 , n179467 );
xor ( n12087 , n179464 , n179468 );
xor ( n12088 , n178916 , n178920 );
xor ( n12089 , n12088 , n179070 );
buf ( n179472 , n12089 );
buf ( n179473 , n179472 );
and ( n12092 , n12087 , n179473 );
and ( n12093 , n179464 , n179468 );
or ( n12094 , n12092 , n12093 );
buf ( n179477 , n12094 );
buf ( n179478 , n179477 );
xor ( n12097 , n178818 , n11466 );
xnor ( n12098 , n12097 , n179074 );
buf ( n179481 , n12098 );
xor ( n12100 , n179478 , n179481 );
buf ( n179483 , n178901 );
not ( n12102 , n179483 );
buf ( n179485 , n177809 );
not ( n12104 , n179485 );
buf ( n179487 , n178909 );
not ( n12106 , n179487 );
and ( n12107 , n12104 , n12106 );
buf ( n179490 , n177809 );
buf ( n179491 , n178909 );
and ( n12110 , n179490 , n179491 );
nor ( n12111 , n12107 , n12110 );
buf ( n179494 , n12111 );
buf ( n179495 , n179494 );
not ( n12114 , n179495 );
and ( n12115 , n12102 , n12114 );
buf ( n179498 , n178901 );
buf ( n179499 , n179494 );
and ( n12118 , n179498 , n179499 );
nor ( n12119 , n12115 , n12118 );
buf ( n179502 , n12119 );
buf ( n179503 , n179502 );
not ( n12122 , n179503 );
buf ( n179505 , n12122 );
buf ( n179506 , n179505 );
not ( n12125 , n179506 );
xor ( n12126 , n179027 , n179040 );
xor ( n12127 , n12126 , n179054 );
buf ( n179510 , n12127 );
buf ( n12129 , n179510 );
buf ( n179512 , n12129 );
buf ( n179513 , n178946 );
not ( n12132 , n179513 );
buf ( n179515 , n178960 );
not ( n12134 , n179515 );
buf ( n179517 , n12134 );
buf ( n179518 , n179517 );
not ( n12137 , n179518 );
or ( n12138 , n12132 , n12137 );
buf ( n179521 , n179517 );
buf ( n179522 , n178946 );
or ( n12141 , n179521 , n179522 );
nand ( n12142 , n12138 , n12141 );
buf ( n179525 , n12142 );
xor ( n12144 , n179525 , n178933 );
buf ( n179527 , n12144 );
or ( n12146 , n179512 , n179527 );
xnor ( n179529 , n178981 , n179009 );
not ( n12148 , n178994 );
and ( n12149 , n179529 , n12148 );
not ( n12150 , n179529 );
and ( n12151 , n12150 , n178994 );
nor ( n179534 , n12149 , n12151 );
buf ( n179535 , n179534 );
nand ( n12154 , n12146 , n179535 );
buf ( n179537 , n12154 );
buf ( n179538 , n179537 );
buf ( n179539 , n12144 );
buf ( n179540 , n12129 );
nand ( n12159 , n179539 , n179540 );
buf ( n179542 , n12159 );
buf ( n179543 , n179542 );
nand ( n12162 , n179538 , n179543 );
buf ( n179545 , n12162 );
buf ( n179546 , n179545 );
not ( n12165 , n179546 );
or ( n12166 , n12125 , n12165 );
buf ( n179549 , n179502 );
not ( n12168 , n179549 );
buf ( n179551 , n179545 );
not ( n12170 , n179551 );
buf ( n179553 , n12170 );
buf ( n179554 , n179553 );
not ( n12173 , n179554 );
or ( n179556 , n12168 , n12173 );
or ( n12175 , n3844 , n3831 );
not ( n12176 , n12175 );
not ( n12177 , n171342 );
or ( n12178 , n12176 , n12177 );
nand ( n12179 , n3850 , n3831 );
nand ( n179562 , n12178 , n12179 );
buf ( n179563 , n179562 );
not ( n12182 , n179563 );
xor ( n12183 , n179327 , n179340 );
xor ( n12184 , n12183 , n179354 );
buf ( n179567 , n12184 );
buf ( n179568 , n179567 );
not ( n12187 , n179568 );
or ( n12188 , n12182 , n12187 );
buf ( n179571 , n179562 );
buf ( n179572 , n179567 );
or ( n12191 , n179571 , n179572 );
xor ( n12192 , n178870 , n178883 );
xor ( n12193 , n12192 , n178897 );
buf ( n179576 , n12193 );
buf ( n179577 , n179576 );
nand ( n12196 , n12191 , n179577 );
buf ( n179579 , n12196 );
buf ( n179580 , n179579 );
nand ( n12199 , n12188 , n179580 );
buf ( n179582 , n12199 );
buf ( n179583 , n179582 );
nand ( n12202 , n179556 , n179583 );
buf ( n179585 , n12202 );
buf ( n179586 , n179585 );
nand ( n12205 , n12166 , n179586 );
buf ( n179588 , n12205 );
not ( n12207 , n179588 );
buf ( n179590 , n178909 );
not ( n12209 , n179590 );
buf ( n179592 , n171500 );
not ( n12211 , n179592 );
buf ( n179594 , n168861 );
not ( n12213 , n179594 );
or ( n12214 , n12211 , n12213 );
buf ( n179597 , n168870 );
buf ( n179598 , n178215 );
nand ( n12217 , n179597 , n179598 );
buf ( n179600 , n12217 );
buf ( n179601 , n179600 );
nand ( n12220 , n12214 , n179601 );
buf ( n179603 , n12220 );
buf ( n179604 , n179603 );
not ( n12223 , n179604 );
buf ( n179606 , n12223 );
buf ( n179607 , n179606 );
not ( n12226 , n179607 );
or ( n12227 , n12209 , n12226 );
xor ( n12228 , n171133 , n171146 );
and ( n12229 , n12228 , n171167 );
and ( n12230 , n171133 , n171146 );
or ( n12231 , n12229 , n12230 );
buf ( n179614 , n12231 );
buf ( n179615 , n179614 );
nand ( n12234 , n12227 , n179615 );
buf ( n179617 , n12234 );
buf ( n179618 , n179617 );
buf ( n179619 , n179603 );
buf ( n179620 , n830 );
nand ( n12239 , n179619 , n179620 );
buf ( n179622 , n12239 );
buf ( n179623 , n179622 );
nand ( n12242 , n179618 , n179623 );
buf ( n179625 , n12242 );
buf ( n179626 , n179625 );
xor ( n12245 , n171558 , n171575 );
and ( n12246 , n12245 , n171590 );
and ( n12247 , n171558 , n171575 );
or ( n12248 , n12246 , n12247 );
buf ( n179631 , n12248 );
buf ( n179632 , n179631 );
xor ( n12251 , n171372 , n171389 );
and ( n12252 , n12251 , n171407 );
and ( n12253 , n171372 , n171389 );
or ( n12254 , n12252 , n12253 );
buf ( n179637 , n12254 );
buf ( n179638 , n179637 );
xor ( n12257 , n179632 , n179638 );
buf ( n179640 , n171250 );
not ( n12259 , n179640 );
buf ( n179642 , n171224 );
not ( n12261 , n179642 );
buf ( n179644 , n12261 );
buf ( n179645 , n179644 );
not ( n12264 , n179645 );
or ( n12265 , n12259 , n12264 );
buf ( n179648 , n171274 );
nand ( n12267 , n12265 , n179648 );
buf ( n179650 , n12267 );
buf ( n179651 , n179650 );
buf ( n179652 , n171224 );
buf ( n179653 , n171247 );
nand ( n12272 , n179652 , n179653 );
buf ( n179655 , n12272 );
buf ( n179656 , n179655 );
nand ( n12275 , n179651 , n179656 );
buf ( n179658 , n12275 );
buf ( n179659 , n179658 );
and ( n12278 , n12257 , n179659 );
and ( n12279 , n179632 , n179638 );
or ( n12280 , n12278 , n12279 );
buf ( n179663 , n12280 );
buf ( n179664 , n179663 );
xor ( n12283 , n179626 , n179664 );
xor ( n12284 , n11623 , n11580 );
xor ( n12285 , n12284 , n179058 );
buf ( n179668 , n12285 );
and ( n12287 , n12283 , n179668 );
and ( n12288 , n179626 , n179664 );
or ( n12289 , n12287 , n12288 );
buf ( n179672 , n12289 );
not ( n12291 , n179672 );
or ( n12292 , n12207 , n12291 );
buf ( n179675 , n179396 );
not ( n12294 , n179675 );
buf ( n179677 , n179418 );
not ( n12296 , n179677 );
or ( n12297 , n12294 , n12296 );
buf ( n179680 , n179418 );
buf ( n179681 , n179396 );
or ( n12300 , n179680 , n179681 );
nand ( n12301 , n12297 , n12300 );
buf ( n179684 , n12301 );
buf ( n179685 , n179684 );
buf ( n12304 , n179371 );
buf ( n179687 , n12304 );
and ( n12306 , n179685 , n179687 );
not ( n12307 , n179685 );
not ( n12308 , n12304 );
buf ( n179691 , n12308 );
and ( n12310 , n12307 , n179691 );
nor ( n12311 , n12306 , n12310 );
buf ( n179694 , n12311 );
not ( n12316 , n179694 );
nor ( n12317 , n179588 , n179672 );
or ( n12318 , n12316 , n12317 );
nand ( n12319 , n12292 , n12318 );
buf ( n179699 , n12319 );
and ( n179700 , n12100 , n179699 );
and ( n12322 , n179478 , n179481 );
or ( n12323 , n179700 , n12322 );
buf ( n179703 , n12323 );
buf ( n179704 , n179703 );
xor ( n12326 , n12064 , n179704 );
buf ( n179706 , n12326 );
buf ( n179707 , n179308 );
not ( n12329 , n179707 );
buf ( n179709 , n12329 );
buf ( n179710 , n179709 );
not ( n12332 , n179710 );
buf ( n179712 , n179430 );
not ( n12334 , n179712 );
and ( n12335 , n12332 , n12334 );
buf ( n179715 , n179430 );
buf ( n179716 , n179709 );
and ( n179717 , n179715 , n179716 );
nor ( n12339 , n12335 , n179717 );
buf ( n179719 , n12339 );
not ( n12341 , n179719 );
xor ( n12342 , n179312 , n12341 );
buf ( n179722 , n12342 );
xor ( n12344 , n179359 , n179363 );
xor ( n12345 , n12344 , n179367 );
buf ( n179725 , n12345 );
xor ( n12347 , n179403 , n179407 );
xor ( n179727 , n12347 , n179414 );
buf ( n179728 , n179727 );
xor ( n12350 , n179725 , n179728 );
buf ( n179730 , n171284 );
not ( n12352 , n179730 );
buf ( n179732 , n3880 );
not ( n12354 , n179732 );
or ( n12355 , n12352 , n12354 );
buf ( n179735 , n171409 );
nand ( n12357 , n12355 , n179735 );
buf ( n179737 , n12357 );
buf ( n179738 , n179737 );
buf ( n179739 , n171284 );
not ( n12361 , n179739 );
buf ( n179741 , n3883 );
nand ( n12363 , n12361 , n179741 );
buf ( n179743 , n12363 );
buf ( n179744 , n179743 );
nand ( n12366 , n179738 , n179744 );
buf ( n179746 , n12366 );
buf ( n179747 , n179746 );
buf ( n179748 , n179603 );
not ( n12370 , n179748 );
buf ( n179750 , n178909 );
not ( n12372 , n179750 );
and ( n12373 , n12370 , n12372 );
buf ( n179753 , n179603 );
buf ( n179754 , n178909 );
and ( n12376 , n179753 , n179754 );
nor ( n12377 , n12373 , n12376 );
buf ( n179757 , n12377 );
xnor ( n12379 , n179614 , n179757 );
buf ( n179759 , n12379 );
or ( n12381 , n179747 , n179759 );
xor ( n12382 , n179632 , n179638 );
xor ( n12383 , n12382 , n179659 );
buf ( n179763 , n12383 );
buf ( n179764 , n179763 );
nand ( n12386 , n12381 , n179764 );
buf ( n179766 , n12386 );
buf ( n179767 , n179766 );
buf ( n179768 , n179746 );
buf ( n179769 , n12379 );
nand ( n12391 , n179768 , n179769 );
buf ( n179771 , n12391 );
buf ( n179772 , n179771 );
nand ( n12394 , n179767 , n179772 );
buf ( n179774 , n12394 );
and ( n12396 , n12350 , n179774 );
and ( n12397 , n179725 , n179728 );
or ( n12398 , n12396 , n12397 );
xor ( n12399 , n179464 , n179468 );
xor ( n12400 , n12399 , n179473 );
buf ( n179780 , n12400 );
xor ( n12402 , n12398 , n179780 );
xor ( n12403 , n179626 , n179664 );
xor ( n12404 , n12403 , n179668 );
buf ( n179784 , n12404 );
not ( n12406 , n179784 );
buf ( n179786 , n171522 );
not ( n12408 , n179786 );
buf ( n179788 , n12408 );
buf ( n179789 , n179788 );
not ( n12411 , n179789 );
buf ( n179791 , n171528 );
not ( n12413 , n179791 );
or ( n12414 , n12411 , n12413 );
buf ( n179794 , n171506 );
nand ( n12416 , n12414 , n179794 );
buf ( n179796 , n12416 );
buf ( n179797 , n179796 );
buf ( n179798 , n171533 );
buf ( n179799 , n171522 );
nand ( n12421 , n179798 , n179799 );
buf ( n179801 , n12421 );
buf ( n179802 , n179801 );
nand ( n12424 , n179797 , n179802 );
buf ( n179804 , n12424 );
not ( n12426 , n179804 );
buf ( n179806 , n171169 );
not ( n12428 , n179806 );
buf ( n179808 , n171184 );
not ( n12430 , n179808 );
or ( n12431 , n12428 , n12430 );
buf ( n179811 , n171184 );
buf ( n179812 , n171169 );
or ( n12434 , n179811 , n179812 );
buf ( n179814 , n12434 );
buf ( n179815 , n179814 );
buf ( n179816 , n171191 );
nand ( n12438 , n179815 , n179816 );
buf ( n179818 , n12438 );
buf ( n179819 , n179818 );
nand ( n12441 , n12431 , n179819 );
buf ( n179821 , n12441 );
not ( n12443 , n179821 );
or ( n12444 , n12426 , n12443 );
not ( n12445 , n179804 );
not ( n12446 , n12445 );
not ( n12447 , n179821 );
not ( n12448 , n12447 );
or ( n12449 , n12446 , n12448 );
buf ( n179829 , n171442 );
not ( n12451 , n179829 );
buf ( n179831 , n12451 );
buf ( n179832 , n179831 );
not ( n12454 , n179832 );
buf ( n179834 , n171459 );
not ( n12456 , n179834 );
or ( n12457 , n12454 , n12456 );
buf ( n179837 , n171465 );
nand ( n12459 , n12457 , n179837 );
buf ( n179839 , n12459 );
buf ( n179840 , n179839 );
buf ( n179841 , n171442 );
buf ( n179842 , n171456 );
nand ( n12464 , n179841 , n179842 );
buf ( n179844 , n12464 );
buf ( n179845 , n179844 );
nand ( n12467 , n179840 , n179845 );
buf ( n179847 , n12467 );
nand ( n12469 , n12449 , n179847 );
nand ( n12470 , n12444 , n12469 );
not ( n12471 , n12470 );
or ( n12472 , n12406 , n12471 );
nor ( n12473 , n179784 , n12470 );
buf ( n179853 , n179502 );
not ( n12475 , n179853 );
buf ( n179855 , n179582 );
not ( n179856 , n179855 );
or ( n12478 , n12475 , n179856 );
buf ( n179858 , n179582 );
buf ( n179859 , n179502 );
or ( n12481 , n179858 , n179859 );
nand ( n179861 , n12478 , n12481 );
buf ( n179862 , n179861 );
buf ( n179863 , n179862 );
buf ( n179864 , n179545 );
buf ( n12486 , n179864 );
buf ( n179866 , n12486 );
buf ( n179867 , n179866 );
xnor ( n12489 , n179863 , n179867 );
buf ( n179869 , n12489 );
or ( n12491 , n12473 , n179869 );
nand ( n12492 , n12472 , n12491 );
and ( n12493 , n12402 , n12492 );
and ( n12494 , n12398 , n179780 );
or ( n12495 , n12493 , n12494 );
buf ( n179875 , n12495 );
xor ( n12497 , n179722 , n179875 );
xor ( n12498 , n179478 , n179481 );
xor ( n179878 , n12498 , n179699 );
buf ( n179879 , n179878 );
buf ( n179880 , n179879 );
and ( n12502 , n12497 , n179880 );
and ( n12503 , n179722 , n179875 );
or ( n12504 , n12502 , n12503 );
buf ( n179884 , n12504 );
xor ( n12506 , n179706 , n179884 );
not ( n12507 , n12506 );
xor ( n12508 , n12445 , n179821 );
not ( n179888 , n179847 );
xnor ( n12510 , n12508 , n179888 );
not ( n12511 , n12510 );
buf ( n179891 , n171127 );
not ( n12513 , n179891 );
buf ( n179893 , n171194 );
not ( n12515 , n179893 );
or ( n12516 , n12513 , n12515 );
buf ( n179896 , n171204 );
nand ( n12518 , n12516 , n179896 );
buf ( n179898 , n12518 );
buf ( n179899 , n171197 );
buf ( n179900 , n171124 );
nand ( n12522 , n179899 , n179900 );
buf ( n179902 , n12522 );
nand ( n12524 , n179898 , n179902 );
not ( n12525 , n12524 );
not ( n12526 , n12525 );
or ( n12527 , n12511 , n12526 );
xor ( n12528 , n179763 , n12379 );
xor ( n12529 , n12528 , n179746 );
nand ( n12530 , n12527 , n12529 );
buf ( n179910 , n12530 );
not ( n12532 , n12510 );
nand ( n12533 , n12524 , n12532 );
buf ( n179913 , n12533 );
nand ( n12535 , n179910 , n179913 );
buf ( n179915 , n12535 );
buf ( n179916 , n179915 );
not ( n12538 , n179916 );
xor ( n12539 , n179725 , n179728 );
xor ( n12540 , n12539 , n179774 );
buf ( n12541 , n12540 );
buf ( n179921 , n12541 );
not ( n12543 , n179921 );
buf ( n179923 , n12543 );
buf ( n179924 , n179923 );
not ( n12546 , n12148 );
not ( n12547 , n179529 );
and ( n12548 , n12546 , n12547 );
and ( n12549 , n12148 , n179529 );
nor ( n12550 , n12548 , n12549 );
not ( n12551 , n12550 );
not ( n12552 , n179510 );
not ( n12553 , n12552 );
or ( n12554 , n12551 , n12553 );
or ( n12555 , n12550 , n12552 );
nand ( n12556 , n12554 , n12555 );
buf ( n179936 , n12556 );
buf ( n179937 , n12144 );
not ( n12559 , n179937 );
buf ( n179939 , n12559 );
buf ( n179940 , n179939 );
and ( n12562 , n179936 , n179940 );
not ( n12563 , n179936 );
buf ( n179943 , n12144 );
and ( n12565 , n12563 , n179943 );
nor ( n12566 , n12562 , n12565 );
buf ( n179946 , n12566 );
buf ( n179947 , n179946 );
not ( n12569 , n179947 );
buf ( n179949 , n12569 );
not ( n12571 , n179949 );
xor ( n12572 , n179562 , n179576 );
xnor ( n12573 , n12572 , n179567 );
buf ( n179953 , n12573 );
not ( n12575 , n179953 );
buf ( n179955 , n12575 );
not ( n12577 , n179955 );
or ( n12578 , n12571 , n12577 );
not ( n12579 , n12573 );
not ( n12580 , n179946 );
or ( n12581 , n12579 , n12580 );
buf ( n179961 , n171488 );
not ( n12583 , n179961 );
buf ( n179963 , n171592 );
not ( n12585 , n179963 );
buf ( n179965 , n4066 );
nand ( n12587 , n12585 , n179965 );
buf ( n179967 , n12587 );
buf ( n179968 , n179967 );
not ( n12590 , n179968 );
or ( n12591 , n12583 , n12590 );
buf ( n179971 , n4066 );
not ( n12593 , n179971 );
buf ( n179973 , n171592 );
nand ( n12595 , n12593 , n179973 );
buf ( n179975 , n12595 );
buf ( n179976 , n179975 );
nand ( n12598 , n12591 , n179976 );
buf ( n179978 , n12598 );
nand ( n12600 , n12581 , n179978 );
nand ( n12601 , n12578 , n12600 );
buf ( n179981 , n12601 );
not ( n12603 , n179981 );
buf ( n179983 , n12603 );
buf ( n179984 , n179983 );
nand ( n12606 , n179924 , n179984 );
buf ( n179986 , n12606 );
buf ( n179987 , n179986 );
not ( n12609 , n179987 );
or ( n12610 , n12538 , n12609 );
buf ( n179990 , n12541 );
buf ( n179991 , n12601 );
nand ( n12613 , n179990 , n179991 );
buf ( n179993 , n12613 );
buf ( n179994 , n179993 );
nand ( n12616 , n12610 , n179994 );
buf ( n179996 , n12616 );
not ( n12618 , n179996 );
xor ( n12619 , n12398 , n179780 );
xor ( n12620 , n12619 , n12492 );
not ( n12621 , n12620 );
and ( n12622 , n12618 , n12621 );
xor ( n12623 , n179588 , n179672 );
and ( n12624 , n12623 , n179694 );
not ( n12625 , n12623 );
and ( n12626 , n12625 , n12316 );
or ( n12627 , n12624 , n12626 );
nor ( n12628 , n12622 , n12627 );
nor ( n12629 , n12618 , n12621 );
nor ( n12630 , n12628 , n12629 );
not ( n12631 , n12630 );
buf ( n180011 , n12631 );
xor ( n12633 , n179722 , n179875 );
xor ( n12634 , n12633 , n179880 );
buf ( n180014 , n12634 );
buf ( n180015 , n180014 );
and ( n12637 , n180011 , n180015 );
buf ( n180017 , n12637 );
not ( n12642 , n180017 );
and ( n12643 , n12507 , n12642 );
and ( n12644 , n12627 , n179996 );
not ( n12645 , n12627 );
not ( n12646 , n179996 );
and ( n180023 , n12645 , n12646 );
nor ( n12648 , n12644 , n180023 );
xor ( n12649 , n12621 , n12648 );
buf ( n180026 , n12649 );
xor ( n12651 , n12470 , n179784 );
buf ( n180028 , n12651 );
buf ( n180029 , n179869 );
not ( n12654 , n180029 );
buf ( n180031 , n12654 );
buf ( n180032 , n180031 );
and ( n12657 , n180028 , n180032 );
not ( n12658 , n180028 );
buf ( n180035 , n179869 );
and ( n12660 , n12658 , n180035 );
nor ( n12661 , n12657 , n12660 );
buf ( n180038 , n12661 );
buf ( n180039 , n180038 );
not ( n12664 , n180039 );
xor ( n12665 , n171420 , n171467 );
and ( n12666 , n12665 , n171474 );
and ( n12667 , n171420 , n171467 );
or ( n12668 , n12666 , n12667 );
buf ( n180045 , n12668 );
buf ( n180046 , n180045 );
buf ( n180047 , n12573 );
buf ( n12672 , n180047 );
buf ( n180049 , n12672 );
buf ( n180050 , n180049 );
buf ( n180051 , n179978 );
not ( n12676 , n180051 );
buf ( n180053 , n179946 );
not ( n12678 , n180053 );
and ( n12679 , n12676 , n12678 );
buf ( n180056 , n179978 );
buf ( n180057 , n179946 );
and ( n12682 , n180056 , n180057 );
nor ( n12683 , n12679 , n12682 );
buf ( n180060 , n12683 );
buf ( n180061 , n180060 );
xor ( n12686 , n180050 , n180061 );
buf ( n180063 , n12686 );
buf ( n180064 , n180063 );
xor ( n12689 , n180046 , n180064 );
xor ( n12690 , n171609 , n171620 );
and ( n12691 , n12690 , n171627 );
and ( n12692 , n171609 , n171620 );
or ( n12693 , n12691 , n12692 );
buf ( n180070 , n12693 );
buf ( n180071 , n180070 );
and ( n12696 , n12689 , n180071 );
and ( n12697 , n180046 , n180064 );
or ( n12698 , n12696 , n12697 );
buf ( n180075 , n12698 );
buf ( n180076 , n180075 );
not ( n12701 , n180076 );
or ( n12702 , n12664 , n12701 );
buf ( n180079 , n180038 );
not ( n12704 , n180079 );
buf ( n180081 , n12704 );
buf ( n180082 , n180081 );
not ( n12707 , n180082 );
buf ( n180084 , n180075 );
not ( n12709 , n180084 );
buf ( n180086 , n12709 );
buf ( n180087 , n180086 );
not ( n12712 , n180087 );
or ( n12713 , n12707 , n12712 );
not ( n12714 , n12601 );
not ( n12715 , n12540 );
not ( n12716 , n12715 );
or ( n12717 , n12714 , n12716 );
nand ( n12718 , n12540 , n179983 );
nand ( n12719 , n12717 , n12718 );
buf ( n180096 , n12719 );
buf ( n180097 , n12530 );
buf ( n180098 , n12533 );
and ( n180099 , n180097 , n180098 );
buf ( n180100 , n180099 );
buf ( n180101 , n180100 );
xor ( n12726 , n180096 , n180101 );
buf ( n180103 , n12726 );
buf ( n180104 , n180103 );
not ( n180105 , n180104 );
buf ( n180106 , n180105 );
buf ( n180107 , n180106 );
nand ( n12732 , n12713 , n180107 );
buf ( n180109 , n12732 );
buf ( n180110 , n180109 );
nand ( n12735 , n12702 , n180110 );
buf ( n180112 , n12735 );
buf ( n180113 , n180112 );
and ( n12738 , n180026 , n180113 );
buf ( n180115 , n12738 );
xor ( n12740 , n180011 , n180015 );
buf ( n180117 , n12740 );
nor ( n12742 , n180115 , n180117 );
nor ( n12743 , n12643 , n12742 );
buf ( n180120 , n12743 );
xor ( n12745 , n178794 , n179445 );
and ( n12746 , n12745 , n179704 );
and ( n12747 , n178794 , n179445 );
or ( n12748 , n12746 , n12747 );
buf ( n180125 , n12748 );
buf ( n180126 , n180125 );
not ( n12751 , n180126 );
buf ( n180128 , n11799 );
not ( n12753 , n180128 );
buf ( n180130 , n11763 );
not ( n12755 , n180130 );
or ( n12756 , n12753 , n12755 );
buf ( n180133 , n179237 );
nand ( n12758 , n12756 , n180133 );
buf ( n180135 , n12758 );
buf ( n180136 , n180135 );
buf ( n180137 , n11799 );
not ( n12762 , n180137 );
not ( n12763 , n11763 );
buf ( n180140 , n12763 );
nand ( n12765 , n12762 , n180140 );
buf ( n180142 , n12765 );
buf ( n180143 , n180142 );
nand ( n12768 , n180136 , n180143 );
buf ( n180145 , n12768 );
buf ( n180146 , n180145 );
not ( n12771 , n179183 );
not ( n12772 , n179161 );
or ( n12773 , n12771 , n12772 );
buf ( n180150 , n179183 );
buf ( n180151 , n179161 );
nor ( n12776 , n180150 , n180151 );
buf ( n180153 , n12776 );
buf ( n180154 , n11772 );
not ( n12779 , n180154 );
buf ( n180156 , n12779 );
or ( n12781 , n180153 , n180156 );
nand ( n12782 , n12773 , n12781 );
buf ( n180159 , n12782 );
buf ( n180160 , n179256 );
not ( n12785 , n180160 );
buf ( n180162 , n168615 );
not ( n12787 , n180162 );
or ( n12788 , n12785 , n12787 );
buf ( n180165 , n168619 );
buf ( n180166 , n783 );
buf ( n180167 , n808 );
xor ( n12792 , n180166 , n180167 );
buf ( n180169 , n12792 );
buf ( n180170 , n180169 );
nand ( n12795 , n180165 , n180170 );
buf ( n180172 , n12795 );
buf ( n180173 , n180172 );
nand ( n12798 , n12788 , n180173 );
buf ( n180175 , n12798 );
buf ( n180176 , n180175 );
buf ( n180177 , n178742 );
not ( n12802 , n180177 );
buf ( n180179 , n1321 );
not ( n12804 , n180179 );
or ( n12805 , n12802 , n12804 );
buf ( n180182 , n168806 );
buf ( n180183 , n773 );
buf ( n180184 , n818 );
xor ( n12809 , n180183 , n180184 );
buf ( n180186 , n12809 );
buf ( n180187 , n180186 );
nand ( n12812 , n180182 , n180187 );
buf ( n180189 , n12812 );
buf ( n180190 , n180189 );
nand ( n12815 , n12805 , n180190 );
buf ( n180192 , n12815 );
buf ( n180193 , n180192 );
xor ( n12818 , n180176 , n180193 );
buf ( n180195 , n178759 );
not ( n12820 , n180195 );
buf ( n180197 , n168977 );
not ( n180198 , n180197 );
buf ( n180199 , n180198 );
buf ( n180200 , n180199 );
not ( n12825 , n180200 );
or ( n12826 , n12820 , n12825 );
buf ( n180203 , n170708 );
buf ( n180204 , n781 );
buf ( n180205 , n810 );
xor ( n12830 , n180204 , n180205 );
buf ( n180207 , n12830 );
buf ( n180208 , n180207 );
nand ( n12833 , n180203 , n180208 );
buf ( n180210 , n12833 );
buf ( n180211 , n180210 );
nand ( n12836 , n12826 , n180211 );
buf ( n180213 , n12836 );
buf ( n180214 , n180213 );
xor ( n12839 , n12818 , n180214 );
buf ( n180216 , n12839 );
buf ( n180217 , n180216 );
xor ( n12842 , n180159 , n180217 );
buf ( n180219 , n793 );
buf ( n180220 , n800 );
and ( n12845 , n180219 , n180220 );
buf ( n180222 , n12845 );
buf ( n180223 , n180222 );
buf ( n180224 , n11768 );
not ( n12849 , n180224 );
buf ( n180226 , n3497 );
not ( n12851 , n180226 );
or ( n12852 , n12849 , n12851 );
buf ( n180229 , n170972 );
buf ( n180230 , n791 );
buf ( n180231 , n800 );
xor ( n12856 , n180230 , n180231 );
buf ( n180233 , n12856 );
buf ( n180234 , n180233 );
nand ( n12859 , n180229 , n180234 );
buf ( n180236 , n12859 );
buf ( n180237 , n180236 );
nand ( n12862 , n12852 , n180237 );
buf ( n180239 , n12862 );
buf ( n180240 , n180239 );
xor ( n12865 , n180223 , n180240 );
buf ( n180242 , n179203 );
not ( n12867 , n180242 );
buf ( n180244 , n2251 );
not ( n12869 , n180244 );
or ( n12870 , n12867 , n12869 );
buf ( n180247 , n771 );
buf ( n180248 , n820 );
xnor ( n12873 , n180247 , n180248 );
buf ( n180250 , n12873 );
buf ( n180251 , n180250 );
not ( n12876 , n180251 );
buf ( n180253 , n168656 );
nand ( n12878 , n12876 , n180253 );
buf ( n180255 , n12878 );
buf ( n180256 , n180255 );
nand ( n12881 , n12870 , n180256 );
buf ( n180258 , n12881 );
buf ( n180259 , n180258 );
xor ( n12884 , n12865 , n180259 );
buf ( n180261 , n12884 );
buf ( n180262 , n180261 );
xor ( n12887 , n12842 , n180262 );
buf ( n180264 , n12887 );
buf ( n180265 , n180264 );
xor ( n12890 , n180146 , n180265 );
xor ( n12891 , n179246 , n179291 );
and ( n12892 , n12891 , n179298 );
and ( n12893 , n179246 , n179291 );
or ( n12894 , n12892 , n12893 );
buf ( n180271 , n12894 );
buf ( n180272 , n180271 );
xor ( n12897 , n12890 , n180272 );
buf ( n180274 , n12897 );
buf ( n180275 , n180274 );
xor ( n12900 , n179098 , n179239 );
and ( n12901 , n12900 , n179301 );
and ( n12902 , n179098 , n179239 );
or ( n12903 , n12901 , n12902 );
buf ( n180280 , n12903 );
buf ( n180281 , n180280 );
xor ( n12906 , n180275 , n180281 );
not ( n12907 , n179221 );
not ( n12908 , n1806 );
or ( n12909 , n12907 , n12908 );
buf ( n180286 , n169169 );
buf ( n180287 , n824 );
nand ( n12912 , n180286 , n180287 );
buf ( n180289 , n12912 );
nand ( n12914 , n12909 , n180289 );
not ( n12915 , n179177 );
not ( n12916 , n3764 );
or ( n12917 , n12915 , n12916 );
buf ( n180294 , n777 );
buf ( n180295 , n814 );
xor ( n12920 , n180294 , n180295 );
buf ( n180297 , n12920 );
nand ( n12922 , n180297 , n169250 );
nand ( n12923 , n12917 , n12922 );
xor ( n12924 , n12914 , n12923 );
buf ( n180301 , n179106 );
not ( n12926 , n180301 );
buf ( n180303 , n178232 );
not ( n12928 , n180303 );
or ( n12929 , n12926 , n12928 );
buf ( n180306 , n168867 );
buf ( n180307 , n789 );
buf ( n180308 , n802 );
xor ( n12933 , n180307 , n180308 );
buf ( n180310 , n12933 );
buf ( n180311 , n180310 );
nand ( n12936 , n180306 , n180311 );
buf ( n180313 , n12936 );
buf ( n180314 , n180313 );
nand ( n12939 , n12929 , n180314 );
buf ( n180316 , n12939 );
xor ( n12941 , n12924 , n180316 );
buf ( n180318 , n12941 );
buf ( n180319 , n11898 );
not ( n12944 , n180319 );
buf ( n180321 , n168713 );
not ( n12946 , n180321 );
or ( n12947 , n12944 , n12946 );
buf ( n180324 , n2823 );
buf ( n180325 , n785 );
buf ( n180326 , n806 );
xor ( n12951 , n180325 , n180326 );
buf ( n180328 , n12951 );
buf ( n180329 , n180328 );
nand ( n12954 , n180324 , n180329 );
buf ( n180331 , n12954 );
buf ( n180332 , n180331 );
nand ( n12957 , n12947 , n180332 );
buf ( n180334 , n12957 );
not ( n12959 , n179141 );
not ( n12960 , n169314 );
or ( n12961 , n12959 , n12960 );
buf ( n180338 , n775 );
buf ( n180339 , n816 );
xor ( n12964 , n180338 , n180339 );
buf ( n180341 , n12964 );
nand ( n12966 , n169845 , n180341 );
nand ( n12967 , n12961 , n12966 );
xor ( n12968 , n180334 , n12967 );
buf ( n180345 , n11738 );
not ( n12970 , n180345 );
buf ( n180347 , n168832 );
not ( n12972 , n180347 );
or ( n12973 , n12970 , n12972 );
buf ( n180350 , n168759 );
xor ( n12975 , n804 , n787 );
buf ( n180352 , n12975 );
nand ( n12977 , n180350 , n180352 );
buf ( n180354 , n12977 );
buf ( n180355 , n180354 );
nand ( n12980 , n12973 , n180355 );
buf ( n180357 , n12980 );
xor ( n12982 , n12968 , n180357 );
buf ( n180359 , n12982 );
xor ( n12984 , n180318 , n180359 );
buf ( n180361 , n178777 );
not ( n12986 , n180361 );
buf ( n180363 , n1907 );
not ( n12988 , n180363 );
or ( n12989 , n12986 , n12988 );
buf ( n180366 , n6287 );
buf ( n180367 , n779 );
buf ( n180368 , n812 );
xor ( n12996 , n180367 , n180368 );
buf ( n180370 , n12996 );
buf ( n180371 , n180370 );
nand ( n12999 , n180366 , n180371 );
buf ( n180373 , n12999 );
buf ( n180374 , n180373 );
nand ( n13002 , n12989 , n180374 );
buf ( n180376 , n13002 );
buf ( n180377 , n180376 );
buf ( n180378 , n11884 );
not ( n13006 , n180378 );
buf ( n180380 , n169411 );
not ( n13008 , n180380 );
or ( n13009 , n13006 , n13008 );
buf ( n180383 , n171055 );
buf ( n180384 , n769 );
buf ( n180385 , n822 );
xor ( n13013 , n180384 , n180385 );
buf ( n180387 , n13013 );
buf ( n180388 , n180387 );
nand ( n13016 , n180383 , n180388 );
buf ( n180390 , n13016 );
buf ( n180391 , n180390 );
nand ( n13019 , n13009 , n180391 );
buf ( n180393 , n13019 );
buf ( n180394 , n180393 );
not ( n13022 , n180394 );
buf ( n180396 , n13022 );
buf ( n180397 , n180396 );
xor ( n13025 , n180377 , n180397 );
buf ( n180399 , n11725 );
not ( n13027 , n180399 );
buf ( n180401 , n13027 );
buf ( n180402 , n180401 );
not ( n13030 , n180402 );
buf ( n180404 , n179129 );
not ( n13032 , n180404 );
or ( n13033 , n13030 , n13032 );
buf ( n180407 , n179147 );
nand ( n13035 , n13033 , n180407 );
buf ( n180409 , n13035 );
buf ( n180410 , n180409 );
nand ( n13038 , n11745 , n11725 );
buf ( n180412 , n13038 );
nand ( n13040 , n180410 , n180412 );
buf ( n180414 , n13040 );
buf ( n180415 , n180414 );
xor ( n13043 , n13025 , n180415 );
buf ( n180417 , n13043 );
buf ( n180418 , n180417 );
xor ( n13046 , n12984 , n180418 );
buf ( n180420 , n13046 );
buf ( n180421 , n180420 );
buf ( n180422 , n178789 );
not ( n13050 , n180422 );
buf ( n180424 , n178614 );
not ( n13052 , n180424 );
or ( n13053 , n13050 , n13052 );
buf ( n180427 , n178614 );
buf ( n180428 , n178789 );
or ( n13056 , n180427 , n180428 );
buf ( n180430 , n178619 );
nand ( n13058 , n13056 , n180430 );
buf ( n180432 , n13058 );
buf ( n180433 , n180432 );
nand ( n13061 , n13053 , n180433 );
buf ( n180435 , n13061 );
buf ( n180436 , n180435 );
xor ( n13064 , n180421 , n180436 );
xor ( n13065 , n178558 , n178605 );
and ( n13066 , n13065 , n178612 );
and ( n13067 , n178558 , n178605 );
or ( n13068 , n13066 , n13067 );
buf ( n180442 , n13068 );
buf ( n180443 , n180442 );
xor ( n13071 , n178671 , n178731 );
and ( n13072 , n13071 , n178787 );
and ( n13073 , n178671 , n178731 );
or ( n13074 , n13072 , n13073 );
buf ( n180448 , n13074 );
buf ( n180449 , n180448 );
xor ( n13077 , n180443 , n180449 );
buf ( n180451 , n179262 );
buf ( n180452 , n179275 );
nand ( n13080 , n180451 , n180452 );
buf ( n180454 , n13080 );
buf ( n180455 , n180454 );
buf ( n180456 , n179262 );
buf ( n180457 , n179275 );
or ( n13085 , n180456 , n180457 );
buf ( n180459 , n179289 );
nand ( n13087 , n13085 , n180459 );
buf ( n180461 , n13087 );
buf ( n180462 , n180461 );
nand ( n13090 , n180455 , n180462 );
buf ( n180464 , n13090 );
buf ( n180465 , n180464 );
buf ( n180466 , n179227 );
not ( n13094 , n180466 );
buf ( n180468 , n179209 );
not ( n13096 , n180468 );
or ( n13097 , n13094 , n13096 );
buf ( n180471 , n179233 );
not ( n13099 , n180471 );
buf ( n180473 , n179209 );
not ( n13101 , n180473 );
buf ( n180475 , n13101 );
buf ( n180476 , n180475 );
not ( n13104 , n180476 );
or ( n13105 , n13099 , n13104 );
buf ( n180479 , n179193 );
nand ( n13107 , n13105 , n180479 );
buf ( n180481 , n13107 );
buf ( n180482 , n180481 );
nand ( n13110 , n13097 , n180482 );
buf ( n180484 , n13110 );
buf ( n180485 , n180484 );
xor ( n13113 , n180465 , n180485 );
xor ( n13114 , n178749 , n178766 );
and ( n13115 , n13114 , n178784 );
and ( n13116 , n178749 , n178766 );
or ( n13117 , n13115 , n13116 );
buf ( n180491 , n13117 );
buf ( n180492 , n180491 );
xor ( n13120 , n13113 , n180492 );
buf ( n180494 , n13120 );
buf ( n180495 , n180494 );
xor ( n13123 , n13077 , n180495 );
buf ( n180497 , n13123 );
buf ( n180498 , n180497 );
xor ( n13126 , n13064 , n180498 );
buf ( n180500 , n13126 );
buf ( n180501 , n180500 );
xor ( n13129 , n12906 , n180501 );
buf ( n180503 , n13129 );
buf ( n180504 , n180503 );
xor ( n13132 , n178109 , n178556 );
and ( n13133 , n13132 , n178791 );
and ( n13134 , n178109 , n178556 );
or ( n13135 , n13133 , n13134 );
buf ( n180509 , n13135 );
buf ( n180510 , n180509 );
not ( n13138 , n180510 );
buf ( n180512 , n13138 );
buf ( n180513 , n180512 );
and ( n13141 , n180504 , n180513 );
not ( n13142 , n180504 );
buf ( n180516 , n180509 );
and ( n13144 , n13142 , n180516 );
nor ( n13145 , n13141 , n13144 );
buf ( n180519 , n13145 );
buf ( n180520 , n180519 );
xor ( n13148 , n179086 , n179304 );
and ( n13149 , n13148 , n179442 );
and ( n13150 , n179086 , n179304 );
or ( n13151 , n13149 , n13150 );
buf ( n180525 , n13151 );
buf ( n180526 , n180525 );
buf ( n13154 , n180526 );
buf ( n180528 , n13154 );
buf ( n180529 , n180528 );
and ( n13157 , n180520 , n180529 );
not ( n180531 , n180520 );
buf ( n180532 , n180528 );
not ( n13160 , n180532 );
buf ( n180534 , n13160 );
buf ( n180535 , n180534 );
and ( n13163 , n180531 , n180535 );
nor ( n13164 , n13157 , n13163 );
buf ( n180538 , n13164 );
not ( n13166 , n180538 );
not ( n13167 , n13166 );
buf ( n180541 , n13167 );
not ( n13169 , n180541 );
or ( n13170 , n12751 , n13169 );
buf ( n180544 , n180125 );
not ( n13172 , n180544 );
buf ( n180546 , n13172 );
buf ( n180547 , n180546 );
buf ( n180548 , n13166 );
nand ( n13176 , n180547 , n180548 );
buf ( n180550 , n13176 );
buf ( n180551 , n180550 );
nand ( n13179 , n13170 , n180551 );
buf ( n180553 , n13179 );
buf ( n180554 , n180553 );
buf ( n180555 , n179706 );
buf ( n180556 , n179884 );
and ( n13184 , n180555 , n180556 );
buf ( n180558 , n13184 );
buf ( n180559 , n180558 );
nor ( n13187 , n180554 , n180559 );
buf ( n180561 , n13187 );
buf ( n180562 , n180561 );
and ( n13190 , n13166 , n180125 );
buf ( n180564 , n13190 );
buf ( n180565 , n180509 );
not ( n13193 , n180565 );
buf ( n180567 , n180525 );
not ( n13195 , n180567 );
or ( n13196 , n13193 , n13195 );
buf ( n180570 , n180512 );
not ( n13198 , n180570 );
buf ( n180572 , n180525 );
not ( n13200 , n180572 );
buf ( n180574 , n13200 );
buf ( n180575 , n180574 );
not ( n13203 , n180575 );
or ( n13204 , n13198 , n13203 );
buf ( n180578 , n180503 );
buf ( n13206 , n180578 );
buf ( n180580 , n13206 );
buf ( n180581 , n180580 );
nand ( n13209 , n13204 , n180581 );
buf ( n180583 , n13209 );
buf ( n180584 , n180583 );
nand ( n13212 , n13196 , n180584 );
buf ( n180586 , n13212 );
not ( n13214 , n180586 );
not ( n13215 , n13214 );
buf ( n180589 , n13215 );
not ( n13217 , n180589 );
xor ( n13218 , n180421 , n180436 );
and ( n13219 , n13218 , n180498 );
and ( n13220 , n180421 , n180436 );
or ( n13221 , n13219 , n13220 );
buf ( n180595 , n13221 );
buf ( n180596 , n180595 );
xor ( n13224 , n180275 , n180281 );
and ( n13225 , n13224 , n180501 );
and ( n13226 , n180275 , n180281 );
or ( n13227 , n13225 , n13226 );
buf ( n180601 , n13227 );
buf ( n180602 , n180601 );
xor ( n13230 , n180596 , n180602 );
xor ( n13231 , n180146 , n180265 );
and ( n13232 , n13231 , n180272 );
and ( n13233 , n180146 , n180265 );
or ( n13234 , n13232 , n13233 );
buf ( n180608 , n13234 );
xor ( n13236 , n180159 , n180217 );
and ( n13237 , n13236 , n180262 );
and ( n13238 , n180159 , n180217 );
or ( n13239 , n13237 , n13238 );
buf ( n180613 , n13239 );
xor ( n13241 , n180223 , n180240 );
and ( n13242 , n13241 , n180259 );
and ( n13243 , n180223 , n180240 );
or ( n13244 , n13242 , n13243 );
buf ( n180618 , n13244 );
buf ( n180619 , n180618 );
buf ( n180620 , n180169 );
not ( n13248 , n180620 );
buf ( n180622 , n169545 );
not ( n13250 , n180622 );
or ( n13251 , n13248 , n13250 );
buf ( n180625 , n168619 );
buf ( n180626 , n782 );
buf ( n180627 , n808 );
xor ( n13255 , n180626 , n180627 );
buf ( n180629 , n13255 );
buf ( n180630 , n180629 );
nand ( n13258 , n180625 , n180630 );
buf ( n180632 , n13258 );
buf ( n180633 , n180632 );
nand ( n13261 , n13251 , n180633 );
buf ( n180635 , n13261 );
buf ( n180636 , n180635 );
buf ( n180637 , n180207 );
not ( n13265 , n180637 );
buf ( n180639 , n169951 );
not ( n13267 , n180639 );
or ( n13268 , n13265 , n13267 );
buf ( n180642 , n168989 );
buf ( n180643 , n780 );
buf ( n180644 , n810 );
xor ( n13272 , n180643 , n180644 );
buf ( n180646 , n13272 );
buf ( n180647 , n180646 );
nand ( n13275 , n180642 , n180647 );
buf ( n180649 , n13275 );
buf ( n180650 , n180649 );
nand ( n13278 , n13268 , n180650 );
buf ( n180652 , n13278 );
buf ( n180653 , n180652 );
xor ( n13281 , n180636 , n180653 );
buf ( n180655 , n7665 );
buf ( n180656 , n180341 );
not ( n13284 , n180656 );
buf ( n180658 , n13284 );
buf ( n180659 , n180658 );
or ( n13287 , n180655 , n180659 );
buf ( n180661 , n169845 );
not ( n13289 , n180661 );
buf ( n180663 , n13289 );
buf ( n180664 , n180663 );
buf ( n180665 , n774 );
buf ( n180666 , n816 );
xor ( n13294 , n180665 , n180666 );
buf ( n180668 , n13294 );
buf ( n180669 , n180668 );
not ( n13297 , n180669 );
buf ( n180671 , n13297 );
buf ( n180672 , n180671 );
or ( n13300 , n180664 , n180672 );
nand ( n13301 , n13287 , n13300 );
buf ( n180675 , n13301 );
buf ( n180676 , n180675 );
xor ( n13304 , n13281 , n180676 );
buf ( n180678 , n13304 );
buf ( n180679 , n180678 );
xor ( n13307 , n180619 , n180679 );
buf ( n180681 , n180186 );
not ( n13309 , n180681 );
buf ( n180683 , n171706 );
not ( n13311 , n180683 );
or ( n13312 , n13309 , n13311 );
buf ( n180686 , n168806 );
buf ( n180687 , n772 );
buf ( n180688 , n818 );
xor ( n13316 , n180687 , n180688 );
buf ( n180690 , n13316 );
buf ( n180691 , n180690 );
nand ( n13319 , n180686 , n180691 );
buf ( n180693 , n13319 );
buf ( n180694 , n180693 );
nand ( n13325 , n13312 , n180694 );
buf ( n180696 , n13325 );
not ( n13327 , n180696 );
buf ( n180698 , n180387 );
not ( n13329 , n180698 );
buf ( n180700 , n169411 );
not ( n13331 , n180700 );
or ( n13332 , n13329 , n13331 );
buf ( n180703 , n171055 );
buf ( n180704 , n768 );
buf ( n180705 , n822 );
xor ( n13336 , n180704 , n180705 );
buf ( n180707 , n13336 );
buf ( n180708 , n180707 );
nand ( n13339 , n180703 , n180708 );
buf ( n180710 , n13339 );
buf ( n180711 , n180710 );
nand ( n13342 , n13332 , n180711 );
buf ( n180713 , n13342 );
not ( n13344 , n180713 );
buf ( n180715 , n170562 );
not ( n13346 , n180715 );
buf ( n180717 , n169151 );
not ( n13348 , n180717 );
or ( n13349 , n13346 , n13348 );
buf ( n180720 , n824 );
nand ( n13351 , n13349 , n180720 );
buf ( n180722 , n13351 );
nand ( n13353 , n13327 , n13344 , n180722 );
not ( n13354 , n180696 );
nor ( n13355 , n13354 , n180722 );
nand ( n13356 , n13344 , n13355 );
nor ( n13357 , n180722 , n180696 );
nand ( n13358 , n180713 , n13357 );
nand ( n13359 , n180722 , n180696 );
not ( n13360 , n13359 );
nand ( n13361 , n13360 , n180713 );
nand ( n13362 , n13353 , n13356 , n13358 , n13361 );
buf ( n180733 , n13362 );
xor ( n13364 , n13307 , n180733 );
buf ( n180735 , n13364 );
xor ( n13366 , n180613 , n180735 );
buf ( n180737 , n180297 );
not ( n13368 , n180737 );
buf ( n180739 , n169241 );
not ( n13370 , n180739 );
or ( n13371 , n13368 , n13370 );
buf ( n180742 , n169250 );
buf ( n180743 , n776 );
buf ( n180744 , n814 );
xor ( n13375 , n180743 , n180744 );
buf ( n180746 , n13375 );
buf ( n180747 , n180746 );
nand ( n13378 , n180742 , n180747 );
buf ( n180749 , n13378 );
buf ( n180750 , n180749 );
nand ( n13381 , n13371 , n180750 );
buf ( n180752 , n13381 );
buf ( n180753 , n180752 );
not ( n13384 , n180753 );
buf ( n180755 , n13384 );
buf ( n180756 , n180755 );
not ( n13387 , n180756 );
buf ( n180758 , n180310 );
not ( n13389 , n180758 );
buf ( n13390 , n1389 );
buf ( n180761 , n13390 );
not ( n13392 , n180761 );
or ( n13393 , n13389 , n13392 );
buf ( n180764 , n168867 );
buf ( n180765 , n788 );
buf ( n180766 , n802 );
xor ( n13397 , n180765 , n180766 );
buf ( n180768 , n13397 );
buf ( n180769 , n180768 );
nand ( n13400 , n180764 , n180769 );
buf ( n180771 , n13400 );
buf ( n180772 , n180771 );
nand ( n13403 , n13393 , n180772 );
buf ( n180774 , n13403 );
buf ( n180775 , n180774 );
not ( n13406 , n180775 );
and ( n13407 , n13387 , n13406 );
buf ( n180778 , n180774 );
buf ( n180779 , n180755 );
and ( n13410 , n180778 , n180779 );
nor ( n13411 , n13407 , n13410 );
buf ( n180782 , n13411 );
buf ( n180783 , n180233 );
not ( n13414 , n180783 );
buf ( n180785 , n3497 );
not ( n13416 , n180785 );
or ( n13417 , n13414 , n13416 );
buf ( n180788 , n170972 );
buf ( n180789 , n790 );
buf ( n180790 , n800 );
xor ( n13421 , n180789 , n180790 );
buf ( n180792 , n13421 );
buf ( n180793 , n180792 );
nand ( n13424 , n180788 , n180793 );
buf ( n180795 , n13424 );
buf ( n180796 , n180795 );
nand ( n13427 , n13417 , n180796 );
buf ( n180798 , n13427 );
and ( n13429 , n180782 , n180798 );
not ( n13430 , n180782 );
buf ( n180801 , n180798 );
not ( n13432 , n180801 );
buf ( n180803 , n13432 );
and ( n13434 , n13430 , n180803 );
nor ( n13435 , n13429 , n13434 );
buf ( n180806 , n180328 );
not ( n13437 , n180806 );
buf ( n180808 , n169635 );
not ( n13439 , n180808 );
or ( n13440 , n13437 , n13439 );
buf ( n180811 , n169641 );
buf ( n180812 , n784 );
buf ( n180813 , n806 );
xor ( n13444 , n180812 , n180813 );
buf ( n180815 , n13444 );
buf ( n180816 , n180815 );
nand ( n13447 , n180811 , n180816 );
buf ( n180818 , n13447 );
buf ( n180819 , n180818 );
nand ( n13450 , n13440 , n180819 );
buf ( n180821 , n13450 );
buf ( n180822 , n180821 );
not ( n13453 , n2251 );
not ( n13454 , n180250 );
not ( n13455 , n13454 );
or ( n13456 , n13453 , n13455 );
buf ( n180827 , n168655 );
xor ( n13458 , n820 , n770 );
buf ( n180829 , n13458 );
nand ( n13460 , n180827 , n180829 );
buf ( n180831 , n13460 );
nand ( n13462 , n13456 , n180831 );
buf ( n180833 , n13462 );
xor ( n13464 , n180822 , n180833 );
buf ( n180835 , n12975 );
not ( n13466 , n180835 );
buf ( n180837 , n168832 );
not ( n13468 , n180837 );
or ( n13469 , n13466 , n13468 );
buf ( n180840 , n178447 );
buf ( n180841 , n786 );
buf ( n180842 , n804 );
xor ( n13473 , n180841 , n180842 );
buf ( n180844 , n13473 );
buf ( n180845 , n180844 );
nand ( n13476 , n180840 , n180845 );
buf ( n180847 , n13476 );
buf ( n180848 , n180847 );
nand ( n13479 , n13469 , n180848 );
buf ( n180850 , n13479 );
buf ( n180851 , n180850 );
xor ( n13482 , n13464 , n180851 );
buf ( n180853 , n13482 );
not ( n13484 , n180853 );
and ( n13485 , n13435 , n13484 );
not ( n13486 , n13435 );
and ( n13487 , n13486 , n180853 );
nor ( n13488 , n13485 , n13487 );
buf ( n180859 , n13488 );
buf ( n180860 , n792 );
buf ( n180861 , n800 );
and ( n13492 , n180860 , n180861 );
buf ( n180863 , n13492 );
buf ( n180864 , n180863 );
buf ( n180865 , n180393 );
xor ( n13496 , n180864 , n180865 );
buf ( n180867 , n180370 );
not ( n13498 , n180867 );
buf ( n180869 , n1907 );
not ( n13500 , n180869 );
or ( n13501 , n13498 , n13500 );
buf ( n180872 , n1535 );
buf ( n180873 , n778 );
buf ( n180874 , n812 );
xor ( n13505 , n180873 , n180874 );
buf ( n180876 , n13505 );
buf ( n180877 , n180876 );
nand ( n13508 , n180872 , n180877 );
buf ( n180879 , n13508 );
buf ( n180880 , n180879 );
nand ( n13511 , n13501 , n180880 );
buf ( n180882 , n13511 );
buf ( n180883 , n180882 );
xor ( n13514 , n13496 , n180883 );
buf ( n180885 , n13514 );
buf ( n180886 , n180885 );
and ( n13517 , n180859 , n180886 );
not ( n13518 , n180859 );
buf ( n180889 , n180885 );
not ( n13520 , n180889 );
buf ( n180891 , n13520 );
buf ( n180892 , n180891 );
and ( n13523 , n13518 , n180892 );
nor ( n13524 , n13517 , n13523 );
buf ( n180895 , n13524 );
xor ( n13526 , n13366 , n180895 );
xor ( n13527 , n180608 , n13526 );
xor ( n13528 , n180318 , n180359 );
and ( n13529 , n13528 , n180418 );
and ( n13530 , n180318 , n180359 );
or ( n13531 , n13529 , n13530 );
buf ( n180902 , n13531 );
buf ( n180903 , n180902 );
xor ( n13534 , n180377 , n180397 );
and ( n13535 , n13534 , n180415 );
and ( n13536 , n180377 , n180397 );
or ( n13537 , n13535 , n13536 );
buf ( n180908 , n13537 );
buf ( n180909 , n180908 );
buf ( n180910 , n12914 );
not ( n13541 , n180910 );
buf ( n180912 , n12923 );
not ( n13543 , n180912 );
or ( n13544 , n13541 , n13543 );
or ( n13545 , n12923 , n12914 );
nand ( n13546 , n13545 , n180316 );
buf ( n180917 , n13546 );
nand ( n13548 , n13544 , n180917 );
buf ( n180919 , n13548 );
buf ( n180920 , n180919 );
buf ( n180921 , n180357 );
not ( n13552 , n180921 );
buf ( n180923 , n180334 );
not ( n13554 , n180923 );
or ( n13555 , n13552 , n13554 );
buf ( n180926 , n180357 );
buf ( n180927 , n180334 );
or ( n13558 , n180926 , n180927 );
buf ( n180929 , n12967 );
nand ( n13560 , n13558 , n180929 );
buf ( n180931 , n13560 );
buf ( n180932 , n180931 );
nand ( n13563 , n13555 , n180932 );
buf ( n180934 , n13563 );
buf ( n180935 , n180934 );
xor ( n13566 , n180920 , n180935 );
xor ( n13567 , n180176 , n180193 );
and ( n13568 , n13567 , n180214 );
and ( n13569 , n180176 , n180193 );
or ( n13570 , n13568 , n13569 );
buf ( n180941 , n13570 );
buf ( n180942 , n180941 );
xor ( n13573 , n13566 , n180942 );
buf ( n180944 , n13573 );
buf ( n180945 , n180944 );
xor ( n13576 , n180909 , n180945 );
xor ( n13577 , n180465 , n180485 );
and ( n13578 , n13577 , n180492 );
and ( n13579 , n180465 , n180485 );
or ( n13580 , n13578 , n13579 );
buf ( n180951 , n13580 );
buf ( n180952 , n180951 );
xor ( n13583 , n13576 , n180952 );
buf ( n180954 , n13583 );
buf ( n180955 , n180954 );
xor ( n13586 , n180903 , n180955 );
xor ( n13587 , n180443 , n180449 );
and ( n13588 , n13587 , n180495 );
and ( n13589 , n180443 , n180449 );
or ( n13590 , n13588 , n13589 );
buf ( n180961 , n13590 );
buf ( n180962 , n180961 );
xor ( n13593 , n13586 , n180962 );
buf ( n180964 , n13593 );
xor ( n13595 , n13527 , n180964 );
buf ( n180966 , n13595 );
xor ( n13597 , n13230 , n180966 );
buf ( n180968 , n13597 );
buf ( n180969 , n180968 );
not ( n13600 , n180969 );
buf ( n180971 , n13600 );
buf ( n180972 , n180971 );
not ( n13603 , n180972 );
or ( n13604 , n13217 , n13603 );
buf ( n180975 , n180968 );
buf ( n180976 , n13214 );
nand ( n13607 , n180975 , n180976 );
buf ( n180978 , n13607 );
buf ( n180979 , n180978 );
nand ( n13610 , n13604 , n180979 );
buf ( n180981 , n13610 );
buf ( n180982 , n180981 );
nor ( n13613 , n180564 , n180982 );
buf ( n180984 , n13613 );
buf ( n180985 , n180984 );
nor ( n13616 , n180562 , n180985 );
buf ( n180987 , n13616 );
buf ( n180988 , n180987 );
nand ( n13619 , n180120 , n180988 );
buf ( n180990 , n13619 );
buf ( n180991 , n180990 );
not ( n13622 , n180991 );
xor ( n13623 , n180103 , n180038 );
and ( n13624 , n13623 , n180075 );
not ( n13625 , n13623 );
and ( n13626 , n13625 , n180086 );
nor ( n13627 , n13624 , n13626 );
not ( n13628 , n13627 );
xor ( n13629 , n12524 , n12510 );
not ( n13630 , n12529 );
and ( n13631 , n13629 , n13630 );
not ( n13632 , n13629 );
and ( n13633 , n13632 , n12529 );
nor ( n13634 , n13631 , n13633 );
xor ( n13635 , n171208 , n171477 );
and ( n13636 , n13635 , n171630 );
and ( n13637 , n171208 , n171477 );
or ( n13638 , n13636 , n13637 );
buf ( n181009 , n13638 );
xor ( n13640 , n13634 , n181009 );
xor ( n13641 , n180046 , n180064 );
xor ( n181012 , n13641 , n180071 );
buf ( n181013 , n181012 );
and ( n13647 , n13640 , n181013 );
and ( n13648 , n13634 , n181009 );
or ( n13649 , n13647 , n13648 );
and ( n13650 , n13628 , n13649 );
not ( n13651 , n13628 );
not ( n13652 , n13649 );
and ( n13653 , n13651 , n13652 );
nor ( n13654 , n13650 , n13653 );
xor ( n13655 , n13634 , n181009 );
xor ( n13656 , n13655 , n181013 );
buf ( n181024 , n13656 );
xor ( n13658 , n171112 , n171118 );
and ( n13659 , n13658 , n171633 );
and ( n13660 , n171112 , n171118 );
or ( n13661 , n13659 , n13660 );
buf ( n181029 , n13661 );
buf ( n181030 , n181029 );
and ( n13664 , n181024 , n181030 );
buf ( n181032 , n13664 );
nor ( n13666 , n13654 , n181032 );
buf ( n181034 , n13628 );
buf ( n181035 , n13649 );
and ( n13669 , n181034 , n181035 );
buf ( n181037 , n13669 );
buf ( n181038 , n181037 );
xor ( n13672 , n12649 , n180112 );
buf ( n181040 , n13672 );
nor ( n13674 , n181038 , n181040 );
buf ( n181042 , n13674 );
nor ( n13676 , n13666 , n181042 );
buf ( n181044 , n13676 );
not ( n13678 , n181044 );
buf ( n181046 , n171654 );
buf ( n181047 , n181029 );
not ( n13681 , n181047 );
not ( n13682 , n13656 );
buf ( n181050 , n13682 );
not ( n13684 , n181050 );
or ( n13685 , n13681 , n13684 );
buf ( n181053 , n13656 );
buf ( n181054 , n181029 );
not ( n13688 , n181054 );
buf ( n181056 , n13688 );
buf ( n181057 , n181056 );
nand ( n13691 , n181053 , n181057 );
buf ( n181059 , n13691 );
buf ( n181060 , n181059 );
nand ( n13694 , n13685 , n181060 );
buf ( n181062 , n13694 );
not ( n13696 , n181062 );
and ( n13697 , n171635 , n171104 );
not ( n13698 , n13697 );
nand ( n13699 , n13696 , n13698 );
buf ( n181067 , n13699 );
nand ( n13701 , n181046 , n181067 );
buf ( n181069 , n13701 );
buf ( n181070 , n181069 );
nor ( n13704 , n13678 , n181070 );
buf ( n181072 , n13704 );
buf ( n181073 , n181072 );
nand ( n13707 , n13622 , n181073 );
buf ( n181075 , n13707 );
buf ( n181076 , n181075 );
not ( n13710 , n181076 );
buf ( n181078 , n13710 );
buf ( n181079 , n181078 );
not ( n13713 , n181079 );
buf ( n181081 , n13713 );
buf ( n181082 , n181081 );
not ( n13716 , n170972 );
buf ( n181084 , n789 );
buf ( n181085 , n800 );
xor ( n13719 , n181084 , n181085 );
buf ( n181087 , n13719 );
not ( n13721 , n181087 );
or ( n13722 , n13716 , n13721 );
nand ( n13723 , n3497 , n180792 );
nand ( n13724 , n13722 , n13723 );
buf ( n181092 , n13724 );
buf ( n181093 , n180707 );
not ( n13727 , n181093 );
buf ( n181095 , n1939 );
not ( n13729 , n181095 );
or ( n13730 , n13727 , n13729 );
buf ( n181098 , n822 );
buf ( n181099 , n171055 );
nand ( n13733 , n181098 , n181099 );
buf ( n181101 , n13733 );
buf ( n181102 , n181101 );
nand ( n13736 , n13730 , n181102 );
buf ( n181104 , n13736 );
buf ( n181105 , n181104 );
xor ( n13739 , n181092 , n181105 );
buf ( n181107 , n180876 );
not ( n13741 , n181107 );
buf ( n181109 , n1907 );
not ( n13743 , n181109 );
or ( n13744 , n13741 , n13743 );
buf ( n181112 , n6287 );
buf ( n181113 , n777 );
buf ( n181114 , n812 );
xor ( n13748 , n181113 , n181114 );
buf ( n181116 , n13748 );
buf ( n181117 , n181116 );
nand ( n13751 , n181112 , n181117 );
buf ( n181119 , n13751 );
buf ( n181120 , n181119 );
nand ( n13754 , n13744 , n181120 );
buf ( n181122 , n13754 );
buf ( n181123 , n181122 );
xor ( n13757 , n13739 , n181123 );
buf ( n181125 , n13757 );
buf ( n181126 , n181125 );
buf ( n181127 , n180815 );
not ( n13761 , n181127 );
buf ( n181129 , n168713 );
not ( n13763 , n181129 );
or ( n13764 , n13761 , n13763 );
buf ( n181132 , n2823 );
buf ( n181133 , n783 );
buf ( n181134 , n806 );
xor ( n13768 , n181133 , n181134 );
buf ( n181136 , n13768 );
buf ( n181137 , n181136 );
nand ( n13771 , n181132 , n181137 );
buf ( n181139 , n13771 );
buf ( n181140 , n181139 );
nand ( n13774 , n13764 , n181140 );
buf ( n181142 , n13774 );
buf ( n181143 , n181142 );
not ( n13777 , n181143 );
buf ( n181145 , n13777 );
buf ( n181146 , n181145 );
not ( n13780 , n181146 );
buf ( n181148 , n180629 );
not ( n13782 , n181148 );
buf ( n181150 , n177984 );
not ( n13784 , n181150 );
or ( n13785 , n13782 , n13784 );
buf ( n181153 , n168619 );
buf ( n181154 , n781 );
buf ( n181155 , n808 );
xor ( n13789 , n181154 , n181155 );
buf ( n181157 , n13789 );
buf ( n181158 , n181157 );
nand ( n13792 , n181153 , n181158 );
buf ( n181160 , n13792 );
buf ( n181161 , n181160 );
nand ( n13795 , n13785 , n181161 );
buf ( n181163 , n13795 );
buf ( n181164 , n180668 );
not ( n13798 , n181164 );
buf ( n181166 , n169314 );
not ( n13800 , n181166 );
or ( n13801 , n13798 , n13800 );
buf ( n181169 , n169320 );
buf ( n181170 , n773 );
buf ( n181171 , n816 );
xor ( n13805 , n181170 , n181171 );
buf ( n181173 , n13805 );
buf ( n181174 , n181173 );
nand ( n13808 , n181169 , n181174 );
buf ( n181176 , n13808 );
buf ( n181177 , n181176 );
nand ( n13811 , n13801 , n181177 );
buf ( n181179 , n13811 );
xor ( n13813 , n181163 , n181179 );
buf ( n181181 , n13813 );
not ( n13815 , n181181 );
or ( n13816 , n13780 , n13815 );
buf ( n181184 , n13813 );
buf ( n181185 , n181145 );
or ( n13819 , n181184 , n181185 );
nand ( n13820 , n13816 , n13819 );
buf ( n181188 , n13820 );
buf ( n181189 , n181188 );
xor ( n13823 , n181126 , n181189 );
buf ( n181191 , n180746 );
not ( n13825 , n181191 );
buf ( n181193 , n169241 );
not ( n13827 , n181193 );
or ( n13828 , n13825 , n13827 );
buf ( n181196 , n169931 );
buf ( n181197 , n775 );
buf ( n181198 , n814 );
xor ( n13832 , n181197 , n181198 );
buf ( n181200 , n13832 );
buf ( n181201 , n181200 );
nand ( n13835 , n181196 , n181201 );
buf ( n181203 , n13835 );
buf ( n181204 , n181203 );
nand ( n13838 , n13828 , n181204 );
buf ( n181206 , n13838 );
buf ( n181207 , n180844 );
not ( n13841 , n181207 );
buf ( n181209 , n168750 );
not ( n13843 , n181209 );
or ( n13844 , n13841 , n13843 );
buf ( n181212 , n168759 );
xor ( n13846 , n804 , n785 );
buf ( n181214 , n13846 );
nand ( n13848 , n181212 , n181214 );
buf ( n181216 , n13848 );
buf ( n181217 , n181216 );
nand ( n13851 , n13844 , n181217 );
buf ( n181219 , n13851 );
buf ( n181220 , n181219 );
not ( n13854 , n181220 );
buf ( n181222 , n13854 );
xor ( n13856 , n181206 , n181222 );
buf ( n181224 , n180768 );
not ( n13858 , n181224 );
buf ( n181226 , n168861 );
not ( n13860 , n181226 );
or ( n13861 , n13858 , n13860 );
buf ( n181229 , n168870 );
xor ( n13863 , n802 , n787 );
buf ( n181231 , n13863 );
nand ( n13865 , n181229 , n181231 );
buf ( n181233 , n13865 );
buf ( n181234 , n181233 );
nand ( n13868 , n13861 , n181234 );
buf ( n181236 , n13868 );
xnor ( n13870 , n13856 , n181236 );
buf ( n181238 , n13870 );
xor ( n13872 , n13823 , n181238 );
buf ( n181240 , n13872 );
buf ( n181241 , n181240 );
xor ( n13875 , n180909 , n180945 );
and ( n13876 , n13875 , n180952 );
and ( n13877 , n180909 , n180945 );
or ( n13878 , n13876 , n13877 );
buf ( n181246 , n13878 );
buf ( n181247 , n181246 );
xor ( n13881 , n181241 , n181247 );
xor ( n13882 , n180864 , n180865 );
and ( n13883 , n13882 , n180883 );
and ( n13884 , n180864 , n180865 );
or ( n13885 , n13883 , n13884 );
buf ( n181253 , n13885 );
buf ( n181254 , n181253 );
xor ( n13888 , n180920 , n180935 );
and ( n13889 , n13888 , n180942 );
and ( n13890 , n180920 , n180935 );
or ( n13891 , n13889 , n13890 );
buf ( n181259 , n13891 );
buf ( n181260 , n181259 );
xor ( n13894 , n181254 , n181260 );
buf ( n181262 , n13458 );
not ( n13896 , n181262 );
buf ( n181264 , n2108 );
not ( n13898 , n181264 );
or ( n13899 , n13896 , n13898 );
buf ( n181267 , n168656 );
buf ( n181268 , n769 );
buf ( n181269 , n820 );
xor ( n13903 , n181268 , n181269 );
buf ( n181271 , n13903 );
buf ( n181272 , n181271 );
nand ( n13906 , n181267 , n181272 );
buf ( n181274 , n13906 );
buf ( n181275 , n181274 );
nand ( n13909 , n13899 , n181275 );
buf ( n181277 , n13909 );
buf ( n181278 , n181277 );
not ( n13912 , n181278 );
buf ( n181280 , n13912 );
buf ( n181281 , n181280 );
xor ( n13915 , n180636 , n180653 );
and ( n13916 , n13915 , n180676 );
and ( n13917 , n180636 , n180653 );
or ( n13918 , n13916 , n13917 );
buf ( n181286 , n13918 );
buf ( n181287 , n181286 );
xor ( n13921 , n181281 , n181287 );
xor ( n13922 , n180822 , n180833 );
and ( n13923 , n13922 , n180851 );
and ( n13924 , n180822 , n180833 );
or ( n13925 , n13923 , n13924 );
buf ( n181293 , n13925 );
buf ( n181294 , n181293 );
xor ( n13928 , n13921 , n181294 );
buf ( n181296 , n13928 );
buf ( n181297 , n181296 );
xor ( n13931 , n13894 , n181297 );
buf ( n181299 , n13931 );
buf ( n181300 , n181299 );
xor ( n13934 , n13881 , n181300 );
buf ( n181302 , n13934 );
buf ( n181303 , n181302 );
buf ( n181304 , n180798 );
not ( n13938 , n181304 );
buf ( n181306 , n180752 );
not ( n13940 , n181306 );
or ( n13941 , n13938 , n13940 );
buf ( n181309 , n180752 );
buf ( n181310 , n180798 );
or ( n13944 , n181309 , n181310 );
buf ( n181312 , n180774 );
nand ( n13946 , n13944 , n181312 );
buf ( n181314 , n13946 );
buf ( n181315 , n181314 );
nand ( n13949 , n13941 , n181315 );
buf ( n181317 , n13949 );
not ( n13951 , n180722 );
nand ( n13952 , n13951 , n13354 );
not ( n13953 , n13952 );
not ( n13954 , n180713 );
or ( n13955 , n13953 , n13954 );
nand ( n13956 , n13955 , n13359 );
and ( n13957 , n181317 , n13956 );
not ( n13958 , n181317 );
and ( n13959 , n180713 , n13952 );
nor ( n13960 , n13959 , n13360 );
and ( n13961 , n13958 , n13960 );
nor ( n13962 , n13957 , n13961 );
buf ( n181330 , n13962 );
buf ( n181331 , n791 );
buf ( n181332 , n800 );
nand ( n13966 , n181331 , n181332 );
buf ( n181334 , n13966 );
buf ( n181335 , n181334 );
not ( n13969 , n181335 );
buf ( n181337 , n13969 );
buf ( n181338 , n181337 );
buf ( n181339 , n180690 );
not ( n13976 , n181339 );
buf ( n181341 , n171706 );
not ( n13978 , n181341 );
or ( n13979 , n13976 , n13978 );
buf ( n181344 , n168806 );
buf ( n181345 , n771 );
buf ( n181346 , n818 );
xor ( n13983 , n181345 , n181346 );
buf ( n181348 , n13983 );
buf ( n181349 , n181348 );
nand ( n13986 , n181344 , n181349 );
buf ( n181351 , n13986 );
buf ( n181352 , n181351 );
nand ( n13989 , n13979 , n181352 );
buf ( n181354 , n13989 );
buf ( n181355 , n181354 );
xor ( n13992 , n181338 , n181355 );
buf ( n181357 , n180646 );
not ( n13994 , n181357 );
buf ( n181359 , n178360 );
not ( n13996 , n181359 );
or ( n13997 , n13994 , n13996 );
buf ( n181362 , n172582 );
buf ( n181363 , n779 );
buf ( n181364 , n810 );
xor ( n14001 , n181363 , n181364 );
buf ( n181366 , n14001 );
buf ( n181367 , n181366 );
nand ( n14004 , n181362 , n181367 );
buf ( n181369 , n14004 );
buf ( n181370 , n181369 );
nand ( n14007 , n13997 , n181370 );
buf ( n181372 , n14007 );
buf ( n181373 , n181372 );
xnor ( n14010 , n13992 , n181373 );
buf ( n181375 , n14010 );
buf ( n181376 , n181375 );
not ( n14013 , n181376 );
buf ( n181378 , n14013 );
buf ( n181379 , n181378 );
and ( n14016 , n181330 , n181379 );
not ( n14017 , n181330 );
buf ( n181382 , n181375 );
and ( n14019 , n14017 , n181382 );
nor ( n14020 , n14016 , n14019 );
buf ( n181385 , n14020 );
buf ( n181386 , n181385 );
buf ( n181387 , n180853 );
buf ( n181388 , n180885 );
or ( n14025 , n181387 , n181388 );
not ( n14026 , n13435 );
buf ( n181391 , n14026 );
nand ( n14028 , n14025 , n181391 );
buf ( n181393 , n14028 );
buf ( n181394 , n181393 );
buf ( n181395 , n180853 );
buf ( n181396 , n180885 );
nand ( n14033 , n181395 , n181396 );
buf ( n181398 , n14033 );
buf ( n181399 , n181398 );
nand ( n14036 , n181394 , n181399 );
buf ( n181401 , n14036 );
buf ( n181402 , n181401 );
xor ( n14039 , n181386 , n181402 );
xor ( n14040 , n180619 , n180679 );
and ( n14041 , n14040 , n180733 );
and ( n14042 , n180619 , n180679 );
or ( n14043 , n14041 , n14042 );
buf ( n181408 , n14043 );
buf ( n181409 , n181408 );
xor ( n14046 , n14039 , n181409 );
buf ( n181411 , n14046 );
xor ( n14048 , n180613 , n180735 );
and ( n14049 , n14048 , n180895 );
and ( n14050 , n180613 , n180735 );
or ( n14051 , n14049 , n14050 );
xor ( n14052 , n181411 , n14051 );
xor ( n14053 , n180903 , n180955 );
and ( n14054 , n14053 , n180962 );
and ( n14055 , n180903 , n180955 );
or ( n14056 , n14054 , n14055 );
buf ( n181421 , n14056 );
xor ( n14058 , n14052 , n181421 );
buf ( n181423 , n14058 );
xor ( n14060 , n181303 , n181423 );
xor ( n14061 , n180608 , n13526 );
and ( n14062 , n14061 , n180964 );
and ( n14063 , n180608 , n13526 );
or ( n14064 , n14062 , n14063 );
buf ( n181429 , n14064 );
xor ( n14066 , n14060 , n181429 );
buf ( n181431 , n14066 );
xor ( n14068 , n180596 , n180602 );
and ( n14069 , n14068 , n180966 );
and ( n14070 , n180596 , n180602 );
or ( n14071 , n14069 , n14070 );
buf ( n181436 , n14071 );
and ( n14073 , n181431 , n181436 );
not ( n14074 , n14073 );
xor ( n14075 , n181254 , n181260 );
and ( n14076 , n14075 , n181297 );
and ( n14077 , n181254 , n181260 );
or ( n14078 , n14076 , n14077 );
buf ( n181443 , n14078 );
buf ( n181444 , n181443 );
not ( n14081 , n181444 );
buf ( n181446 , n13846 );
not ( n14083 , n181446 );
buf ( n181448 , n1578 );
not ( n14085 , n181448 );
or ( n14086 , n14083 , n14085 );
buf ( n181451 , n168759 );
xor ( n14088 , n804 , n784 );
buf ( n181453 , n14088 );
nand ( n14090 , n181451 , n181453 );
buf ( n181455 , n14090 );
buf ( n181456 , n181455 );
nand ( n14093 , n14086 , n181456 );
buf ( n181458 , n14093 );
buf ( n181459 , n13863 );
not ( n14096 , n181459 );
buf ( n181461 , n178232 );
not ( n14098 , n181461 );
or ( n14099 , n14096 , n14098 );
buf ( n181464 , n168867 );
xor ( n14101 , n802 , n786 );
buf ( n181466 , n14101 );
nand ( n14103 , n181464 , n181466 );
buf ( n181468 , n14103 );
buf ( n181469 , n181468 );
nand ( n14106 , n14099 , n181469 );
buf ( n181471 , n14106 );
xor ( n14108 , n181458 , n181471 );
buf ( n181473 , n181348 );
not ( n14110 , n181473 );
buf ( n181475 , n1321 );
not ( n14112 , n181475 );
or ( n14113 , n14110 , n14112 );
buf ( n181478 , n168806 );
buf ( n181479 , n770 );
buf ( n181480 , n818 );
xor ( n14117 , n181479 , n181480 );
buf ( n181482 , n14117 );
buf ( n181483 , n181482 );
nand ( n14120 , n181478 , n181483 );
buf ( n181485 , n14120 );
buf ( n181486 , n181485 );
nand ( n14123 , n14113 , n181486 );
buf ( n181488 , n14123 );
not ( n14125 , n181488 );
xor ( n14126 , n14108 , n14125 );
buf ( n181491 , n181271 );
not ( n14128 , n181491 );
buf ( n181493 , n2251 );
not ( n14130 , n181493 );
or ( n14131 , n14128 , n14130 );
buf ( n181496 , n768 );
buf ( n181497 , n820 );
xor ( n14134 , n181496 , n181497 );
buf ( n181499 , n14134 );
buf ( n181500 , n181499 );
buf ( n181501 , n168656 );
nand ( n14138 , n181500 , n181501 );
buf ( n181503 , n14138 );
buf ( n181504 , n181503 );
nand ( n14141 , n14131 , n181504 );
buf ( n181506 , n14141 );
buf ( n181507 , n169420 );
not ( n14144 , n181507 );
buf ( n181509 , n2418 );
not ( n14146 , n181509 );
buf ( n181511 , n14146 );
buf ( n181512 , n181511 );
not ( n14149 , n181512 );
or ( n14150 , n14144 , n14149 );
buf ( n181515 , n822 );
nand ( n14152 , n14150 , n181515 );
buf ( n181517 , n14152 );
xor ( n14154 , n181506 , n181517 );
buf ( n181519 , n181173 );
not ( n14156 , n181519 );
buf ( n181521 , n169836 );
not ( n14158 , n181521 );
or ( n14159 , n14156 , n14158 );
buf ( n181524 , n169320 );
buf ( n181525 , n772 );
buf ( n181526 , n816 );
xor ( n14163 , n181525 , n181526 );
buf ( n181528 , n14163 );
buf ( n181529 , n181528 );
nand ( n14166 , n181524 , n181529 );
buf ( n181531 , n14166 );
buf ( n181532 , n181531 );
nand ( n14169 , n14159 , n181532 );
buf ( n181534 , n14169 );
xor ( n14171 , n14154 , n181534 );
xor ( n14172 , n14126 , n14171 );
buf ( n181537 , n181157 );
not ( n14174 , n181537 );
buf ( n181539 , n177984 );
not ( n14176 , n181539 );
or ( n14177 , n14174 , n14176 );
buf ( n181542 , n168619 );
buf ( n181543 , n780 );
buf ( n181544 , n808 );
xor ( n14181 , n181543 , n181544 );
buf ( n181546 , n14181 );
buf ( n181547 , n181546 );
nand ( n14184 , n181542 , n181547 );
buf ( n181549 , n14184 );
buf ( n181550 , n181549 );
nand ( n14187 , n14177 , n181550 );
buf ( n181552 , n14187 );
buf ( n181553 , n181552 );
not ( n14190 , n181553 );
buf ( n181555 , n14190 );
buf ( n181556 , n181555 );
buf ( n181557 , n181200 );
not ( n14194 , n181557 );
buf ( n181559 , n169922 );
not ( n14196 , n181559 );
or ( n14197 , n14194 , n14196 );
buf ( n181562 , n169250 );
buf ( n181563 , n774 );
buf ( n181564 , n814 );
xor ( n14201 , n181563 , n181564 );
buf ( n181566 , n14201 );
buf ( n181567 , n181566 );
nand ( n14204 , n181562 , n181567 );
buf ( n181569 , n14204 );
buf ( n181570 , n181569 );
nand ( n14207 , n14197 , n181570 );
buf ( n181572 , n14207 );
buf ( n181573 , n181572 );
and ( n14210 , n181556 , n181573 );
not ( n14211 , n181556 );
buf ( n181576 , n181572 );
not ( n14213 , n181576 );
buf ( n181578 , n14213 );
buf ( n181579 , n181578 );
and ( n14216 , n14211 , n181579 );
or ( n14217 , n14210 , n14216 );
buf ( n181582 , n14217 );
buf ( n181583 , n181582 );
buf ( n181584 , n181136 );
not ( n14221 , n181584 );
buf ( n181586 , n168713 );
buf ( n14223 , n181586 );
buf ( n181588 , n14223 );
buf ( n181589 , n181588 );
not ( n14226 , n181589 );
or ( n14227 , n14221 , n14226 );
buf ( n181592 , n2823 );
buf ( n14229 , n181592 );
buf ( n181594 , n14229 );
buf ( n181595 , n181594 );
buf ( n181596 , n782 );
buf ( n181597 , n806 );
xor ( n14234 , n181596 , n181597 );
buf ( n181599 , n14234 );
buf ( n181600 , n181599 );
nand ( n14237 , n181595 , n181600 );
buf ( n181602 , n14237 );
buf ( n181603 , n181602 );
nand ( n14240 , n14227 , n181603 );
buf ( n181605 , n14240 );
buf ( n181606 , n181605 );
xnor ( n14243 , n181583 , n181606 );
buf ( n181608 , n14243 );
xnor ( n14245 , n14172 , n181608 );
buf ( n181610 , n14245 );
not ( n14247 , n181610 );
and ( n14248 , n14081 , n14247 );
buf ( n181613 , n181443 );
buf ( n181614 , n14245 );
and ( n14251 , n181613 , n181614 );
nor ( n14252 , n14248 , n14251 );
buf ( n181617 , n14252 );
buf ( n181618 , n181617 );
buf ( n181619 , n790 );
buf ( n181620 , n800 );
and ( n14257 , n181619 , n181620 );
buf ( n181622 , n14257 );
buf ( n181623 , n181622 );
buf ( n181624 , n181087 );
not ( n14261 , n181624 );
buf ( n181626 , n3497 );
not ( n14263 , n181626 );
or ( n14264 , n14261 , n14263 );
xor ( n14265 , n800 , n788 );
nand ( n14266 , n170972 , n14265 );
buf ( n181631 , n14266 );
nand ( n14268 , n14264 , n181631 );
buf ( n181633 , n14268 );
buf ( n181634 , n181633 );
xor ( n14271 , n181623 , n181634 );
buf ( n181636 , n181116 );
not ( n14273 , n181636 );
buf ( n181638 , n1907 );
not ( n14275 , n181638 );
or ( n14276 , n14273 , n14275 );
buf ( n14277 , n1534 );
buf ( n181642 , n14277 );
buf ( n181643 , n776 );
buf ( n181644 , n812 );
xor ( n14281 , n181643 , n181644 );
buf ( n181646 , n14281 );
buf ( n181647 , n181646 );
nand ( n14284 , n181642 , n181647 );
buf ( n181649 , n14284 );
buf ( n181650 , n181649 );
nand ( n14287 , n14276 , n181650 );
buf ( n181652 , n14287 );
buf ( n181653 , n181652 );
xor ( n14290 , n14271 , n181653 );
buf ( n181655 , n14290 );
buf ( n181656 , n181219 );
not ( n14293 , n181656 );
buf ( n181658 , n181206 );
not ( n14298 , n181658 );
or ( n14299 , n14293 , n14298 );
buf ( n181661 , n181222 );
not ( n14301 , n181661 );
buf ( n181663 , n181206 );
not ( n14303 , n181663 );
buf ( n181665 , n14303 );
buf ( n181666 , n181665 );
not ( n14306 , n181666 );
or ( n14307 , n14301 , n14306 );
buf ( n181669 , n181236 );
nand ( n14309 , n14307 , n181669 );
buf ( n181671 , n14309 );
buf ( n181672 , n181671 );
nand ( n14312 , n14299 , n181672 );
buf ( n181674 , n14312 );
buf ( n181675 , n181674 );
not ( n14315 , n181675 );
buf ( n181677 , n181277 );
not ( n14317 , n181677 );
buf ( n181679 , n181366 );
not ( n14319 , n181679 );
buf ( n181681 , n169951 );
not ( n14321 , n181681 );
or ( n14322 , n14319 , n14321 );
buf ( n181684 , n170708 );
buf ( n181685 , n778 );
buf ( n181686 , n810 );
xor ( n14326 , n181685 , n181686 );
buf ( n181688 , n14326 );
buf ( n181689 , n181688 );
nand ( n14329 , n181684 , n181689 );
buf ( n181691 , n14329 );
buf ( n181692 , n181691 );
nand ( n14332 , n14322 , n181692 );
buf ( n181694 , n14332 );
buf ( n181695 , n181694 );
not ( n14335 , n181695 );
buf ( n181697 , n14335 );
buf ( n181698 , n181697 );
not ( n14338 , n181698 );
and ( n14339 , n14317 , n14338 );
buf ( n181701 , n181277 );
buf ( n181702 , n181697 );
and ( n14342 , n181701 , n181702 );
nor ( n14343 , n14339 , n14342 );
buf ( n181705 , n14343 );
buf ( n181706 , n181705 );
not ( n14346 , n181706 );
and ( n14347 , n14315 , n14346 );
buf ( n181709 , n181674 );
buf ( n181710 , n181705 );
and ( n14350 , n181709 , n181710 );
nor ( n14351 , n14347 , n14350 );
buf ( n181713 , n14351 );
xor ( n14353 , n181655 , n181713 );
xor ( n14354 , n181281 , n181287 );
and ( n14355 , n14354 , n181294 );
and ( n14356 , n181281 , n181287 );
or ( n14357 , n14355 , n14356 );
buf ( n181719 , n14357 );
xor ( n14359 , n14353 , n181719 );
not ( n14360 , n14359 );
buf ( n14361 , n14360 );
not ( n14362 , n14361 );
buf ( n181724 , n14362 );
and ( n14364 , n181618 , n181724 );
not ( n14365 , n181618 );
buf ( n181727 , n14361 );
and ( n14367 , n14365 , n181727 );
nor ( n14368 , n14364 , n14367 );
buf ( n181730 , n14368 );
buf ( n181731 , n181730 );
not ( n14371 , n181378 );
not ( n14372 , n13956 );
or ( n14373 , n14371 , n14372 );
not ( n14374 , n181375 );
not ( n14375 , n13960 );
or ( n14376 , n14374 , n14375 );
nand ( n14377 , n14376 , n181317 );
nand ( n14378 , n14373 , n14377 );
buf ( n181740 , n14378 );
not ( n14380 , n181354 );
nand ( n14381 , n14380 , n181334 );
not ( n14382 , n14381 );
not ( n14383 , n181372 );
or ( n14384 , n14382 , n14383 );
buf ( n181746 , n181354 );
buf ( n181747 , n181337 );
nand ( n14387 , n181746 , n181747 );
buf ( n181749 , n14387 );
nand ( n14389 , n14384 , n181749 );
buf ( n181751 , n14389 );
buf ( n181752 , n181163 );
buf ( n181753 , n181142 );
or ( n14393 , n181752 , n181753 );
buf ( n181755 , n181179 );
nand ( n14395 , n14393 , n181755 );
buf ( n181757 , n14395 );
buf ( n181758 , n181757 );
buf ( n181759 , n181163 );
buf ( n181760 , n181142 );
nand ( n14400 , n181759 , n181760 );
buf ( n181762 , n14400 );
buf ( n181763 , n181762 );
nand ( n14403 , n181758 , n181763 );
buf ( n181765 , n14403 );
buf ( n181766 , n181765 );
xor ( n14406 , n181751 , n181766 );
xor ( n14407 , n181092 , n181105 );
and ( n14408 , n14407 , n181123 );
and ( n14409 , n181092 , n181105 );
or ( n14410 , n14408 , n14409 );
buf ( n181772 , n14410 );
buf ( n181773 , n181772 );
xor ( n14413 , n14406 , n181773 );
buf ( n181775 , n14413 );
buf ( n181776 , n181775 );
xor ( n14416 , n181740 , n181776 );
xor ( n14417 , n181126 , n181189 );
and ( n14418 , n14417 , n181238 );
and ( n14419 , n181126 , n181189 );
or ( n14420 , n14418 , n14419 );
buf ( n181782 , n14420 );
buf ( n181783 , n181782 );
xor ( n14423 , n14416 , n181783 );
buf ( n181785 , n14423 );
buf ( n181786 , n181785 );
xor ( n14426 , n181386 , n181402 );
and ( n14427 , n14426 , n181409 );
and ( n14428 , n181386 , n181402 );
or ( n14429 , n14427 , n14428 );
buf ( n181791 , n14429 );
buf ( n181792 , n181791 );
xor ( n14432 , n181786 , n181792 );
xor ( n14433 , n181241 , n181247 );
and ( n14434 , n14433 , n181300 );
and ( n14435 , n181241 , n181247 );
or ( n14436 , n14434 , n14435 );
buf ( n181798 , n14436 );
buf ( n181799 , n181798 );
xor ( n14439 , n14432 , n181799 );
buf ( n181801 , n14439 );
buf ( n181802 , n181801 );
xor ( n14442 , n181731 , n181802 );
xor ( n14443 , n181411 , n14051 );
and ( n14444 , n14443 , n181421 );
and ( n14445 , n181411 , n14051 );
or ( n14446 , n14444 , n14445 );
buf ( n181808 , n14446 );
xor ( n14448 , n14442 , n181808 );
buf ( n181810 , n14448 );
buf ( n181811 , n181810 );
not ( n14451 , n181811 );
buf ( n181813 , n14451 );
buf ( n181814 , n181813 );
not ( n14454 , n181814 );
xor ( n14455 , n181303 , n181423 );
and ( n14456 , n14455 , n181429 );
and ( n14457 , n181303 , n181423 );
or ( n14458 , n14456 , n14457 );
buf ( n181820 , n14458 );
buf ( n181821 , n181820 );
not ( n14461 , n181821 );
or ( n14462 , n14454 , n14461 );
buf ( n181824 , n181820 );
not ( n14464 , n181824 );
buf ( n181826 , n14464 );
buf ( n181827 , n181826 );
buf ( n181828 , n181810 );
nand ( n14468 , n181827 , n181828 );
buf ( n181830 , n14468 );
buf ( n181831 , n181830 );
nand ( n14471 , n14462 , n181831 );
buf ( n181833 , n14471 );
not ( n14473 , n181833 );
and ( n14474 , n14074 , n14473 );
buf ( n181836 , n181436 );
not ( n14476 , n181836 );
not ( n14477 , n181431 );
buf ( n181839 , n14477 );
not ( n14479 , n181839 );
or ( n14480 , n14476 , n14479 );
buf ( n181842 , n181436 );
not ( n14482 , n181842 );
buf ( n181844 , n14482 );
buf ( n181845 , n181844 );
buf ( n181846 , n181431 );
nand ( n14486 , n181845 , n181846 );
buf ( n181848 , n14486 );
buf ( n181849 , n181848 );
nand ( n14489 , n14480 , n181849 );
buf ( n181851 , n14489 );
buf ( n181852 , n181851 );
buf ( n181853 , n180968 );
buf ( n181854 , n13215 );
and ( n14494 , n181853 , n181854 );
buf ( n181856 , n14494 );
buf ( n181857 , n181856 );
nor ( n14497 , n181852 , n181857 );
buf ( n181859 , n14497 );
nor ( n14499 , n14474 , n181859 );
buf ( n181861 , n14499 );
buf ( n181862 , n14101 );
not ( n14502 , n181862 );
buf ( n181864 , n168861 );
not ( n14504 , n181864 );
or ( n14505 , n14502 , n14504 );
buf ( n181867 , n168870 );
buf ( n181868 , n785 );
buf ( n181869 , n802 );
xor ( n14509 , n181868 , n181869 );
buf ( n181871 , n14509 );
buf ( n181872 , n181871 );
nand ( n14512 , n181867 , n181872 );
buf ( n181874 , n14512 );
buf ( n181875 , n181874 );
nand ( n14515 , n14505 , n181875 );
buf ( n181877 , n14515 );
buf ( n181878 , n181877 );
not ( n14518 , n14265 );
not ( n14519 , n177819 );
or ( n14520 , n14518 , n14519 );
buf ( n181882 , n170972 );
buf ( n181883 , n787 );
buf ( n181884 , n800 );
xor ( n14524 , n181883 , n181884 );
buf ( n181886 , n14524 );
buf ( n181887 , n181886 );
nand ( n14527 , n181882 , n181887 );
buf ( n181889 , n14527 );
nand ( n14529 , n14520 , n181889 );
buf ( n181891 , n14529 );
xor ( n14531 , n181878 , n181891 );
buf ( n181893 , n181646 );
not ( n14533 , n181893 );
buf ( n181895 , n1907 );
not ( n14535 , n181895 );
or ( n14536 , n14533 , n14535 );
not ( n14537 , n1535 );
not ( n14538 , n14537 );
buf ( n181900 , n14538 );
buf ( n181901 , n775 );
buf ( n181902 , n812 );
xor ( n14542 , n181901 , n181902 );
buf ( n181904 , n14542 );
buf ( n181905 , n181904 );
nand ( n14545 , n181900 , n181905 );
buf ( n181907 , n14545 );
buf ( n181908 , n181907 );
nand ( n14548 , n14536 , n181908 );
buf ( n181910 , n14548 );
buf ( n181911 , n181910 );
xor ( n14551 , n14531 , n181911 );
buf ( n181913 , n14551 );
buf ( n181914 , n181913 );
buf ( n181915 , n181546 );
not ( n14555 , n181915 );
buf ( n181917 , n177984 );
not ( n14557 , n181917 );
or ( n14558 , n14555 , n14557 );
buf ( n181920 , n168619 );
buf ( n181921 , n779 );
buf ( n181922 , n808 );
xor ( n14562 , n181921 , n181922 );
buf ( n181924 , n14562 );
buf ( n181925 , n181924 );
nand ( n14565 , n181920 , n181925 );
buf ( n181927 , n14565 );
buf ( n181928 , n181927 );
nand ( n14568 , n14558 , n181928 );
buf ( n181930 , n14568 );
buf ( n181931 , n181930 );
buf ( n181932 , n181688 );
not ( n14572 , n181932 );
buf ( n181934 , n180199 );
not ( n14574 , n181934 );
or ( n14575 , n14572 , n14574 );
buf ( n181937 , n172582 );
buf ( n181938 , n777 );
buf ( n181939 , n810 );
xor ( n14579 , n181938 , n181939 );
buf ( n181941 , n14579 );
buf ( n181942 , n181941 );
nand ( n14582 , n181937 , n181942 );
buf ( n181944 , n14582 );
buf ( n181945 , n181944 );
nand ( n14585 , n14575 , n181945 );
buf ( n181947 , n14585 );
buf ( n181948 , n181947 );
xor ( n14588 , n181931 , n181948 );
buf ( n181950 , n181482 );
not ( n14590 , n181950 );
buf ( n181952 , n1321 );
not ( n14592 , n181952 );
or ( n14593 , n14590 , n14592 );
buf ( n181955 , n168806 );
buf ( n181956 , n769 );
buf ( n181957 , n818 );
xor ( n14597 , n181956 , n181957 );
buf ( n181959 , n14597 );
buf ( n181960 , n181959 );
nand ( n14600 , n181955 , n181960 );
buf ( n181962 , n14600 );
buf ( n181963 , n181962 );
nand ( n14603 , n14593 , n181963 );
buf ( n181965 , n14603 );
buf ( n181966 , n181965 );
not ( n14606 , n181966 );
buf ( n181968 , n14606 );
buf ( n181969 , n181968 );
xor ( n14612 , n14588 , n181969 );
buf ( n181971 , n14612 );
buf ( n181972 , n181971 );
xor ( n14615 , n181914 , n181972 );
xor ( n14616 , n181751 , n181766 );
and ( n14617 , n14616 , n181773 );
and ( n14618 , n181751 , n181766 );
or ( n14619 , n14617 , n14618 );
buf ( n181978 , n14619 );
buf ( n181979 , n181978 );
xor ( n14622 , n14615 , n181979 );
buf ( n181981 , n14622 );
buf ( n181982 , n181981 );
buf ( n14625 , n181982 );
buf ( n181984 , n14625 );
buf ( n181985 , n181984 );
not ( n14628 , n181985 );
buf ( n181987 , n181655 );
not ( n14630 , n181987 );
buf ( n181989 , n181713 );
not ( n14632 , n181989 );
buf ( n181991 , n14632 );
buf ( n181992 , n181991 );
not ( n14635 , n181992 );
or ( n14636 , n14630 , n14635 );
buf ( n181995 , n181655 );
not ( n14638 , n181995 );
buf ( n181997 , n14638 );
buf ( n181998 , n181997 );
not ( n14641 , n181998 );
buf ( n182000 , n181713 );
not ( n14643 , n182000 );
or ( n14644 , n14641 , n14643 );
buf ( n182003 , n181719 );
nand ( n14646 , n14644 , n182003 );
buf ( n182005 , n14646 );
buf ( n182006 , n182005 );
nand ( n14649 , n14636 , n182006 );
buf ( n182008 , n14649 );
buf ( n182009 , n182008 );
not ( n14652 , n182009 );
not ( n14653 , n181552 );
not ( n14654 , n181572 );
or ( n14655 , n14653 , n14654 );
buf ( n182014 , n181555 );
not ( n14657 , n182014 );
buf ( n182016 , n181578 );
not ( n14659 , n182016 );
or ( n14660 , n14657 , n14659 );
buf ( n182019 , n181605 );
nand ( n14662 , n14660 , n182019 );
buf ( n182021 , n14662 );
nand ( n14664 , n14655 , n182021 );
not ( n14665 , n14664 );
buf ( n182024 , n789 );
buf ( n182025 , n800 );
and ( n14668 , n182024 , n182025 );
buf ( n182027 , n14668 );
buf ( n182028 , n182027 );
buf ( n182029 , n181528 );
not ( n14672 , n182029 );
buf ( n182031 , n169836 );
not ( n14674 , n182031 );
or ( n14675 , n14672 , n14674 );
buf ( n182034 , n169320 );
buf ( n182035 , n771 );
buf ( n182036 , n816 );
xor ( n14679 , n182035 , n182036 );
buf ( n182038 , n14679 );
buf ( n182039 , n182038 );
nand ( n14682 , n182034 , n182039 );
buf ( n182041 , n14682 );
buf ( n182042 , n182041 );
nand ( n14685 , n14675 , n182042 );
buf ( n182044 , n14685 );
buf ( n182045 , n182044 );
xor ( n14688 , n182028 , n182045 );
buf ( n182047 , n181499 );
not ( n14690 , n182047 );
buf ( n182049 , n2251 );
not ( n14692 , n182049 );
or ( n14693 , n14690 , n14692 );
buf ( n182052 , n820 );
buf ( n182053 , n2513 );
nand ( n14696 , n182052 , n182053 );
buf ( n182055 , n14696 );
buf ( n182056 , n182055 );
nand ( n14699 , n14693 , n182056 );
buf ( n182058 , n14699 );
buf ( n182059 , n182058 );
xor ( n14702 , n14688 , n182059 );
buf ( n182061 , n14702 );
buf ( n182062 , n182061 );
not ( n14705 , n182062 );
buf ( n182064 , n14705 );
not ( n14707 , n182064 );
or ( n14708 , n14665 , n14707 );
not ( n14709 , n14664 );
nand ( n14710 , n14709 , n182061 );
nand ( n14711 , n14708 , n14710 );
not ( n14712 , n14088 );
not ( n14713 , n168832 );
or ( n14714 , n14712 , n14713 );
buf ( n182073 , n168838 );
buf ( n182074 , n783 );
buf ( n182075 , n804 );
xor ( n14718 , n182074 , n182075 );
buf ( n182077 , n14718 );
buf ( n182078 , n182077 );
nand ( n14721 , n182073 , n182078 );
buf ( n182080 , n14721 );
nand ( n14723 , n14714 , n182080 );
buf ( n182082 , n181599 );
not ( n14725 , n182082 );
buf ( n182084 , n168713 );
not ( n14727 , n182084 );
or ( n14728 , n14725 , n14727 );
buf ( n182087 , n2823 );
buf ( n182088 , n781 );
buf ( n182089 , n806 );
xor ( n14732 , n182088 , n182089 );
buf ( n182091 , n14732 );
buf ( n182092 , n182091 );
nand ( n14735 , n182087 , n182092 );
buf ( n182094 , n14735 );
buf ( n182095 , n182094 );
nand ( n14738 , n14728 , n182095 );
buf ( n182097 , n14738 );
xor ( n14740 , n14723 , n182097 );
buf ( n182099 , n181566 );
not ( n14742 , n182099 );
buf ( n182101 , n171013 );
not ( n14744 , n182101 );
or ( n14745 , n14742 , n14744 );
buf ( n182104 , n169250 );
buf ( n182105 , n773 );
buf ( n182106 , n814 );
xor ( n14749 , n182105 , n182106 );
buf ( n182108 , n14749 );
buf ( n182109 , n182108 );
nand ( n14752 , n182104 , n182109 );
buf ( n182111 , n14752 );
buf ( n182112 , n182111 );
nand ( n14755 , n14745 , n182112 );
buf ( n182114 , n14755 );
not ( n14757 , n182114 );
xor ( n14758 , n14740 , n14757 );
and ( n14759 , n14711 , n14758 );
not ( n14760 , n14711 );
not ( n182119 , n14758 );
and ( n14762 , n14760 , n182119 );
nor ( n14763 , n14759 , n14762 );
buf ( n182122 , n14763 );
not ( n14765 , n182122 );
and ( n14766 , n14652 , n14765 );
buf ( n182125 , n182008 );
buf ( n182126 , n14763 );
and ( n14769 , n182125 , n182126 );
nor ( n14770 , n14766 , n14769 );
buf ( n182129 , n14770 );
buf ( n182130 , n182129 );
not ( n14773 , n182130 );
or ( n14774 , n14628 , n14773 );
buf ( n182133 , n182129 );
buf ( n182134 , n181984 );
or ( n14777 , n182133 , n182134 );
nand ( n14778 , n14774 , n14777 );
buf ( n182137 , n14778 );
buf ( n182138 , n182137 );
xor ( n14781 , n181786 , n181792 );
and ( n14782 , n14781 , n181799 );
and ( n14783 , n181786 , n181792 );
or ( n14784 , n14782 , n14783 );
buf ( n182143 , n14784 );
buf ( n182144 , n182143 );
xor ( n14787 , n182138 , n182144 );
xor ( n14788 , n181740 , n181776 );
and ( n14789 , n14788 , n181783 );
and ( n14790 , n181740 , n181776 );
or ( n14791 , n14789 , n14790 );
buf ( n182150 , n14791 );
buf ( n182151 , n182150 );
buf ( n182152 , n181280 );
buf ( n182153 , n181697 );
nand ( n14796 , n182152 , n182153 );
buf ( n182155 , n14796 );
buf ( n182156 , n182155 );
not ( n14799 , n182156 );
buf ( n182158 , n181674 );
not ( n14801 , n182158 );
or ( n14802 , n14799 , n14801 );
buf ( n182161 , n181694 );
buf ( n182162 , n181277 );
nand ( n14805 , n182161 , n182162 );
buf ( n182164 , n14805 );
buf ( n182165 , n182164 );
nand ( n14808 , n14802 , n182165 );
buf ( n182167 , n14808 );
buf ( n182168 , n182167 );
not ( n14811 , n181488 );
buf ( n182170 , n181458 );
buf ( n182171 , n181471 );
or ( n14814 , n182170 , n182171 );
buf ( n182173 , n14814 );
not ( n14816 , n182173 );
or ( n14817 , n14811 , n14816 );
buf ( n182176 , n181458 );
buf ( n182177 , n181471 );
nand ( n14820 , n182176 , n182177 );
buf ( n182179 , n14820 );
nand ( n14822 , n14817 , n182179 );
buf ( n182181 , n14822 );
buf ( n182182 , n181517 );
not ( n14825 , n182182 );
buf ( n182184 , n181506 );
not ( n14827 , n182184 );
or ( n14828 , n14825 , n14827 );
buf ( n182187 , n181506 );
buf ( n182188 , n181517 );
or ( n14831 , n182187 , n182188 );
buf ( n182190 , n181534 );
nand ( n14833 , n14831 , n182190 );
buf ( n182192 , n14833 );
buf ( n182193 , n182192 );
nand ( n14836 , n14828 , n182193 );
buf ( n182195 , n14836 );
buf ( n182196 , n182195 );
xor ( n14839 , n182181 , n182196 );
xor ( n14840 , n181623 , n181634 );
and ( n14841 , n14840 , n181653 );
and ( n14842 , n181623 , n181634 );
or ( n14843 , n14841 , n14842 );
buf ( n182202 , n14843 );
buf ( n182203 , n182202 );
xor ( n14846 , n14839 , n182203 );
buf ( n182205 , n14846 );
buf ( n182206 , n182205 );
xor ( n14849 , n182168 , n182206 );
not ( n14850 , n14171 );
buf ( n182209 , n14126 );
not ( n14852 , n182209 );
buf ( n182211 , n14852 );
not ( n14854 , n182211 );
or ( n14855 , n14850 , n14854 );
buf ( n182214 , n14171 );
buf ( n182215 , n182211 );
nor ( n14858 , n182214 , n182215 );
buf ( n182217 , n14858 );
or ( n14860 , n181608 , n182217 );
nand ( n14861 , n14855 , n14860 );
buf ( n182220 , n14861 );
xor ( n14863 , n14849 , n182220 );
buf ( n182222 , n14863 );
buf ( n182223 , n182222 );
xor ( n14866 , n182151 , n182223 );
buf ( n182225 , n14245 );
not ( n14868 , n182225 );
buf ( n182227 , n14359 );
not ( n14870 , n182227 );
or ( n14871 , n14868 , n14870 );
buf ( n182230 , n181443 );
nand ( n14873 , n14871 , n182230 );
buf ( n182232 , n14873 );
buf ( n182233 , n182232 );
buf ( n182234 , n14360 );
buf ( n182235 , n14245 );
not ( n14878 , n182235 );
buf ( n182237 , n14878 );
buf ( n182238 , n182237 );
nand ( n14881 , n182234 , n182238 );
buf ( n182240 , n14881 );
buf ( n182241 , n182240 );
nand ( n14884 , n182233 , n182241 );
buf ( n182243 , n14884 );
buf ( n182244 , n182243 );
xor ( n14887 , n14866 , n182244 );
buf ( n182246 , n14887 );
buf ( n182247 , n182246 );
and ( n14890 , n14787 , n182247 );
and ( n14891 , n182138 , n182144 );
or ( n14892 , n14890 , n14891 );
buf ( n182251 , n14892 );
buf ( n182252 , n182251 );
not ( n14895 , n182252 );
buf ( n182254 , n14895 );
buf ( n182255 , n182254 );
not ( n14898 , n182255 );
buf ( n182257 , n182108 );
not ( n14900 , n182257 );
buf ( n182259 , n169241 );
not ( n14902 , n182259 );
or ( n14903 , n14900 , n14902 );
buf ( n182262 , n169250 );
buf ( n182263 , n772 );
buf ( n182264 , n814 );
xor ( n14907 , n182263 , n182264 );
buf ( n182266 , n14907 );
buf ( n182267 , n182266 );
nand ( n182268 , n182262 , n182267 );
buf ( n182269 , n182268 );
buf ( n182270 , n182269 );
nand ( n14916 , n14903 , n182270 );
buf ( n182272 , n14916 );
buf ( n182273 , n182272 );
buf ( n182274 , n181959 );
not ( n14920 , n182274 );
buf ( n182276 , n1321 );
not ( n14922 , n182276 );
or ( n14923 , n14920 , n14922 );
buf ( n182279 , n168806 );
buf ( n182280 , n768 );
buf ( n182281 , n818 );
xor ( n14927 , n182280 , n182281 );
buf ( n182283 , n14927 );
buf ( n182284 , n182283 );
nand ( n14930 , n182279 , n182284 );
buf ( n182286 , n14930 );
buf ( n182287 , n182286 );
nand ( n14933 , n14923 , n182287 );
buf ( n182289 , n14933 );
buf ( n182290 , n182289 );
xor ( n14936 , n182273 , n182290 );
buf ( n182292 , n2512 );
not ( n14938 , n182292 );
buf ( n182294 , n2251 );
not ( n14940 , n182294 );
buf ( n182296 , n14940 );
buf ( n182297 , n182296 );
not ( n14943 , n182297 );
or ( n14944 , n14938 , n14943 );
buf ( n182300 , n820 );
nand ( n14946 , n14944 , n182300 );
buf ( n182302 , n14946 );
buf ( n182303 , n182302 );
xor ( n14949 , n14936 , n182303 );
buf ( n182305 , n14949 );
buf ( n182306 , n182305 );
xor ( n14952 , n181931 , n181948 );
and ( n14953 , n14952 , n181969 );
and ( n14954 , n181931 , n181948 );
or ( n14955 , n14953 , n14954 );
buf ( n182311 , n14955 );
buf ( n182312 , n182311 );
xor ( n14958 , n182306 , n182312 );
not ( n14959 , n182077 );
not ( n14960 , n1578 );
or ( n14961 , n14959 , n14960 );
buf ( n182317 , n168838 );
buf ( n182318 , n782 );
buf ( n182319 , n804 );
xor ( n14965 , n182318 , n182319 );
buf ( n182321 , n14965 );
buf ( n182322 , n182321 );
nand ( n14968 , n182317 , n182322 );
buf ( n182324 , n14968 );
nand ( n14970 , n14961 , n182324 );
not ( n14971 , n182091 );
not ( n14972 , n168713 );
or ( n14973 , n14971 , n14972 );
buf ( n182329 , n168719 );
buf ( n182330 , n780 );
buf ( n182331 , n806 );
xor ( n14977 , n182330 , n182331 );
buf ( n182333 , n14977 );
buf ( n182334 , n182333 );
nand ( n14980 , n182329 , n182334 );
buf ( n182336 , n14980 );
nand ( n14982 , n14973 , n182336 );
xor ( n14983 , n14970 , n14982 );
not ( n14984 , n181904 );
not ( n14985 , n2757 );
or ( n14986 , n14984 , n14985 );
buf ( n182342 , n6287 );
buf ( n182343 , n774 );
buf ( n182344 , n812 );
xor ( n14990 , n182343 , n182344 );
buf ( n182346 , n14990 );
buf ( n182347 , n182346 );
nand ( n14993 , n182342 , n182347 );
buf ( n182349 , n14993 );
nand ( n14995 , n14986 , n182349 );
xor ( n14996 , n14983 , n14995 );
buf ( n182352 , n14996 );
xor ( n14998 , n14958 , n182352 );
buf ( n182354 , n14998 );
buf ( n182355 , n181941 );
not ( n15001 , n182355 );
buf ( n182357 , n178360 );
not ( n15003 , n182357 );
or ( n15004 , n15001 , n15003 );
buf ( n182360 , n172582 );
buf ( n182361 , n776 );
buf ( n182362 , n810 );
xor ( n15008 , n182361 , n182362 );
buf ( n182364 , n15008 );
buf ( n182365 , n182364 );
nand ( n15011 , n182360 , n182365 );
buf ( n182367 , n15011 );
buf ( n182368 , n182367 );
nand ( n15014 , n15004 , n182368 );
buf ( n182370 , n15014 );
buf ( n182371 , n182370 );
buf ( n182372 , n788 );
buf ( n182373 , n800 );
and ( n15019 , n182372 , n182373 );
buf ( n182375 , n15019 );
buf ( n182376 , n182375 );
and ( n15022 , n182371 , n182376 );
not ( n15023 , n182371 );
buf ( n182379 , n788 );
buf ( n182380 , n800 );
nand ( n15026 , n182379 , n182380 );
buf ( n182382 , n15026 );
buf ( n182383 , n182382 );
and ( n15029 , n15023 , n182383 );
nor ( n15030 , n15022 , n15029 );
buf ( n182386 , n15030 );
buf ( n182387 , n182386 );
buf ( n182388 , n181924 );
not ( n15034 , n182388 );
buf ( n182390 , n177984 );
not ( n15036 , n182390 );
or ( n15037 , n15034 , n15036 );
buf ( n182393 , n168619 );
buf ( n182394 , n778 );
buf ( n182395 , n808 );
xor ( n15041 , n182394 , n182395 );
buf ( n182397 , n15041 );
buf ( n182398 , n182397 );
nand ( n15044 , n182393 , n182398 );
buf ( n182400 , n15044 );
buf ( n182401 , n182400 );
nand ( n15047 , n15037 , n182401 );
buf ( n182403 , n15047 );
buf ( n182404 , n182403 );
not ( n15050 , n182404 );
buf ( n182406 , n15050 );
buf ( n182407 , n182406 );
and ( n15053 , n182387 , n182407 );
not ( n15054 , n182387 );
buf ( n182410 , n182403 );
and ( n15056 , n15054 , n182410 );
nor ( n15057 , n15053 , n15056 );
buf ( n182413 , n15057 );
buf ( n182414 , n182413 );
not ( n15060 , n182414 );
xor ( n15061 , n181878 , n181891 );
and ( n15062 , n15061 , n181911 );
and ( n15063 , n181878 , n181891 );
or ( n15064 , n15062 , n15063 );
buf ( n182420 , n15064 );
buf ( n182421 , n182420 );
not ( n15067 , n182421 );
or ( n15068 , n15060 , n15067 );
buf ( n182424 , n182420 );
buf ( n182425 , n182413 );
or ( n15071 , n182424 , n182425 );
nand ( n15072 , n15068 , n15071 );
buf ( n182428 , n15072 );
buf ( n182429 , n182428 );
buf ( n182430 , n182038 );
not ( n15076 , n182430 );
buf ( n182432 , n169836 );
not ( n15078 , n182432 );
or ( n15079 , n15076 , n15078 );
buf ( n182435 , n169845 );
xor ( n15081 , n816 , n770 );
buf ( n182437 , n15081 );
nand ( n15083 , n182435 , n182437 );
buf ( n182439 , n15083 );
buf ( n182440 , n182439 );
nand ( n15086 , n15079 , n182440 );
buf ( n182442 , n15086 );
buf ( n182443 , n181871 );
not ( n15089 , n182443 );
buf ( n182445 , n168861 );
not ( n15091 , n182445 );
or ( n15092 , n15089 , n15091 );
buf ( n182448 , n168870 );
buf ( n182449 , n784 );
buf ( n182450 , n802 );
xor ( n15096 , n182449 , n182450 );
buf ( n182452 , n15096 );
buf ( n182453 , n182452 );
nand ( n15099 , n182448 , n182453 );
buf ( n182455 , n15099 );
buf ( n182456 , n182455 );
nand ( n15102 , n15092 , n182456 );
buf ( n182458 , n15102 );
xor ( n15104 , n182442 , n182458 );
buf ( n182460 , n181886 );
not ( n15106 , n182460 );
buf ( n182462 , n3497 );
not ( n15108 , n182462 );
or ( n15109 , n15106 , n15108 );
buf ( n182465 , n170972 );
buf ( n182466 , n786 );
buf ( n182467 , n800 );
xor ( n15113 , n182466 , n182467 );
buf ( n182469 , n15113 );
buf ( n182470 , n182469 );
nand ( n15116 , n182465 , n182470 );
buf ( n182472 , n15116 );
buf ( n182473 , n182472 );
nand ( n15119 , n15109 , n182473 );
buf ( n182475 , n15119 );
xor ( n15121 , n15104 , n182475 );
buf ( n182477 , n15121 );
not ( n15123 , n182477 );
buf ( n182479 , n15123 );
buf ( n182480 , n182479 );
and ( n15126 , n182429 , n182480 );
not ( n15127 , n182429 );
buf ( n182483 , n15121 );
and ( n15129 , n15127 , n182483 );
nor ( n15130 , n15126 , n15129 );
buf ( n182486 , n15130 );
xor ( n15132 , n182354 , n182486 );
xor ( n15133 , n181914 , n181972 );
and ( n15134 , n15133 , n181979 );
and ( n15135 , n181914 , n181972 );
or ( n15136 , n15134 , n15135 );
buf ( n182492 , n15136 );
buf ( n182493 , n182492 );
not ( n15139 , n182493 );
buf ( n182495 , n15139 );
and ( n15141 , n15132 , n182495 );
not ( n15142 , n15132 );
and ( n15143 , n15142 , n182492 );
nor ( n15144 , n15141 , n15143 );
buf ( n182500 , n15144 );
xor ( n15146 , n182151 , n182223 );
and ( n15147 , n15146 , n182244 );
and ( n15148 , n182151 , n182223 );
or ( n15149 , n15147 , n15148 );
buf ( n182505 , n15149 );
buf ( n182506 , n182505 );
xor ( n15152 , n182500 , n182506 );
xor ( n15153 , n182168 , n182206 );
and ( n15154 , n15153 , n182220 );
and ( n15155 , n182168 , n182206 );
or ( n15156 , n15154 , n15155 );
buf ( n182512 , n15156 );
buf ( n182513 , n182512 );
xor ( n15159 , n182181 , n182196 );
and ( n15160 , n15159 , n182203 );
and ( n15161 , n182181 , n182196 );
or ( n15162 , n15160 , n15161 );
buf ( n182518 , n15162 );
buf ( n182519 , n182518 );
buf ( n182520 , n181965 );
xor ( n15166 , n182028 , n182045 );
and ( n15167 , n15166 , n182059 );
and ( n15168 , n182028 , n182045 );
or ( n15169 , n15167 , n15168 );
buf ( n182525 , n15169 );
buf ( n182526 , n182525 );
xor ( n15172 , n182520 , n182526 );
or ( n15173 , n14723 , n182114 );
nand ( n15174 , n15173 , n182097 );
buf ( n182530 , n15174 );
buf ( n182531 , n182114 );
buf ( n182532 , n14723 );
nand ( n15178 , n182531 , n182532 );
buf ( n182534 , n15178 );
buf ( n182535 , n182534 );
nand ( n15181 , n182530 , n182535 );
buf ( n182537 , n15181 );
buf ( n182538 , n182537 );
xor ( n15184 , n15172 , n182538 );
buf ( n182540 , n15184 );
buf ( n182541 , n182540 );
xor ( n15187 , n182519 , n182541 );
not ( n15188 , n14709 );
not ( n15189 , n182064 );
or ( n15190 , n15188 , n15189 );
nand ( n15191 , n15190 , n182119 );
buf ( n182547 , n15191 );
buf ( n182548 , n14709 );
not ( n15194 , n182548 );
buf ( n182550 , n182061 );
nand ( n15196 , n15194 , n182550 );
buf ( n182552 , n15196 );
buf ( n182553 , n182552 );
nand ( n15199 , n182547 , n182553 );
buf ( n182555 , n15199 );
buf ( n182556 , n182555 );
xor ( n15202 , n15187 , n182556 );
buf ( n182558 , n15202 );
buf ( n182559 , n182558 );
xor ( n15208 , n182513 , n182559 );
not ( n15209 , n14763 );
nor ( n15210 , n15209 , n181981 );
buf ( n182563 , n15210 );
buf ( n182564 , n182008 );
not ( n15213 , n182564 );
buf ( n182566 , n15213 );
buf ( n182567 , n182566 );
or ( n15216 , n182563 , n182567 );
buf ( n182569 , n181981 );
buf ( n182570 , n15209 );
nand ( n15219 , n182569 , n182570 );
buf ( n182572 , n15219 );
buf ( n182573 , n182572 );
nand ( n15222 , n15216 , n182573 );
buf ( n182575 , n15222 );
buf ( n182576 , n182575 );
xor ( n15225 , n15208 , n182576 );
buf ( n182578 , n15225 );
buf ( n182579 , n182578 );
xor ( n15228 , n15152 , n182579 );
buf ( n182581 , n15228 );
buf ( n182582 , n182581 );
not ( n15231 , n182582 );
or ( n15232 , n14898 , n15231 );
buf ( n182585 , n182254 );
buf ( n182586 , n182581 );
or ( n15235 , n182585 , n182586 );
nand ( n15236 , n15232 , n15235 );
buf ( n182589 , n15236 );
buf ( n182590 , n182589 );
not ( n15239 , n182590 );
xor ( n15240 , n182138 , n182144 );
xor ( n15241 , n15240 , n182247 );
buf ( n182594 , n15241 );
buf ( n182595 , n182594 );
xor ( n15244 , n181731 , n181802 );
and ( n15245 , n15244 , n181808 );
and ( n15246 , n181731 , n181802 );
or ( n15247 , n15245 , n15246 );
buf ( n182600 , n15247 );
buf ( n182601 , n182600 );
nand ( n15250 , n182595 , n182601 );
buf ( n182603 , n15250 );
buf ( n182604 , n182603 );
nand ( n15253 , n15239 , n182604 );
buf ( n182606 , n15253 );
buf ( n182607 , n182606 );
not ( n15256 , n182607 );
buf ( n182609 , n15256 );
buf ( n182610 , n182609 );
buf ( n182611 , n181820 );
buf ( n182612 , n181810 );
and ( n15261 , n182611 , n182612 );
buf ( n182614 , n15261 );
buf ( n182615 , n182614 );
buf ( n182616 , n182600 );
buf ( n182617 , n182594 );
and ( n15266 , n182616 , n182617 );
not ( n15267 , n182616 );
buf ( n182620 , n182594 );
not ( n15269 , n182620 );
buf ( n182622 , n15269 );
buf ( n182623 , n182622 );
and ( n15272 , n15267 , n182623 );
nor ( n15273 , n15266 , n15272 );
buf ( n182626 , n15273 );
buf ( n182627 , n182626 );
nor ( n15276 , n182615 , n182627 );
buf ( n182629 , n15276 );
buf ( n182630 , n182629 );
nor ( n15279 , n182610 , n182630 );
buf ( n182632 , n15279 );
buf ( n182633 , n182632 );
nand ( n15282 , n181861 , n182633 );
buf ( n182635 , n15282 );
buf ( n182636 , n182635 );
not ( n15285 , n182636 );
xor ( n15286 , n182500 , n182506 );
and ( n15287 , n15286 , n182579 );
and ( n15288 , n182500 , n182506 );
or ( n15289 , n15287 , n15288 );
buf ( n182642 , n15289 );
buf ( n182643 , n15121 );
buf ( n182644 , n182413 );
not ( n15293 , n182644 );
buf ( n182646 , n15293 );
buf ( n182647 , n182646 );
or ( n15296 , n182643 , n182647 );
buf ( n182649 , n182420 );
nand ( n15298 , n15296 , n182649 );
buf ( n182651 , n15298 );
buf ( n182652 , n182651 );
buf ( n182653 , n15121 );
buf ( n182654 , n182646 );
nand ( n15303 , n182653 , n182654 );
buf ( n182656 , n15303 );
buf ( n182657 , n182656 );
nand ( n15306 , n182652 , n182657 );
buf ( n182659 , n15306 );
buf ( n182660 , n182659 );
xor ( n15309 , n182306 , n182312 );
and ( n15310 , n15309 , n182352 );
and ( n15311 , n182306 , n182312 );
or ( n15312 , n15310 , n15311 );
buf ( n182665 , n15312 );
buf ( n182666 , n182665 );
xor ( n15315 , n182660 , n182666 );
buf ( n182668 , n787 );
buf ( n182669 , n800 );
and ( n15318 , n182668 , n182669 );
buf ( n182671 , n15318 );
buf ( n182672 , n182671 );
buf ( n182673 , n182364 );
not ( n15322 , n182673 );
buf ( n182675 , n178360 );
not ( n15324 , n182675 );
or ( n15325 , n15322 , n15324 );
buf ( n182678 , n170708 );
buf ( n182679 , n775 );
buf ( n182680 , n810 );
xor ( n15329 , n182679 , n182680 );
buf ( n182682 , n15329 );
buf ( n182683 , n182682 );
nand ( n15332 , n182678 , n182683 );
buf ( n182685 , n15332 );
buf ( n182686 , n182685 );
nand ( n15335 , n15325 , n182686 );
buf ( n182688 , n15335 );
buf ( n182689 , n182688 );
xor ( n15338 , n182672 , n182689 );
buf ( n182691 , n182469 );
not ( n15340 , n182691 );
buf ( n182693 , n3497 );
not ( n15342 , n182693 );
or ( n15343 , n15340 , n15342 );
buf ( n182696 , n170972 );
buf ( n182697 , n785 );
buf ( n182698 , n800 );
xor ( n182699 , n182697 , n182698 );
buf ( n182700 , n182699 );
buf ( n182701 , n182700 );
nand ( n15350 , n182696 , n182701 );
buf ( n182703 , n15350 );
buf ( n182704 , n182703 );
nand ( n15353 , n15343 , n182704 );
buf ( n182706 , n15353 );
buf ( n182707 , n182706 );
xor ( n15356 , n15338 , n182707 );
buf ( n182709 , n15356 );
buf ( n182710 , n182452 );
not ( n15359 , n182710 );
buf ( n182712 , n1389 );
not ( n15361 , n182712 );
or ( n15362 , n15359 , n15361 );
buf ( n182715 , n168867 );
buf ( n182716 , n783 );
buf ( n182717 , n802 );
xor ( n15366 , n182716 , n182717 );
buf ( n182719 , n15366 );
buf ( n182720 , n182719 );
nand ( n15369 , n182715 , n182720 );
buf ( n182722 , n15369 );
buf ( n182723 , n182722 );
nand ( n15372 , n15362 , n182723 );
buf ( n182725 , n15372 );
buf ( n182726 , n182725 );
buf ( n182727 , n182321 );
not ( n15376 , n182727 );
buf ( n182729 , n168750 );
not ( n15378 , n182729 );
or ( n15379 , n15376 , n15378 );
buf ( n182732 , n178447 );
buf ( n182733 , n781 );
buf ( n182734 , n804 );
xor ( n15383 , n182733 , n182734 );
buf ( n182736 , n15383 );
buf ( n182737 , n182736 );
nand ( n15386 , n182732 , n182737 );
buf ( n182739 , n15386 );
buf ( n182740 , n182739 );
nand ( n15389 , n15379 , n182740 );
buf ( n182742 , n15389 );
buf ( n182743 , n182742 );
xor ( n15392 , n182726 , n182743 );
buf ( n182745 , n182346 );
not ( n15394 , n182745 );
buf ( n182747 , n1907 );
not ( n15396 , n182747 );
or ( n15397 , n15394 , n15396 );
buf ( n182750 , n14277 );
buf ( n182751 , n773 );
buf ( n182752 , n812 );
xor ( n15401 , n182751 , n182752 );
buf ( n182754 , n15401 );
buf ( n182755 , n182754 );
nand ( n15404 , n182750 , n182755 );
buf ( n182757 , n15404 );
buf ( n182758 , n182757 );
nand ( n15407 , n15397 , n182758 );
buf ( n182760 , n15407 );
buf ( n182761 , n182760 );
xor ( n15410 , n15392 , n182761 );
buf ( n182763 , n15410 );
xor ( n15412 , n182709 , n182763 );
buf ( n182765 , n182266 );
not ( n15414 , n182765 );
buf ( n182767 , n171013 );
not ( n15416 , n182767 );
or ( n15417 , n15414 , n15416 );
buf ( n182770 , n169931 );
buf ( n182771 , n771 );
buf ( n182772 , n814 );
xor ( n15421 , n182771 , n182772 );
buf ( n182774 , n15421 );
buf ( n182775 , n182774 );
nand ( n15424 , n182770 , n182775 );
buf ( n182777 , n15424 );
buf ( n182778 , n182777 );
nand ( n15427 , n15417 , n182778 );
buf ( n182780 , n15427 );
buf ( n182781 , n182780 );
buf ( n182782 , n182397 );
not ( n15431 , n182782 );
buf ( n182784 , n177984 );
not ( n15433 , n182784 );
or ( n15434 , n15431 , n15433 );
buf ( n182787 , n2554 );
buf ( n182788 , n777 );
buf ( n182789 , n808 );
xor ( n15438 , n182788 , n182789 );
buf ( n182791 , n15438 );
buf ( n182792 , n182791 );
nand ( n15441 , n182787 , n182792 );
buf ( n182794 , n15441 );
buf ( n182795 , n182794 );
nand ( n15444 , n15434 , n182795 );
buf ( n182797 , n15444 );
buf ( n182798 , n182797 );
xor ( n15447 , n182781 , n182798 );
buf ( n182800 , n182283 );
not ( n15449 , n182800 );
buf ( n182802 , n2566 );
not ( n15451 , n182802 );
or ( n15452 , n15449 , n15451 );
buf ( n182805 , n818 );
buf ( n182806 , n168806 );
nand ( n15455 , n182805 , n182806 );
buf ( n182808 , n15455 );
buf ( n182809 , n182808 );
nand ( n15458 , n15452 , n182809 );
buf ( n182811 , n15458 );
buf ( n182812 , n182811 );
xor ( n15461 , n15447 , n182812 );
buf ( n182814 , n15461 );
xor ( n15463 , n15412 , n182814 );
buf ( n182816 , n15463 );
xor ( n15465 , n15315 , n182816 );
buf ( n182818 , n15465 );
buf ( n182819 , n182818 );
xor ( n15468 , n182513 , n182559 );
and ( n15469 , n15468 , n182576 );
and ( n15470 , n182513 , n182559 );
or ( n15471 , n15469 , n15470 );
buf ( n182824 , n15471 );
buf ( n182825 , n182824 );
xor ( n15474 , n182819 , n182825 );
buf ( n182827 , n182333 );
not ( n15476 , n182827 );
buf ( n182829 , n168713 );
not ( n15478 , n182829 );
or ( n15479 , n15476 , n15478 );
buf ( n182832 , n2823 );
xor ( n15481 , n806 , n779 );
buf ( n182834 , n15481 );
nand ( n15483 , n182832 , n182834 );
buf ( n182836 , n15483 );
buf ( n182837 , n182836 );
nand ( n182838 , n15479 , n182837 );
buf ( n182839 , n182838 );
not ( n15491 , n15081 );
not ( n15492 , n169836 );
or ( n15493 , n15491 , n15492 );
buf ( n182843 , n169320 );
buf ( n182844 , n769 );
buf ( n182845 , n816 );
xor ( n15497 , n182844 , n182845 );
buf ( n182847 , n15497 );
buf ( n182848 , n182847 );
nand ( n15500 , n182843 , n182848 );
buf ( n182850 , n15500 );
nand ( n15502 , n15493 , n182850 );
xor ( n15503 , n182839 , n15502 );
buf ( n182853 , n182458 );
not ( n15505 , n182853 );
buf ( n182855 , n182475 );
not ( n15507 , n182855 );
or ( n15508 , n15505 , n15507 );
buf ( n182858 , n182475 );
buf ( n182859 , n182458 );
or ( n15511 , n182858 , n182859 );
buf ( n182861 , n182442 );
nand ( n15513 , n15511 , n182861 );
buf ( n182863 , n15513 );
buf ( n182864 , n182863 );
nand ( n15516 , n15508 , n182864 );
buf ( n182866 , n15516 );
xnor ( n15518 , n15503 , n182866 );
buf ( n182868 , n15518 );
xor ( n15520 , n182520 , n182526 );
and ( n15521 , n15520 , n182538 );
and ( n15522 , n182520 , n182526 );
or ( n15523 , n15521 , n15522 );
buf ( n182873 , n15523 );
buf ( n182874 , n182873 );
xor ( n15526 , n182868 , n182874 );
or ( n15527 , n14970 , n14982 );
nand ( n15528 , n15527 , n14995 );
buf ( n182878 , n15528 );
buf ( n182879 , n14982 );
buf ( n182880 , n14970 );
nand ( n15532 , n182879 , n182880 );
buf ( n182882 , n15532 );
buf ( n182883 , n182882 );
nand ( n15535 , n182878 , n182883 );
buf ( n182885 , n15535 );
buf ( n182886 , n182885 );
buf ( n182887 , n182403 );
buf ( n182888 , n182375 );
or ( n15540 , n182887 , n182888 );
buf ( n182890 , n182370 );
nand ( n15542 , n15540 , n182890 );
buf ( n182892 , n15542 );
buf ( n182893 , n182892 );
buf ( n182894 , n182403 );
buf ( n182895 , n182375 );
nand ( n15547 , n182894 , n182895 );
buf ( n182897 , n15547 );
buf ( n182898 , n182897 );
nand ( n15550 , n182893 , n182898 );
buf ( n182900 , n15550 );
buf ( n182901 , n182900 );
xor ( n15553 , n182886 , n182901 );
xor ( n15554 , n182273 , n182290 );
and ( n15555 , n15554 , n182303 );
and ( n15556 , n182273 , n182290 );
or ( n15557 , n15555 , n15556 );
buf ( n182907 , n15557 );
buf ( n182908 , n182907 );
xor ( n15560 , n15553 , n182908 );
buf ( n182910 , n15560 );
buf ( n182911 , n182910 );
xor ( n15563 , n15526 , n182911 );
buf ( n182913 , n15563 );
buf ( n182914 , n182913 );
xor ( n15566 , n182519 , n182541 );
and ( n15567 , n15566 , n182556 );
and ( n15568 , n182519 , n182541 );
or ( n15569 , n15567 , n15568 );
buf ( n182919 , n15569 );
buf ( n182920 , n182919 );
xor ( n15572 , n182914 , n182920 );
buf ( n182922 , n182354 );
not ( n15574 , n182922 );
buf ( n182924 , n182492 );
not ( n15576 , n182924 );
or ( n15577 , n15574 , n15576 );
buf ( n182927 , n182492 );
buf ( n182928 , n182354 );
or ( n15580 , n182927 , n182928 );
buf ( n182930 , n182486 );
not ( n15582 , n182930 );
buf ( n182932 , n15582 );
buf ( n182933 , n182932 );
nand ( n15585 , n15580 , n182933 );
buf ( n182935 , n15585 );
buf ( n182936 , n182935 );
nand ( n15588 , n15577 , n182936 );
buf ( n182938 , n15588 );
buf ( n182939 , n182938 );
xor ( n15591 , n15572 , n182939 );
buf ( n182941 , n15591 );
buf ( n182942 , n182941 );
xor ( n15594 , n15474 , n182942 );
buf ( n182944 , n15594 );
xor ( n15596 , n182642 , n182944 );
buf ( n182946 , n15596 );
not ( n15598 , n182946 );
buf ( n182948 , n15598 );
not ( n15600 , n182948 );
buf ( n182950 , n182581 );
buf ( n182951 , n182251 );
nand ( n15603 , n182950 , n182951 );
buf ( n182953 , n15603 );
not ( n15605 , n182953 );
or ( n15606 , n15600 , n15605 );
xor ( n15607 , n182819 , n182825 );
and ( n15608 , n15607 , n182942 );
and ( n15609 , n182819 , n182825 );
or ( n15610 , n15608 , n15609 );
buf ( n182960 , n15610 );
buf ( n182961 , n182960 );
not ( n15613 , n182961 );
xor ( n15614 , n182660 , n182666 );
and ( n15615 , n15614 , n182816 );
and ( n15616 , n182660 , n182666 );
or ( n15617 , n15615 , n15616 );
buf ( n182967 , n15617 );
buf ( n182968 , n182967 );
xor ( n15620 , n182914 , n182920 );
and ( n15621 , n15620 , n182939 );
and ( n15622 , n182914 , n182920 );
or ( n15623 , n15621 , n15622 );
buf ( n182973 , n15623 );
buf ( n182974 , n182973 );
xor ( n15626 , n182968 , n182974 );
xor ( n15627 , n182868 , n182874 );
and ( n15628 , n15627 , n182911 );
and ( n15629 , n182868 , n182874 );
or ( n15630 , n15628 , n15629 );
buf ( n182980 , n15630 );
buf ( n182981 , n182980 );
not ( n15633 , n15481 );
not ( n15634 , n181588 );
or ( n15635 , n15633 , n15634 );
buf ( n182985 , n181594 );
buf ( n182986 , n778 );
buf ( n182987 , n806 );
xor ( n15639 , n182986 , n182987 );
buf ( n182989 , n15639 );
buf ( n182990 , n182989 );
nand ( n15642 , n182985 , n182990 );
buf ( n182992 , n15642 );
nand ( n15644 , n15635 , n182992 );
xor ( n15645 , n15502 , n15644 );
not ( n15646 , n182791 );
not ( n15647 , n170019 );
or ( n15648 , n15646 , n15647 );
buf ( n182998 , n2554 );
buf ( n182999 , n776 );
buf ( n183000 , n808 );
xor ( n15652 , n182999 , n183000 );
buf ( n183002 , n15652 );
buf ( n183003 , n183002 );
nand ( n15655 , n182998 , n183003 );
buf ( n183005 , n15655 );
nand ( n15657 , n15648 , n183005 );
xor ( n15658 , n15645 , n15657 );
buf ( n183008 , n15658 );
buf ( n183009 , n182839 );
not ( n15661 , n183009 );
buf ( n183011 , n15502 );
nand ( n15663 , n15661 , n183011 );
buf ( n183013 , n15663 );
buf ( n183014 , n183013 );
not ( n15666 , n183014 );
buf ( n183016 , n182866 );
not ( n15668 , n183016 );
or ( n15669 , n15666 , n15668 );
buf ( n183019 , n15502 );
not ( n15671 , n183019 );
buf ( n183021 , n182839 );
nand ( n15673 , n15671 , n183021 );
buf ( n183023 , n15673 );
buf ( n183024 , n183023 );
nand ( n15676 , n15669 , n183024 );
buf ( n183026 , n15676 );
buf ( n183027 , n183026 );
xor ( n15679 , n183008 , n183027 );
xor ( n15680 , n182886 , n182901 );
and ( n15681 , n15680 , n182908 );
and ( n15682 , n182886 , n182901 );
or ( n15683 , n15681 , n15682 );
buf ( n183033 , n15683 );
buf ( n183034 , n183033 );
xor ( n15686 , n15679 , n183034 );
buf ( n183036 , n15686 );
buf ( n183037 , n183036 );
xor ( n15689 , n182981 , n183037 );
not ( n15690 , n182814 );
not ( n15691 , n182763 );
or ( n15692 , n15690 , n15691 );
buf ( n183042 , n182814 );
buf ( n183043 , n182763 );
or ( n15695 , n183042 , n183043 );
buf ( n183045 , n182709 );
nand ( n15697 , n15695 , n183045 );
buf ( n183047 , n15697 );
nand ( n15699 , n15692 , n183047 );
buf ( n183049 , n15699 );
xor ( n15701 , n182672 , n182689 );
and ( n15702 , n15701 , n182707 );
and ( n15703 , n182672 , n182689 );
or ( n15704 , n15702 , n15703 );
buf ( n183054 , n15704 );
buf ( n183055 , n183054 );
xor ( n15707 , n182726 , n182743 );
and ( n15708 , n15707 , n182761 );
and ( n15709 , n182726 , n182743 );
or ( n15710 , n15708 , n15709 );
buf ( n183060 , n15710 );
buf ( n183061 , n183060 );
xor ( n15713 , n183055 , n183061 );
xor ( n15714 , n182781 , n182798 );
and ( n15715 , n15714 , n182812 );
and ( n15716 , n182781 , n182798 );
or ( n15717 , n15715 , n15716 );
buf ( n183067 , n15717 );
buf ( n183068 , n183067 );
xor ( n15720 , n15713 , n183068 );
buf ( n183070 , n15720 );
buf ( n183071 , n183070 );
xor ( n15723 , n183049 , n183071 );
buf ( n183073 , n786 );
buf ( n183074 , n800 );
and ( n15726 , n183073 , n183074 );
buf ( n183076 , n15726 );
buf ( n183077 , n183076 );
buf ( n183078 , n182700 );
not ( n15730 , n183078 );
buf ( n183080 , n3497 );
not ( n15732 , n183080 );
or ( n15733 , n15730 , n15732 );
buf ( n183083 , n170972 );
buf ( n183084 , n784 );
buf ( n183085 , n800 );
xor ( n15737 , n183084 , n183085 );
buf ( n183087 , n15737 );
buf ( n183088 , n183087 );
nand ( n15740 , n183083 , n183088 );
buf ( n183090 , n15740 );
buf ( n183091 , n183090 );
nand ( n15743 , n15733 , n183091 );
buf ( n183093 , n15743 );
buf ( n183094 , n183093 );
xor ( n15746 , n183077 , n183094 );
buf ( n183096 , n182774 );
not ( n15748 , n183096 );
buf ( n183098 , n169922 );
buf ( n15750 , n183098 );
buf ( n183100 , n15750 );
buf ( n183101 , n183100 );
not ( n15753 , n183101 );
or ( n15754 , n15748 , n15753 );
buf ( n183104 , n169250 );
buf ( n183105 , n770 );
buf ( n183106 , n814 );
xor ( n15758 , n183105 , n183106 );
buf ( n183108 , n15758 );
buf ( n183109 , n183108 );
nand ( n15764 , n183104 , n183109 );
buf ( n183111 , n15764 );
buf ( n183112 , n183111 );
nand ( n15767 , n15754 , n183112 );
buf ( n183114 , n15767 );
buf ( n183115 , n183114 );
xor ( n15770 , n15746 , n183115 );
buf ( n183117 , n15770 );
buf ( n183118 , n183117 );
not ( n15773 , n182754 );
not ( n15774 , n2757 );
or ( n15775 , n15773 , n15774 );
buf ( n183122 , n3220 );
buf ( n183123 , n772 );
buf ( n183124 , n812 );
xor ( n15779 , n183123 , n183124 );
buf ( n183126 , n15779 );
buf ( n183127 , n183126 );
nand ( n15782 , n183122 , n183127 );
buf ( n183129 , n15782 );
nand ( n15784 , n15775 , n183129 );
buf ( n183131 , n168806 );
not ( n15786 , n183131 );
buf ( n183133 , n15786 );
buf ( n183134 , n183133 );
not ( n15789 , n183134 );
buf ( n183136 , n168793 );
not ( n15791 , n183136 );
or ( n15792 , n15789 , n15791 );
buf ( n183139 , n818 );
nand ( n15794 , n15792 , n183139 );
buf ( n183141 , n15794 );
xor ( n15796 , n15784 , n183141 );
buf ( n183143 , n182847 );
not ( n15798 , n183143 );
buf ( n183145 , n171029 );
not ( n15800 , n183145 );
or ( n15801 , n15798 , n15800 );
buf ( n183148 , n169320 );
buf ( n183149 , n768 );
buf ( n183150 , n816 );
xor ( n15805 , n183149 , n183150 );
buf ( n183152 , n15805 );
buf ( n183153 , n183152 );
nand ( n15808 , n183148 , n183153 );
buf ( n183155 , n15808 );
buf ( n183156 , n183155 );
nand ( n15811 , n15801 , n183156 );
buf ( n183158 , n15811 );
xor ( n15813 , n15796 , n183158 );
buf ( n183160 , n15813 );
xor ( n15815 , n183118 , n183160 );
buf ( n183162 , n182719 );
not ( n15817 , n183162 );
buf ( n183164 , n168861 );
not ( n15819 , n183164 );
or ( n15820 , n15817 , n15819 );
buf ( n183167 , n168870 );
buf ( n183168 , n782 );
buf ( n183169 , n802 );
xor ( n15824 , n183168 , n183169 );
buf ( n183171 , n15824 );
buf ( n183172 , n183171 );
nand ( n15827 , n183167 , n183172 );
buf ( n183174 , n15827 );
buf ( n183175 , n183174 );
nand ( n15830 , n15820 , n183175 );
buf ( n183177 , n15830 );
buf ( n183178 , n183177 );
buf ( n183179 , n182736 );
not ( n15834 , n183179 );
buf ( n183181 , n168750 );
buf ( n15836 , n183181 );
buf ( n183183 , n15836 );
buf ( n183184 , n183183 );
not ( n15839 , n183184 );
or ( n15840 , n15834 , n15839 );
buf ( n183187 , n178447 );
buf ( n183188 , n780 );
buf ( n183189 , n804 );
xor ( n15844 , n183188 , n183189 );
buf ( n183191 , n15844 );
buf ( n183192 , n183191 );
nand ( n15847 , n183187 , n183192 );
buf ( n183194 , n15847 );
buf ( n183195 , n183194 );
nand ( n15850 , n15840 , n183195 );
buf ( n183197 , n15850 );
buf ( n183198 , n183197 );
xor ( n15853 , n183178 , n183198 );
buf ( n183200 , n182682 );
not ( n15855 , n183200 );
buf ( n183202 , n180199 );
not ( n15857 , n183202 );
or ( n15858 , n15855 , n15857 );
buf ( n183205 , n172582 );
buf ( n183206 , n774 );
buf ( n183207 , n810 );
xor ( n15862 , n183206 , n183207 );
buf ( n183209 , n15862 );
buf ( n183210 , n183209 );
nand ( n15865 , n183205 , n183210 );
buf ( n183212 , n15865 );
buf ( n183213 , n183212 );
nand ( n15868 , n15858 , n183213 );
buf ( n183215 , n15868 );
buf ( n183216 , n183215 );
xor ( n15871 , n15853 , n183216 );
buf ( n183218 , n15871 );
buf ( n183219 , n183218 );
xor ( n15874 , n15815 , n183219 );
buf ( n183221 , n15874 );
buf ( n183222 , n183221 );
xor ( n15877 , n15723 , n183222 );
buf ( n183224 , n15877 );
buf ( n183225 , n183224 );
xor ( n15880 , n15689 , n183225 );
buf ( n183227 , n15880 );
buf ( n183228 , n183227 );
xor ( n15883 , n15626 , n183228 );
buf ( n183230 , n15883 );
buf ( n183231 , n183230 );
not ( n15886 , n183231 );
buf ( n183233 , n15886 );
buf ( n183234 , n183233 );
not ( n15889 , n183234 );
or ( n15890 , n15613 , n15889 );
buf ( n183237 , n183230 );
buf ( n183238 , n182960 );
not ( n183239 , n183238 );
buf ( n183240 , n183239 );
buf ( n183241 , n183240 );
nand ( n15896 , n183237 , n183241 );
buf ( n183243 , n15896 );
buf ( n183244 , n183243 );
nand ( n15899 , n15890 , n183244 );
buf ( n183246 , n15899 );
not ( n15901 , n183246 );
buf ( n183248 , n182642 );
buf ( n183249 , n182944 );
and ( n15904 , n183248 , n183249 );
buf ( n183251 , n15904 );
not ( n15906 , n183251 );
nand ( n15907 , n15901 , n15906 );
nand ( n15908 , n15606 , n15907 );
not ( n15909 , n15908 );
buf ( n183256 , n15909 );
buf ( n183257 , n183230 );
buf ( n15912 , n183257 );
buf ( n183259 , n15912 );
and ( n15914 , n183259 , n182960 );
buf ( n183261 , n15914 );
xor ( n15916 , n182968 , n182974 );
and ( n15917 , n15916 , n183228 );
and ( n15918 , n182968 , n182974 );
or ( n15919 , n15917 , n15918 );
buf ( n183266 , n15919 );
xor ( n15921 , n183077 , n183094 );
and ( n15922 , n15921 , n183115 );
and ( n15923 , n183077 , n183094 );
or ( n15924 , n15922 , n15923 );
buf ( n183271 , n15924 );
buf ( n183272 , n183271 );
buf ( n183273 , n183171 );
not ( n15928 , n183273 );
buf ( n183275 , n168861 );
not ( n15930 , n183275 );
or ( n15931 , n15928 , n15930 );
buf ( n183278 , n168870 );
buf ( n183279 , n781 );
buf ( n183280 , n802 );
xor ( n15935 , n183279 , n183280 );
buf ( n183282 , n15935 );
buf ( n183283 , n183282 );
nand ( n15938 , n183278 , n183283 );
buf ( n183285 , n15938 );
buf ( n183286 , n183285 );
nand ( n15941 , n15931 , n183286 );
buf ( n183288 , n15941 );
buf ( n183289 , n183288 );
buf ( n183290 , n183087 );
not ( n15945 , n183290 );
buf ( n183292 , n177819 );
not ( n15947 , n183292 );
or ( n15948 , n15945 , n15947 );
buf ( n183295 , n170972 );
buf ( n183296 , n783 );
buf ( n183297 , n800 );
xor ( n15952 , n183296 , n183297 );
buf ( n183299 , n15952 );
buf ( n183300 , n183299 );
nand ( n15955 , n183295 , n183300 );
buf ( n183302 , n15955 );
buf ( n183303 , n183302 );
nand ( n15958 , n15948 , n183303 );
buf ( n183305 , n15958 );
buf ( n183306 , n183305 );
xor ( n15961 , n183289 , n183306 );
buf ( n183308 , n180199 );
not ( n15963 , n183308 );
buf ( n183310 , n15963 );
buf ( n183311 , n183310 );
buf ( n183312 , n183209 );
not ( n15967 , n183312 );
buf ( n183314 , n15967 );
buf ( n183315 , n183314 );
or ( n15970 , n183311 , n183315 );
buf ( n183317 , n172582 );
not ( n15972 , n183317 );
buf ( n183319 , n15972 );
buf ( n183320 , n183319 );
buf ( n183321 , n773 );
buf ( n183322 , n810 );
xor ( n15977 , n183321 , n183322 );
buf ( n183324 , n15977 );
buf ( n183325 , n183324 );
not ( n15980 , n183325 );
buf ( n183327 , n15980 );
buf ( n183328 , n183327 );
or ( n15983 , n183320 , n183328 );
nand ( n15984 , n15970 , n15983 );
buf ( n183331 , n15984 );
buf ( n183332 , n183331 );
xor ( n15987 , n15961 , n183332 );
buf ( n183334 , n15987 );
buf ( n183335 , n183334 );
xor ( n15990 , n183272 , n183335 );
buf ( n183337 , n785 );
buf ( n183338 , n800 );
and ( n15993 , n183337 , n183338 );
buf ( n183340 , n15993 );
buf ( n183341 , n183340 );
buf ( n183342 , n183002 );
not ( n15997 , n183342 );
buf ( n183344 , n170019 );
not ( n15999 , n183344 );
or ( n16000 , n15997 , n15999 );
buf ( n183347 , n2554 );
buf ( n183348 , n775 );
buf ( n183349 , n808 );
xor ( n16004 , n183348 , n183349 );
buf ( n183351 , n16004 );
buf ( n183352 , n183351 );
nand ( n16007 , n183347 , n183352 );
buf ( n183354 , n16007 );
buf ( n183355 , n183354 );
nand ( n16010 , n16000 , n183355 );
buf ( n183357 , n16010 );
buf ( n183358 , n183357 );
xor ( n16013 , n183341 , n183358 );
buf ( n183360 , n183108 );
not ( n16015 , n183360 );
buf ( n183362 , n183100 );
not ( n16017 , n183362 );
or ( n16018 , n16015 , n16017 );
buf ( n183365 , n169250 );
buf ( n183366 , n769 );
buf ( n183367 , n814 );
xor ( n183368 , n183366 , n183367 );
buf ( n183369 , n183368 );
buf ( n183370 , n183369 );
nand ( n16028 , n183365 , n183370 );
buf ( n183372 , n16028 );
buf ( n183373 , n183372 );
nand ( n16031 , n16018 , n183373 );
buf ( n183375 , n16031 );
buf ( n183376 , n183375 );
xor ( n16034 , n16013 , n183376 );
buf ( n183378 , n16034 );
buf ( n183379 , n183378 );
xor ( n16037 , n15990 , n183379 );
buf ( n183381 , n16037 );
buf ( n183382 , n183152 );
not ( n16040 , n183382 );
buf ( n183384 , n174938 );
not ( n16042 , n183384 );
or ( n16043 , n16040 , n16042 );
buf ( n183387 , n169320 );
buf ( n183388 , n816 );
nand ( n16046 , n183387 , n183388 );
buf ( n183390 , n16046 );
buf ( n183391 , n183390 );
nand ( n16049 , n16043 , n183391 );
buf ( n183393 , n16049 );
buf ( n183394 , n183141 );
not ( n16052 , n183394 );
buf ( n183396 , n183158 );
not ( n16054 , n183396 );
or ( n16055 , n16052 , n16054 );
buf ( n183399 , n183158 );
buf ( n183400 , n183141 );
or ( n16058 , n183399 , n183400 );
buf ( n183402 , n15784 );
nand ( n16060 , n16058 , n183402 );
buf ( n183404 , n16060 );
buf ( n183405 , n183404 );
nand ( n16063 , n16055 , n183405 );
buf ( n183407 , n16063 );
xor ( n16065 , n183393 , n183407 );
xor ( n16066 , n183178 , n183198 );
and ( n16067 , n16066 , n183216 );
and ( n16068 , n183178 , n183198 );
or ( n16069 , n16067 , n16068 );
buf ( n183413 , n16069 );
xor ( n16071 , n16065 , n183413 );
buf ( n183415 , n16071 );
not ( n16073 , n183415 );
xor ( n16074 , n183118 , n183160 );
and ( n16075 , n16074 , n183219 );
and ( n16076 , n183118 , n183160 );
or ( n16077 , n16075 , n16076 );
buf ( n183421 , n16077 );
buf ( n183422 , n183421 );
not ( n16080 , n183422 );
or ( n16081 , n16073 , n16080 );
buf ( n183425 , n183421 );
buf ( n183426 , n16071 );
or ( n16084 , n183425 , n183426 );
nand ( n16085 , n16081 , n16084 );
buf ( n183429 , n16085 );
xor ( n16087 , n183381 , n183429 );
buf ( n183431 , n16087 );
xor ( n16089 , n15502 , n15644 );
and ( n16090 , n16089 , n15657 );
and ( n16091 , n15502 , n15644 );
or ( n16092 , n16090 , n16091 );
buf ( n183436 , n16092 );
buf ( n183437 , n183191 );
not ( n16095 , n183437 );
buf ( n183439 , n183183 );
not ( n16097 , n183439 );
or ( n16098 , n16095 , n16097 );
buf ( n183442 , n178447 );
buf ( n183443 , n779 );
buf ( n183444 , n804 );
xor ( n16102 , n183443 , n183444 );
buf ( n183446 , n16102 );
buf ( n183447 , n183446 );
nand ( n16105 , n183442 , n183447 );
buf ( n183449 , n16105 );
buf ( n183450 , n183449 );
nand ( n16108 , n16098 , n183450 );
buf ( n183452 , n16108 );
buf ( n183453 , n183452 );
buf ( n183454 , n183126 );
not ( n16112 , n183454 );
buf ( n183456 , n1907 );
not ( n16114 , n183456 );
or ( n16115 , n16112 , n16114 );
buf ( n183459 , n14277 );
buf ( n183460 , n771 );
buf ( n183461 , n812 );
xor ( n16119 , n183460 , n183461 );
buf ( n183463 , n16119 );
buf ( n183464 , n183463 );
nand ( n16122 , n183459 , n183464 );
buf ( n183466 , n16122 );
buf ( n183467 , n183466 );
nand ( n16125 , n16115 , n183467 );
buf ( n183469 , n16125 );
buf ( n183470 , n183469 );
xor ( n16128 , n183453 , n183470 );
buf ( n183472 , n182989 );
not ( n16130 , n183472 );
buf ( n183474 , n181588 );
not ( n16132 , n183474 );
or ( n16133 , n16130 , n16132 );
buf ( n183477 , n181594 );
buf ( n183478 , n777 );
buf ( n183479 , n806 );
xor ( n16137 , n183478 , n183479 );
buf ( n183481 , n16137 );
buf ( n183482 , n183481 );
nand ( n16140 , n183477 , n183482 );
buf ( n183484 , n16140 );
buf ( n183485 , n183484 );
nand ( n16143 , n16133 , n183485 );
buf ( n183487 , n16143 );
buf ( n183488 , n183487 );
xor ( n16146 , n16128 , n183488 );
buf ( n183490 , n16146 );
buf ( n183491 , n183490 );
xor ( n16149 , n183436 , n183491 );
xor ( n16150 , n183055 , n183061 );
and ( n183494 , n16150 , n183068 );
and ( n16152 , n183055 , n183061 );
or ( n16153 , n183494 , n16152 );
buf ( n183497 , n16153 );
buf ( n183498 , n183497 );
xor ( n16156 , n16149 , n183498 );
buf ( n183500 , n16156 );
buf ( n183501 , n183500 );
xor ( n16159 , n183008 , n183027 );
and ( n16160 , n16159 , n183034 );
and ( n16161 , n183008 , n183027 );
or ( n16162 , n16160 , n16161 );
buf ( n183506 , n16162 );
buf ( n183507 , n183506 );
xor ( n16165 , n183501 , n183507 );
xor ( n16166 , n183049 , n183071 );
and ( n16167 , n16166 , n183222 );
and ( n16168 , n183049 , n183071 );
or ( n16169 , n16167 , n16168 );
buf ( n183513 , n16169 );
buf ( n183514 , n183513 );
xor ( n16172 , n16165 , n183514 );
buf ( n183516 , n16172 );
buf ( n183517 , n183516 );
xor ( n16175 , n183431 , n183517 );
xor ( n16176 , n182981 , n183037 );
and ( n16177 , n16176 , n183225 );
and ( n16178 , n182981 , n183037 );
or ( n16179 , n16177 , n16178 );
buf ( n183523 , n16179 );
buf ( n183524 , n183523 );
xor ( n16182 , n16175 , n183524 );
buf ( n183526 , n16182 );
xor ( n16184 , n183266 , n183526 );
buf ( n183528 , n16184 );
nor ( n16186 , n183261 , n183528 );
buf ( n183530 , n16186 );
buf ( n183531 , n183530 );
not ( n16189 , n183531 );
buf ( n183533 , n16189 );
buf ( n183534 , n183533 );
and ( n16192 , n183256 , n183534 );
buf ( n183536 , n16192 );
buf ( n183537 , n183536 );
nand ( n16195 , n15285 , n183537 );
buf ( n183539 , n16195 );
buf ( n183540 , n183539 );
nor ( n16198 , n181082 , n183540 );
buf ( n183542 , n16198 );
buf ( n183543 , n183542 );
not ( n16201 , n183543 );
buf ( n183545 , n177727 );
not ( n16203 , n183545 );
or ( n16204 , n16201 , n16203 );
buf ( n183548 , n183539 );
not ( n16206 , n183548 );
buf ( n183550 , n16206 );
buf ( n183551 , n183550 );
not ( n16209 , n183551 );
buf ( n183553 , n180553 );
buf ( n183554 , n180558 );
nand ( n16212 , n183553 , n183554 );
buf ( n183556 , n16212 );
not ( n16214 , n183556 );
not ( n16215 , n180984 );
and ( n16216 , n16214 , n16215 );
buf ( n183560 , n180981 );
buf ( n16218 , n183560 );
buf ( n183562 , n16218 );
and ( n16220 , n183562 , n13190 );
nor ( n16221 , n16216 , n16220 );
buf ( n183565 , n16221 );
buf ( n16223 , n183565 );
buf ( n183567 , n16223 );
nand ( n16225 , n180117 , n180115 );
not ( n16226 , n16225 );
buf ( n183570 , n16226 );
not ( n16228 , n183570 );
buf ( n183572 , n12506 );
not ( n16230 , n183572 );
buf ( n183574 , n16230 );
buf ( n183575 , n183574 );
buf ( n183576 , n180017 );
not ( n16234 , n183576 );
buf ( n183578 , n16234 );
buf ( n183579 , n183578 );
nand ( n16237 , n183575 , n183579 );
buf ( n183581 , n16237 );
buf ( n183582 , n183581 );
not ( n16240 , n183582 );
or ( n16241 , n16228 , n16240 );
buf ( n183585 , n12506 );
buf ( n183586 , n180017 );
nand ( n16244 , n183585 , n183586 );
buf ( n183588 , n16244 );
buf ( n183589 , n183588 );
nand ( n16247 , n16241 , n183589 );
buf ( n183591 , n16247 );
buf ( n183592 , n183591 );
buf ( n183593 , n180987 );
nand ( n16251 , n183592 , n183593 );
buf ( n183595 , n16251 );
nand ( n16253 , n183567 , n183595 );
not ( n16254 , n16253 );
buf ( n183598 , n180990 );
not ( n16256 , n183598 );
buf ( n183600 , n16256 );
nor ( n16258 , n181062 , n13697 );
or ( n16259 , n4190 , n16258 );
nand ( n16260 , n13697 , n181062 );
nand ( n16261 , n16259 , n16260 );
not ( n16262 , n16261 );
nor ( n16263 , n181042 , n13666 );
not ( n16264 , n16263 );
or ( n16265 , n16262 , n16264 );
not ( n16266 , n181042 );
nand ( n16267 , n13654 , n181032 );
not ( n16268 , n16267 );
and ( n16269 , n16266 , n16268 );
buf ( n183613 , n13672 );
buf ( n183614 , n181037 );
nand ( n16272 , n183613 , n183614 );
buf ( n183616 , n16272 );
buf ( n183617 , n183616 );
not ( n16275 , n183617 );
buf ( n183619 , n16275 );
nor ( n16280 , n16269 , n183619 );
nand ( n16281 , n16265 , n16280 );
nand ( n16282 , n183600 , n16281 );
nand ( n16283 , n16254 , n16282 );
buf ( n183624 , n16283 );
not ( n16285 , n183624 );
or ( n16286 , n16209 , n16285 );
buf ( n183627 , n181833 );
not ( n16288 , n183627 );
buf ( n183629 , n16288 );
buf ( n183630 , n183629 );
buf ( n183631 , n14073 );
not ( n16292 , n183631 );
buf ( n183633 , n16292 );
buf ( n183634 , n183633 );
nand ( n16295 , n183630 , n183634 );
buf ( n183636 , n16295 );
not ( n16297 , n183636 );
nand ( n16298 , n181851 , n181856 );
not ( n16299 , n16298 );
not ( n16300 , n16299 );
or ( n16301 , n16297 , n16300 );
nand ( n16302 , n181833 , n14073 );
nand ( n16303 , n16301 , n16302 );
buf ( n183644 , n16303 );
buf ( n183645 , n182609 );
buf ( n183646 , n182629 );
nor ( n16307 , n183645 , n183646 );
buf ( n183648 , n16307 );
buf ( n183649 , n183648 );
nand ( n16310 , n183644 , n183649 );
buf ( n183651 , n16310 );
buf ( n183652 , n183651 );
buf ( n183653 , n182626 );
not ( n16314 , n183653 );
buf ( n183655 , n16314 );
buf ( n183656 , n183655 );
buf ( n183657 , n182614 );
not ( n16318 , n183657 );
buf ( n183659 , n16318 );
buf ( n183660 , n183659 );
nor ( n16321 , n183656 , n183660 );
buf ( n183662 , n16321 );
buf ( n183663 , n183662 );
not ( n16324 , n183663 );
buf ( n183665 , n182606 );
not ( n16326 , n183665 );
or ( n16327 , n16324 , n16326 );
not ( n16328 , n182603 );
nand ( n16329 , n16328 , n182589 );
buf ( n183670 , n16329 );
nand ( n16331 , n16327 , n183670 );
buf ( n183672 , n16331 );
buf ( n183673 , n183672 );
not ( n16334 , n183673 );
buf ( n183675 , n16334 );
buf ( n183676 , n183675 );
nand ( n16337 , n183652 , n183676 );
buf ( n183678 , n16337 );
and ( n16339 , n183536 , n183678 );
buf ( n183680 , n183533 );
not ( n16341 , n183680 );
buf ( n183682 , n182953 );
buf ( n183683 , n182948 );
nor ( n16344 , n183682 , n183683 );
buf ( n183685 , n16344 );
buf ( n183686 , n183685 );
not ( n16347 , n183686 );
buf ( n183688 , n15901 );
buf ( n183689 , n15906 );
nand ( n16350 , n183688 , n183689 );
buf ( n183691 , n16350 );
buf ( n183692 , n183691 );
not ( n16353 , n183692 );
or ( n16354 , n16347 , n16353 );
buf ( n183695 , n183246 );
buf ( n183696 , n183251 );
nand ( n16357 , n183695 , n183696 );
buf ( n183698 , n16357 );
buf ( n183699 , n183698 );
nand ( n16360 , n16354 , n183699 );
buf ( n183701 , n16360 );
buf ( n183702 , n183701 );
buf ( n16363 , n183702 );
buf ( n183704 , n16363 );
buf ( n183705 , n183704 );
not ( n16366 , n183705 );
or ( n16367 , n16341 , n16366 );
buf ( n183708 , n15914 );
buf ( n183709 , n16184 );
nand ( n16370 , n183708 , n183709 );
buf ( n183711 , n16370 );
buf ( n183712 , n183711 );
nand ( n16373 , n16367 , n183712 );
buf ( n183714 , n16373 );
nor ( n16375 , n16339 , n183714 );
buf ( n183716 , n16375 );
nand ( n16377 , n16286 , n183716 );
buf ( n183718 , n16377 );
buf ( n183719 , n183718 );
not ( n16380 , n183719 );
buf ( n183721 , n16380 );
buf ( n183722 , n183721 );
nand ( n16383 , n16204 , n183722 );
buf ( n183724 , n16383 );
buf ( n183725 , n183724 );
buf ( n183726 , n183526 );
buf ( n183727 , n183266 );
and ( n16388 , n183726 , n183727 );
buf ( n183729 , n16388 );
buf ( n183730 , n183729 );
not ( n16391 , n183413 );
buf ( n183732 , n183393 );
not ( n16393 , n183732 );
buf ( n183734 , n16393 );
not ( n16395 , n183734 );
or ( n16396 , n16391 , n16395 );
buf ( n183737 , n183413 );
buf ( n183738 , n183734 );
nor ( n183739 , n183737 , n183738 );
buf ( n183740 , n183739 );
buf ( n183741 , n183407 );
not ( n16402 , n183741 );
buf ( n183743 , n16402 );
or ( n16404 , n183740 , n183743 );
nand ( n16405 , n16396 , n16404 );
buf ( n183746 , n16405 );
xor ( n16407 , n183272 , n183335 );
and ( n16408 , n16407 , n183379 );
and ( n16409 , n183272 , n183335 );
or ( n16410 , n16408 , n16409 );
buf ( n183751 , n16410 );
buf ( n183752 , n183751 );
xor ( n16413 , n183746 , n183752 );
xor ( n16414 , n183341 , n183358 );
and ( n16415 , n16414 , n183376 );
and ( n16416 , n183341 , n183358 );
or ( n16417 , n16415 , n16416 );
buf ( n183758 , n16417 );
buf ( n183759 , n183758 );
xor ( n16420 , n183453 , n183470 );
and ( n16421 , n16420 , n183488 );
and ( n16422 , n183453 , n183470 );
or ( n16423 , n16421 , n16422 );
buf ( n183764 , n16423 );
buf ( n183765 , n183764 );
xor ( n16426 , n183759 , n183765 );
buf ( n183767 , n784 );
buf ( n183768 , n800 );
and ( n16429 , n183767 , n183768 );
buf ( n183770 , n16429 );
buf ( n183771 , n183770 );
buf ( n183772 , n183481 );
not ( n16433 , n183772 );
buf ( n183774 , n181588 );
not ( n16435 , n183774 );
or ( n16436 , n16433 , n16435 );
buf ( n183777 , n181594 );
buf ( n183778 , n776 );
buf ( n183779 , n806 );
xor ( n16440 , n183778 , n183779 );
buf ( n183781 , n16440 );
buf ( n183782 , n183781 );
nand ( n16443 , n183777 , n183782 );
buf ( n183784 , n16443 );
buf ( n183785 , n183784 );
nand ( n16446 , n16436 , n183785 );
buf ( n183787 , n16446 );
buf ( n183788 , n183787 );
xor ( n16449 , n183771 , n183788 );
buf ( n183790 , n183463 );
not ( n16451 , n183790 );
buf ( n183792 , n1907 );
not ( n16453 , n183792 );
or ( n16454 , n16451 , n16453 );
not ( n16455 , n14537 );
buf ( n183796 , n16455 );
buf ( n183797 , n770 );
buf ( n183798 , n812 );
xor ( n16459 , n183797 , n183798 );
buf ( n183800 , n16459 );
buf ( n183801 , n183800 );
nand ( n16462 , n183796 , n183801 );
buf ( n183803 , n16462 );
buf ( n183804 , n183803 );
nand ( n16465 , n16454 , n183804 );
buf ( n183806 , n16465 );
buf ( n183807 , n183806 );
xor ( n16468 , n16449 , n183807 );
buf ( n183809 , n16468 );
buf ( n183810 , n183809 );
xor ( n16471 , n16426 , n183810 );
buf ( n183812 , n16471 );
buf ( n183813 , n183812 );
xor ( n16474 , n16413 , n183813 );
buf ( n183815 , n16474 );
buf ( n183816 , n183815 );
buf ( n183817 , n183351 );
not ( n16478 , n183817 );
buf ( n183819 , n170019 );
not ( n16480 , n183819 );
or ( n16481 , n16478 , n16480 );
buf ( n183822 , n2554 );
buf ( n183823 , n774 );
buf ( n183824 , n808 );
xor ( n16485 , n183823 , n183824 );
buf ( n183826 , n16485 );
buf ( n183827 , n183826 );
nand ( n16488 , n183822 , n183827 );
buf ( n183829 , n16488 );
buf ( n183830 , n183829 );
nand ( n16491 , n16481 , n183830 );
buf ( n183832 , n16491 );
buf ( n183833 , n183832 );
buf ( n183834 , n183282 );
not ( n16495 , n183834 );
buf ( n183836 , n170419 );
not ( n16497 , n183836 );
or ( n16498 , n16495 , n16497 );
buf ( n183839 , n168870 );
buf ( n183840 , n780 );
buf ( n183841 , n802 );
xor ( n16502 , n183840 , n183841 );
buf ( n183843 , n16502 );
buf ( n183844 , n183843 );
nand ( n16505 , n183839 , n183844 );
buf ( n183846 , n16505 );
buf ( n183847 , n183846 );
nand ( n16508 , n16498 , n183847 );
buf ( n183849 , n16508 );
buf ( n183850 , n183849 );
xor ( n16511 , n183833 , n183850 );
buf ( n183852 , n183299 );
not ( n16513 , n183852 );
buf ( n183854 , n177819 );
not ( n16515 , n183854 );
or ( n16516 , n16513 , n16515 );
buf ( n183857 , n170972 );
buf ( n183858 , n782 );
buf ( n183859 , n800 );
xor ( n16523 , n183858 , n183859 );
buf ( n183861 , n16523 );
buf ( n183862 , n183861 );
nand ( n16526 , n183857 , n183862 );
buf ( n183864 , n16526 );
buf ( n183865 , n183864 );
nand ( n16529 , n16516 , n183865 );
buf ( n183867 , n16529 );
buf ( n183868 , n183867 );
xor ( n16532 , n16511 , n183868 );
buf ( n183870 , n16532 );
buf ( n183871 , n183870 );
buf ( n183872 , n183369 );
not ( n16536 , n183872 );
buf ( n183874 , n183100 );
not ( n16538 , n183874 );
or ( n16539 , n16536 , n16538 );
buf ( n183877 , n169250 );
buf ( n183878 , n768 );
buf ( n183879 , n814 );
xor ( n16543 , n183878 , n183879 );
buf ( n183881 , n16543 );
buf ( n183882 , n183881 );
nand ( n16546 , n183877 , n183882 );
buf ( n183884 , n16546 );
buf ( n183885 , n183884 );
nand ( n16549 , n16539 , n183885 );
buf ( n183887 , n16549 );
buf ( n183888 , n183887 );
buf ( n183889 , n169842 );
buf ( n183890 , n174938 );
or ( n16554 , n183889 , n183890 );
buf ( n183892 , n816 );
nand ( n16556 , n16554 , n183892 );
buf ( n183894 , n16556 );
buf ( n183895 , n183894 );
xor ( n16559 , n183888 , n183895 );
buf ( n183897 , n183324 );
not ( n16561 , n183897 );
buf ( n183899 , n180199 );
not ( n16563 , n183899 );
or ( n16564 , n16561 , n16563 );
buf ( n183902 , n183319 );
not ( n16566 , n183902 );
buf ( n183904 , n16566 );
buf ( n183905 , n183904 );
buf ( n183906 , n772 );
buf ( n183907 , n810 );
xor ( n16571 , n183906 , n183907 );
buf ( n183909 , n16571 );
buf ( n183910 , n183909 );
nand ( n16574 , n183905 , n183910 );
buf ( n183912 , n16574 );
buf ( n183913 , n183912 );
nand ( n16577 , n16564 , n183913 );
buf ( n183915 , n16577 );
buf ( n183916 , n183915 );
xor ( n16580 , n16559 , n183916 );
buf ( n183918 , n16580 );
buf ( n183919 , n183918 );
xor ( n16583 , n183871 , n183919 );
buf ( n183921 , n183393 );
buf ( n183922 , n183446 );
not ( n16586 , n183922 );
buf ( n183924 , n183183 );
not ( n16588 , n183924 );
or ( n16589 , n16586 , n16588 );
buf ( n183927 , n178447 );
buf ( n183928 , n778 );
buf ( n183929 , n804 );
xor ( n16593 , n183928 , n183929 );
buf ( n183931 , n16593 );
buf ( n183932 , n183931 );
nand ( n16596 , n183927 , n183932 );
buf ( n183934 , n16596 );
buf ( n183935 , n183934 );
nand ( n16599 , n16589 , n183935 );
buf ( n183937 , n16599 );
buf ( n183938 , n183937 );
xor ( n16602 , n183921 , n183938 );
xor ( n16603 , n183289 , n183306 );
and ( n16604 , n16603 , n183332 );
and ( n16605 , n183289 , n183306 );
or ( n16606 , n16604 , n16605 );
buf ( n183944 , n16606 );
buf ( n183945 , n183944 );
xor ( n16609 , n16602 , n183945 );
buf ( n183947 , n16609 );
buf ( n183948 , n183947 );
xor ( n16612 , n16583 , n183948 );
buf ( n183950 , n16612 );
buf ( n183951 , n183950 );
xor ( n16615 , n183436 , n183491 );
and ( n16616 , n16615 , n183498 );
and ( n16617 , n183436 , n183491 );
or ( n16618 , n16616 , n16617 );
buf ( n183956 , n16618 );
buf ( n183957 , n183956 );
xor ( n16621 , n183951 , n183957 );
buf ( n183959 , n183421 );
buf ( n183960 , n16071 );
not ( n16624 , n183960 );
buf ( n183962 , n16624 );
buf ( n183963 , n183962 );
or ( n16627 , n183959 , n183963 );
buf ( n183965 , n183381 );
nand ( n16629 , n16627 , n183965 );
buf ( n183967 , n16629 );
buf ( n183968 , n183967 );
buf ( n183969 , n183421 );
buf ( n183970 , n183962 );
nand ( n16634 , n183969 , n183970 );
buf ( n183972 , n16634 );
buf ( n183973 , n183972 );
nand ( n183974 , n183968 , n183973 );
buf ( n183975 , n183974 );
buf ( n183976 , n183975 );
xor ( n16640 , n16621 , n183976 );
buf ( n183978 , n16640 );
buf ( n183979 , n183978 );
xor ( n16643 , n183816 , n183979 );
xor ( n16644 , n183501 , n183507 );
and ( n16645 , n16644 , n183514 );
and ( n16646 , n183501 , n183507 );
or ( n16647 , n16645 , n16646 );
buf ( n183985 , n16647 );
buf ( n183986 , n183985 );
xor ( n16650 , n16643 , n183986 );
buf ( n183988 , n16650 );
buf ( n183989 , n183988 );
xor ( n16653 , n183431 , n183517 );
and ( n16654 , n16653 , n183524 );
and ( n16655 , n183431 , n183517 );
or ( n16656 , n16654 , n16655 );
buf ( n183994 , n16656 );
buf ( n183995 , n183994 );
xor ( n16659 , n183989 , n183995 );
buf ( n183997 , n16659 );
buf ( n183998 , n183997 );
nand ( n16662 , n183730 , n183998 );
buf ( n184000 , n16662 );
buf ( n184001 , n184000 );
not ( n16665 , n184001 );
buf ( n184003 , n183729 );
buf ( n184004 , n183997 );
nor ( n16668 , n184003 , n184004 );
buf ( n184006 , n16668 );
buf ( n184007 , n184006 );
nor ( n16671 , n16665 , n184007 );
buf ( n184009 , n16671 );
buf ( n184010 , n184009 );
and ( n16674 , n183725 , n184010 );
not ( n16675 , n183725 );
buf ( n184013 , n184009 );
not ( n16677 , n184013 );
buf ( n184015 , n16677 );
buf ( n184016 , n184015 );
and ( n16680 , n16675 , n184016 );
nor ( n16681 , n16674 , n16680 );
buf ( n184019 , n16681 );
buf ( n16683 , n184019 );
buf ( n184021 , n181078 );
not ( n16685 , n184021 );
buf ( n184023 , n16685 );
buf ( n184024 , n184023 );
buf ( n184025 , n182635 );
not ( n16689 , n184025 );
not ( n16690 , n15596 );
nand ( n16691 , n16690 , n182953 );
buf ( n184029 , n16691 );
nand ( n16693 , n16689 , n184029 );
buf ( n184031 , n16693 );
buf ( n184032 , n184031 );
nor ( n16696 , n184024 , n184032 );
buf ( n184034 , n16696 );
buf ( n184035 , n184034 );
not ( n16699 , n184035 );
buf ( n184037 , n177737 );
not ( n16701 , n184037 );
or ( n16702 , n16699 , n16701 );
buf ( n184040 , n184031 );
not ( n16704 , n184040 );
buf ( n184042 , n16704 );
buf ( n184043 , n184042 );
not ( n16707 , n184043 );
not ( n16708 , n16253 );
nand ( n16709 , n16708 , n16282 );
buf ( n184047 , n16709 );
not ( n16711 , n184047 );
or ( n16712 , n16707 , n16711 );
buf ( n184050 , n16691 );
not ( n16714 , n184050 );
buf ( n184052 , n183678 );
not ( n16716 , n184052 );
or ( n16717 , n16714 , n16716 );
not ( n16718 , n183685 );
buf ( n184056 , n16718 );
nand ( n16720 , n16717 , n184056 );
buf ( n184058 , n16720 );
buf ( n184059 , n184058 );
not ( n16723 , n184059 );
buf ( n184061 , n16723 );
buf ( n184062 , n184061 );
nand ( n16726 , n16712 , n184062 );
buf ( n184064 , n16726 );
buf ( n184065 , n184064 );
not ( n16729 , n184065 );
buf ( n184067 , n16729 );
buf ( n184068 , n184067 );
nand ( n16732 , n16702 , n184068 );
buf ( n184070 , n16732 );
buf ( n184071 , n184070 );
buf ( n16735 , n183691 );
buf ( n184073 , n16735 );
buf ( n184074 , n183698 );
and ( n16738 , n184073 , n184074 );
buf ( n184076 , n16738 );
buf ( n184077 , n184076 );
and ( n16741 , n184071 , n184077 );
not ( n16742 , n184071 );
buf ( n184080 , n184076 );
not ( n16744 , n184080 );
buf ( n184082 , n16744 );
buf ( n184083 , n184082 );
and ( n16747 , n16742 , n184083 );
nor ( n16748 , n16741 , n16747 );
buf ( n184086 , n16748 );
buf ( n16750 , n184086 );
buf ( n184088 , n183530 );
buf ( n184089 , n184006 );
nor ( n16756 , n184088 , n184089 );
buf ( n184091 , n16756 );
nand ( n16758 , n184091 , n15909 );
not ( n16759 , n16758 );
nand ( n16760 , n182632 , n14499 , n16759 );
not ( n16761 , n16760 );
not ( n16762 , n183651 );
not ( n16763 , n16758 );
and ( n16764 , n16762 , n16763 );
buf ( n184099 , n183672 );
not ( n16766 , n184099 );
buf ( n184101 , n16759 );
not ( n16768 , n184101 );
or ( n16769 , n16766 , n16768 );
not ( n16770 , n184091 );
not ( n16771 , n183701 );
or ( n16772 , n16770 , n16771 );
not ( n16773 , n183711 );
not ( n16774 , n184006 );
and ( n16775 , n16773 , n16774 );
buf ( n184110 , n184000 );
not ( n16777 , n184110 );
buf ( n184112 , n16777 );
nor ( n16779 , n16775 , n184112 );
nand ( n16780 , n16772 , n16779 );
buf ( n184115 , n16780 );
not ( n16782 , n184115 );
buf ( n184117 , n16782 );
buf ( n184118 , n184117 );
nand ( n16785 , n16769 , n184118 );
buf ( n184120 , n16785 );
nor ( n16787 , n16764 , n184120 );
not ( n16788 , n16787 );
or ( n16789 , n16761 , n16788 );
buf ( n184124 , n183595 );
buf ( n184125 , n184117 );
nand ( n16792 , n184124 , n184125 );
buf ( n184127 , n16792 );
not ( n16794 , n184127 );
buf ( n184129 , n183651 );
not ( n16796 , n184129 );
buf ( n184131 , n16221 );
buf ( n184132 , n183675 );
nand ( n16799 , n184131 , n184132 );
buf ( n184134 , n16799 );
buf ( n184135 , n184134 );
nor ( n16802 , n16796 , n184135 );
buf ( n184137 , n16802 );
nand ( n16804 , n183600 , n16281 );
nand ( n16805 , n16794 , n184137 , n16804 );
nand ( n16806 , n16789 , n16805 );
buf ( n184141 , n16806 );
not ( n16808 , n184141 );
buf ( n184143 , n16808 );
buf ( n184144 , n184143 );
buf ( n184145 , n775 );
buf ( n184146 , n804 );
xor ( n16813 , n184145 , n184146 );
buf ( n184148 , n16813 );
buf ( n184149 , n184148 );
not ( n16816 , n184149 );
buf ( n184151 , n183183 );
not ( n16818 , n184151 );
or ( n16819 , n16816 , n16818 );
buf ( n184154 , n178447 );
buf ( n184155 , n774 );
buf ( n184156 , n804 );
xor ( n16823 , n184155 , n184156 );
buf ( n184158 , n16823 );
buf ( n184159 , n184158 );
nand ( n16826 , n184154 , n184159 );
buf ( n184161 , n16826 );
buf ( n184162 , n184161 );
nand ( n16829 , n16819 , n184162 );
buf ( n184164 , n16829 );
buf ( n184165 , n184164 );
buf ( n184166 , n800 );
buf ( n184167 , n780 );
and ( n16834 , n184166 , n184167 );
buf ( n184169 , n16834 );
buf ( n184170 , n184169 );
xor ( n16837 , n184165 , n184170 );
buf ( n184172 , n16837 );
buf ( n184173 , n184172 );
buf ( n184174 , n771 );
buf ( n184175 , n808 );
xor ( n16842 , n184174 , n184175 );
buf ( n184177 , n16842 );
buf ( n184178 , n184177 );
not ( n16845 , n184178 );
buf ( n184180 , n170019 );
not ( n16847 , n184180 );
or ( n16848 , n16845 , n16847 );
buf ( n184183 , n2554 );
xor ( n16850 , n808 , n770 );
buf ( n184185 , n16850 );
nand ( n16852 , n184183 , n184185 );
buf ( n184187 , n16852 );
buf ( n184188 , n184187 );
nand ( n16855 , n16848 , n184188 );
buf ( n184190 , n16855 );
buf ( n184191 , n184190 );
xor ( n16858 , n184173 , n184191 );
buf ( n184193 , n16858 );
buf ( n184194 , n184193 );
buf ( n184195 , n768 );
buf ( n184196 , n812 );
xor ( n16863 , n184195 , n184196 );
buf ( n184198 , n16863 );
buf ( n184199 , n184198 );
not ( n16866 , n184199 );
buf ( n184201 , n1907 );
not ( n16868 , n184201 );
or ( n16869 , n16866 , n16868 );
buf ( n184204 , n14277 );
buf ( n184205 , n812 );
nand ( n16872 , n184204 , n184205 );
buf ( n184207 , n16872 );
buf ( n184208 , n184207 );
nand ( n16875 , n16869 , n184208 );
buf ( n184210 , n16875 );
buf ( n184211 , n184210 );
not ( n16878 , n184211 );
buf ( n184213 , n16878 );
buf ( n184214 , n184213 );
xor ( n16881 , n184166 , n184167 );
buf ( n184216 , n16881 );
buf ( n184217 , n184216 );
not ( n16884 , n184217 );
buf ( n184219 , n177819 );
not ( n16886 , n184219 );
or ( n16887 , n16884 , n16886 );
buf ( n184222 , n170972 );
buf ( n184223 , n800 );
buf ( n184224 , n779 );
xor ( n16891 , n184223 , n184224 );
buf ( n184226 , n16891 );
buf ( n184227 , n184226 );
nand ( n16894 , n184222 , n184227 );
buf ( n184229 , n16894 );
buf ( n184230 , n184229 );
nand ( n16897 , n16887 , n184230 );
buf ( n184232 , n16897 );
buf ( n184233 , n184232 );
xor ( n16900 , n184214 , n184233 );
buf ( n184235 , n183100 );
not ( n16902 , n184235 );
buf ( n184237 , n16902 );
buf ( n184238 , n184237 );
buf ( n184239 , n169250 );
not ( n16906 , n184239 );
buf ( n184241 , n16906 );
buf ( n184242 , n184241 );
and ( n16909 , n184238 , n184242 );
buf ( n184244 , n814 );
not ( n16911 , n184244 );
buf ( n184246 , n16911 );
buf ( n184247 , n184246 );
nor ( n16914 , n16909 , n184247 );
buf ( n184249 , n16914 );
buf ( n184250 , n184249 );
not ( n16917 , n184250 );
buf ( n184252 , n170019 );
buf ( n184253 , n773 );
buf ( n184254 , n808 );
xor ( n16921 , n184253 , n184254 );
buf ( n184256 , n16921 );
buf ( n184257 , n184256 );
and ( n16924 , n184252 , n184257 );
buf ( n184259 , n2554 );
xor ( n16926 , n808 , n772 );
buf ( n184261 , n16926 );
and ( n16928 , n184259 , n184261 );
nor ( n16929 , n16924 , n16928 );
buf ( n184264 , n16929 );
buf ( n184265 , n184264 );
not ( n16932 , n184265 );
or ( n16933 , n16917 , n16932 );
buf ( n184268 , n769 );
buf ( n184269 , n812 );
xor ( n16936 , n184268 , n184269 );
buf ( n184271 , n16936 );
buf ( n184272 , n184271 );
not ( n16939 , n184272 );
buf ( n184274 , n1907 );
not ( n16941 , n184274 );
or ( n16942 , n16939 , n16941 );
buf ( n184277 , n16455 );
buf ( n184278 , n184198 );
nand ( n16945 , n184277 , n184278 );
buf ( n184280 , n16945 );
buf ( n184281 , n184280 );
nand ( n16948 , n16942 , n184281 );
buf ( n184283 , n16948 );
buf ( n184284 , n184283 );
nand ( n16951 , n16933 , n184284 );
buf ( n184286 , n16951 );
buf ( n184287 , n184286 );
buf ( n184288 , n184249 );
not ( n16955 , n184288 );
buf ( n184290 , n184264 );
not ( n16957 , n184290 );
buf ( n184292 , n16957 );
buf ( n184293 , n184292 );
nand ( n16960 , n16955 , n184293 );
buf ( n184295 , n16960 );
buf ( n184296 , n184295 );
nand ( n16963 , n184287 , n184296 );
buf ( n184298 , n16963 );
buf ( n184299 , n184298 );
and ( n16966 , n16900 , n184299 );
and ( n16967 , n184214 , n184233 );
or ( n16968 , n16966 , n16967 );
buf ( n184303 , n16968 );
buf ( n184304 , n184303 );
xor ( n16971 , n184194 , n184304 );
buf ( n184306 , n777 );
buf ( n184307 , n802 );
xor ( n184308 , n184306 , n184307 );
buf ( n184309 , n184308 );
buf ( n184310 , n184309 );
not ( n16980 , n184310 );
buf ( n184312 , n170419 );
not ( n16982 , n184312 );
or ( n16983 , n16980 , n16982 );
buf ( n184315 , n168870 );
xor ( n16985 , n802 , n776 );
buf ( n184317 , n16985 );
nand ( n16987 , n184315 , n184317 );
buf ( n184319 , n16987 );
buf ( n184320 , n184319 );
nand ( n16990 , n16983 , n184320 );
buf ( n184322 , n16990 );
buf ( n184323 , n184226 );
not ( n16993 , n184323 );
buf ( n184325 , n177819 );
not ( n16995 , n184325 );
or ( n16996 , n16993 , n16995 );
buf ( n184328 , n170972 );
buf ( n184329 , n800 );
buf ( n184330 , n778 );
xor ( n17000 , n184329 , n184330 );
buf ( n184332 , n17000 );
buf ( n184333 , n184332 );
nand ( n17003 , n184328 , n184333 );
buf ( n184335 , n17003 );
buf ( n184336 , n184335 );
nand ( n17006 , n16996 , n184336 );
buf ( n184338 , n17006 );
xor ( n17008 , n184322 , n184338 );
buf ( n184340 , n17008 );
buf ( n184341 , n184210 );
and ( n17011 , n184340 , n184341 );
not ( n17012 , n184340 );
buf ( n184344 , n184213 );
and ( n17014 , n17012 , n184344 );
nor ( n17015 , n17011 , n17014 );
buf ( n184347 , n17015 );
buf ( n184348 , n184347 );
xor ( n17018 , n16971 , n184348 );
buf ( n184350 , n17018 );
buf ( n184351 , n184350 );
buf ( n184352 , n16926 );
not ( n17022 , n184352 );
buf ( n184354 , n170019 );
not ( n17024 , n184354 );
or ( n17025 , n17022 , n17024 );
buf ( n184357 , n2554 );
buf ( n184358 , n184177 );
nand ( n17028 , n184357 , n184358 );
buf ( n184360 , n17028 );
buf ( n184361 , n184360 );
nand ( n17031 , n17025 , n184361 );
buf ( n184363 , n17031 );
buf ( n184364 , n776 );
buf ( n184365 , n804 );
xor ( n17035 , n184364 , n184365 );
buf ( n184367 , n17035 );
buf ( n184368 , n184367 );
not ( n17038 , n184368 );
buf ( n184370 , n183183 );
not ( n17040 , n184370 );
or ( n17041 , n17038 , n17040 );
buf ( n184373 , n178447 );
buf ( n184374 , n184148 );
nand ( n17044 , n184373 , n184374 );
buf ( n184376 , n17044 );
buf ( n184377 , n184376 );
nand ( n17047 , n17041 , n184377 );
buf ( n184379 , n17047 );
buf ( n17049 , n184379 );
xor ( n17050 , n184363 , n17049 );
buf ( n184382 , n778 );
buf ( n184383 , n802 );
xor ( n17053 , n184382 , n184383 );
buf ( n184385 , n17053 );
buf ( n184386 , n184385 );
not ( n17056 , n184386 );
buf ( n184388 , n170419 );
not ( n17058 , n184388 );
or ( n17059 , n17056 , n17058 );
buf ( n184391 , n168870 );
buf ( n184392 , n184309 );
nand ( n17062 , n184391 , n184392 );
buf ( n184394 , n17062 );
buf ( n184395 , n184394 );
nand ( n17065 , n17059 , n184395 );
buf ( n184397 , n17065 );
not ( n17067 , n184397 );
xor ( n17068 , n17050 , n17067 );
not ( n17069 , n17068 );
not ( n17070 , n17069 );
buf ( n184402 , n777 );
buf ( n184403 , n804 );
xor ( n17073 , n184402 , n184403 );
buf ( n184405 , n17073 );
buf ( n184406 , n184405 );
not ( n17076 , n184406 );
buf ( n184408 , n183183 );
not ( n17078 , n184408 );
or ( n17079 , n17076 , n17078 );
buf ( n184411 , n178447 );
buf ( n184412 , n184367 );
nand ( n17082 , n184411 , n184412 );
buf ( n184414 , n17082 );
buf ( n184415 , n184414 );
nand ( n17085 , n17079 , n184415 );
buf ( n184417 , n17085 );
buf ( n184418 , n184417 );
buf ( n184419 , n779 );
buf ( n184420 , n802 );
xor ( n17090 , n184419 , n184420 );
buf ( n184422 , n17090 );
buf ( n184423 , n184422 );
not ( n17093 , n184423 );
buf ( n184425 , n170419 );
not ( n17095 , n184425 );
or ( n17096 , n17093 , n17095 );
buf ( n184428 , n168870 );
buf ( n184429 , n184385 );
nand ( n17099 , n184428 , n184429 );
buf ( n184431 , n17099 );
buf ( n184432 , n184431 );
nand ( n17102 , n17096 , n184432 );
buf ( n184434 , n17102 );
buf ( n184435 , n184434 );
xor ( n17105 , n184418 , n184435 );
xor ( n17106 , n810 , n771 );
buf ( n184438 , n17106 );
not ( n17108 , n184438 );
buf ( n184440 , n180199 );
not ( n17110 , n184440 );
or ( n17111 , n17108 , n17110 );
buf ( n184443 , n183904 );
buf ( n184444 , n770 );
buf ( n184445 , n810 );
xor ( n17115 , n184444 , n184445 );
buf ( n184447 , n17115 );
buf ( n184448 , n184447 );
nand ( n17118 , n184443 , n184448 );
buf ( n184450 , n17118 );
buf ( n184451 , n184450 );
nand ( n17121 , n17111 , n184451 );
buf ( n184453 , n17121 );
buf ( n184454 , n184453 );
and ( n17124 , n17105 , n184454 );
and ( n17125 , n184418 , n184435 );
or ( n17126 , n17124 , n17125 );
buf ( n184458 , n17126 );
buf ( n17128 , n184458 );
not ( n17129 , n17128 );
buf ( n184461 , n782 );
buf ( n184462 , n800 );
and ( n17132 , n184461 , n184462 );
buf ( n184464 , n17132 );
buf ( n184465 , n184464 );
buf ( n184466 , n781 );
buf ( n184467 , n800 );
xor ( n17137 , n184466 , n184467 );
buf ( n184469 , n17137 );
buf ( n184470 , n184469 );
not ( n17140 , n184470 );
buf ( n184472 , n177819 );
not ( n17142 , n184472 );
or ( n17143 , n17140 , n17142 );
buf ( n184475 , n170972 );
buf ( n184476 , n184216 );
nand ( n17146 , n184475 , n184476 );
buf ( n184478 , n17146 );
buf ( n184479 , n184478 );
nand ( n17149 , n17143 , n184479 );
buf ( n184481 , n17149 );
buf ( n184482 , n184481 );
xor ( n17152 , n184465 , n184482 );
xor ( n17153 , n806 , n775 );
buf ( n184485 , n17153 );
not ( n17155 , n184485 );
buf ( n184487 , n181588 );
not ( n17157 , n184487 );
or ( n17158 , n17155 , n17157 );
buf ( n184490 , n181594 );
buf ( n184491 , n774 );
buf ( n184492 , n806 );
xor ( n17162 , n184491 , n184492 );
buf ( n184494 , n17162 );
buf ( n184495 , n184494 );
nand ( n17165 , n184490 , n184495 );
buf ( n184497 , n17165 );
buf ( n184498 , n184497 );
nand ( n17168 , n17158 , n184498 );
buf ( n184500 , n17168 );
buf ( n184501 , n184500 );
and ( n17171 , n17152 , n184501 );
and ( n17172 , n184465 , n184482 );
or ( n17173 , n17171 , n17172 );
buf ( n184505 , n17173 );
buf ( n17175 , n184505 );
not ( n17176 , n17175 );
nand ( n17177 , n17129 , n17176 );
not ( n17178 , n17177 );
or ( n17179 , n17070 , n17178 );
nand ( n17180 , n17175 , n17128 );
nand ( n17181 , n17179 , n17180 );
buf ( n184513 , n17181 );
not ( n17183 , n184363 );
not ( n17184 , n17183 );
not ( n17185 , n17067 );
or ( n17186 , n17184 , n17185 );
nand ( n17187 , n17186 , n17049 );
or ( n184519 , n17067 , n17183 );
nand ( n17192 , n17187 , n184519 );
buf ( n184521 , n781 );
buf ( n184522 , n800 );
and ( n17195 , n184521 , n184522 );
buf ( n184524 , n17195 );
buf ( n184525 , n184524 );
buf ( n184526 , n184494 );
not ( n17199 , n184526 );
buf ( n184528 , n168713 );
not ( n17201 , n184528 );
or ( n17202 , n17199 , n17201 );
buf ( n184531 , n181594 );
buf ( n184532 , n773 );
buf ( n184533 , n806 );
xor ( n17206 , n184532 , n184533 );
buf ( n184535 , n17206 );
buf ( n184536 , n184535 );
nand ( n17209 , n184531 , n184536 );
buf ( n184538 , n17209 );
buf ( n184539 , n184538 );
nand ( n17212 , n17202 , n184539 );
buf ( n184541 , n17212 );
buf ( n184542 , n184541 );
xor ( n17215 , n184525 , n184542 );
buf ( n184544 , n184447 );
not ( n17217 , n184544 );
buf ( n184546 , n180199 );
not ( n17219 , n184546 );
or ( n17220 , n17217 , n17219 );
buf ( n184549 , n183904 );
buf ( n184550 , n769 );
buf ( n184551 , n810 );
xor ( n17224 , n184550 , n184551 );
buf ( n184553 , n17224 );
buf ( n184554 , n184553 );
nand ( n17227 , n184549 , n184554 );
buf ( n184556 , n17227 );
buf ( n184557 , n184556 );
nand ( n17230 , n17220 , n184557 );
buf ( n184559 , n17230 );
buf ( n184560 , n184559 );
and ( n17233 , n17215 , n184560 );
and ( n17234 , n184525 , n184542 );
or ( n17235 , n17233 , n17234 );
buf ( n184564 , n17235 );
buf ( n17237 , n184564 );
xor ( n17238 , n17192 , n17237 );
not ( n17239 , n1554 );
not ( n17240 , n14537 );
or ( n17241 , n17239 , n17240 );
nand ( n17242 , n17241 , n812 );
buf ( n184571 , n17242 );
buf ( n184572 , n184553 );
not ( n17245 , n184572 );
buf ( n184574 , n180199 );
not ( n17247 , n184574 );
or ( n17248 , n17245 , n17247 );
buf ( n184577 , n183904 );
buf ( n184578 , n768 );
buf ( n184579 , n810 );
xor ( n17252 , n184578 , n184579 );
buf ( n184581 , n17252 );
buf ( n184582 , n184581 );
nand ( n17255 , n184577 , n184582 );
buf ( n184584 , n17255 );
buf ( n184585 , n184584 );
nand ( n17258 , n17248 , n184585 );
buf ( n184587 , n17258 );
buf ( n184588 , n184587 );
xor ( n17261 , n184571 , n184588 );
buf ( n184590 , n184535 );
not ( n17263 , n184590 );
buf ( n184592 , n181588 );
not ( n17265 , n184592 );
or ( n17266 , n17263 , n17265 );
buf ( n184595 , n181594 );
xor ( n17268 , n806 , n772 );
buf ( n184597 , n17268 );
nand ( n17270 , n184595 , n184597 );
buf ( n184599 , n17270 );
buf ( n184600 , n184599 );
nand ( n17273 , n17266 , n184600 );
buf ( n184602 , n17273 );
buf ( n184603 , n184602 );
xor ( n17276 , n17261 , n184603 );
buf ( n184605 , n17276 );
xor ( n17278 , n17238 , n184605 );
buf ( n184607 , n17278 );
xor ( n17280 , n184513 , n184607 );
xor ( n17281 , n184525 , n184542 );
xor ( n17282 , n17281 , n184560 );
buf ( n184611 , n17282 );
buf ( n184612 , n184611 );
xor ( n17285 , n184214 , n184233 );
xor ( n17286 , n17285 , n184299 );
buf ( n184615 , n17286 );
buf ( n184616 , n184615 );
xor ( n17289 , n184612 , n184616 );
buf ( n184618 , n183881 );
not ( n184619 , n184618 );
buf ( n184620 , n183100 );
not ( n17293 , n184620 );
or ( n17294 , n184619 , n17293 );
buf ( n184623 , n184241 );
not ( n17296 , n184623 );
buf ( n184625 , n814 );
nand ( n17298 , n17296 , n184625 );
buf ( n184627 , n17298 );
buf ( n184628 , n184627 );
nand ( n17301 , n17294 , n184628 );
buf ( n184630 , n17301 );
buf ( n184631 , n184630 );
buf ( n184632 , n183781 );
not ( n17305 , n184632 );
buf ( n184634 , n181588 );
not ( n17307 , n184634 );
or ( n17308 , n17305 , n17307 );
buf ( n184637 , n181594 );
buf ( n184638 , n17153 );
nand ( n17311 , n184637 , n184638 );
buf ( n184640 , n17311 );
buf ( n184641 , n184640 );
nand ( n17314 , n17308 , n184641 );
buf ( n184643 , n17314 );
buf ( n184644 , n184643 );
not ( n17317 , n184644 );
not ( n17318 , n183904 );
not ( n17319 , n17106 );
or ( n17320 , n17318 , n17319 );
nand ( n17321 , n183909 , n180199 );
nand ( n17322 , n17320 , n17321 );
buf ( n184651 , n17322 );
not ( n17324 , n184651 );
or ( n17325 , n17317 , n17324 );
buf ( n184654 , n17322 );
buf ( n184655 , n184643 );
or ( n17328 , n184654 , n184655 );
buf ( n184657 , n183800 );
not ( n17330 , n184657 );
buf ( n184659 , n2757 );
not ( n17332 , n184659 );
or ( n17333 , n17330 , n17332 );
buf ( n184662 , n14538 );
buf ( n184663 , n184271 );
nand ( n17336 , n184662 , n184663 );
buf ( n184665 , n17336 );
buf ( n184666 , n184665 );
nand ( n17339 , n17333 , n184666 );
buf ( n184668 , n17339 );
buf ( n184669 , n184668 );
nand ( n17342 , n17328 , n184669 );
buf ( n184671 , n17342 );
buf ( n184672 , n184671 );
nand ( n17345 , n17325 , n184672 );
buf ( n184674 , n17345 );
buf ( n184675 , n184674 );
xor ( n17348 , n184631 , n184675 );
buf ( n184677 , n783 );
buf ( n184678 , n800 );
and ( n17351 , n184677 , n184678 );
buf ( n184680 , n17351 );
buf ( n184681 , n184680 );
buf ( n184682 , n183826 );
not ( n17355 , n184682 );
buf ( n184684 , n170019 );
not ( n17357 , n184684 );
or ( n17358 , n17355 , n17357 );
buf ( n184687 , n2554 );
buf ( n184688 , n184256 );
nand ( n17361 , n184687 , n184688 );
buf ( n184690 , n17361 );
buf ( n184691 , n184690 );
nand ( n17364 , n17358 , n184691 );
buf ( n184693 , n17364 );
buf ( n184694 , n184693 );
xor ( n17367 , n184681 , n184694 );
buf ( n184696 , n183861 );
not ( n17369 , n184696 );
buf ( n184698 , n177819 );
not ( n17371 , n184698 );
or ( n17372 , n17369 , n17371 );
buf ( n184701 , n170972 );
buf ( n184702 , n184469 );
nand ( n17375 , n184701 , n184702 );
buf ( n184704 , n17375 );
buf ( n184705 , n184704 );
nand ( n17378 , n17372 , n184705 );
buf ( n184707 , n17378 );
buf ( n184708 , n184707 );
and ( n17381 , n17367 , n184708 );
and ( n17382 , n184681 , n184694 );
or ( n17383 , n17381 , n17382 );
buf ( n184712 , n17383 );
buf ( n184713 , n184712 );
and ( n17386 , n17348 , n184713 );
and ( n17387 , n184631 , n184675 );
or ( n17388 , n17386 , n17387 );
buf ( n184717 , n17388 );
buf ( n184718 , n184717 );
and ( n17394 , n17289 , n184718 );
and ( n17395 , n184612 , n184616 );
or ( n17396 , n17394 , n17395 );
buf ( n184722 , n17396 );
buf ( n184723 , n184722 );
xor ( n17399 , n17280 , n184723 );
buf ( n184725 , n17399 );
buf ( n184726 , n184725 );
xor ( n17402 , n184351 , n184726 );
xor ( n17403 , n184465 , n184482 );
xor ( n17404 , n17403 , n184501 );
buf ( n184730 , n17404 );
buf ( n184731 , n184730 );
xor ( n17407 , n184418 , n184435 );
xor ( n17408 , n17407 , n184454 );
buf ( n184734 , n17408 );
buf ( n184735 , n184734 );
xor ( n17411 , n184731 , n184735 );
xor ( n17412 , n184249 , n184283 );
buf ( n184738 , n17412 );
buf ( n184739 , n184264 );
and ( n17415 , n184738 , n184739 );
not ( n17416 , n184738 );
buf ( n184742 , n184292 );
and ( n17418 , n17416 , n184742 );
nor ( n17419 , n17415 , n17418 );
buf ( n184745 , n17419 );
buf ( n184746 , n184745 );
and ( n17422 , n17411 , n184746 );
and ( n17423 , n184731 , n184735 );
or ( n17424 , n17422 , n17423 );
buf ( n184750 , n17424 );
buf ( n184751 , n184750 );
and ( n17427 , n17128 , n17176 , n17068 );
not ( n17428 , n17427 );
nand ( n17429 , n17175 , n17128 , n17069 );
nand ( n17430 , n17176 , n17129 , n17069 );
not ( n17431 , n17128 );
nand ( n17432 , n17431 , n17175 , n17068 );
nand ( n17433 , n17428 , n17429 , n17430 , n17432 );
buf ( n184759 , n17433 );
xor ( n17435 , n184751 , n184759 );
xor ( n17436 , n184612 , n184616 );
xor ( n17437 , n17436 , n184718 );
buf ( n184763 , n17437 );
buf ( n184764 , n184763 );
and ( n17440 , n17435 , n184764 );
and ( n17441 , n184751 , n184759 );
or ( n17442 , n17440 , n17441 );
buf ( n184768 , n17442 );
buf ( n184769 , n184768 );
xor ( n17445 , n17402 , n184769 );
buf ( n184771 , n17445 );
buf ( n184772 , n184771 );
buf ( n184773 , n183931 );
not ( n17449 , n184773 );
buf ( n184775 , n183183 );
not ( n17451 , n184775 );
or ( n17452 , n17449 , n17451 );
buf ( n184778 , n178447 );
buf ( n184779 , n184405 );
nand ( n17455 , n184778 , n184779 );
buf ( n184781 , n17455 );
buf ( n184782 , n184781 );
nand ( n17458 , n17452 , n184782 );
buf ( n184784 , n17458 );
buf ( n184785 , n184784 );
buf ( n184786 , n183843 );
not ( n17462 , n184786 );
buf ( n184788 , n170419 );
not ( n17464 , n184788 );
or ( n17465 , n17462 , n17464 );
buf ( n184791 , n168870 );
buf ( n184792 , n184422 );
nand ( n17468 , n184791 , n184792 );
buf ( n184794 , n17468 );
buf ( n184795 , n184794 );
nand ( n17471 , n17465 , n184795 );
buf ( n184797 , n17471 );
buf ( n184798 , n184797 );
xor ( n17474 , n184785 , n184798 );
buf ( n184800 , n184630 );
not ( n17476 , n184800 );
buf ( n184802 , n17476 );
buf ( n184803 , n184802 );
and ( n17479 , n17474 , n184803 );
and ( n17480 , n184785 , n184798 );
or ( n17481 , n17479 , n17480 );
buf ( n184807 , n17481 );
buf ( n184808 , n184807 );
xor ( n17484 , n184631 , n184675 );
xor ( n17485 , n17484 , n184713 );
buf ( n184811 , n17485 );
buf ( n184812 , n184811 );
xor ( n17488 , n184808 , n184812 );
xor ( n184814 , n183771 , n183788 );
and ( n17490 , n184814 , n183807 );
and ( n17491 , n183771 , n183788 );
or ( n17492 , n17490 , n17491 );
buf ( n184818 , n17492 );
buf ( n184819 , n184818 );
xor ( n17495 , n183833 , n183850 );
and ( n17496 , n17495 , n183868 );
and ( n17497 , n183833 , n183850 );
or ( n17498 , n17496 , n17497 );
buf ( n184824 , n17498 );
buf ( n184825 , n184824 );
xor ( n17501 , n184819 , n184825 );
xor ( n17502 , n183888 , n183895 );
and ( n17503 , n17502 , n183916 );
and ( n17504 , n183888 , n183895 );
or ( n17505 , n17503 , n17504 );
buf ( n184831 , n17505 );
buf ( n184832 , n184831 );
and ( n17508 , n17501 , n184832 );
and ( n17509 , n184819 , n184825 );
or ( n17510 , n17508 , n17509 );
buf ( n184836 , n17510 );
buf ( n184837 , n184836 );
and ( n17513 , n17488 , n184837 );
and ( n17514 , n184808 , n184812 );
or ( n17515 , n17513 , n17514 );
buf ( n184841 , n17515 );
buf ( n184842 , n184841 );
xor ( n17518 , n184751 , n184759 );
xor ( n17519 , n17518 , n184764 );
buf ( n184845 , n17519 );
buf ( n184846 , n184845 );
xor ( n17522 , n184842 , n184846 );
xor ( n17523 , n184681 , n184694 );
xor ( n17524 , n17523 , n184708 );
buf ( n184850 , n17524 );
buf ( n184851 , n184850 );
xor ( n17527 , n17322 , n184643 );
xor ( n17528 , n17527 , n184668 );
buf ( n184854 , n17528 );
xor ( n17530 , n184851 , n184854 );
xor ( n17531 , n184785 , n184798 );
xor ( n17532 , n17531 , n184803 );
buf ( n184858 , n17532 );
buf ( n184859 , n184858 );
and ( n17535 , n17530 , n184859 );
and ( n17536 , n184851 , n184854 );
or ( n17537 , n17535 , n17536 );
buf ( n184863 , n17537 );
buf ( n184864 , n184863 );
xor ( n17540 , n184731 , n184735 );
xor ( n17541 , n17540 , n184746 );
buf ( n184867 , n17541 );
buf ( n184868 , n184867 );
xor ( n17544 , n184864 , n184868 );
xor ( n17545 , n183921 , n183938 );
and ( n17546 , n17545 , n183945 );
and ( n17547 , n183921 , n183938 );
or ( n17548 , n17546 , n17547 );
buf ( n184874 , n17548 );
buf ( n184875 , n184874 );
xor ( n17551 , n183759 , n183765 );
and ( n17552 , n17551 , n183810 );
and ( n17553 , n183759 , n183765 );
or ( n17554 , n17552 , n17553 );
buf ( n184880 , n17554 );
buf ( n184881 , n184880 );
xor ( n17557 , n184875 , n184881 );
xor ( n17558 , n184819 , n184825 );
xor ( n17559 , n17558 , n184832 );
buf ( n184885 , n17559 );
buf ( n184886 , n184885 );
and ( n17562 , n17557 , n184886 );
and ( n17563 , n184875 , n184881 );
or ( n17564 , n17562 , n17563 );
buf ( n184890 , n17564 );
buf ( n184891 , n184890 );
and ( n17567 , n17544 , n184891 );
and ( n17568 , n184864 , n184868 );
or ( n17569 , n17567 , n17568 );
buf ( n184895 , n17569 );
buf ( n184896 , n184895 );
and ( n17572 , n17522 , n184896 );
and ( n17573 , n184842 , n184846 );
or ( n17574 , n17572 , n17573 );
buf ( n184900 , n17574 );
buf ( n184901 , n184900 );
xor ( n17577 , n184772 , n184901 );
buf ( n184903 , n17577 );
buf ( n184904 , n184903 );
not ( n17580 , n184904 );
buf ( n184906 , n17580 );
buf ( n184907 , n184906 );
xor ( n17583 , n184842 , n184846 );
xor ( n184909 , n17583 , n184896 );
buf ( n184910 , n184909 );
buf ( n184911 , n184910 );
xor ( n17590 , n184808 , n184812 );
xor ( n17591 , n17590 , n184837 );
buf ( n184914 , n17591 );
buf ( n184915 , n184914 );
xor ( n17594 , n183871 , n183919 );
and ( n17595 , n17594 , n183948 );
and ( n17596 , n183871 , n183919 );
or ( n17597 , n17595 , n17596 );
buf ( n184920 , n17597 );
buf ( n184921 , n184920 );
xor ( n17600 , n184851 , n184854 );
xor ( n17601 , n17600 , n184859 );
buf ( n184924 , n17601 );
buf ( n184925 , n184924 );
xor ( n17604 , n184921 , n184925 );
xor ( n17605 , n183746 , n183752 );
and ( n17606 , n17605 , n183813 );
and ( n17607 , n183746 , n183752 );
or ( n17608 , n17606 , n17607 );
buf ( n184931 , n17608 );
buf ( n184932 , n184931 );
and ( n17611 , n17604 , n184932 );
and ( n17612 , n184921 , n184925 );
or ( n17613 , n17611 , n17612 );
buf ( n184936 , n17613 );
buf ( n184937 , n184936 );
xor ( n17616 , n184915 , n184937 );
xor ( n17617 , n184864 , n184868 );
xor ( n17618 , n17617 , n184891 );
buf ( n184941 , n17618 );
buf ( n184942 , n184941 );
and ( n17621 , n17616 , n184942 );
and ( n17622 , n184915 , n184937 );
or ( n17623 , n17621 , n17622 );
buf ( n184946 , n17623 );
buf ( n184947 , n184946 );
and ( n17626 , n184911 , n184947 );
buf ( n184949 , n17626 );
buf ( n184950 , n184949 );
not ( n17629 , n184950 );
buf ( n184952 , n17629 );
buf ( n184953 , n184952 );
nand ( n17632 , n184907 , n184953 );
buf ( n184955 , n17632 );
buf ( n184956 , n184955 );
xor ( n17635 , n184915 , n184937 );
xor ( n17636 , n17635 , n184942 );
buf ( n184959 , n17636 );
buf ( n184960 , n184959 );
xor ( n17639 , n184875 , n184881 );
xor ( n17640 , n17639 , n184886 );
buf ( n184963 , n17640 );
buf ( n184964 , n184963 );
xor ( n17643 , n184921 , n184925 );
xor ( n17644 , n17643 , n184932 );
buf ( n184967 , n17644 );
buf ( n184968 , n184967 );
xor ( n17647 , n184964 , n184968 );
xor ( n17648 , n183951 , n183957 );
and ( n17649 , n17648 , n183976 );
and ( n17650 , n183951 , n183957 );
or ( n17651 , n17649 , n17650 );
buf ( n184974 , n17651 );
buf ( n184975 , n184974 );
and ( n17654 , n17647 , n184975 );
and ( n17655 , n184964 , n184968 );
or ( n17656 , n17654 , n17655 );
buf ( n184979 , n17656 );
buf ( n184980 , n184979 );
and ( n17659 , n184960 , n184980 );
buf ( n184982 , n17659 );
buf ( n184983 , n184982 );
not ( n17662 , n184983 );
xor ( n17663 , n184911 , n184947 );
buf ( n184986 , n17663 );
buf ( n184987 , n184986 );
not ( n17666 , n184987 );
buf ( n184989 , n17666 );
buf ( n184990 , n184989 );
nand ( n17669 , n17662 , n184990 );
buf ( n184992 , n17669 );
buf ( n184993 , n184992 );
and ( n17672 , n184956 , n184993 );
buf ( n184995 , n17672 );
buf ( n184996 , n184995 );
xor ( n17675 , n183816 , n183979 );
and ( n17676 , n17675 , n183986 );
and ( n184999 , n183816 , n183979 );
or ( n17678 , n17676 , n184999 );
buf ( n185001 , n17678 );
xor ( n17680 , n184964 , n184968 );
xor ( n17681 , n17680 , n184975 );
buf ( n185004 , n17681 );
xor ( n17683 , n185001 , n185004 );
buf ( n185006 , n17683 );
and ( n17685 , n183989 , n183995 );
buf ( n185008 , n17685 );
buf ( n185009 , n185008 );
nor ( n17688 , n185006 , n185009 );
buf ( n185011 , n17688 );
buf ( n185012 , n185011 );
buf ( n185013 , n185004 );
buf ( n185014 , n185001 );
and ( n17693 , n185013 , n185014 );
buf ( n185016 , n17693 );
buf ( n185017 , n185016 );
buf ( n185018 , n184979 );
not ( n17697 , n185018 );
buf ( n185020 , n184959 );
not ( n17699 , n185020 );
buf ( n185022 , n17699 );
buf ( n185023 , n185022 );
not ( n17702 , n185023 );
or ( n17703 , n17697 , n17702 );
buf ( n185026 , n184979 );
not ( n17705 , n185026 );
buf ( n185028 , n184959 );
nand ( n17707 , n17705 , n185028 );
buf ( n185030 , n17707 );
buf ( n185031 , n185030 );
nand ( n17710 , n17703 , n185031 );
buf ( n185033 , n17710 );
buf ( n185034 , n185033 );
nor ( n17713 , n185017 , n185034 );
buf ( n185036 , n17713 );
buf ( n185037 , n185036 );
nor ( n17716 , n185012 , n185037 );
buf ( n185039 , n17716 );
buf ( n185040 , n185039 );
nand ( n17719 , n184996 , n185040 );
buf ( n185042 , n17719 );
buf ( n185043 , n185042 );
buf ( n17722 , n185043 );
buf ( n185045 , n17722 );
buf ( n185046 , n185045 );
not ( n17725 , n185046 );
buf ( n185048 , n17725 );
buf ( n185049 , n185048 );
and ( n17728 , n184772 , n184901 );
buf ( n185051 , n17728 );
buf ( n185052 , n185051 );
not ( n17731 , n185052 );
xor ( n17732 , n184351 , n184726 );
and ( n17733 , n17732 , n184769 );
and ( n17734 , n184351 , n184726 );
or ( n17735 , n17733 , n17734 );
buf ( n185058 , n17735 );
buf ( n185059 , n185058 );
xor ( n17738 , n184194 , n184304 );
and ( n17739 , n17738 , n184348 );
and ( n17740 , n184194 , n184304 );
or ( n17741 , n17739 , n17740 );
buf ( n185064 , n17741 );
buf ( n185065 , n185064 );
xor ( n17744 , n184513 , n184607 );
and ( n17745 , n17744 , n184723 );
and ( n17746 , n184513 , n184607 );
or ( n17747 , n17745 , n17746 );
buf ( n185070 , n17747 );
buf ( n185071 , n185070 );
xor ( n17750 , n185065 , n185071 );
buf ( n185073 , n184581 );
not ( n17752 , n185073 );
buf ( n185075 , n178360 );
not ( n17754 , n185075 );
or ( n17755 , n17752 , n17754 );
buf ( n185078 , n183904 );
buf ( n185079 , n810 );
nand ( n17758 , n185078 , n185079 );
buf ( n185081 , n17758 );
buf ( n185082 , n185081 );
nand ( n17761 , n17755 , n185082 );
buf ( n185084 , n17761 );
buf ( n185085 , n185084 );
not ( n17764 , n185085 );
buf ( n185087 , n17764 );
buf ( n185088 , n185087 );
buf ( n185089 , n184190 );
buf ( n185090 , n184169 );
or ( n17772 , n185089 , n185090 );
buf ( n185092 , n184164 );
nand ( n17774 , n17772 , n185092 );
buf ( n185094 , n17774 );
buf ( n185095 , n185094 );
buf ( n185096 , n184169 );
buf ( n185097 , n184190 );
nand ( n17779 , n185096 , n185097 );
buf ( n185099 , n17779 );
buf ( n185100 , n185099 );
nand ( n17782 , n185095 , n185100 );
buf ( n185102 , n17782 );
buf ( n185103 , n185102 );
xor ( n17785 , n185088 , n185103 );
xor ( n17786 , n184571 , n184588 );
and ( n17787 , n17786 , n184603 );
and ( n17788 , n184571 , n184588 );
or ( n17789 , n17787 , n17788 );
buf ( n185109 , n17789 );
buf ( n185110 , n185109 );
xor ( n17792 , n17785 , n185110 );
buf ( n185112 , n17792 );
buf ( n185113 , n185112 );
not ( n17795 , n184605 );
or ( n17796 , n17192 , n17237 );
not ( n17797 , n17796 );
or ( n17798 , n17795 , n17797 );
nand ( n17799 , n17237 , n17192 );
nand ( n17800 , n17798 , n17799 );
buf ( n185120 , n17800 );
xor ( n17802 , n185113 , n185120 );
buf ( n185122 , n184322 );
buf ( n185123 , n184338 );
or ( n17805 , n185122 , n185123 );
buf ( n185125 , n184210 );
nand ( n17807 , n17805 , n185125 );
buf ( n185127 , n17807 );
buf ( n185128 , n185127 );
buf ( n185129 , n184338 );
buf ( n185130 , n184322 );
nand ( n17812 , n185129 , n185130 );
buf ( n185132 , n17812 );
buf ( n185133 , n185132 );
nand ( n17815 , n185128 , n185133 );
buf ( n185135 , n17815 );
buf ( n185136 , n185135 );
buf ( n185137 , n184158 );
not ( n17819 , n185137 );
buf ( n185139 , n183183 );
not ( n17821 , n185139 );
or ( n17822 , n17819 , n17821 );
buf ( n185142 , n178447 );
buf ( n185143 , n773 );
buf ( n185144 , n804 );
xor ( n17826 , n185143 , n185144 );
buf ( n185146 , n17826 );
buf ( n185147 , n185146 );
nand ( n17829 , n185142 , n185147 );
buf ( n185149 , n17829 );
buf ( n185150 , n185149 );
nand ( n17832 , n17822 , n185150 );
buf ( n185152 , n17832 );
buf ( n185153 , n185152 );
buf ( n185154 , n16985 );
not ( n17836 , n185154 );
buf ( n185156 , n170419 );
not ( n17838 , n185156 );
or ( n17839 , n17836 , n17838 );
buf ( n185159 , n168870 );
xor ( n17841 , n802 , n775 );
buf ( n185161 , n17841 );
nand ( n17843 , n185159 , n185161 );
buf ( n185163 , n17843 );
buf ( n185164 , n185163 );
nand ( n17846 , n17839 , n185164 );
buf ( n185166 , n17846 );
buf ( n185167 , n185166 );
xor ( n17849 , n185153 , n185167 );
buf ( n185169 , n16850 );
not ( n17851 , n185169 );
buf ( n185171 , n170019 );
not ( n17853 , n185171 );
or ( n17854 , n17851 , n17853 );
buf ( n185174 , n2554 );
buf ( n185175 , n769 );
buf ( n185176 , n808 );
xor ( n17858 , n185175 , n185176 );
buf ( n185178 , n17858 );
buf ( n185179 , n185178 );
nand ( n17861 , n185174 , n185179 );
buf ( n185181 , n17861 );
buf ( n185182 , n185181 );
nand ( n17864 , n17854 , n185182 );
buf ( n185184 , n17864 );
buf ( n185185 , n185184 );
xor ( n17867 , n17849 , n185185 );
buf ( n185187 , n17867 );
buf ( n185188 , n185187 );
xor ( n17870 , n185136 , n185188 );
and ( n17871 , n184223 , n184224 );
buf ( n185191 , n17871 );
buf ( n185192 , n17268 );
not ( n17874 , n185192 );
buf ( n185194 , n181588 );
not ( n17876 , n185194 );
or ( n17877 , n17874 , n17876 );
buf ( n185197 , n181594 );
xor ( n17879 , n806 , n771 );
buf ( n185199 , n17879 );
nand ( n17881 , n185197 , n185199 );
buf ( n185201 , n17881 );
buf ( n185202 , n185201 );
nand ( n17884 , n17877 , n185202 );
buf ( n185204 , n17884 );
xor ( n17886 , n185191 , n185204 );
buf ( n185206 , n184332 );
not ( n17888 , n185206 );
buf ( n185208 , n177819 );
not ( n17890 , n185208 );
or ( n17891 , n17888 , n17890 );
buf ( n185211 , n170972 );
buf ( n185212 , n800 );
buf ( n185213 , n777 );
xor ( n17895 , n185212 , n185213 );
buf ( n185215 , n17895 );
buf ( n185216 , n185215 );
nand ( n17898 , n185211 , n185216 );
buf ( n185218 , n17898 );
buf ( n185219 , n185218 );
nand ( n17901 , n17891 , n185219 );
buf ( n185221 , n17901 );
xor ( n17903 , n17886 , n185221 );
buf ( n185223 , n17903 );
xor ( n17905 , n17870 , n185223 );
buf ( n185225 , n17905 );
buf ( n185226 , n185225 );
xor ( n17908 , n17802 , n185226 );
buf ( n185228 , n17908 );
buf ( n185229 , n185228 );
xor ( n17911 , n17750 , n185229 );
buf ( n185231 , n17911 );
buf ( n185232 , n185231 );
xor ( n17914 , n185059 , n185232 );
buf ( n185234 , n17914 );
buf ( n185235 , n185234 );
not ( n17917 , n185235 );
buf ( n185237 , n17917 );
buf ( n185238 , n185237 );
nand ( n17920 , n17731 , n185238 );
buf ( n185240 , n17920 );
buf ( n185241 , n185240 );
and ( n17923 , n185059 , n185232 );
buf ( n185243 , n17923 );
nand ( n17925 , n185191 , n185204 );
nand ( n17926 , n185191 , n185221 );
nand ( n17927 , n185204 , n185221 );
nand ( n17928 , n17925 , n17926 , n17927 );
buf ( n185248 , n17928 );
buf ( n185249 , n185178 );
not ( n17931 , n185249 );
buf ( n185251 , n170019 );
not ( n17933 , n185251 );
or ( n17934 , n17931 , n17933 );
buf ( n185254 , n2554 );
buf ( n185255 , n768 );
buf ( n185256 , n808 );
xor ( n17938 , n185255 , n185256 );
buf ( n185258 , n17938 );
buf ( n185259 , n185258 );
nand ( n17944 , n185254 , n185259 );
buf ( n185261 , n17944 );
buf ( n185262 , n185261 );
nand ( n17947 , n17934 , n185262 );
buf ( n185264 , n17947 );
buf ( n185265 , n185264 );
buf ( n185266 , n183319 );
not ( n17951 , n185266 );
buf ( n185268 , n183310 );
not ( n17953 , n185268 );
or ( n17954 , n17951 , n17953 );
buf ( n185271 , n810 );
nand ( n17956 , n17954 , n185271 );
buf ( n185273 , n17956 );
buf ( n185274 , n185273 );
xor ( n17959 , n185265 , n185274 );
buf ( n185276 , n185146 );
not ( n17961 , n185276 );
buf ( n185278 , n183183 );
not ( n17963 , n185278 );
or ( n17964 , n17961 , n17963 );
buf ( n185281 , n178447 );
buf ( n185282 , n772 );
buf ( n185283 , n804 );
xor ( n17968 , n185282 , n185283 );
buf ( n185285 , n17968 );
buf ( n185286 , n185285 );
nand ( n17971 , n185281 , n185286 );
buf ( n185288 , n17971 );
buf ( n185289 , n185288 );
nand ( n17974 , n17964 , n185289 );
buf ( n185291 , n17974 );
buf ( n185292 , n185291 );
xor ( n17977 , n17959 , n185292 );
buf ( n185294 , n17977 );
buf ( n185295 , n185294 );
xor ( n17980 , n185248 , n185295 );
buf ( n185297 , n185215 );
not ( n17982 , n185297 );
buf ( n185299 , n177819 );
not ( n17984 , n185299 );
or ( n17985 , n17982 , n17984 );
buf ( n185302 , n170972 );
buf ( n185303 , n800 );
buf ( n185304 , n776 );
xor ( n17989 , n185303 , n185304 );
buf ( n185306 , n17989 );
buf ( n185307 , n185306 );
nand ( n17992 , n185302 , n185307 );
buf ( n185309 , n17992 );
buf ( n185310 , n185309 );
nand ( n17995 , n17985 , n185310 );
buf ( n185312 , n17995 );
buf ( n185313 , n185312 );
buf ( n185314 , n17841 );
not ( n17999 , n185314 );
buf ( n185316 , n170419 );
not ( n18001 , n185316 );
or ( n18002 , n17999 , n18001 );
buf ( n185319 , n168870 );
buf ( n185320 , n802 );
buf ( n185321 , n774 );
xor ( n18006 , n185320 , n185321 );
buf ( n185323 , n18006 );
buf ( n185324 , n185323 );
nand ( n18009 , n185319 , n185324 );
buf ( n185326 , n18009 );
buf ( n185327 , n185326 );
nand ( n18012 , n18002 , n185327 );
buf ( n185329 , n18012 );
buf ( n185330 , n185329 );
xor ( n18015 , n185313 , n185330 );
buf ( n185332 , n17879 );
not ( n18017 , n185332 );
buf ( n185334 , n181588 );
not ( n18019 , n185334 );
or ( n18020 , n18017 , n18019 );
buf ( n185337 , n181594 );
buf ( n185338 , n770 );
buf ( n185339 , n806 );
xor ( n18024 , n185338 , n185339 );
buf ( n185341 , n18024 );
buf ( n185342 , n185341 );
nand ( n18027 , n185337 , n185342 );
buf ( n185344 , n18027 );
buf ( n185345 , n185344 );
nand ( n18030 , n18020 , n185345 );
buf ( n185347 , n18030 );
buf ( n185348 , n185347 );
xor ( n18033 , n18015 , n185348 );
buf ( n185350 , n18033 );
buf ( n185351 , n185350 );
xor ( n18036 , n17980 , n185351 );
buf ( n185353 , n18036 );
buf ( n185354 , n185353 );
and ( n18039 , n184329 , n184330 );
buf ( n185356 , n18039 );
buf ( n185357 , n185356 );
buf ( n185358 , n185084 );
xor ( n18043 , n185357 , n185358 );
xor ( n18044 , n185153 , n185167 );
and ( n18045 , n18044 , n185185 );
and ( n18046 , n185153 , n185167 );
or ( n18047 , n18045 , n18046 );
buf ( n185364 , n18047 );
buf ( n185365 , n185364 );
xor ( n18050 , n18043 , n185365 );
buf ( n185367 , n18050 );
buf ( n185368 , n185367 );
xor ( n18053 , n185088 , n185103 );
and ( n18054 , n18053 , n185110 );
and ( n18055 , n185088 , n185103 );
or ( n18056 , n18054 , n18055 );
buf ( n185373 , n18056 );
buf ( n185374 , n185373 );
xor ( n18059 , n185368 , n185374 );
xor ( n18060 , n185136 , n185188 );
and ( n18061 , n18060 , n185223 );
and ( n18062 , n185136 , n185188 );
or ( n18063 , n18061 , n18062 );
buf ( n185380 , n18063 );
buf ( n185381 , n185380 );
xor ( n18066 , n18059 , n185381 );
buf ( n185383 , n18066 );
buf ( n185384 , n185383 );
xor ( n18069 , n185354 , n185384 );
xor ( n18070 , n185113 , n185120 );
and ( n18071 , n18070 , n185226 );
and ( n18072 , n185113 , n185120 );
or ( n18073 , n18071 , n18072 );
buf ( n185390 , n18073 );
buf ( n185391 , n185390 );
xor ( n18076 , n18069 , n185391 );
buf ( n185393 , n18076 );
buf ( n185394 , n185393 );
xor ( n18079 , n185065 , n185071 );
and ( n18080 , n18079 , n185229 );
and ( n18081 , n185065 , n185071 );
or ( n18082 , n18080 , n18081 );
buf ( n185399 , n18082 );
buf ( n185400 , n185399 );
xor ( n18085 , n185394 , n185400 );
buf ( n185402 , n18085 );
or ( n18087 , n185243 , n185402 );
buf ( n185404 , n18087 );
and ( n18089 , n185241 , n185404 );
buf ( n185406 , n18089 );
buf ( n185407 , n185406 );
nand ( n18092 , n185049 , n185407 );
buf ( n185409 , n18092 );
buf ( n185410 , n185409 );
not ( n18095 , n185410 );
buf ( n185412 , n18095 );
buf ( n185413 , n185412 );
nand ( n18098 , n184144 , n185413 );
buf ( n185415 , n18098 );
buf ( n185416 , n177727 );
nand ( n18101 , n14499 , n182632 );
buf ( n185418 , n18101 );
not ( n18106 , n185418 );
buf ( n185420 , n13676 );
buf ( n185421 , n180987 );
and ( n18109 , n185420 , n185421 );
buf ( n185423 , n18109 );
buf ( n185424 , n185423 );
buf ( n185425 , n184091 );
buf ( n185426 , n15909 );
buf ( n185427 , n183581 );
buf ( n18115 , n185427 );
buf ( n185429 , n18115 );
buf ( n185430 , n185429 );
and ( n18118 , n185425 , n185426 , n185430 );
buf ( n185432 , n18118 );
buf ( n185433 , n185432 );
buf ( n185434 , n181069 );
buf ( n185435 , n12742 );
nor ( n18123 , n185434 , n185435 );
buf ( n185437 , n18123 );
buf ( n185438 , n185437 );
nand ( n18126 , n18106 , n185424 , n185433 , n185438 );
buf ( n185440 , n18126 );
buf ( n185441 , n185440 );
not ( n18129 , n185441 );
buf ( n185443 , n18129 );
buf ( n185444 , n185443 );
not ( n18132 , n185444 );
buf ( n185446 , n18132 );
buf ( n185447 , n185446 );
buf ( n185448 , n185409 );
nor ( n18136 , n185447 , n185448 );
buf ( n185450 , n18136 );
buf ( n185451 , n185450 );
nand ( n18139 , n185416 , n185451 );
buf ( n185453 , n18139 );
buf ( n185454 , n185406 );
not ( n18142 , n185454 );
buf ( n185456 , n184995 );
not ( n18144 , n185456 );
buf ( n185458 , n17683 );
buf ( n185459 , n185008 );
nand ( n18147 , n185458 , n185459 );
buf ( n185461 , n18147 );
not ( n18149 , n185461 );
not ( n18150 , n18149 );
not ( n18151 , n185036 );
not ( n18152 , n18151 );
or ( n18153 , n18150 , n18152 );
nand ( n18154 , n185016 , n185033 );
nand ( n18155 , n18153 , n18154 );
buf ( n185469 , n18155 );
not ( n18157 , n185469 );
or ( n18158 , n18144 , n18157 );
buf ( n185472 , n184955 );
buf ( n185473 , n184982 );
buf ( n185474 , n184986 );
nand ( n18162 , n185473 , n185474 );
buf ( n185476 , n18162 );
buf ( n185477 , n185476 );
not ( n18165 , n185477 );
buf ( n185479 , n18165 );
buf ( n185480 , n185479 );
and ( n18168 , n185472 , n185480 );
buf ( n185482 , n184906 );
buf ( n185483 , n184952 );
nor ( n18171 , n185482 , n185483 );
buf ( n185485 , n18171 );
buf ( n185486 , n185485 );
nor ( n18174 , n18168 , n185486 );
buf ( n185488 , n18174 );
buf ( n185489 , n185488 );
nand ( n18177 , n18158 , n185489 );
buf ( n185491 , n18177 );
buf ( n185492 , n185491 );
buf ( n18180 , n185492 );
buf ( n185494 , n18180 );
buf ( n185495 , n185494 );
not ( n18183 , n185495 );
or ( n18184 , n18142 , n18183 );
buf ( n185498 , n18087 );
not ( n18186 , n185498 );
buf ( n185500 , n185051 );
buf ( n18188 , n185500 );
buf ( n185502 , n18188 );
buf ( n185503 , n185502 );
buf ( n185504 , n185234 );
nand ( n18192 , n185503 , n185504 );
buf ( n185506 , n18192 );
buf ( n185507 , n185506 );
not ( n18195 , n185507 );
buf ( n185509 , n18195 );
buf ( n185510 , n185509 );
not ( n18198 , n185510 );
or ( n18199 , n18186 , n18198 );
buf ( n185513 , n185243 );
buf ( n185514 , n185402 );
nand ( n18202 , n185513 , n185514 );
buf ( n185516 , n18202 );
buf ( n185517 , n185516 );
nand ( n18205 , n18199 , n185517 );
buf ( n185519 , n18205 );
buf ( n185520 , n185519 );
not ( n18208 , n185520 );
buf ( n185522 , n18208 );
buf ( n185523 , n185522 );
nand ( n18211 , n18184 , n185523 );
buf ( n185525 , n18211 );
buf ( n185526 , n185525 );
not ( n18214 , n185526 );
buf ( n185528 , n18214 );
nand ( n18216 , n185415 , n185453 , n185528 );
and ( n18217 , n185394 , n185400 );
buf ( n185531 , n18217 );
buf ( n185532 , n185531 );
xor ( n18220 , n185265 , n185274 );
and ( n18221 , n18220 , n185292 );
and ( n18222 , n185265 , n185274 );
or ( n18223 , n18221 , n18222 );
buf ( n185537 , n18223 );
buf ( n185538 , n185537 );
xor ( n18226 , n185313 , n185330 );
and ( n18227 , n18226 , n185348 );
and ( n18228 , n185313 , n185330 );
or ( n18229 , n18227 , n18228 );
buf ( n185543 , n18229 );
buf ( n185544 , n185543 );
xor ( n18232 , n185538 , n185544 );
buf ( n185546 , n185306 );
not ( n18234 , n185546 );
buf ( n185548 , n177819 );
not ( n18236 , n185548 );
or ( n18237 , n18234 , n18236 );
buf ( n185551 , n170972 );
buf ( n185552 , n775 );
buf ( n185553 , n800 );
xor ( n18241 , n185552 , n185553 );
buf ( n185555 , n18241 );
buf ( n185556 , n185555 );
nand ( n18244 , n185551 , n185556 );
buf ( n185558 , n18244 );
buf ( n185559 , n185558 );
nand ( n18247 , n18237 , n185559 );
buf ( n185561 , n18247 );
buf ( n185562 , n185258 );
not ( n18250 , n185562 );
buf ( n185564 , n170019 );
not ( n18252 , n185564 );
or ( n18253 , n18250 , n18252 );
buf ( n185567 , n2554 );
buf ( n185568 , n808 );
nand ( n185569 , n185567 , n185568 );
buf ( n185570 , n185569 );
buf ( n185571 , n185570 );
nand ( n18262 , n18253 , n185571 );
buf ( n185573 , n18262 );
xor ( n18264 , n185561 , n185573 );
buf ( n185575 , n185323 );
not ( n18266 , n185575 );
buf ( n185577 , n170419 );
not ( n18268 , n185577 );
or ( n18269 , n18266 , n18268 );
buf ( n185580 , n168870 );
buf ( n185581 , n802 );
buf ( n185582 , n773 );
xor ( n18273 , n185581 , n185582 );
buf ( n185584 , n18273 );
buf ( n185585 , n185584 );
nand ( n18276 , n185580 , n185585 );
buf ( n185587 , n18276 );
buf ( n185588 , n185587 );
nand ( n18279 , n18269 , n185588 );
buf ( n185590 , n18279 );
xor ( n18281 , n18264 , n185590 );
buf ( n185592 , n18281 );
xor ( n18283 , n18232 , n185592 );
buf ( n185594 , n18283 );
buf ( n185595 , n185594 );
and ( n18286 , n185212 , n185213 );
buf ( n185597 , n18286 );
buf ( n185598 , n185597 );
buf ( n185599 , n185285 );
not ( n18290 , n185599 );
buf ( n185601 , n183183 );
not ( n18292 , n185601 );
or ( n18293 , n18290 , n18292 );
buf ( n185604 , n178447 );
buf ( n185605 , n771 );
buf ( n185606 , n804 );
xor ( n18297 , n185605 , n185606 );
buf ( n185608 , n18297 );
buf ( n185609 , n185608 );
nand ( n18300 , n185604 , n185609 );
buf ( n185611 , n18300 );
buf ( n185612 , n185611 );
nand ( n18303 , n18293 , n185612 );
buf ( n185614 , n18303 );
buf ( n185615 , n185614 );
xor ( n18306 , n185598 , n185615 );
buf ( n185617 , n185341 );
not ( n18308 , n185617 );
buf ( n185619 , n181588 );
not ( n18310 , n185619 );
or ( n18311 , n18308 , n18310 );
buf ( n185622 , n181594 );
xor ( n18313 , n806 , n769 );
buf ( n185624 , n18313 );
nand ( n18315 , n185622 , n185624 );
buf ( n185626 , n18315 );
buf ( n185627 , n185626 );
nand ( n18318 , n18311 , n185627 );
buf ( n185629 , n18318 );
buf ( n185630 , n185629 );
not ( n18321 , n185630 );
buf ( n185632 , n18321 );
buf ( n185633 , n185632 );
xor ( n18324 , n18306 , n185633 );
buf ( n185635 , n18324 );
buf ( n185636 , n185635 );
xor ( n18327 , n185357 , n185358 );
and ( n18328 , n18327 , n185365 );
and ( n185639 , n185357 , n185358 );
or ( n18330 , n18328 , n185639 );
buf ( n185641 , n18330 );
buf ( n185642 , n185641 );
xor ( n18333 , n185636 , n185642 );
xor ( n18334 , n185248 , n185295 );
and ( n18335 , n18334 , n185351 );
and ( n18336 , n185248 , n185295 );
or ( n18337 , n18335 , n18336 );
buf ( n185648 , n18337 );
buf ( n185649 , n185648 );
xor ( n18340 , n18333 , n185649 );
buf ( n185651 , n18340 );
buf ( n185652 , n185651 );
xor ( n18343 , n185595 , n185652 );
xor ( n18344 , n185368 , n185374 );
and ( n18345 , n18344 , n185381 );
and ( n18346 , n185368 , n185374 );
or ( n18347 , n18345 , n18346 );
buf ( n185658 , n18347 );
buf ( n185659 , n185658 );
xor ( n18350 , n18343 , n185659 );
buf ( n185661 , n18350 );
buf ( n185662 , n185661 );
xor ( n18353 , n185354 , n185384 );
and ( n18354 , n18353 , n185391 );
and ( n18355 , n185354 , n185384 );
or ( n18356 , n18354 , n18355 );
buf ( n185667 , n18356 );
buf ( n185668 , n185667 );
xor ( n18359 , n185662 , n185668 );
buf ( n185670 , n18359 );
buf ( n185671 , n185670 );
nor ( n18362 , n185532 , n185671 );
buf ( n185673 , n18362 );
buf ( n185674 , n185673 );
not ( n18365 , n185674 );
buf ( n185676 , n18365 );
buf ( n185677 , n185531 );
buf ( n185678 , n185670 );
nand ( n18369 , n185677 , n185678 );
buf ( n185680 , n18369 );
nand ( n18371 , n185676 , n185680 );
not ( n18372 , n18371 );
and ( n18373 , n18216 , n18372 );
not ( n18374 , n18216 );
and ( n18375 , n18374 , n18371 );
nor ( n18376 , n18373 , n18375 );
buf ( n18377 , n18376 );
buf ( n185688 , n181081 );
buf ( n185689 , n182635 );
nor ( n18380 , n185688 , n185689 );
buf ( n185691 , n18380 );
buf ( n185692 , n185691 );
not ( n18383 , n185692 );
buf ( n185694 , n177727 );
not ( n18385 , n185694 );
or ( n18386 , n18383 , n18385 );
buf ( n185697 , n182635 );
not ( n18388 , n185697 );
buf ( n185699 , n18388 );
buf ( n185700 , n185699 );
not ( n18391 , n185700 );
buf ( n185702 , n16283 );
not ( n18393 , n185702 );
or ( n18394 , n18391 , n18393 );
buf ( n185705 , n183678 );
not ( n18396 , n185705 );
buf ( n185707 , n18396 );
buf ( n185708 , n185707 );
nand ( n18402 , n18394 , n185708 );
buf ( n185710 , n18402 );
buf ( n185711 , n185710 );
not ( n18405 , n185711 );
buf ( n185713 , n18405 );
buf ( n185714 , n185713 );
nand ( n18408 , n18386 , n185714 );
buf ( n185716 , n18408 );
buf ( n185717 , n185716 );
buf ( n185718 , n16691 );
buf ( n185719 , n16718 );
nand ( n18413 , n185718 , n185719 );
buf ( n185721 , n18413 );
buf ( n185722 , n185721 );
not ( n18416 , n185722 );
buf ( n185724 , n18416 );
buf ( n185725 , n185724 );
and ( n18419 , n185717 , n185725 );
not ( n18420 , n185717 );
buf ( n185728 , n185721 );
and ( n18422 , n18420 , n185728 );
nor ( n18423 , n18419 , n18422 );
buf ( n185731 , n18423 );
buf ( n18425 , n185731 );
buf ( n185733 , n177669 );
not ( n18427 , n185733 );
nor ( n18428 , n175266 , n175037 );
nor ( n18429 , n176201 , n18428 );
buf ( n185737 , n18429 );
not ( n18431 , n185737 );
or ( n18432 , n18427 , n18431 );
not ( n18433 , n18428 );
not ( n18434 , n18433 );
not ( n18435 , n8687 );
or ( n18436 , n18434 , n18435 );
nand ( n18437 , n175266 , n175037 );
nand ( n18438 , n18436 , n18437 );
buf ( n185746 , n18438 );
not ( n18440 , n185746 );
buf ( n185748 , n18440 );
buf ( n185749 , n185748 );
nand ( n18443 , n18432 , n185749 );
buf ( n185751 , n18443 );
buf ( n185752 , n185751 );
buf ( n185753 , n8709 );
buf ( n185754 , n8714 );
and ( n18448 , n185753 , n185754 );
buf ( n185756 , n18448 );
buf ( n185757 , n185756 );
and ( n18451 , n185752 , n185757 );
not ( n18452 , n185752 );
buf ( n185760 , n185756 );
not ( n18454 , n185760 );
buf ( n185762 , n18454 );
buf ( n185763 , n185762 );
and ( n18457 , n18452 , n185763 );
nor ( n18458 , n18451 , n18457 );
buf ( n185766 , n18458 );
buf ( n18460 , n185766 );
buf ( n185768 , n171657 );
not ( n18462 , n185768 );
buf ( n185770 , n177727 );
not ( n18464 , n185770 );
or ( n18465 , n18462 , n18464 );
buf ( n185773 , n171662 );
nand ( n185774 , n18465 , n185773 );
buf ( n185775 , n185774 );
buf ( n185776 , n185775 );
nand ( n18470 , n13699 , n16260 );
buf ( n185778 , n18470 );
not ( n18472 , n185778 );
buf ( n185780 , n18472 );
buf ( n185781 , n185780 );
and ( n18475 , n185776 , n185781 );
not ( n18476 , n185776 );
buf ( n185784 , n18470 );
and ( n18478 , n18476 , n185784 );
nor ( n18479 , n18475 , n18478 );
buf ( n185787 , n18479 );
buf ( n18481 , n185787 );
buf ( n185789 , n181072 );
buf ( n18483 , n185789 );
buf ( n185791 , n18483 );
buf ( n185792 , n185791 );
not ( n18486 , n185792 );
buf ( n185794 , n18486 );
buf ( n185795 , n185794 );
buf ( n185796 , n12743 );
buf ( n18490 , n185796 );
buf ( n185798 , n18490 );
buf ( n185799 , n185798 );
buf ( n185800 , n180561 );
not ( n18494 , n185800 );
buf ( n185802 , n18494 );
buf ( n185803 , n185802 );
nand ( n18497 , n185799 , n185803 );
buf ( n185805 , n18497 );
buf ( n185806 , n185805 );
nor ( n18500 , n185795 , n185806 );
buf ( n185808 , n18500 );
buf ( n185809 , n185808 );
not ( n18503 , n185809 );
buf ( n185811 , n177737 );
not ( n18505 , n185811 );
or ( n18506 , n18503 , n18505 );
buf ( n18507 , n16281 );
buf ( n185815 , n18507 );
not ( n18509 , n185815 );
buf ( n185817 , n185805 );
not ( n18511 , n185817 );
buf ( n185819 , n18511 );
buf ( n185820 , n185819 );
not ( n18514 , n185820 );
or ( n18515 , n18509 , n18514 );
buf ( n185823 , n185802 );
not ( n18517 , n185823 );
buf ( n185825 , n183591 );
buf ( n18519 , n185825 );
buf ( n185827 , n18519 );
buf ( n185828 , n185827 );
not ( n18522 , n185828 );
or ( n18523 , n18517 , n18522 );
buf ( n185831 , n183556 );
nand ( n18525 , n18523 , n185831 );
buf ( n185833 , n18525 );
buf ( n185834 , n185833 );
not ( n18528 , n185834 );
buf ( n185836 , n18528 );
buf ( n185837 , n185836 );
nand ( n18531 , n18515 , n185837 );
buf ( n185839 , n18531 );
not ( n18536 , n185839 );
buf ( n185841 , n18536 );
nand ( n18538 , n18506 , n185841 );
buf ( n185843 , n18538 );
buf ( n185844 , n180984 );
and ( n18541 , n183562 , n13190 );
buf ( n185846 , n18541 );
or ( n18543 , n185844 , n185846 );
buf ( n185848 , n18543 );
xnor ( n18545 , n185843 , n185848 );
buf ( n18546 , n18545 );
not ( n18547 , n10214 );
buf ( n185852 , n176677 );
not ( n18549 , n185852 );
buf ( n185854 , n18549 );
buf ( n185855 , n185854 );
buf ( n185856 , n177629 );
nand ( n18553 , n185855 , n185856 );
buf ( n185858 , n18553 );
not ( n18555 , n185858 );
or ( n18556 , n18547 , n18555 );
not ( n18557 , n185858 );
nand ( n18558 , n18557 , n10163 , n177616 );
nand ( n18559 , n18556 , n18558 );
buf ( n18560 , n18559 );
buf ( n18561 , n184992 );
buf ( n185866 , n18561 );
buf ( n18563 , n185866 );
buf ( n185868 , n18563 );
buf ( n185869 , n185868 );
not ( n18566 , n185869 );
buf ( n185871 , n18155 );
not ( n18568 , n185871 );
or ( n18569 , n18566 , n18568 );
buf ( n185874 , n185476 );
nand ( n18571 , n18569 , n185874 );
buf ( n185876 , n18571 );
not ( n18573 , n185876 );
buf ( n185878 , n177740 );
buf ( n185879 , n185440 );
not ( n18576 , n185879 );
buf ( n185881 , n18576 );
buf ( n185882 , n185881 );
buf ( n185883 , n185039 );
buf ( n185884 , n185868 );
and ( n18581 , n185883 , n185884 );
buf ( n185886 , n18581 );
buf ( n185887 , n185886 );
and ( n18584 , n185882 , n185887 );
buf ( n185889 , n18584 );
buf ( n185890 , n185889 );
nand ( n18587 , n185878 , n185890 );
buf ( n185892 , n18587 );
buf ( n185893 , n16806 );
not ( n18590 , n185893 );
buf ( n185895 , n18590 );
buf ( n185896 , n185895 );
buf ( n185897 , n185886 );
nand ( n18594 , n185896 , n185897 );
buf ( n185899 , n18594 );
nand ( n18596 , n18573 , n185892 , n185899 );
buf ( n185901 , n18596 );
buf ( n185902 , n184955 );
not ( n18599 , n185902 );
buf ( n185904 , n185485 );
nor ( n18601 , n18599 , n185904 );
buf ( n185906 , n18601 );
buf ( n185907 , n185906 );
and ( n18604 , n185901 , n185907 );
not ( n18605 , n185901 );
buf ( n185910 , n185906 );
not ( n18607 , n185910 );
buf ( n185912 , n18607 );
buf ( n185913 , n185912 );
and ( n18610 , n18605 , n185913 );
nor ( n18611 , n18604 , n18610 );
buf ( n185916 , n18611 );
buf ( n18613 , n185916 );
buf ( n185918 , n185798 );
not ( n18615 , n185918 );
buf ( n185920 , n185794 );
nor ( n18617 , n18615 , n185920 );
buf ( n185922 , n18617 );
buf ( n185923 , n185922 );
not ( n18620 , n185923 );
buf ( n185925 , n177737 );
not ( n18622 , n185925 );
or ( n18623 , n18620 , n18622 );
buf ( n185928 , n185798 );
buf ( n185929 , n18507 );
and ( n18626 , n185928 , n185929 );
buf ( n185931 , n185827 );
nor ( n18628 , n18626 , n185931 );
buf ( n185933 , n18628 );
buf ( n185934 , n185933 );
nand ( n18631 , n18623 , n185934 );
buf ( n185936 , n18631 );
buf ( n185937 , n185936 );
buf ( n185938 , n185802 );
buf ( n185939 , n183556 );
nand ( n18636 , n185938 , n185939 );
buf ( n185941 , n18636 );
buf ( n185942 , n185941 );
not ( n18639 , n185942 );
buf ( n185944 , n18639 );
buf ( n185945 , n185944 );
and ( n18642 , n185937 , n185945 );
not ( n18643 , n185937 );
buf ( n185948 , n185941 );
and ( n18645 , n18643 , n185948 );
nor ( n18646 , n18642 , n18645 );
buf ( n185951 , n18646 );
buf ( n18648 , n185951 );
buf ( n185953 , n185791 );
not ( n18650 , n185953 );
buf ( n185955 , n177727 );
not ( n18652 , n185955 );
or ( n18653 , n18650 , n18652 );
buf ( n185958 , n18507 );
not ( n18658 , n185958 );
buf ( n185960 , n18658 );
buf ( n185961 , n185960 );
nand ( n18661 , n18653 , n185961 );
buf ( n185963 , n18661 );
buf ( n185964 , n185963 );
or ( n18664 , n180117 , n180115 );
buf ( n185966 , n18664 );
buf ( n185967 , n16225 );
nand ( n18667 , n185966 , n185967 );
buf ( n185969 , n18667 );
buf ( n185970 , n185969 );
not ( n18670 , n185970 );
buf ( n185972 , n18670 );
buf ( n185973 , n185972 );
and ( n18673 , n185964 , n185973 );
not ( n18674 , n185964 );
buf ( n185976 , n185969 );
and ( n18676 , n18674 , n185976 );
nor ( n18677 , n18673 , n18676 );
buf ( n185979 , n18677 );
buf ( n18679 , n185979 );
buf ( n185981 , n181069 );
buf ( n18681 , n185981 );
buf ( n185983 , n18681 );
buf ( n185984 , n185983 );
buf ( n185985 , n13666 );
buf ( n18685 , n185985 );
buf ( n185987 , n18685 );
buf ( n185988 , n185987 );
nor ( n18688 , n185984 , n185988 );
buf ( n185990 , n18688 );
nand ( n18690 , n185990 , n177727 );
not ( n18691 , n18690 );
buf ( n18692 , n16261 );
not ( n18693 , n18692 );
nor ( n18694 , n18693 , n185987 );
nand ( n18695 , n16266 , n183616 );
buf ( n185997 , n16267 );
buf ( n18697 , n185997 );
buf ( n185999 , n18697 );
buf ( n186000 , n185999 );
not ( n18700 , n186000 );
buf ( n186002 , n18700 );
nor ( n18702 , n18694 , n18695 , n186002 );
not ( n18703 , n18702 );
or ( n18704 , n18691 , n18703 );
nor ( n18705 , n18694 , n186002 );
not ( n18706 , n18705 );
not ( n18707 , n18690 );
or ( n18708 , n18706 , n18707 );
nand ( n18709 , n18708 , n18695 );
nand ( n18710 , n18704 , n18709 );
buf ( n18711 , n18710 );
buf ( n186013 , n185011 );
buf ( n186014 , n16760 );
nor ( n18714 , n186013 , n186014 );
buf ( n186016 , n18714 );
not ( n18716 , n186016 );
not ( n18717 , n16283 );
buf ( n186019 , n8751 );
buf ( n186020 , n174167 );
and ( n18720 , n186019 , n186020 );
buf ( n186022 , n18720 );
buf ( n186023 , n186022 );
buf ( n18723 , n186023 );
buf ( n186025 , n18723 );
buf ( n186026 , n186025 );
not ( n18726 , n186026 );
buf ( n186028 , n8688 );
buf ( n186029 , n176164 );
not ( n18729 , n186029 );
buf ( n186031 , n18729 );
buf ( n186032 , n186031 );
nand ( n18732 , n186028 , n186032 );
buf ( n186034 , n18732 );
buf ( n186035 , n186034 );
not ( n18735 , n186035 );
buf ( n186037 , n177669 );
not ( n18737 , n186037 );
nand ( n18738 , n8784 , n176198 );
buf ( n186040 , n18738 );
nor ( n18740 , n18737 , n186040 );
buf ( n186042 , n18740 );
buf ( n186043 , n186042 );
not ( n18743 , n186043 );
buf ( n186045 , n18743 );
buf ( n186046 , n186045 );
nand ( n18746 , n18735 , n186046 );
buf ( n186048 , n18746 );
buf ( n186049 , n186048 );
not ( n18749 , n186049 );
or ( n18750 , n18726 , n18749 );
buf ( n186052 , n177718 );
buf ( n18752 , n186052 );
buf ( n186054 , n18752 );
buf ( n186055 , n186054 );
not ( n18755 , n6725 );
not ( n18756 , n8751 );
or ( n18757 , n18755 , n18756 );
not ( n18758 , n6194 );
nand ( n18759 , n18757 , n18758 );
buf ( n186061 , n18759 );
buf ( n18761 , n186061 );
buf ( n186063 , n18761 );
buf ( n186064 , n186063 );
nor ( n18764 , n186055 , n186064 );
buf ( n186066 , n18764 );
buf ( n186067 , n186066 );
nand ( n18767 , n18750 , n186067 );
buf ( n186069 , n18767 );
buf ( n186070 , n186069 );
buf ( n186071 , n173197 );
not ( n18774 , n186071 );
buf ( n186073 , n186054 );
nor ( n18776 , n18774 , n186073 );
buf ( n186075 , n18776 );
buf ( n186076 , n186075 );
buf ( n186077 , n181075 );
nor ( n18780 , n186076 , n186077 );
buf ( n186079 , n18780 );
buf ( n186080 , n186079 );
nand ( n18783 , n186070 , n186080 );
buf ( n186082 , n18783 );
nand ( n18785 , n18717 , n186082 );
not ( n18786 , n18785 );
or ( n18787 , n18716 , n18786 );
buf ( n186086 , n16759 );
not ( n18789 , n186086 );
buf ( n186088 , n183678 );
not ( n18791 , n186088 );
or ( n18792 , n18789 , n18791 );
buf ( n186091 , n184117 );
nand ( n18794 , n18792 , n186091 );
buf ( n186093 , n18794 );
buf ( n186094 , n186093 );
buf ( n186095 , n185011 );
not ( n18798 , n186095 );
buf ( n186097 , n18798 );
buf ( n186098 , n186097 );
nand ( n18801 , n186094 , n186098 );
buf ( n186100 , n18801 );
buf ( n186101 , n186100 );
buf ( n186102 , n185461 );
and ( n18805 , n186101 , n186102 );
buf ( n186104 , n18805 );
nand ( n18807 , n18787 , n186104 );
and ( n18808 , n18154 , n18151 );
and ( n18809 , n18807 , n18808 );
not ( n18810 , n18807 );
not ( n18811 , n18808 );
and ( n18812 , n18810 , n18811 );
nor ( n18813 , n18809 , n18812 );
buf ( n18814 , n18813 );
not ( n18815 , n8773 );
not ( n18816 , n10214 );
not ( n18817 , n176681 );
or ( n18818 , n18816 , n18817 );
nand ( n18819 , n18818 , n10266 );
not ( n18820 , n18819 );
or ( n186119 , n18815 , n18820 );
buf ( n186120 , n176082 );
buf ( n18823 , n186120 );
buf ( n186122 , n18823 );
not ( n18825 , n186122 );
nand ( n18826 , n186119 , n18825 );
buf ( n186125 , n18826 );
buf ( n186126 , n176098 );
not ( n18829 , n186126 );
buf ( n186128 , n176185 );
buf ( n18831 , n186128 );
buf ( n186130 , n18831 );
buf ( n186131 , n186130 );
nand ( n18834 , n18829 , n186131 );
buf ( n186133 , n18834 );
buf ( n186134 , n186133 );
not ( n18837 , n186134 );
buf ( n186136 , n18837 );
buf ( n186137 , n186136 );
and ( n18840 , n186125 , n186137 );
not ( n18841 , n186125 );
buf ( n186140 , n186133 );
and ( n18843 , n18841 , n186140 );
nor ( n18844 , n18840 , n18843 );
buf ( n186143 , n18844 );
buf ( n18846 , n186143 );
buf ( n186145 , n832 );
buf ( n186146 , n880 );
xor ( n18849 , n186145 , n186146 );
buf ( n186148 , n18849 );
buf ( n186149 , n186148 );
not ( n18852 , n186149 );
not ( n18853 , n880 );
not ( n18854 , n881 );
or ( n18855 , n18853 , n18854 );
not ( n18856 , n880 );
not ( n18857 , n881 );
nand ( n18858 , n18856 , n18857 );
nand ( n18859 , n18855 , n18858 );
xor ( n18860 , n881 , n882 );
nor ( n18861 , n18859 , n18860 );
buf ( n18862 , n18861 );
buf ( n186161 , n18862 );
not ( n18864 , n186161 );
or ( n18865 , n18852 , n18864 );
not ( n18866 , n882 );
not ( n18867 , n881 );
not ( n18868 , n18867 );
or ( n18869 , n18866 , n18868 );
not ( n186168 , n882 );
nand ( n18874 , n186168 , n881 );
nand ( n18875 , n18869 , n18874 );
buf ( n186171 , n18875 );
buf ( n186172 , n880 );
nand ( n18878 , n186171 , n186172 );
buf ( n186174 , n18878 );
buf ( n186175 , n186174 );
nand ( n18881 , n18865 , n186175 );
buf ( n186177 , n18881 );
buf ( n186178 , n186177 );
buf ( n186179 , n843 );
buf ( n186180 , n868 );
xor ( n18886 , n186179 , n186180 );
buf ( n186182 , n18886 );
buf ( n186183 , n186182 );
not ( n18889 , n186183 );
xor ( n18890 , n869 , n870 );
not ( n18891 , n18890 );
buf ( n186187 , n18891 );
buf ( n186188 , n868 );
buf ( n186189 , n869 );
xor ( n18895 , n186188 , n186189 );
buf ( n186191 , n18895 );
buf ( n186192 , n186191 );
and ( n18898 , n186187 , n186192 );
buf ( n186194 , n18898 );
buf ( n186195 , n186194 );
buf ( n18901 , n186195 );
buf ( n186197 , n18901 );
buf ( n186198 , n186197 );
not ( n18904 , n186198 );
or ( n18905 , n18889 , n18904 );
not ( n18906 , n18890 );
not ( n18907 , n18906 );
buf ( n186203 , n18907 );
not ( n18909 , n186203 );
buf ( n186205 , n18909 );
buf ( n186206 , n186205 );
not ( n18912 , n186206 );
buf ( n186208 , n18912 );
buf ( n186209 , n186208 );
buf ( n186210 , n842 );
buf ( n186211 , n868 );
xor ( n18917 , n186210 , n186211 );
buf ( n186213 , n18917 );
buf ( n186214 , n186213 );
nand ( n18920 , n186209 , n186214 );
buf ( n186216 , n18920 );
buf ( n186217 , n186216 );
nand ( n18923 , n18905 , n186217 );
buf ( n186219 , n18923 );
buf ( n186220 , n186219 );
xor ( n18926 , n186178 , n186220 );
buf ( n186222 , n846 );
buf ( n186223 , n866 );
xor ( n18929 , n186222 , n186223 );
buf ( n186225 , n18929 );
buf ( n186226 , n186225 );
not ( n18932 , n186226 );
and ( n18933 , n867 , n866 );
not ( n18934 , n867 );
not ( n18935 , n866 );
and ( n18936 , n18934 , n18935 );
nor ( n18937 , n18933 , n18936 );
not ( n18938 , n18937 );
buf ( n186234 , n867 );
buf ( n186235 , n868 );
xor ( n18941 , n186234 , n186235 );
buf ( n186237 , n18941 );
nor ( n18943 , n18938 , n186237 );
buf ( n186239 , n18943 );
buf ( n18945 , n186239 );
buf ( n186241 , n18945 );
buf ( n186242 , n186241 );
not ( n18948 , n186242 );
or ( n18949 , n18932 , n18948 );
buf ( n186245 , n867 );
buf ( n186246 , n868 );
xor ( n18952 , n186245 , n186246 );
buf ( n186248 , n18952 );
buf ( n186249 , n186248 );
not ( n18955 , n186249 );
buf ( n186251 , n18955 );
buf ( n186252 , n186251 );
not ( n18958 , n186252 );
buf ( n186254 , n18958 );
buf ( n186255 , n186254 );
buf ( n186256 , n845 );
buf ( n186257 , n866 );
xor ( n18963 , n186256 , n186257 );
buf ( n186259 , n18963 );
buf ( n186260 , n186259 );
nand ( n18969 , n186255 , n186260 );
buf ( n186262 , n18969 );
buf ( n186263 , n186262 );
nand ( n18972 , n18949 , n186263 );
buf ( n186265 , n18972 );
buf ( n186266 , n186265 );
buf ( n186267 , n838 );
buf ( n186268 , n874 );
xor ( n18977 , n186267 , n186268 );
buf ( n186270 , n18977 );
buf ( n186271 , n186270 );
not ( n18980 , n186271 );
buf ( n186273 , n875 );
not ( n18982 , n186273 );
buf ( n186275 , n876 );
nand ( n18984 , n18982 , n186275 );
buf ( n186277 , n18984 );
buf ( n186278 , n876 );
not ( n18987 , n186278 );
buf ( n186280 , n875 );
nand ( n18989 , n18987 , n186280 );
buf ( n186282 , n18989 );
xor ( n18991 , n874 , n875 );
and ( n18992 , n186277 , n186282 , n18991 );
buf ( n186285 , n18992 );
buf ( n18994 , n186285 );
buf ( n186287 , n18994 );
buf ( n186288 , n186287 );
not ( n18997 , n186288 );
or ( n18998 , n18980 , n18997 );
xor ( n18999 , n876 , n875 );
buf ( n186292 , n18999 );
not ( n19001 , n186292 );
buf ( n186294 , n19001 );
buf ( n186295 , n186294 );
not ( n19004 , n186295 );
buf ( n186297 , n19004 );
buf ( n186298 , n186297 );
buf ( n186299 , n837 );
buf ( n186300 , n874 );
xor ( n19009 , n186299 , n186300 );
buf ( n186302 , n19009 );
buf ( n186303 , n186302 );
nand ( n19012 , n186298 , n186303 );
buf ( n186305 , n19012 );
buf ( n186306 , n186305 );
nand ( n19015 , n18998 , n186306 );
buf ( n186308 , n19015 );
buf ( n186309 , n186308 );
xor ( n19018 , n186266 , n186309 );
not ( n19019 , n865 );
not ( n19020 , n864 );
not ( n19021 , n19020 );
or ( n19022 , n19019 , n19021 );
nand ( n19023 , n19022 , n866 );
not ( n19024 , n864 );
not ( n19025 , n865 );
not ( n19026 , n19025 );
or ( n19027 , n19024 , n19026 );
not ( n19028 , n866 );
nand ( n19029 , n19027 , n19028 );
nand ( n19030 , n19023 , n19029 );
not ( n19031 , n19030 );
buf ( n186324 , n19031 );
not ( n19033 , n186324 );
buf ( n186326 , n19033 );
buf ( n186327 , n186326 );
buf ( n186328 , n848 );
buf ( n186329 , n864 );
xnor ( n19038 , n186328 , n186329 );
buf ( n186331 , n19038 );
buf ( n186332 , n186331 );
or ( n19041 , n186327 , n186332 );
buf ( n186334 , n865 );
buf ( n186335 , n866 );
xor ( n19044 , n186334 , n186335 );
buf ( n186337 , n19044 );
buf ( n186338 , n186337 );
buf ( n19050 , n186338 );
buf ( n186340 , n19050 );
buf ( n186341 , n186340 );
not ( n19053 , n186341 );
buf ( n186343 , n19053 );
buf ( n186344 , n186343 );
buf ( n186345 , n847 );
buf ( n186346 , n864 );
xor ( n19058 , n186345 , n186346 );
buf ( n186348 , n19058 );
buf ( n186349 , n186348 );
not ( n19061 , n186349 );
buf ( n186351 , n19061 );
buf ( n186352 , n186351 );
or ( n19064 , n186344 , n186352 );
nand ( n19065 , n19041 , n19064 );
buf ( n186355 , n19065 );
buf ( n186356 , n186355 );
and ( n19068 , n19018 , n186356 );
and ( n19069 , n186266 , n186309 );
or ( n19070 , n19068 , n19069 );
buf ( n186360 , n19070 );
buf ( n186361 , n186360 );
and ( n19073 , n18926 , n186361 );
and ( n19074 , n186178 , n186220 );
or ( n19075 , n19073 , n19074 );
buf ( n186365 , n19075 );
buf ( n186366 , n186365 );
buf ( n186367 , n848 );
buf ( n186368 , n864 );
and ( n19080 , n186367 , n186368 );
buf ( n186370 , n19080 );
not ( n19082 , n186370 );
buf ( n186372 , n835 );
buf ( n186373 , n876 );
xor ( n186374 , n186372 , n186373 );
buf ( n186375 , n186374 );
buf ( n186376 , n186375 );
not ( n19088 , n186376 );
not ( n19089 , n876 );
not ( n19090 , n19089 );
nand ( n19091 , n877 , n878 );
not ( n19092 , n19091 );
or ( n19093 , n19090 , n19092 );
or ( n19094 , n877 , n878 );
nand ( n19095 , n19094 , n876 );
nand ( n19096 , n19093 , n19095 );
not ( n19097 , n19096 );
buf ( n19098 , n19097 );
buf ( n186388 , n19098 );
not ( n19100 , n186388 );
or ( n19101 , n19088 , n19100 );
xor ( n19102 , n877 , n878 );
buf ( n19103 , n19102 );
buf ( n186393 , n19103 );
buf ( n19105 , n186393 );
buf ( n186395 , n19105 );
buf ( n186396 , n186395 );
buf ( n186397 , n834 );
buf ( n186398 , n876 );
xor ( n19110 , n186397 , n186398 );
buf ( n186400 , n19110 );
buf ( n186401 , n186400 );
nand ( n19113 , n186396 , n186401 );
buf ( n186403 , n19113 );
buf ( n186404 , n186403 );
nand ( n19116 , n19101 , n186404 );
buf ( n186406 , n19116 );
not ( n19118 , n186406 );
xor ( n19119 , n19082 , n19118 );
buf ( n186409 , n841 );
buf ( n186410 , n870 );
xor ( n19125 , n186409 , n186410 );
buf ( n186412 , n19125 );
buf ( n186413 , n186412 );
not ( n19128 , n186413 );
not ( n19129 , n871 );
not ( n19130 , n872 );
not ( n19131 , n19130 );
or ( n19132 , n19129 , n19131 );
buf ( n186419 , n871 );
not ( n19134 , n186419 );
buf ( n186421 , n872 );
nand ( n19136 , n19134 , n186421 );
buf ( n186423 , n19136 );
nand ( n19138 , n19132 , n186423 );
buf ( n186425 , n19138 );
xnor ( n19140 , n870 , n871 );
buf ( n186427 , n19140 );
nor ( n19142 , n186425 , n186427 );
buf ( n186429 , n19142 );
buf ( n186430 , n186429 );
buf ( n19145 , n186430 );
buf ( n186432 , n19145 );
buf ( n186433 , n186432 );
buf ( n19148 , n186433 );
buf ( n186435 , n19148 );
buf ( n186436 , n186435 );
not ( n19151 , n186436 );
or ( n19152 , n19128 , n19151 );
buf ( n186439 , n19138 );
buf ( n19154 , n186439 );
buf ( n186441 , n19154 );
buf ( n186442 , n186441 );
buf ( n19157 , n186442 );
buf ( n186444 , n19157 );
buf ( n186445 , n186444 );
buf ( n186446 , n840 );
buf ( n186447 , n870 );
xor ( n19162 , n186446 , n186447 );
buf ( n186449 , n19162 );
buf ( n186450 , n186449 );
nand ( n19165 , n186445 , n186450 );
buf ( n186452 , n19165 );
buf ( n186453 , n186452 );
nand ( n19168 , n19152 , n186453 );
buf ( n186455 , n19168 );
xor ( n19170 , n19119 , n186455 );
buf ( n186457 , n836 );
buf ( n186458 , n876 );
xor ( n19173 , n186457 , n186458 );
buf ( n186460 , n19173 );
buf ( n186461 , n186460 );
not ( n19176 , n186461 );
buf ( n19177 , n19097 );
buf ( n186464 , n19177 );
not ( n19179 , n186464 );
or ( n19180 , n19176 , n19179 );
buf ( n186467 , n186395 );
buf ( n186468 , n186375 );
nand ( n19186 , n186467 , n186468 );
buf ( n186470 , n19186 );
buf ( n186471 , n186470 );
nand ( n19189 , n19180 , n186471 );
buf ( n186473 , n19189 );
not ( n19191 , n186473 );
buf ( n186475 , n844 );
buf ( n186476 , n868 );
xor ( n19194 , n186475 , n186476 );
buf ( n186478 , n19194 );
buf ( n186479 , n186478 );
not ( n19197 , n186479 );
buf ( n186481 , n186197 );
not ( n19199 , n186481 );
or ( n19200 , n19197 , n19199 );
buf ( n19201 , n18907 );
buf ( n186485 , n19201 );
buf ( n186486 , n186182 );
nand ( n19204 , n186485 , n186486 );
buf ( n186488 , n19204 );
buf ( n186489 , n186488 );
nand ( n19207 , n19200 , n186489 );
buf ( n186491 , n19207 );
buf ( n186492 , n186491 );
not ( n19210 , n186492 );
buf ( n186494 , n19210 );
nand ( n19212 , n19191 , n186494 );
not ( n19213 , n19212 );
buf ( n186497 , n842 );
buf ( n186498 , n870 );
xor ( n19216 , n186497 , n186498 );
buf ( n186500 , n19216 );
buf ( n186501 , n186500 );
not ( n19219 , n186501 );
buf ( n186503 , n186435 );
not ( n19221 , n186503 );
or ( n19222 , n19219 , n19221 );
buf ( n186506 , n186444 );
buf ( n186507 , n186412 );
nand ( n19225 , n186506 , n186507 );
buf ( n186509 , n19225 );
buf ( n186510 , n186509 );
nand ( n19228 , n19222 , n186510 );
buf ( n186512 , n19228 );
not ( n19230 , n186512 );
or ( n19231 , n19213 , n19230 );
buf ( n186515 , n186473 );
buf ( n186516 , n186491 );
nand ( n19234 , n186515 , n186516 );
buf ( n186518 , n19234 );
nand ( n186519 , n19231 , n186518 );
or ( n19240 , n19170 , n186519 );
buf ( n186521 , n849 );
buf ( n186522 , n864 );
and ( n19243 , n186521 , n186522 );
buf ( n186524 , n19243 );
buf ( n186525 , n840 );
buf ( n186526 , n872 );
xor ( n19247 , n186525 , n186526 );
buf ( n186528 , n19247 );
buf ( n186529 , n186528 );
not ( n19250 , n186529 );
xor ( n19251 , n873 , n874 );
buf ( n186532 , n19251 );
not ( n19253 , n186532 );
buf ( n186534 , n19253 );
buf ( n186535 , n872 );
buf ( n186536 , n873 );
xor ( n19257 , n186535 , n186536 );
buf ( n186538 , n19257 );
nand ( n186539 , n186534 , n186538 );
not ( n19260 , n186539 );
buf ( n186541 , n19260 );
not ( n19262 , n186541 );
or ( n19263 , n19250 , n19262 );
buf ( n19264 , n19251 );
buf ( n19265 , n19264 );
buf ( n186546 , n19265 );
buf ( n186547 , n839 );
buf ( n186548 , n872 );
xor ( n19269 , n186547 , n186548 );
buf ( n186550 , n19269 );
buf ( n186551 , n186550 );
nand ( n19272 , n186546 , n186551 );
buf ( n186553 , n19272 );
buf ( n186554 , n186553 );
nand ( n19275 , n19263 , n186554 );
buf ( n186556 , n19275 );
xor ( n19277 , n186524 , n186556 );
buf ( n186558 , n834 );
buf ( n186559 , n878 );
xor ( n186560 , n186558 , n186559 );
buf ( n186561 , n186560 );
buf ( n186562 , n186561 );
not ( n186563 , n186562 );
xnor ( n186564 , n879 , n878 );
xor ( n186565 , n879 , n880 );
nor ( n186566 , n186564 , n186565 );
buf ( n186567 , n186566 );
buf ( n186568 , n186567 );
buf ( n186569 , n186568 );
buf ( n186570 , n186569 );
not ( n186571 , n186570 );
or ( n186572 , n186563 , n186571 );
buf ( n186573 , n186565 );
buf ( n186574 , n186573 );
buf ( n186575 , n186574 );
buf ( n186576 , n186575 );
buf ( n186577 , n833 );
buf ( n186578 , n878 );
xor ( n186579 , n186577 , n186578 );
buf ( n186580 , n186579 );
buf ( n186581 , n186580 );
nand ( n186582 , n186576 , n186581 );
buf ( n186583 , n186582 );
buf ( n186584 , n186583 );
nand ( n186585 , n186572 , n186584 );
buf ( n186586 , n186585 );
and ( n186587 , n19277 , n186586 );
and ( n186588 , n186524 , n186556 );
or ( n186589 , n186587 , n186588 );
nand ( n186590 , n19240 , n186589 );
nand ( n186591 , n186519 , n19170 );
nand ( n186592 , n186590 , n186591 );
buf ( n186593 , n186592 );
xor ( n186594 , n186366 , n186593 );
buf ( n186595 , n186370 );
not ( n186596 , n186595 );
buf ( n186597 , n186406 );
not ( n186598 , n186597 );
or ( n186599 , n186596 , n186598 );
buf ( n186600 , n186406 );
buf ( n186601 , n186370 );
or ( n186602 , n186600 , n186601 );
buf ( n186603 , n186455 );
nand ( n186604 , n186602 , n186603 );
buf ( n186605 , n186604 );
buf ( n186606 , n186605 );
nand ( n186607 , n186599 , n186606 );
buf ( n186608 , n186607 );
buf ( n186609 , n186608 );
buf ( n186610 , n186259 );
not ( n186611 , n186610 );
buf ( n186612 , n186241 );
not ( n186613 , n186612 );
or ( n186614 , n186611 , n186613 );
buf ( n186615 , n186254 );
buf ( n186616 , n844 );
buf ( n186617 , n866 );
xor ( n186618 , n186616 , n186617 );
buf ( n186619 , n186618 );
buf ( n186620 , n186619 );
nand ( n186621 , n186615 , n186620 );
buf ( n186622 , n186621 );
buf ( n186623 , n186622 );
nand ( n186624 , n186614 , n186623 );
buf ( n186625 , n186624 );
buf ( n186626 , n186625 );
not ( n186627 , n19265 );
buf ( n186628 , n838 );
buf ( n186629 , n872 );
xor ( n186630 , n186628 , n186629 );
buf ( n186631 , n186630 );
not ( n186632 , n186631 );
or ( n186633 , n186627 , n186632 );
nand ( n186634 , n186550 , n19260 );
nand ( n186635 , n186633 , n186634 );
buf ( n186636 , n186635 );
xor ( n186637 , n186626 , n186636 );
buf ( n186638 , n186348 );
not ( n186639 , n186638 );
buf ( n186640 , n19031 );
buf ( n186641 , n186640 );
not ( n186642 , n186641 );
or ( n186643 , n186639 , n186642 );
buf ( n186644 , n186340 );
xor ( n186645 , n864 , n846 );
buf ( n186646 , n186645 );
nand ( n186647 , n186644 , n186646 );
buf ( n186648 , n186647 );
buf ( n186649 , n186648 );
nand ( n186650 , n186643 , n186649 );
buf ( n186651 , n186650 );
buf ( n186652 , n186651 );
and ( n186653 , n186637 , n186652 );
and ( n186654 , n186626 , n186636 );
or ( n186655 , n186653 , n186654 );
buf ( n186656 , n186655 );
buf ( n186657 , n186656 );
xor ( n186658 , n186609 , n186657 );
buf ( n186659 , n186580 );
not ( n186660 , n186659 );
buf ( n186661 , n186569 );
not ( n186662 , n186661 );
or ( n186663 , n186660 , n186662 );
buf ( n186664 , n186575 );
buf ( n186665 , n832 );
buf ( n186666 , n878 );
xor ( n186667 , n186665 , n186666 );
buf ( n186668 , n186667 );
buf ( n186669 , n186668 );
nand ( n186670 , n186664 , n186669 );
buf ( n186671 , n186670 );
buf ( n186672 , n186671 );
nand ( n186673 , n186663 , n186672 );
buf ( n186674 , n186673 );
buf ( n186675 , n186674 );
buf ( n186676 , n18875 );
buf ( n186677 , n18862 );
or ( n186678 , n186676 , n186677 );
buf ( n186679 , n880 );
nand ( n186680 , n186678 , n186679 );
buf ( n186681 , n186680 );
buf ( n186682 , n186681 );
xor ( n186683 , n186675 , n186682 );
buf ( n186684 , n186302 );
not ( n186685 , n186684 );
buf ( n186686 , n186287 );
not ( n186687 , n186686 );
or ( n19411 , n186685 , n186687 );
buf ( n186689 , n186297 );
buf ( n186690 , n836 );
buf ( n186691 , n874 );
xor ( n19415 , n186690 , n186691 );
buf ( n186693 , n19415 );
buf ( n186694 , n186693 );
nand ( n19418 , n186689 , n186694 );
buf ( n186696 , n19418 );
buf ( n186697 , n186696 );
nand ( n19421 , n19411 , n186697 );
buf ( n186699 , n19421 );
buf ( n186700 , n186699 );
and ( n19424 , n186683 , n186700 );
and ( n19425 , n186675 , n186682 );
or ( n19426 , n19424 , n19425 );
buf ( n186704 , n19426 );
buf ( n186705 , n186704 );
xor ( n19429 , n186658 , n186705 );
buf ( n186707 , n19429 );
buf ( n186708 , n186707 );
xor ( n19432 , n186594 , n186708 );
buf ( n186710 , n19432 );
buf ( n186711 , n186710 );
buf ( n186712 , n847 );
buf ( n186713 , n864 );
and ( n19437 , n186712 , n186713 );
buf ( n186715 , n19437 );
buf ( n186716 , n186715 );
buf ( n186717 , n186645 );
not ( n19441 , n186717 );
buf ( n186719 , n19031 );
not ( n19443 , n186719 );
or ( n19444 , n19441 , n19443 );
buf ( n186722 , n186340 );
xor ( n19446 , n864 , n845 );
buf ( n186724 , n19446 );
nand ( n19448 , n186722 , n186724 );
buf ( n186726 , n19448 );
buf ( n186727 , n186726 );
nand ( n19451 , n19444 , n186727 );
buf ( n186729 , n19451 );
buf ( n186730 , n186729 );
xor ( n19454 , n186716 , n186730 );
buf ( n186732 , n186631 );
not ( n19456 , n186732 );
buf ( n186734 , n19260 );
not ( n19458 , n186734 );
or ( n19459 , n19456 , n19458 );
buf ( n186737 , n19265 );
xor ( n19461 , n872 , n837 );
buf ( n186739 , n19461 );
nand ( n19463 , n186737 , n186739 );
buf ( n186741 , n19463 );
buf ( n186742 , n186741 );
nand ( n19466 , n19459 , n186742 );
buf ( n186744 , n19466 );
buf ( n186745 , n186744 );
xor ( n19469 , n19454 , n186745 );
buf ( n186747 , n19469 );
buf ( n186748 , n186747 );
buf ( n186749 , n186619 );
not ( n19473 , n186749 );
buf ( n186751 , n186241 );
not ( n19475 , n186751 );
or ( n19476 , n19473 , n19475 );
buf ( n186754 , n186254 );
buf ( n186755 , n843 );
buf ( n186756 , n866 );
xor ( n19480 , n186755 , n186756 );
buf ( n186758 , n19480 );
buf ( n186759 , n186758 );
nand ( n19483 , n186754 , n186759 );
buf ( n186761 , n19483 );
buf ( n186762 , n186761 );
nand ( n19486 , n19476 , n186762 );
buf ( n186764 , n19486 );
buf ( n186765 , n186764 );
buf ( n186766 , n186213 );
not ( n19490 , n186766 );
buf ( n186768 , n186197 );
not ( n19492 , n186768 );
or ( n19493 , n19490 , n19492 );
buf ( n19494 , n18907 );
buf ( n186772 , n19494 );
buf ( n186773 , n841 );
buf ( n186774 , n868 );
xor ( n19498 , n186773 , n186774 );
buf ( n186776 , n19498 );
buf ( n186777 , n186776 );
nand ( n19501 , n186772 , n186777 );
buf ( n186779 , n19501 );
buf ( n186780 , n186779 );
nand ( n19504 , n19493 , n186780 );
buf ( n186782 , n19504 );
buf ( n186783 , n186782 );
xor ( n19507 , n186765 , n186783 );
buf ( n186785 , n186668 );
not ( n19509 , n186785 );
buf ( n186787 , n186569 );
buf ( n19511 , n186787 );
buf ( n186789 , n19511 );
buf ( n186790 , n186789 );
not ( n19514 , n186790 );
or ( n19515 , n19509 , n19514 );
buf ( n186793 , n186575 );
buf ( n186794 , n878 );
nand ( n19518 , n186793 , n186794 );
buf ( n186796 , n19518 );
buf ( n186797 , n186796 );
nand ( n19521 , n19515 , n186797 );
buf ( n186799 , n19521 );
buf ( n186800 , n186799 );
not ( n19524 , n186800 );
buf ( n186802 , n19524 );
buf ( n186803 , n186802 );
xor ( n19527 , n19507 , n186803 );
buf ( n186805 , n19527 );
buf ( n186806 , n186805 );
xor ( n19530 , n186748 , n186806 );
buf ( n186808 , n186449 );
not ( n19532 , n186808 );
buf ( n186810 , n186435 );
not ( n19534 , n186810 );
or ( n19535 , n19532 , n19534 );
buf ( n186813 , n186444 );
xor ( n19537 , n870 , n839 );
buf ( n186815 , n19537 );
nand ( n19539 , n186813 , n186815 );
buf ( n186817 , n19539 );
buf ( n186818 , n186817 );
nand ( n19542 , n19535 , n186818 );
buf ( n186820 , n19542 );
buf ( n186821 , n186820 );
buf ( n186822 , n186693 );
not ( n19546 , n186822 );
buf ( n186824 , n186287 );
not ( n19548 , n186824 );
or ( n19549 , n19546 , n19548 );
buf ( n186827 , n186297 );
xor ( n19551 , n874 , n835 );
buf ( n186829 , n19551 );
nand ( n19553 , n186827 , n186829 );
buf ( n186831 , n19553 );
buf ( n186832 , n186831 );
nand ( n19556 , n19549 , n186832 );
buf ( n186834 , n19556 );
buf ( n186835 , n186834 );
xor ( n19559 , n186821 , n186835 );
buf ( n186837 , n186400 );
not ( n19561 , n186837 );
buf ( n186839 , n19177 );
not ( n19563 , n186839 );
or ( n19564 , n19561 , n19563 );
buf ( n186842 , n186395 );
xor ( n19566 , n876 , n833 );
buf ( n186844 , n19566 );
nand ( n19568 , n186842 , n186844 );
buf ( n186846 , n19568 );
buf ( n186847 , n186846 );
nand ( n19571 , n19564 , n186847 );
buf ( n186849 , n19571 );
buf ( n186850 , n186849 );
xor ( n19574 , n19559 , n186850 );
buf ( n186852 , n19574 );
buf ( n186853 , n186852 );
xor ( n19577 , n19530 , n186853 );
buf ( n186855 , n19577 );
buf ( n186856 , n186855 );
xor ( n19580 , n186626 , n186636 );
xor ( n19581 , n19580 , n186652 );
buf ( n186859 , n19581 );
buf ( n186860 , n186859 );
xor ( n19584 , n186675 , n186682 );
xor ( n19585 , n19584 , n186700 );
buf ( n186863 , n19585 );
buf ( n186864 , n186863 );
xor ( n19588 , n186860 , n186864 );
xor ( n19589 , n186178 , n186220 );
xor ( n19590 , n19589 , n186361 );
buf ( n186868 , n19590 );
buf ( n186869 , n186868 );
and ( n19593 , n19588 , n186869 );
and ( n19594 , n186860 , n186864 );
or ( n19595 , n19593 , n19594 );
buf ( n186873 , n19595 );
buf ( n186874 , n186873 );
xor ( n19598 , n186856 , n186874 );
buf ( n186876 , n186177 );
not ( n19600 , n186876 );
xor ( n19601 , n883 , n884 );
not ( n19602 , n19601 );
buf ( n186880 , n19602 );
not ( n19604 , n186880 );
and ( n19605 , n883 , n882 );
not ( n19606 , n883 );
not ( n19607 , n882 );
and ( n19608 , n19606 , n19607 );
nor ( n19609 , n19605 , n19608 );
not ( n19610 , n19609 );
xor ( n19611 , n883 , n884 );
nor ( n19612 , n19610 , n19611 );
buf ( n19613 , n19612 );
buf ( n186891 , n19613 );
not ( n19615 , n186891 );
buf ( n186893 , n19615 );
buf ( n186894 , n186893 );
not ( n19618 , n186894 );
or ( n19619 , n19604 , n19618 );
buf ( n186897 , n882 );
nand ( n19621 , n19619 , n186897 );
buf ( n186899 , n19621 );
buf ( n186900 , n186899 );
buf ( n186901 , n837 );
buf ( n186902 , n876 );
xor ( n19626 , n186901 , n186902 );
buf ( n186904 , n19626 );
buf ( n186905 , n186904 );
not ( n19629 , n186905 );
buf ( n186907 , n19098 );
not ( n19631 , n186907 );
or ( n19632 , n19629 , n19631 );
buf ( n186910 , n186395 );
buf ( n186911 , n186460 );
nand ( n19635 , n186910 , n186911 );
buf ( n186913 , n19635 );
buf ( n186914 , n186913 );
nand ( n19638 , n19632 , n186914 );
buf ( n186916 , n19638 );
buf ( n186917 , n186916 );
xor ( n19641 , n186900 , n186917 );
xor ( n19642 , n880 , n833 );
buf ( n186920 , n19642 );
not ( n19644 , n186920 );
buf ( n186922 , n18862 );
buf ( n19646 , n186922 );
buf ( n186924 , n19646 );
buf ( n186925 , n186924 );
not ( n19649 , n186925 );
or ( n19650 , n19644 , n19649 );
buf ( n186928 , n18875 );
buf ( n186929 , n186148 );
nand ( n19653 , n186928 , n186929 );
buf ( n186931 , n19653 );
buf ( n186932 , n186931 );
nand ( n19656 , n19650 , n186932 );
buf ( n186934 , n19656 );
buf ( n186935 , n186934 );
and ( n19659 , n19641 , n186935 );
and ( n19660 , n186900 , n186917 );
or ( n19661 , n19659 , n19660 );
buf ( n186939 , n19661 );
buf ( n186940 , n186939 );
not ( n19664 , n186940 );
buf ( n186942 , n19664 );
buf ( n186943 , n186942 );
not ( n19667 , n186943 );
or ( n19668 , n19600 , n19667 );
xor ( n19669 , n868 , n845 );
buf ( n186947 , n19669 );
not ( n19671 , n186947 );
buf ( n186949 , n186197 );
not ( n19673 , n186949 );
or ( n19674 , n19671 , n19673 );
buf ( n186952 , n18907 );
buf ( n186953 , n186478 );
nand ( n19677 , n186952 , n186953 );
buf ( n186955 , n19677 );
buf ( n186956 , n186955 );
nand ( n19680 , n19674 , n186956 );
buf ( n186958 , n19680 );
buf ( n186959 , n186958 );
not ( n19683 , n186959 );
buf ( n186961 , n847 );
buf ( n186962 , n866 );
xor ( n19686 , n186961 , n186962 );
buf ( n186964 , n19686 );
buf ( n186965 , n186964 );
not ( n19689 , n186965 );
buf ( n186967 , n186241 );
not ( n19691 , n186967 );
or ( n19692 , n19689 , n19691 );
buf ( n186970 , n186254 );
buf ( n186971 , n186225 );
nand ( n19695 , n186970 , n186971 );
buf ( n186973 , n19695 );
buf ( n186974 , n186973 );
nand ( n19698 , n19692 , n186974 );
buf ( n186976 , n19698 );
buf ( n186977 , n186976 );
not ( n19701 , n186977 );
or ( n19702 , n19683 , n19701 );
buf ( n186980 , n186958 );
not ( n19704 , n186980 );
buf ( n186982 , n19704 );
buf ( n186983 , n186982 );
not ( n19707 , n186983 );
buf ( n186985 , n186976 );
not ( n19709 , n186985 );
buf ( n186987 , n19709 );
buf ( n186988 , n186987 );
not ( n19712 , n186988 );
or ( n19713 , n19707 , n19712 );
buf ( n186991 , n839 );
buf ( n186992 , n874 );
xor ( n19716 , n186991 , n186992 );
buf ( n186994 , n19716 );
buf ( n186995 , n186994 );
not ( n19719 , n186995 );
buf ( n186997 , n186287 );
not ( n19721 , n186997 );
or ( n19722 , n19719 , n19721 );
buf ( n187000 , n186297 );
buf ( n187001 , n186270 );
nand ( n19725 , n187000 , n187001 );
buf ( n187003 , n19725 );
buf ( n187004 , n187003 );
nand ( n19728 , n19722 , n187004 );
buf ( n187006 , n19728 );
buf ( n187007 , n187006 );
nand ( n19731 , n19713 , n187007 );
buf ( n187009 , n19731 );
buf ( n187010 , n187009 );
nand ( n19734 , n19702 , n187010 );
buf ( n187012 , n19734 );
buf ( n187013 , n187012 );
nand ( n19737 , n19668 , n187013 );
buf ( n187015 , n19737 );
buf ( n187016 , n187015 );
buf ( n187017 , n186177 );
not ( n19741 , n187017 );
buf ( n187019 , n186939 );
nand ( n19743 , n19741 , n187019 );
buf ( n187021 , n19743 );
buf ( n187022 , n187021 );
nand ( n19746 , n187016 , n187022 );
buf ( n187024 , n19746 );
buf ( n187025 , n187024 );
xor ( n19749 , n186524 , n186556 );
xor ( n19750 , n19749 , n186586 );
not ( n19751 , n19750 );
not ( n19752 , n19751 );
xor ( n19753 , n186266 , n186309 );
xor ( n19754 , n19753 , n186356 );
buf ( n187032 , n19754 );
not ( n19756 , n187032 );
not ( n19757 , n19756 );
or ( n19758 , n19752 , n19757 );
and ( n19759 , n850 , n864 );
buf ( n187037 , n849 );
buf ( n187038 , n864 );
xor ( n19762 , n187037 , n187038 );
buf ( n187040 , n19762 );
not ( n19764 , n187040 );
not ( n19765 , n19031 );
or ( n19766 , n19764 , n19765 );
buf ( n187044 , n186331 );
not ( n19768 , n187044 );
buf ( n187046 , n186340 );
nand ( n19770 , n19768 , n187046 );
buf ( n187048 , n19770 );
nand ( n19772 , n19766 , n187048 );
xor ( n19773 , n19759 , n19772 );
not ( n19774 , n186789 );
buf ( n187052 , n835 );
buf ( n187053 , n878 );
xor ( n19777 , n187052 , n187053 );
buf ( n187055 , n19777 );
not ( n19779 , n187055 );
or ( n19780 , n19774 , n19779 );
buf ( n187058 , n186575 );
buf ( n187059 , n186561 );
nand ( n19783 , n187058 , n187059 );
buf ( n187061 , n19783 );
nand ( n19785 , n19780 , n187061 );
and ( n19786 , n19773 , n19785 );
and ( n19787 , n19759 , n19772 );
or ( n19788 , n19786 , n19787 );
nand ( n19789 , n19758 , n19788 );
not ( n19790 , n19756 );
nand ( n19791 , n19790 , n19750 );
nand ( n19792 , n19789 , n19791 );
buf ( n187070 , n19792 );
xor ( n19794 , n187025 , n187070 );
nand ( n19795 , n186519 , n19170 , n186589 );
not ( n19796 , n186519 );
xor ( n19797 , n19082 , n19118 );
xnor ( n19798 , n19797 , n186455 );
nand ( n19799 , n19796 , n19798 , n186589 );
nor ( n19800 , n19798 , n186589 );
nand ( n19801 , n19800 , n19796 );
not ( n19802 , n186589 );
nand ( n19803 , n19802 , n186519 , n19798 );
nand ( n19804 , n19795 , n19799 , n19801 , n19803 );
buf ( n187082 , n19804 );
and ( n19806 , n19794 , n187082 );
and ( n19807 , n187025 , n187070 );
or ( n19808 , n19806 , n19807 );
buf ( n187086 , n19808 );
buf ( n187087 , n187086 );
xor ( n19811 , n19598 , n187087 );
buf ( n187089 , n19811 );
buf ( n187090 , n187089 );
xor ( n19814 , n186711 , n187090 );
xor ( n19815 , n186860 , n186864 );
xor ( n19816 , n19815 , n186869 );
buf ( n187094 , n19816 );
buf ( n187095 , n187094 );
buf ( n187096 , n186924 );
buf ( n187097 , n834 );
buf ( n187098 , n880 );
xor ( n19822 , n187097 , n187098 );
buf ( n187100 , n19822 );
buf ( n187101 , n187100 );
and ( n19825 , n187096 , n187101 );
buf ( n187103 , n18875 );
buf ( n187104 , n19642 );
and ( n19828 , n187103 , n187104 );
nor ( n19829 , n19825 , n19828 );
buf ( n187107 , n19829 );
buf ( n187108 , n187107 );
not ( n19832 , n187108 );
buf ( n187110 , n19832 );
buf ( n187111 , n187110 );
xor ( n19835 , n870 , n843 );
buf ( n187113 , n19835 );
not ( n19837 , n187113 );
buf ( n187115 , n186435 );
not ( n19839 , n187115 );
or ( n19840 , n19837 , n19839 );
buf ( n187118 , n186444 );
buf ( n187119 , n186500 );
nand ( n19843 , n187118 , n187119 );
buf ( n187121 , n19843 );
buf ( n187122 , n187121 );
nand ( n19846 , n19840 , n187122 );
buf ( n187124 , n19846 );
buf ( n187125 , n187124 );
xor ( n19849 , n187111 , n187125 );
buf ( n187127 , n841 );
buf ( n187128 , n872 );
xor ( n19852 , n187127 , n187128 );
buf ( n187130 , n19852 );
buf ( n187131 , n187130 );
not ( n19855 , n187131 );
buf ( n187133 , n19260 );
not ( n19857 , n187133 );
or ( n19858 , n19855 , n19857 );
buf ( n187136 , n19265 );
buf ( n187137 , n186528 );
nand ( n19861 , n187136 , n187137 );
buf ( n187139 , n19861 );
buf ( n187140 , n187139 );
nand ( n19864 , n19858 , n187140 );
buf ( n187142 , n19864 );
buf ( n187143 , n187142 );
and ( n19867 , n19849 , n187143 );
and ( n19868 , n187111 , n187125 );
or ( n19869 , n19867 , n19868 );
buf ( n187147 , n19869 );
buf ( n187148 , n187147 );
xor ( n19872 , n186494 , n186473 );
xnor ( n19873 , n19872 , n186512 );
buf ( n187151 , n19873 );
xor ( n19875 , n187148 , n187151 );
buf ( n187153 , n848 );
buf ( n187154 , n866 );
xor ( n19878 , n187153 , n187154 );
buf ( n187156 , n19878 );
buf ( n187157 , n187156 );
not ( n19881 , n187157 );
buf ( n187159 , n186241 );
not ( n19883 , n187159 );
or ( n19884 , n19881 , n19883 );
buf ( n187162 , n186254 );
buf ( n187163 , n186964 );
nand ( n19887 , n187162 , n187163 );
buf ( n187165 , n19887 );
buf ( n187166 , n187165 );
nand ( n19890 , n19884 , n187166 );
buf ( n187168 , n19890 );
buf ( n187169 , n187168 );
xor ( n19893 , n868 , n846 );
buf ( n187171 , n19893 );
not ( n19895 , n187171 );
buf ( n187173 , n186197 );
not ( n19897 , n187173 );
or ( n19898 , n19895 , n19897 );
buf ( n187176 , n19494 );
buf ( n187177 , n19669 );
nand ( n19901 , n187176 , n187177 );
buf ( n187179 , n19901 );
buf ( n187180 , n187179 );
nand ( n19904 , n19898 , n187180 );
buf ( n187182 , n19904 );
buf ( n187183 , n187182 );
xor ( n19907 , n187169 , n187183 );
xor ( n19908 , n876 , n838 );
buf ( n187186 , n19908 );
not ( n19910 , n187186 );
buf ( n187188 , n19177 );
not ( n19912 , n187188 );
or ( n19913 , n19910 , n19912 );
buf ( n187191 , n186395 );
buf ( n187192 , n186904 );
nand ( n19916 , n187191 , n187192 );
buf ( n187194 , n19916 );
buf ( n187195 , n187194 );
nand ( n19919 , n19913 , n187195 );
buf ( n187197 , n19919 );
buf ( n187198 , n187197 );
and ( n19922 , n19907 , n187198 );
and ( n19923 , n187169 , n187183 );
or ( n19924 , n19922 , n19923 );
buf ( n187202 , n19924 );
buf ( n187203 , n187202 );
buf ( n187204 , n832 );
buf ( n187205 , n882 );
xor ( n19929 , n187204 , n187205 );
buf ( n187207 , n19929 );
buf ( n187208 , n187207 );
not ( n19932 , n187208 );
buf ( n187210 , n19613 );
not ( n19934 , n187210 );
or ( n19935 , n19932 , n19934 );
not ( n19936 , n883 );
not ( n19937 , n884 );
not ( n19938 , n19937 );
or ( n19939 , n19936 , n19938 );
not ( n19940 , n883 );
nand ( n19941 , n19940 , n884 );
nand ( n19942 , n19939 , n19941 );
buf ( n19943 , n19942 );
buf ( n187221 , n19943 );
buf ( n187222 , n882 );
nand ( n19946 , n187221 , n187222 );
buf ( n187224 , n19946 );
buf ( n187225 , n187224 );
nand ( n19949 , n19935 , n187225 );
buf ( n187227 , n19949 );
buf ( n187228 , n187227 );
buf ( n187229 , n842 );
buf ( n187230 , n872 );
xor ( n19954 , n187229 , n187230 );
buf ( n187232 , n19954 );
buf ( n187233 , n187232 );
not ( n19957 , n187233 );
buf ( n187235 , n19260 );
not ( n19959 , n187235 );
or ( n19960 , n19957 , n19959 );
buf ( n187238 , n19265 );
buf ( n187239 , n187130 );
nand ( n19963 , n187238 , n187239 );
buf ( n187241 , n19963 );
buf ( n187242 , n187241 );
nand ( n19966 , n19960 , n187242 );
buf ( n187244 , n19966 );
buf ( n187245 , n187244 );
xor ( n19969 , n187228 , n187245 );
buf ( n187247 , n836 );
buf ( n187248 , n878 );
xor ( n19972 , n187247 , n187248 );
buf ( n187250 , n19972 );
buf ( n187251 , n187250 );
not ( n19975 , n187251 );
buf ( n187253 , n186789 );
not ( n19977 , n187253 );
or ( n19978 , n19975 , n19977 );
buf ( n187256 , n186575 );
buf ( n187257 , n187055 );
nand ( n19981 , n187256 , n187257 );
buf ( n187259 , n19981 );
buf ( n187260 , n187259 );
nand ( n19984 , n19978 , n187260 );
buf ( n187262 , n19984 );
buf ( n187263 , n187262 );
and ( n19987 , n19969 , n187263 );
and ( n19988 , n187228 , n187245 );
or ( n19989 , n19987 , n19988 );
buf ( n187267 , n19989 );
buf ( n187268 , n187267 );
xor ( n19992 , n187203 , n187268 );
buf ( n187270 , n851 );
buf ( n187271 , n864 );
and ( n19995 , n187270 , n187271 );
buf ( n187273 , n19995 );
buf ( n187274 , n187273 );
buf ( n187275 , n850 );
buf ( n187276 , n864 );
xor ( n20000 , n187275 , n187276 );
buf ( n187278 , n20000 );
buf ( n187279 , n187278 );
not ( n20003 , n187279 );
buf ( n187281 , n19031 );
not ( n20005 , n187281 );
or ( n20006 , n20003 , n20005 );
buf ( n187284 , n186340 );
buf ( n187285 , n187040 );
nand ( n20009 , n187284 , n187285 );
buf ( n187287 , n20009 );
buf ( n187288 , n187287 );
nand ( n20012 , n20006 , n187288 );
buf ( n187290 , n20012 );
buf ( n187291 , n187290 );
xor ( n20015 , n187274 , n187291 );
buf ( n187293 , n840 );
buf ( n187294 , n874 );
xor ( n20018 , n187293 , n187294 );
buf ( n187296 , n20018 );
buf ( n187297 , n187296 );
not ( n20021 , n187297 );
buf ( n187299 , n186287 );
not ( n20023 , n187299 );
or ( n20024 , n20021 , n20023 );
buf ( n187302 , n186297 );
buf ( n187303 , n186994 );
nand ( n20027 , n187302 , n187303 );
buf ( n187305 , n20027 );
buf ( n187306 , n187305 );
nand ( n20030 , n20024 , n187306 );
buf ( n187308 , n20030 );
buf ( n187309 , n187308 );
and ( n20033 , n20015 , n187309 );
and ( n20034 , n187274 , n187291 );
or ( n20035 , n20033 , n20034 );
buf ( n187313 , n20035 );
buf ( n187314 , n187313 );
and ( n20038 , n19992 , n187314 );
and ( n20039 , n187203 , n187268 );
or ( n20040 , n20038 , n20039 );
buf ( n187318 , n20040 );
buf ( n187319 , n187318 );
and ( n20043 , n19875 , n187319 );
and ( n20044 , n187148 , n187151 );
or ( n20045 , n20043 , n20044 );
buf ( n187323 , n20045 );
buf ( n187324 , n187323 );
xor ( n20048 , n187095 , n187324 );
xor ( n20049 , n19759 , n19772 );
xor ( n20050 , n20049 , n19785 );
xor ( n20051 , n186900 , n186917 );
xor ( n20052 , n20051 , n186935 );
buf ( n187330 , n20052 );
xor ( n20054 , n20050 , n187330 );
buf ( n187332 , n187006 );
not ( n20056 , n187332 );
buf ( n187334 , n186982 );
not ( n20058 , n187334 );
buf ( n187336 , n186976 );
not ( n20060 , n187336 );
and ( n20061 , n20058 , n20060 );
buf ( n187339 , n186976 );
buf ( n187340 , n186982 );
and ( n20064 , n187339 , n187340 );
nor ( n20065 , n20061 , n20064 );
buf ( n187343 , n20065 );
buf ( n187344 , n187343 );
not ( n20068 , n187344 );
or ( n20069 , n20056 , n20068 );
buf ( n187347 , n187343 );
buf ( n187348 , n187006 );
or ( n20072 , n187347 , n187348 );
nand ( n20073 , n20069 , n20072 );
buf ( n187351 , n20073 );
and ( n20075 , n20054 , n187351 );
and ( n20076 , n20050 , n187330 );
or ( n20077 , n20075 , n20076 );
buf ( n187355 , n20077 );
and ( n20079 , n19788 , n19750 );
not ( n20080 , n19788 );
and ( n20081 , n20080 , n19751 );
nor ( n20082 , n20079 , n20081 );
and ( n20083 , n20082 , n19790 );
not ( n20084 , n20082 );
and ( n20085 , n20084 , n19756 );
nor ( n20086 , n20083 , n20085 );
buf ( n187364 , n20086 );
or ( n20088 , n187355 , n187364 );
buf ( n187366 , n187012 );
not ( n20090 , n187366 );
buf ( n187368 , n186177 );
not ( n20092 , n187368 );
and ( n20093 , n20090 , n20092 );
buf ( n187371 , n187012 );
buf ( n187372 , n186177 );
and ( n20096 , n187371 , n187372 );
nor ( n20097 , n20093 , n20096 );
buf ( n187375 , n20097 );
buf ( n187376 , n187375 );
buf ( n187377 , n186939 );
and ( n20101 , n187376 , n187377 );
not ( n20102 , n187376 );
buf ( n187380 , n186942 );
and ( n20104 , n20102 , n187380 );
nor ( n20105 , n20101 , n20104 );
buf ( n187383 , n20105 );
buf ( n187384 , n187383 );
not ( n20108 , n187384 );
buf ( n187386 , n20108 );
buf ( n187387 , n187386 );
nand ( n20111 , n20088 , n187387 );
buf ( n187389 , n20111 );
buf ( n187390 , n187389 );
buf ( n187391 , n20086 );
buf ( n187392 , n20077 );
nand ( n20116 , n187391 , n187392 );
buf ( n187394 , n20116 );
buf ( n187395 , n187394 );
nand ( n20119 , n187390 , n187395 );
buf ( n187397 , n20119 );
buf ( n187398 , n187397 );
and ( n20122 , n20048 , n187398 );
and ( n20123 , n187095 , n187324 );
or ( n20124 , n20122 , n20123 );
buf ( n187402 , n20124 );
buf ( n187403 , n187402 );
xor ( n20127 , n19814 , n187403 );
buf ( n187405 , n20127 );
buf ( n20129 , n187405 );
buf ( n187407 , n894 );
buf ( n187408 , n859 );
buf ( n187409 , n866 );
xor ( n20133 , n187408 , n187409 );
buf ( n187411 , n20133 );
buf ( n187412 , n187411 );
not ( n20136 , n187412 );
buf ( n187414 , n186241 );
not ( n20138 , n187414 );
or ( n20139 , n20136 , n20138 );
buf ( n187417 , n186254 );
buf ( n187418 , n858 );
buf ( n187419 , n866 );
xor ( n20143 , n187418 , n187419 );
buf ( n187421 , n20143 );
buf ( n187422 , n187421 );
nand ( n20146 , n187417 , n187422 );
buf ( n187424 , n20146 );
buf ( n187425 , n187424 );
nand ( n20149 , n20139 , n187425 );
buf ( n187427 , n20149 );
buf ( n187428 , n187427 );
xor ( n20152 , n187407 , n187428 );
buf ( n187430 , n863 );
buf ( n187431 , n864 );
and ( n20155 , n187430 , n187431 );
buf ( n187433 , n20155 );
buf ( n187434 , n187433 );
and ( n20158 , n832 , n894 );
not ( n20159 , n832 );
not ( n20160 , n894 );
and ( n20161 , n20159 , n20160 );
nor ( n20162 , n20158 , n20161 );
not ( n20163 , n20162 );
not ( n20164 , n894 );
nor ( n20165 , n20164 , n895 );
not ( n20166 , n20165 );
or ( n20167 , n20163 , n20166 );
nand ( n20168 , n894 , n895 );
nand ( n20169 , n20167 , n20168 );
buf ( n187447 , n20169 );
xor ( n20171 , n187434 , n187447 );
buf ( n187449 , n834 );
buf ( n187450 , n892 );
xor ( n20174 , n187449 , n187450 );
buf ( n187452 , n20174 );
buf ( n187453 , n187452 );
not ( n20177 , n187453 );
and ( n20178 , n893 , n20160 );
not ( n20179 , n893 );
and ( n20180 , n20179 , n894 );
nor ( n20181 , n20178 , n20180 );
not ( n20182 , n892 );
not ( n20183 , n893 );
not ( n20184 , n20183 );
or ( n20185 , n20182 , n20184 );
not ( n20186 , n892 );
nand ( n20187 , n20186 , n893 );
nand ( n20188 , n20185 , n20187 );
nand ( n20189 , n20181 , n20188 );
buf ( n187467 , n20189 );
not ( n20191 , n187467 );
buf ( n187469 , n20191 );
buf ( n187470 , n187469 );
not ( n20194 , n187470 );
or ( n20195 , n20177 , n20194 );
xor ( n20196 , n893 , n894 );
not ( n20197 , n20196 );
buf ( n187475 , n20197 );
not ( n20199 , n187475 );
buf ( n187477 , n20199 );
buf ( n187478 , n187477 );
xor ( n20202 , n892 , n833 );
buf ( n187480 , n20202 );
nand ( n20204 , n187478 , n187480 );
buf ( n187482 , n20204 );
buf ( n187483 , n187482 );
nand ( n20207 , n20195 , n187483 );
buf ( n187485 , n20207 );
buf ( n187486 , n187485 );
and ( n20210 , n20171 , n187486 );
and ( n20211 , n187434 , n187447 );
or ( n20212 , n20210 , n20211 );
buf ( n187490 , n20212 );
buf ( n187491 , n187490 );
and ( n20215 , n20152 , n187491 );
and ( n20216 , n187407 , n187428 );
or ( n20217 , n20215 , n20216 );
buf ( n187495 , n20217 );
buf ( n187496 , n187495 );
not ( n20220 , n187496 );
xor ( n20221 , n882 , n844 );
not ( n20222 , n20221 );
buf ( n187500 , n882 );
buf ( n187501 , n883 );
xnor ( n20225 , n187500 , n187501 );
buf ( n187503 , n20225 );
buf ( n187504 , n187503 );
buf ( n187505 , n19601 );
nor ( n20229 , n187504 , n187505 );
buf ( n187507 , n20229 );
not ( n20231 , n187507 );
or ( n20232 , n20222 , n20231 );
buf ( n187510 , n19601 );
xor ( n20234 , n882 , n843 );
buf ( n187512 , n20234 );
nand ( n20236 , n187510 , n187512 );
buf ( n187514 , n20236 );
nand ( n20238 , n20232 , n187514 );
not ( n20239 , n20238 );
xor ( n20240 , n872 , n854 );
not ( n20241 , n20240 );
xnor ( n20242 , n873 , n874 );
nand ( n20243 , n20242 , n186538 );
not ( n20244 , n20243 );
not ( n20245 , n20244 );
or ( n20246 , n20241 , n20245 );
buf ( n187524 , n19264 );
xor ( n20248 , n872 , n853 );
buf ( n187526 , n20248 );
nand ( n20250 , n187524 , n187526 );
buf ( n187528 , n20250 );
nand ( n20252 , n20246 , n187528 );
not ( n20253 , n20252 );
or ( n20254 , n20239 , n20253 );
or ( n20255 , n20252 , n20238 );
and ( n20256 , n871 , n872 );
not ( n20257 , n871 );
and ( n20258 , n20257 , n19130 );
nor ( n20259 , n20256 , n20258 );
not ( n20260 , n20259 );
buf ( n187538 , n855 );
buf ( n187539 , n870 );
xor ( n20263 , n187538 , n187539 );
buf ( n187541 , n20263 );
not ( n20265 , n187541 );
or ( n20266 , n20260 , n20265 );
not ( n20267 , n20259 );
not ( n20268 , n19140 );
xor ( n20269 , n856 , n870 );
nand ( n20270 , n20267 , n20268 , n20269 );
nand ( n20271 , n20266 , n20270 );
nand ( n20272 , n20255 , n20271 );
nand ( n20273 , n20254 , n20272 );
xor ( n20274 , n876 , n850 );
not ( n20275 , n20274 );
not ( n20276 , n19096 );
not ( n20277 , n20276 );
or ( n20278 , n20275 , n20277 );
buf ( n20279 , n19102 );
buf ( n187557 , n20279 );
xor ( n20281 , n876 , n849 );
buf ( n187559 , n20281 );
nand ( n20283 , n187557 , n187559 );
buf ( n187561 , n20283 );
nand ( n20285 , n20278 , n187561 );
buf ( n187563 , n20285 );
not ( n20287 , n187563 );
xor ( n20288 , n887 , n888 );
not ( n20289 , n20288 );
xor ( n20290 , n886 , n839 );
not ( n20291 , n20290 );
or ( n20292 , n20289 , n20291 );
xor ( n20293 , n887 , n888 );
not ( n20294 , n20293 );
xor ( n20295 , n887 , n886 );
and ( n20296 , n840 , n886 );
not ( n20297 , n840 );
not ( n20298 , n886 );
and ( n20299 , n20297 , n20298 );
nor ( n20300 , n20296 , n20299 );
nand ( n20301 , n20294 , n20295 , n20300 );
nand ( n20302 , n20292 , n20301 );
buf ( n187580 , n20302 );
not ( n20304 , n187580 );
or ( n20305 , n20287 , n20304 );
buf ( n187583 , n20302 );
buf ( n187584 , n20285 );
or ( n20308 , n187583 , n187584 );
buf ( n187586 , n847 );
buf ( n187587 , n878 );
xor ( n20311 , n187586 , n187587 );
buf ( n187589 , n20311 );
not ( n20313 , n187589 );
not ( n20314 , n186575 );
or ( n20315 , n20313 , n20314 );
buf ( n187593 , n848 );
buf ( n187594 , n878 );
xor ( n20318 , n187593 , n187594 );
buf ( n187596 , n20318 );
nand ( n20320 , n187596 , n186566 );
nand ( n20321 , n20315 , n20320 );
buf ( n187599 , n20321 );
nand ( n20323 , n20308 , n187599 );
buf ( n187601 , n20323 );
buf ( n187602 , n187601 );
nand ( n20326 , n20305 , n187602 );
buf ( n187604 , n20326 );
xor ( n20328 , n20273 , n187604 );
buf ( n187606 , n862 );
buf ( n187607 , n864 );
xor ( n20331 , n187606 , n187607 );
buf ( n187609 , n20331 );
buf ( n187610 , n187609 );
not ( n20334 , n187610 );
not ( n20335 , n19030 );
buf ( n187613 , n20335 );
not ( n20337 , n187613 );
or ( n20338 , n20334 , n20337 );
xor ( n20339 , n861 , n864 );
nand ( n20340 , n186337 , n20339 );
buf ( n187618 , n20340 );
nand ( n20342 , n20338 , n187618 );
buf ( n187620 , n20342 );
buf ( n187621 , n187620 );
not ( n20345 , n187621 );
buf ( n187623 , n20345 );
buf ( n187624 , n187623 );
not ( n20348 , n187624 );
buf ( n187626 , n846 );
buf ( n187627 , n880 );
xor ( n20351 , n187626 , n187627 );
buf ( n187629 , n20351 );
buf ( n187630 , n187629 );
not ( n20354 , n187630 );
buf ( n187632 , n18862 );
not ( n20356 , n187632 );
or ( n20357 , n20354 , n20356 );
xor ( n20358 , n881 , n882 );
buf ( n187636 , n20358 );
buf ( n187637 , n845 );
buf ( n187638 , n880 );
xor ( n20362 , n187637 , n187638 );
buf ( n187640 , n20362 );
buf ( n187641 , n187640 );
nand ( n20365 , n187636 , n187641 );
buf ( n187643 , n20365 );
buf ( n187644 , n187643 );
nand ( n20368 , n20357 , n187644 );
buf ( n187646 , n20368 );
buf ( n187647 , n187646 );
not ( n20371 , n187647 );
buf ( n187649 , n20371 );
buf ( n187650 , n187649 );
not ( n20374 , n187650 );
or ( n20375 , n20348 , n20374 );
buf ( n187653 , n838 );
buf ( n187654 , n888 );
xor ( n20378 , n187653 , n187654 );
buf ( n187656 , n20378 );
buf ( n187657 , n187656 );
not ( n20381 , n187657 );
not ( n20382 , n888 );
not ( n20383 , n20382 );
nand ( n20384 , n889 , n890 );
not ( n20385 , n20384 );
not ( n20386 , n20385 );
or ( n20387 , n20383 , n20386 );
nor ( n20388 , n889 , n890 );
nand ( n20389 , n888 , n20388 );
nand ( n20390 , n20387 , n20389 );
buf ( n20391 , n20390 );
buf ( n187669 , n20391 );
not ( n20393 , n187669 );
or ( n20394 , n20381 , n20393 );
xor ( n20395 , n889 , n890 );
buf ( n20396 , n20395 );
buf ( n187674 , n20396 );
xor ( n20398 , n888 , n837 );
buf ( n187676 , n20398 );
nand ( n20400 , n187674 , n187676 );
buf ( n187678 , n20400 );
buf ( n187679 , n187678 );
nand ( n20403 , n20394 , n187679 );
buf ( n187681 , n20403 );
buf ( n187682 , n187681 );
nand ( n20406 , n20375 , n187682 );
buf ( n187684 , n20406 );
buf ( n187685 , n187684 );
buf ( n187686 , n187620 );
buf ( n187687 , n187646 );
nand ( n20411 , n187686 , n187687 );
buf ( n187689 , n20411 );
buf ( n187690 , n187689 );
nand ( n20414 , n187685 , n187690 );
buf ( n187692 , n20414 );
and ( n20416 , n20328 , n187692 );
and ( n20417 , n20273 , n187604 );
or ( n20418 , n20416 , n20417 );
not ( n20419 , n20418 );
not ( n20420 , n20419 );
buf ( n187698 , n20420 );
not ( n20422 , n187698 );
or ( n20423 , n20220 , n20422 );
buf ( n187701 , n187495 );
not ( n20425 , n187701 );
buf ( n187703 , n20425 );
buf ( n187704 , n187703 );
not ( n20428 , n187704 );
buf ( n187706 , n20419 );
not ( n20430 , n187706 );
or ( n20431 , n20428 , n20430 );
xor ( n20432 , n890 , n835 );
buf ( n187710 , n20432 );
not ( n20434 , n187710 );
xnor ( n20435 , n891 , n890 );
xor ( n20436 , n891 , n892 );
nor ( n20437 , n20435 , n20436 );
buf ( n187715 , n20437 );
not ( n20439 , n187715 );
or ( n20440 , n20434 , n20439 );
xor ( n20441 , n890 , n834 );
buf ( n187719 , n20441 );
buf ( n187720 , n20436 );
nand ( n20444 , n187719 , n187720 );
buf ( n187722 , n20444 );
buf ( n187723 , n187722 );
nand ( n20447 , n20440 , n187723 );
buf ( n187725 , n20447 );
buf ( n187726 , n187725 );
xor ( n20450 , n884 , n841 );
buf ( n187728 , n20450 );
not ( n20452 , n187728 );
buf ( n187730 , n885 );
buf ( n187731 , n886 );
xor ( n20455 , n187730 , n187731 );
buf ( n187733 , n20455 );
and ( n20457 , n885 , n884 );
not ( n20458 , n885 );
not ( n20459 , n884 );
and ( n20460 , n20458 , n20459 );
nor ( n20461 , n20457 , n20460 );
not ( n20462 , n20461 );
nor ( n20463 , n187733 , n20462 );
buf ( n187741 , n20463 );
not ( n20465 , n187741 );
or ( n20466 , n20452 , n20465 );
buf ( n187744 , n187733 );
xor ( n20468 , n884 , n840 );
buf ( n187746 , n20468 );
nand ( n20470 , n187744 , n187746 );
buf ( n187748 , n20470 );
buf ( n187749 , n187748 );
nand ( n20473 , n20466 , n187749 );
buf ( n187751 , n20473 );
buf ( n187752 , n187751 );
or ( n20476 , n187726 , n187752 );
buf ( n187754 , n20248 );
not ( n20478 , n187754 );
buf ( n187756 , n20244 );
not ( n20480 , n187756 );
or ( n20481 , n20478 , n20480 );
buf ( n187759 , n19264 );
buf ( n187760 , n852 );
buf ( n187761 , n872 );
xor ( n20485 , n187760 , n187761 );
buf ( n187763 , n20485 );
buf ( n187764 , n187763 );
nand ( n20488 , n187759 , n187764 );
buf ( n187766 , n20488 );
buf ( n187767 , n187766 );
nand ( n20491 , n20481 , n187767 );
buf ( n187769 , n20491 );
buf ( n187770 , n187769 );
nand ( n20494 , n20476 , n187770 );
buf ( n187772 , n20494 );
buf ( n187773 , n187772 );
buf ( n187774 , n187725 );
buf ( n187775 , n187751 );
nand ( n20499 , n187774 , n187775 );
buf ( n187777 , n20499 );
buf ( n187778 , n187777 );
nand ( n20502 , n187773 , n187778 );
buf ( n187780 , n20502 );
buf ( n187781 , n187780 );
buf ( n187782 , n20202 );
not ( n20506 , n187782 );
buf ( n187784 , n187469 );
not ( n20508 , n187784 );
or ( n20509 , n20506 , n20508 );
buf ( n187787 , n187477 );
xor ( n20511 , n892 , n832 );
buf ( n187789 , n20511 );
nand ( n20513 , n187787 , n187789 );
buf ( n187791 , n20513 );
buf ( n187792 , n187791 );
nand ( n20516 , n20509 , n187792 );
buf ( n187794 , n20516 );
buf ( n187795 , n20398 );
not ( n20519 , n187795 );
buf ( n187797 , n20391 );
not ( n20521 , n187797 );
or ( n20522 , n20519 , n20521 );
buf ( n187800 , n20396 );
buf ( n187801 , n836 );
buf ( n187802 , n888 );
xor ( n20526 , n187801 , n187802 );
buf ( n187804 , n20526 );
buf ( n187805 , n187804 );
nand ( n20529 , n187800 , n187805 );
buf ( n187807 , n20529 );
buf ( n187808 , n187807 );
nand ( n20532 , n20522 , n187808 );
buf ( n187810 , n20532 );
xor ( n20534 , n187794 , n187810 );
buf ( n187812 , n187589 );
not ( n20536 , n187812 );
buf ( n187814 , n186569 );
not ( n20538 , n187814 );
or ( n20539 , n20536 , n20538 );
xnor ( n20540 , n878 , n846 );
not ( n20541 , n20540 );
nand ( n20542 , n20541 , n186575 );
buf ( n187820 , n20542 );
nand ( n20544 , n20539 , n187820 );
buf ( n187822 , n20544 );
and ( n20546 , n20534 , n187822 );
and ( n20547 , n187794 , n187810 );
or ( n20548 , n20546 , n20547 );
buf ( n187826 , n20548 );
xor ( n20550 , n187781 , n187826 );
buf ( n187828 , n20290 );
not ( n20552 , n187828 );
nand ( n20553 , n20294 , n20295 );
not ( n20554 , n20553 );
buf ( n187832 , n20554 );
not ( n20556 , n187832 );
or ( n20557 , n20552 , n20556 );
buf ( n20558 , n20288 );
buf ( n187836 , n20558 );
buf ( n187837 , n838 );
buf ( n187838 , n886 );
xor ( n20562 , n187837 , n187838 );
buf ( n187840 , n20562 );
buf ( n187841 , n187840 );
nand ( n20565 , n187836 , n187841 );
buf ( n187843 , n20565 );
buf ( n187844 , n187843 );
nand ( n20568 , n20557 , n187844 );
buf ( n187846 , n20568 );
not ( n20570 , n187846 );
buf ( n187848 , n851 );
buf ( n187849 , n874 );
xor ( n20573 , n187848 , n187849 );
buf ( n187851 , n20573 );
buf ( n187852 , n187851 );
not ( n20576 , n187852 );
buf ( n187854 , n876 );
not ( n20578 , n187854 );
buf ( n187856 , n875 );
nand ( n20580 , n20578 , n187856 );
buf ( n187858 , n20580 );
and ( n20582 , n187858 , n186277 , n18991 );
buf ( n187860 , n20582 );
not ( n20584 , n187860 );
or ( n20585 , n20576 , n20584 );
buf ( n187863 , n186294 );
not ( n20587 , n187863 );
buf ( n187865 , n20587 );
buf ( n187866 , n187865 );
xor ( n20590 , n874 , n850 );
buf ( n187868 , n20590 );
nand ( n20592 , n187866 , n187868 );
buf ( n187870 , n20592 );
buf ( n187871 , n187870 );
nand ( n20595 , n20585 , n187871 );
buf ( n187873 , n20595 );
not ( n20597 , n187873 );
buf ( n187875 , n20281 );
not ( n20599 , n187875 );
buf ( n187877 , n19177 );
not ( n20601 , n187877 );
or ( n20602 , n20599 , n20601 );
buf ( n187880 , n19103 );
xor ( n20604 , n876 , n848 );
buf ( n187882 , n20604 );
nand ( n20606 , n187880 , n187882 );
buf ( n187884 , n20606 );
buf ( n187885 , n187884 );
nand ( n20609 , n20602 , n187885 );
buf ( n187887 , n20609 );
not ( n20611 , n187887 );
nand ( n20612 , n20597 , n20611 );
not ( n20613 , n20612 );
or ( n20614 , n20570 , n20613 );
nand ( n20615 , n187887 , n187873 );
nand ( n20616 , n20614 , n20615 );
buf ( n187894 , n20616 );
xor ( n20618 , n20550 , n187894 );
buf ( n187896 , n20618 );
buf ( n187897 , n187896 );
nand ( n20621 , n20431 , n187897 );
buf ( n187899 , n20621 );
buf ( n187900 , n187899 );
nand ( n20624 , n20423 , n187900 );
buf ( n187902 , n20624 );
buf ( n187903 , n187902 );
buf ( n187904 , n894 );
not ( n20628 , n187904 );
buf ( n187906 , n20628 );
buf ( n187907 , n187906 );
not ( n20631 , n20511 );
not ( n20632 , n20189 );
not ( n20633 , n20632 );
or ( n20634 , n20631 , n20633 );
buf ( n20635 , n187477 );
buf ( n187913 , n20635 );
buf ( n187914 , n892 );
nand ( n20638 , n187913 , n187914 );
buf ( n187916 , n20638 );
nand ( n20640 , n20634 , n187916 );
not ( n20641 , n20640 );
buf ( n187919 , n20641 );
xor ( n20643 , n187907 , n187919 );
buf ( n187921 , n862 );
buf ( n187922 , n864 );
nand ( n20646 , n187921 , n187922 );
buf ( n187924 , n20646 );
buf ( n187925 , n187924 );
not ( n20649 , n187925 );
buf ( n187927 , n20649 );
buf ( n187928 , n187927 );
not ( n20652 , n187928 );
buf ( n187930 , n20339 );
not ( n20654 , n187930 );
buf ( n187932 , n19031 );
not ( n20656 , n187932 );
or ( n20657 , n20654 , n20656 );
buf ( n187935 , n186337 );
xor ( n20659 , n864 , n860 );
buf ( n187937 , n20659 );
nand ( n20661 , n187935 , n187937 );
buf ( n187939 , n20661 );
buf ( n187940 , n187939 );
nand ( n20664 , n20657 , n187940 );
buf ( n187942 , n20664 );
buf ( n187943 , n187942 );
not ( n20667 , n187943 );
or ( n20668 , n20652 , n20667 );
buf ( n187946 , n187640 );
not ( n20670 , n187946 );
nand ( n20671 , n18867 , n882 );
nand ( n20672 , n18856 , n18857 );
nand ( n20673 , n880 , n881 );
nand ( n20674 , n20671 , n20672 , n18874 , n20673 );
not ( n20675 , n20674 );
buf ( n187953 , n20675 );
not ( n20677 , n187953 );
or ( n20678 , n20670 , n20677 );
not ( n20679 , n18874 );
not ( n20680 , n20671 );
or ( n20681 , n20679 , n20680 );
xor ( n20682 , n880 , n844 );
nand ( n20683 , n20681 , n20682 );
buf ( n187961 , n20683 );
nand ( n20685 , n20678 , n187961 );
buf ( n187963 , n20685 );
buf ( n187964 , n187963 );
buf ( n187965 , n19031 );
buf ( n187966 , n20339 );
nand ( n20690 , n187965 , n187966 );
buf ( n187968 , n20690 );
buf ( n187969 , n187968 );
buf ( n187970 , n187939 );
buf ( n187971 , n187924 );
nand ( n20695 , n187969 , n187970 , n187971 );
buf ( n187973 , n20695 );
buf ( n187974 , n187973 );
nand ( n20698 , n187964 , n187974 );
buf ( n187976 , n20698 );
buf ( n187977 , n187976 );
nand ( n20701 , n20668 , n187977 );
buf ( n187979 , n20701 );
buf ( n187980 , n187979 );
xor ( n20704 , n20643 , n187980 );
buf ( n187982 , n20704 );
buf ( n20706 , n187982 );
buf ( n187984 , n20706 );
not ( n20708 , n187984 );
buf ( n187986 , n187924 );
buf ( n187987 , n187963 );
xor ( n20711 , n187986 , n187987 );
buf ( n187989 , n187942 );
xor ( n20713 , n20711 , n187989 );
buf ( n187991 , n20713 );
buf ( n187992 , n187991 );
not ( n20716 , n187992 );
buf ( n187994 , n20716 );
not ( n20718 , n187994 );
buf ( n187996 , n842 );
buf ( n187997 , n884 );
xor ( n20721 , n187996 , n187997 );
buf ( n187999 , n20721 );
buf ( n188000 , n187999 );
not ( n20724 , n188000 );
xnor ( n20725 , n885 , n884 );
nor ( n20726 , n20725 , n187733 );
buf ( n20727 , n20726 );
buf ( n188005 , n20727 );
not ( n20729 , n188005 );
or ( n20730 , n20724 , n20729 );
buf ( n188008 , n187733 );
buf ( n20732 , n188008 );
buf ( n188010 , n20732 );
buf ( n188011 , n188010 );
buf ( n188012 , n20450 );
nand ( n20736 , n188011 , n188012 );
buf ( n188014 , n20736 );
buf ( n188015 , n188014 );
nand ( n20739 , n20730 , n188015 );
buf ( n188017 , n20739 );
not ( n20741 , n188017 );
buf ( n188019 , n836 );
buf ( n188020 , n890 );
xor ( n20744 , n188019 , n188020 );
buf ( n188022 , n20744 );
buf ( n188023 , n188022 );
not ( n20747 , n188023 );
buf ( n188025 , n20437 );
not ( n20749 , n188025 );
or ( n20750 , n20747 , n20749 );
buf ( n188028 , n20432 );
buf ( n188029 , n20436 );
nand ( n20753 , n188028 , n188029 );
buf ( n188031 , n20753 );
buf ( n188032 , n188031 );
nand ( n20756 , n20750 , n188032 );
buf ( n188034 , n20756 );
buf ( n188035 , n188034 );
not ( n20759 , n188035 );
buf ( n188037 , n20759 );
nand ( n20761 , n20741 , n188037 );
not ( n20762 , n20761 );
buf ( n188040 , n852 );
buf ( n188041 , n874 );
xor ( n20765 , n188040 , n188041 );
buf ( n188043 , n20765 );
buf ( n188044 , n188043 );
not ( n20768 , n188044 );
and ( n20769 , n18991 , n186277 , n187858 );
buf ( n188047 , n20769 );
not ( n20771 , n188047 );
or ( n20772 , n20768 , n20771 );
buf ( n188050 , n18999 );
buf ( n188051 , n187851 );
nand ( n20775 , n188050 , n188051 );
buf ( n188053 , n20775 );
buf ( n188054 , n188053 );
nand ( n20778 , n20772 , n188054 );
buf ( n188056 , n20778 );
not ( n20780 , n188056 );
or ( n20781 , n20762 , n20780 );
buf ( n188059 , n188034 );
buf ( n188060 , n188017 );
nand ( n20784 , n188059 , n188060 );
buf ( n188062 , n20784 );
nand ( n20786 , n20781 , n188062 );
not ( n20787 , n20786 );
or ( n20788 , n20718 , n20787 );
not ( n20789 , n187991 );
buf ( n188067 , n20786 );
not ( n20791 , n188067 );
buf ( n188069 , n20791 );
not ( n20793 , n188069 );
or ( n20794 , n20789 , n20793 );
not ( n20795 , n20234 );
not ( n20796 , n19609 );
nor ( n20797 , n20796 , n19942 );
not ( n20798 , n20797 );
or ( n20799 , n20795 , n20798 );
not ( n20800 , n19602 );
buf ( n188078 , n20800 );
buf ( n188079 , n842 );
buf ( n188080 , n882 );
xor ( n20804 , n188079 , n188080 );
buf ( n188082 , n20804 );
buf ( n188083 , n188082 );
nand ( n20807 , n188078 , n188083 );
buf ( n188085 , n20807 );
nand ( n20809 , n20799 , n188085 );
not ( n20810 , n186191 );
nor ( n20811 , n20810 , n18890 );
not ( n20812 , n20811 );
buf ( n188090 , n857 );
buf ( n188091 , n868 );
xor ( n20815 , n188090 , n188091 );
buf ( n188093 , n20815 );
not ( n20817 , n188093 );
or ( n20818 , n20812 , n20817 );
not ( n20819 , n18906 );
buf ( n188097 , n20819 );
buf ( n188098 , n856 );
buf ( n188099 , n868 );
xor ( n20823 , n188098 , n188099 );
buf ( n188101 , n20823 );
buf ( n188102 , n188101 );
nand ( n20826 , n188097 , n188102 );
buf ( n188104 , n20826 );
nand ( n20828 , n20818 , n188104 );
xor ( n20829 , n20809 , n20828 );
buf ( n188107 , n186441 );
buf ( n188108 , n854 );
buf ( n188109 , n870 );
xor ( n20833 , n188108 , n188109 );
buf ( n188111 , n20833 );
buf ( n188112 , n188111 );
nand ( n20836 , n188107 , n188112 );
buf ( n188114 , n20836 );
nor ( n20838 , n20259 , n19140 );
nand ( n20839 , n187541 , n20838 );
nand ( n20840 , n188114 , n20839 );
xor ( n20841 , n20829 , n20840 );
nand ( n20842 , n20794 , n20841 );
nand ( n20843 , n20788 , n20842 );
buf ( n188121 , n20843 );
not ( n20845 , n188121 );
or ( n20846 , n20708 , n20845 );
or ( n20847 , n20843 , n187982 );
xor ( n20848 , n187794 , n187810 );
xor ( n20849 , n20848 , n187822 );
xor ( n20850 , n187751 , n187725 );
and ( n20851 , n20850 , n187769 );
not ( n20852 , n20850 );
not ( n20853 , n187769 );
and ( n20854 , n20852 , n20853 );
nor ( n20855 , n20851 , n20854 );
buf ( n20856 , n20855 );
or ( n20857 , n20849 , n20856 );
xor ( n20858 , n187873 , n20611 );
xnor ( n20859 , n20858 , n187846 );
nand ( n20860 , n20857 , n20859 );
nand ( n20861 , n20849 , n20856 );
nand ( n20862 , n20860 , n20861 );
nand ( n20863 , n20847 , n20862 );
buf ( n188141 , n20863 );
nand ( n20865 , n20846 , n188141 );
buf ( n188143 , n20865 );
buf ( n188144 , n188143 );
xor ( n20868 , n187903 , n188144 );
buf ( n188146 , n20868 );
buf ( n188147 , n188146 );
buf ( n188148 , n861 );
buf ( n188149 , n864 );
and ( n20873 , n188148 , n188149 );
buf ( n188151 , n20873 );
buf ( n188152 , n187840 );
not ( n20876 , n188152 );
and ( n20877 , n20294 , n20295 );
buf ( n188155 , n20877 );
not ( n20879 , n188155 );
or ( n20880 , n20876 , n20879 );
buf ( n188158 , n20288 );
buf ( n188159 , n837 );
buf ( n188160 , n886 );
xor ( n20884 , n188159 , n188160 );
buf ( n188162 , n20884 );
buf ( n188163 , n188162 );
nand ( n20887 , n188158 , n188163 );
buf ( n188165 , n20887 );
buf ( n188166 , n188165 );
nand ( n20890 , n20880 , n188166 );
buf ( n188168 , n20890 );
xor ( n20892 , n188151 , n188168 );
buf ( n188170 , n20441 );
not ( n20894 , n188170 );
buf ( n188172 , n20437 );
not ( n20896 , n188172 );
or ( n20897 , n20894 , n20896 );
buf ( n188175 , n833 );
buf ( n188176 , n890 );
xor ( n20900 , n188175 , n188176 );
buf ( n188178 , n20900 );
buf ( n20902 , n20436 );
nand ( n20903 , n188178 , n20902 );
buf ( n188181 , n20903 );
nand ( n20905 , n20897 , n188181 );
buf ( n188183 , n20905 );
xor ( n20907 , n20892 , n188183 );
buf ( n188185 , n20907 );
not ( n20909 , n188185 );
not ( n20910 , n187804 );
not ( n20911 , n20390 );
or ( n20912 , n20910 , n20911 );
buf ( n188190 , n20396 );
buf ( n188191 , n835 );
buf ( n188192 , n888 );
xor ( n20916 , n188191 , n188192 );
buf ( n188194 , n20916 );
buf ( n188195 , n188194 );
nand ( n20919 , n188190 , n188195 );
buf ( n188197 , n20919 );
nand ( n20921 , n20912 , n188197 );
not ( n20922 , n20921 );
buf ( n188200 , n20590 );
not ( n20924 , n188200 );
buf ( n188202 , n20769 );
not ( n20926 , n188202 );
or ( n20927 , n20924 , n20926 );
xor ( n20928 , n874 , n849 );
nand ( n20929 , n18999 , n20928 );
buf ( n188207 , n20929 );
nand ( n20931 , n20927 , n188207 );
buf ( n188209 , n20931 );
not ( n20933 , n188209 );
buf ( n188211 , n187763 );
not ( n20935 , n188211 );
buf ( n188213 , n186534 );
buf ( n188214 , n186538 );
and ( n20938 , n188213 , n188214 );
buf ( n188216 , n20938 );
buf ( n188217 , n188216 );
not ( n20941 , n188217 );
or ( n20942 , n20935 , n20941 );
buf ( n188220 , n19264 );
buf ( n188221 , n851 );
buf ( n188222 , n872 );
xor ( n20946 , n188221 , n188222 );
buf ( n188224 , n20946 );
buf ( n188225 , n188224 );
nand ( n20949 , n188220 , n188225 );
buf ( n188227 , n20949 );
buf ( n188228 , n188227 );
nand ( n20952 , n20942 , n188228 );
buf ( n188230 , n20952 );
nand ( n20954 , n20933 , n188230 );
buf ( n188232 , n187763 );
not ( n20956 , n188232 );
buf ( n188234 , n188216 );
not ( n20958 , n188234 );
or ( n20959 , n20956 , n20958 );
buf ( n188237 , n188227 );
nand ( n20961 , n20959 , n188237 );
buf ( n188239 , n20961 );
buf ( n188240 , n188239 );
not ( n20964 , n188240 );
buf ( n188242 , n20964 );
buf ( n188243 , n188242 );
buf ( n188244 , n188209 );
nand ( n20968 , n188243 , n188244 );
buf ( n188246 , n20968 );
nand ( n20970 , n20954 , n188246 );
not ( n20971 , n20970 );
or ( n20972 , n20922 , n20971 );
buf ( n188250 , n20921 );
not ( n20974 , n188250 );
buf ( n188252 , n20974 );
nand ( n20976 , n20954 , n188246 , n188252 );
nand ( n20977 , n20972 , n20976 );
buf ( n188255 , n20977 );
not ( n20979 , n188255 );
buf ( n188257 , n20979 );
buf ( n188258 , n188257 );
not ( n20982 , n188258 );
or ( n20983 , n20909 , n20982 );
buf ( n188261 , n20977 );
not ( n20985 , n188261 );
not ( n20986 , n20907 );
buf ( n188264 , n20986 );
not ( n20988 , n188264 );
or ( n20989 , n20985 , n20988 );
not ( n20990 , n20811 );
not ( n20991 , n188101 );
or ( n20992 , n20990 , n20991 );
buf ( n20993 , n18890 );
xor ( n20994 , n855 , n868 );
nand ( n20995 , n20993 , n20994 );
nand ( n20996 , n20992 , n20995 );
not ( n20997 , n20838 );
not ( n20998 , n188111 );
or ( n20999 , n20997 , n20998 );
buf ( n188277 , n186441 );
buf ( n188278 , n853 );
buf ( n188279 , n870 );
xor ( n21003 , n188278 , n188279 );
buf ( n188281 , n21003 );
buf ( n188282 , n188281 );
nand ( n21006 , n188277 , n188282 );
buf ( n188284 , n21006 );
nand ( n21008 , n20999 , n188284 );
xor ( n21009 , n20996 , n21008 );
not ( n21010 , n188082 );
not ( n21011 , n187507 );
or ( n21012 , n21010 , n21011 );
buf ( n188290 , n19601 );
buf ( n188291 , n841 );
buf ( n188292 , n882 );
xor ( n21016 , n188291 , n188292 );
buf ( n188294 , n21016 );
buf ( n188295 , n188294 );
nand ( n21019 , n188290 , n188295 );
buf ( n188297 , n21019 );
nand ( n21021 , n21012 , n188297 );
xor ( n21022 , n21009 , n21021 );
buf ( n188300 , n21022 );
nand ( n21024 , n20989 , n188300 );
buf ( n188302 , n21024 );
buf ( n188303 , n188302 );
nand ( n21027 , n20983 , n188303 );
buf ( n188305 , n21027 );
not ( n21029 , n188305 );
or ( n21030 , n20809 , n20828 );
nand ( n21031 , n21030 , n20840 );
buf ( n188309 , n20809 );
buf ( n188310 , n20828 );
nand ( n21034 , n188309 , n188310 );
buf ( n188312 , n21034 );
nand ( n21036 , n21031 , n188312 );
not ( n21037 , n21036 );
and ( n21038 , n879 , n878 );
not ( n21039 , n879 );
not ( n21040 , n878 );
and ( n21041 , n21039 , n21040 );
nor ( n21042 , n21038 , n21041 );
not ( n21043 , n21042 );
not ( n21044 , n21043 );
not ( n21045 , n186565 );
nand ( n21046 , n21044 , n21045 );
not ( n21047 , n21046 );
not ( n21048 , n20540 );
and ( n21049 , n21047 , n21048 );
xor ( n21050 , n878 , n845 );
not ( n21051 , n21050 );
nor ( n21052 , n21051 , n21045 );
nor ( n21053 , n21049 , n21052 );
not ( n21054 , n21053 );
not ( n21055 , n21054 );
buf ( n188333 , n20604 );
not ( n21057 , n188333 );
buf ( n188335 , n20276 );
not ( n21059 , n188335 );
or ( n21060 , n21057 , n21059 );
buf ( n188338 , n20279 );
xor ( n21062 , n876 , n847 );
buf ( n188340 , n21062 );
nand ( n21064 , n188338 , n188340 );
buf ( n188342 , n21064 );
buf ( n188343 , n188342 );
nand ( n21067 , n21060 , n188343 );
buf ( n188345 , n21067 );
not ( n21069 , n188345 );
not ( n21070 , n21069 );
or ( n21071 , n21055 , n21070 );
nand ( n21072 , n21053 , n188345 );
nand ( n21073 , n21071 , n21072 );
not ( n21074 , n20468 );
not ( n21075 , n20463 );
or ( n21076 , n21074 , n21075 );
buf ( n188354 , n187733 );
xor ( n21078 , n884 , n839 );
buf ( n188356 , n21078 );
nand ( n21080 , n188354 , n188356 );
buf ( n188358 , n21080 );
nand ( n21082 , n21076 , n188358 );
not ( n21083 , n21082 );
and ( n21084 , n21073 , n21083 );
not ( n21085 , n21073 );
and ( n21086 , n21085 , n21082 );
nor ( n21087 , n21084 , n21086 );
not ( n21088 , n21087 );
not ( n21089 , n21088 );
or ( n21090 , n21037 , n21089 );
buf ( n188368 , n21036 );
not ( n21092 , n188368 );
buf ( n188370 , n21092 );
not ( n21094 , n188370 );
not ( n21095 , n21087 );
or ( n21096 , n21094 , n21095 );
buf ( n188374 , n187421 );
not ( n21098 , n188374 );
buf ( n188376 , n18943 );
not ( n21100 , n188376 );
or ( n21101 , n21098 , n21100 );
buf ( n188379 , n186248 );
buf ( n188380 , n857 );
buf ( n188381 , n866 );
xor ( n21105 , n188380 , n188381 );
buf ( n188383 , n21105 );
buf ( n188384 , n188383 );
nand ( n21108 , n188379 , n188384 );
buf ( n188386 , n21108 );
buf ( n188387 , n188386 );
nand ( n21111 , n21101 , n188387 );
buf ( n188389 , n21111 );
buf ( n188390 , n188389 );
not ( n21114 , n188390 );
and ( n21115 , n20675 , n20682 );
nand ( n21116 , n18874 , n20671 );
xor ( n21117 , n880 , n843 );
and ( n21118 , n21116 , n21117 );
nor ( n21119 , n21115 , n21118 );
buf ( n188397 , n21119 );
not ( n21121 , n188397 );
or ( n21122 , n21114 , n21121 );
buf ( n188400 , n21119 );
buf ( n188401 , n188389 );
or ( n21125 , n188400 , n188401 );
nand ( n21126 , n21122 , n21125 );
buf ( n188404 , n21126 );
buf ( n188405 , n188404 );
buf ( n188406 , n20659 );
not ( n21130 , n188406 );
buf ( n188408 , n19031 );
not ( n21132 , n188408 );
or ( n21133 , n21130 , n21132 );
buf ( n188411 , n186337 );
buf ( n188412 , n859 );
buf ( n188413 , n864 );
xor ( n21137 , n188412 , n188413 );
buf ( n188415 , n21137 );
buf ( n188416 , n188415 );
nand ( n21140 , n188411 , n188416 );
buf ( n188418 , n21140 );
buf ( n188419 , n188418 );
nand ( n21143 , n21133 , n188419 );
buf ( n188421 , n21143 );
buf ( n188422 , n188421 );
not ( n21146 , n188422 );
buf ( n188424 , n21146 );
buf ( n188425 , n188424 );
and ( n21149 , n188405 , n188425 );
not ( n21150 , n188405 );
buf ( n188428 , n188421 );
and ( n21152 , n21150 , n188428 );
nor ( n21153 , n21149 , n21152 );
buf ( n188431 , n21153 );
buf ( n188432 , n188431 );
not ( n21156 , n188432 );
buf ( n188434 , n21156 );
nand ( n21158 , n21096 , n188434 );
nand ( n21159 , n21090 , n21158 );
not ( n21160 , n21159 );
not ( n21161 , n21160 );
and ( n21162 , n21029 , n21161 );
and ( n21163 , n21160 , n188305 );
nor ( n21164 , n21162 , n21163 );
buf ( n188442 , n188242 );
not ( n21166 , n188442 );
buf ( n188444 , n188252 );
not ( n21168 , n188444 );
or ( n21169 , n21166 , n21168 );
buf ( n188447 , n188209 );
nand ( n21171 , n21169 , n188447 );
buf ( n188449 , n21171 );
buf ( n188450 , n188449 );
buf ( n188451 , n20921 );
buf ( n188452 , n188239 );
nand ( n21176 , n188451 , n188452 );
buf ( n188454 , n21176 );
buf ( n188455 , n188454 );
nand ( n21179 , n188450 , n188455 );
buf ( n188457 , n21179 );
not ( n21181 , n21082 );
not ( n21182 , n188345 );
or ( n21183 , n21181 , n21182 );
or ( n21184 , n21082 , n188345 );
nand ( n21185 , n21184 , n21054 );
nand ( n21186 , n21183 , n21185 );
and ( n21187 , n188457 , n21186 );
not ( n21188 , n188457 );
buf ( n188466 , n21186 );
not ( n21190 , n188466 );
buf ( n188468 , n21190 );
and ( n21192 , n21188 , n188468 );
nor ( n21193 , n21187 , n21192 );
or ( n21194 , n20996 , n21021 );
nand ( n21195 , n21194 , n21008 );
nand ( n21196 , n20996 , n21021 );
nand ( n21197 , n21195 , n21196 );
not ( n21198 , n21197 );
and ( n21199 , n21193 , n21198 );
not ( n21200 , n21193 );
and ( n21201 , n21200 , n21197 );
nor ( n21202 , n21199 , n21201 );
buf ( n21203 , n21202 );
and ( n21204 , n21164 , n21203 );
not ( n21205 , n21164 );
buf ( n188483 , n21202 );
not ( n21207 , n188483 );
buf ( n188485 , n21207 );
and ( n21209 , n21205 , n188485 );
nor ( n21210 , n21204 , n21209 );
buf ( n188488 , n21210 );
and ( n21212 , n188147 , n188488 );
not ( n21213 , n188147 );
buf ( n188491 , n21210 );
not ( n21215 , n188491 );
buf ( n188493 , n21215 );
buf ( n188494 , n188493 );
and ( n21218 , n21213 , n188494 );
nor ( n21219 , n21212 , n21218 );
buf ( n188497 , n21219 );
buf ( n188498 , n188497 );
not ( n21222 , n188498 );
buf ( n188500 , n21222 );
buf ( n188501 , n188500 );
not ( n21225 , n188501 );
xor ( n21226 , n20855 , n20849 );
xor ( n21227 , n21226 , n20859 );
not ( n21228 , n21227 );
buf ( n188506 , n188069 );
not ( n21230 , n188506 );
buf ( n188508 , n187994 );
not ( n21232 , n188508 );
or ( n21233 , n21230 , n21232 );
buf ( n188511 , n187991 );
buf ( n188512 , n20786 );
nand ( n21236 , n188511 , n188512 );
buf ( n188514 , n21236 );
buf ( n188515 , n188514 );
nand ( n21239 , n21233 , n188515 );
buf ( n188517 , n21239 );
buf ( n188518 , n188517 );
buf ( n188519 , n20841 );
not ( n21243 , n188519 );
buf ( n188521 , n21243 );
buf ( n188522 , n188521 );
and ( n21246 , n188518 , n188522 );
not ( n21247 , n188518 );
buf ( n188525 , n20841 );
and ( n21249 , n21247 , n188525 );
nor ( n21250 , n21246 , n21249 );
buf ( n188528 , n21250 );
buf ( n188529 , n188528 );
not ( n21253 , n188529 );
buf ( n188531 , n21253 );
not ( n21255 , n188531 );
or ( n21256 , n21228 , n21255 );
nor ( n21257 , n21227 , n188531 );
and ( n21258 , n187681 , n187620 );
not ( n21259 , n187681 );
and ( n21260 , n21259 , n187623 );
nor ( n21261 , n21258 , n21260 );
buf ( n188539 , n21261 );
buf ( n188540 , n187649 );
and ( n21264 , n188539 , n188540 );
not ( n21265 , n188539 );
buf ( n188543 , n187646 );
and ( n21267 , n21265 , n188543 );
or ( n21268 , n21264 , n21267 );
buf ( n188546 , n21268 );
buf ( n188547 , n188546 );
buf ( n188548 , n860 );
buf ( n188549 , n866 );
xor ( n21273 , n188548 , n188549 );
buf ( n188551 , n21273 );
buf ( n188552 , n188551 );
not ( n21276 , n188552 );
buf ( n188554 , n186241 );
not ( n21278 , n188554 );
or ( n21279 , n21276 , n21278 );
buf ( n188557 , n186248 );
buf ( n21281 , n188557 );
buf ( n188559 , n21281 );
buf ( n188560 , n188559 );
buf ( n188561 , n187411 );
nand ( n21285 , n188560 , n188561 );
buf ( n188563 , n21285 );
buf ( n188564 , n188563 );
nand ( n21288 , n21279 , n188564 );
buf ( n188566 , n21288 );
buf ( n188567 , n188566 );
buf ( n188568 , n858 );
buf ( n188569 , n868 );
xor ( n21293 , n188568 , n188569 );
buf ( n188571 , n21293 );
buf ( n188572 , n188571 );
not ( n21296 , n188572 );
buf ( n188574 , n186197 );
not ( n21298 , n188574 );
or ( n21299 , n21296 , n21298 );
buf ( n188577 , n19494 );
buf ( n188578 , n188093 );
nand ( n21302 , n188577 , n188578 );
buf ( n188580 , n21302 );
buf ( n188581 , n188580 );
nand ( n21305 , n21299 , n188581 );
buf ( n188583 , n21305 );
buf ( n188584 , n188583 );
xor ( n21308 , n188567 , n188584 );
buf ( n188586 , n863 );
buf ( n188587 , n865 );
or ( n21311 , n188586 , n188587 );
buf ( n188589 , n866 );
nand ( n21313 , n21311 , n188589 );
buf ( n188591 , n21313 );
buf ( n188592 , n188591 );
buf ( n188593 , n863 );
buf ( n188594 , n865 );
nand ( n21318 , n188593 , n188594 );
buf ( n188596 , n21318 );
buf ( n188597 , n188596 );
buf ( n188598 , n864 );
and ( n21322 , n188592 , n188597 , n188598 );
buf ( n188600 , n21322 );
buf ( n188601 , n188600 );
xor ( n21325 , n894 , n833 );
buf ( n188603 , n21325 );
not ( n21327 , n188603 );
not ( n21328 , n895 );
nand ( n21329 , n21328 , n894 );
not ( n21330 , n21329 );
buf ( n188608 , n21330 );
not ( n21332 , n188608 );
or ( n21333 , n21327 , n21332 );
buf ( n188611 , n20162 );
buf ( n188612 , n895 );
nand ( n21336 , n188611 , n188612 );
buf ( n188614 , n21336 );
buf ( n188615 , n188614 );
nand ( n21339 , n21333 , n188615 );
buf ( n188617 , n21339 );
buf ( n188618 , n188617 );
and ( n21342 , n188601 , n188618 );
buf ( n188620 , n21342 );
buf ( n188621 , n188620 );
xor ( n21345 , n21308 , n188621 );
buf ( n188623 , n21345 );
buf ( n188624 , n188623 );
xor ( n21348 , n188547 , n188624 );
buf ( n188626 , n860 );
buf ( n188627 , n868 );
xor ( n21351 , n188626 , n188627 );
buf ( n188629 , n21351 );
buf ( n188630 , n188629 );
not ( n21354 , n188630 );
buf ( n188632 , n20811 );
not ( n21356 , n188632 );
or ( n21357 , n21354 , n21356 );
buf ( n188635 , n20819 );
buf ( n188636 , n859 );
buf ( n188637 , n868 );
xor ( n21361 , n188636 , n188637 );
buf ( n188639 , n21361 );
buf ( n188640 , n188639 );
nand ( n21364 , n188635 , n188640 );
buf ( n188642 , n21364 );
buf ( n188643 , n188642 );
nand ( n21367 , n21357 , n188643 );
buf ( n188645 , n21367 );
buf ( n188646 , n188645 );
not ( n21370 , n188646 );
buf ( n188648 , n21370 );
buf ( n188649 , n188648 );
not ( n21373 , n188649 );
buf ( n188651 , n846 );
buf ( n188652 , n882 );
xor ( n21376 , n188651 , n188652 );
buf ( n188654 , n21376 );
buf ( n188655 , n188654 );
not ( n21379 , n188655 );
buf ( n188657 , n187507 );
not ( n21381 , n188657 );
or ( n21382 , n21379 , n21381 );
buf ( n188660 , n19942 );
buf ( n188661 , n845 );
buf ( n188662 , n882 );
xor ( n21386 , n188661 , n188662 );
buf ( n188664 , n21386 );
buf ( n188665 , n188664 );
nand ( n21389 , n188660 , n188665 );
buf ( n188667 , n21389 );
buf ( n188668 , n188667 );
nand ( n21392 , n21382 , n188668 );
buf ( n188670 , n21392 );
buf ( n188671 , n188670 );
not ( n21395 , n188671 );
buf ( n188673 , n21395 );
buf ( n188674 , n188673 );
not ( n21398 , n188674 );
or ( n21399 , n21373 , n21398 );
xor ( n21400 , n870 , n858 );
buf ( n188678 , n21400 );
not ( n21402 , n188678 );
buf ( n188680 , n186432 );
not ( n21404 , n188680 );
or ( n21405 , n21402 , n21404 );
buf ( n188683 , n186441 );
buf ( n188684 , n857 );
buf ( n188685 , n870 );
xor ( n21409 , n188684 , n188685 );
buf ( n188687 , n21409 );
buf ( n188688 , n188687 );
nand ( n21412 , n188683 , n188688 );
buf ( n188690 , n21412 );
buf ( n188691 , n188690 );
nand ( n21415 , n21405 , n188691 );
buf ( n188693 , n21415 );
buf ( n188694 , n188693 );
nand ( n21418 , n21399 , n188694 );
buf ( n188696 , n21418 );
buf ( n188697 , n188696 );
buf ( n188698 , n188670 );
buf ( n188699 , n188645 );
nand ( n21423 , n188698 , n188699 );
buf ( n188701 , n21423 );
buf ( n188702 , n188701 );
nand ( n21426 , n188697 , n188702 );
buf ( n188704 , n21426 );
buf ( n188705 , n188704 );
buf ( n188706 , n844 );
buf ( n188707 , n884 );
xor ( n21431 , n188706 , n188707 );
buf ( n188709 , n21431 );
not ( n21433 , n188709 );
not ( n21434 , n20463 );
or ( n21435 , n21433 , n21434 );
buf ( n188713 , n187733 );
buf ( n188714 , n843 );
buf ( n188715 , n884 );
xor ( n21439 , n188714 , n188715 );
buf ( n188717 , n21439 );
buf ( n188718 , n188717 );
nand ( n21442 , n188713 , n188718 );
buf ( n188720 , n21442 );
nand ( n21444 , n21435 , n188720 );
buf ( n188722 , n856 );
buf ( n188723 , n872 );
xor ( n21447 , n188722 , n188723 );
buf ( n188725 , n21447 );
not ( n21449 , n188725 );
not ( n21450 , n20244 );
or ( n21451 , n21449 , n21450 );
buf ( n188729 , n19264 );
buf ( n188730 , n855 );
buf ( n188731 , n872 );
xor ( n21455 , n188730 , n188731 );
buf ( n188733 , n21455 );
buf ( n188734 , n188733 );
nand ( n21458 , n188729 , n188734 );
buf ( n188736 , n21458 );
nand ( n21460 , n21451 , n188736 );
xor ( n21461 , n21444 , n21460 );
buf ( n188739 , n838 );
buf ( n188740 , n890 );
xor ( n21464 , n188739 , n188740 );
buf ( n188742 , n21464 );
not ( n21466 , n188742 );
nor ( n21467 , n890 , n891 );
not ( n21468 , n21467 );
nand ( n21469 , n890 , n891 );
nand ( n21470 , n21468 , n21469 );
nor ( n21471 , n20436 , n21470 );
buf ( n188749 , n21471 );
buf ( n21473 , n188749 );
buf ( n188751 , n21473 );
not ( n21475 , n188751 );
or ( n21476 , n21466 , n21475 );
buf ( n188754 , n20902 );
buf ( n188755 , n837 );
buf ( n188756 , n890 );
xor ( n21480 , n188755 , n188756 );
buf ( n188758 , n21480 );
buf ( n188759 , n188758 );
nand ( n21483 , n188754 , n188759 );
buf ( n188761 , n21483 );
nand ( n21485 , n21476 , n188761 );
and ( n21486 , n21461 , n21485 );
and ( n21487 , n21444 , n21460 );
or ( n21488 , n21486 , n21487 );
buf ( n188766 , n21488 );
or ( n21490 , n188705 , n188766 );
buf ( n188768 , n852 );
buf ( n188769 , n876 );
xor ( n21493 , n188768 , n188769 );
buf ( n188771 , n21493 );
buf ( n188772 , n188771 );
not ( n21496 , n188772 );
buf ( n188774 , n20276 );
not ( n21498 , n188774 );
or ( n21499 , n21496 , n21498 );
buf ( n188777 , n19103 );
buf ( n188778 , n851 );
buf ( n188779 , n876 );
xor ( n21503 , n188778 , n188779 );
buf ( n188781 , n21503 );
buf ( n188782 , n188781 );
nand ( n21506 , n188777 , n188782 );
buf ( n188784 , n21506 );
buf ( n188785 , n188784 );
nand ( n21509 , n21499 , n188785 );
buf ( n188787 , n21509 );
not ( n21511 , n188787 );
not ( n21512 , n20288 );
buf ( n188790 , n841 );
buf ( n188791 , n886 );
xor ( n21515 , n188790 , n188791 );
buf ( n188793 , n21515 );
not ( n21517 , n188793 );
or ( n21518 , n21512 , n21517 );
buf ( n21519 , n20294 );
and ( n21520 , n842 , n886 );
not ( n21521 , n842 );
and ( n21522 , n21521 , n20298 );
nor ( n21523 , n21520 , n21522 );
nand ( n21524 , n20295 , n21519 , n21523 );
nand ( n21525 , n21518 , n21524 );
not ( n21526 , n21525 );
or ( n21527 , n21511 , n21526 );
buf ( n188805 , n188787 );
not ( n21529 , n188805 );
buf ( n188807 , n21529 );
not ( n21531 , n188807 );
not ( n21532 , n21525 );
not ( n21533 , n21532 );
or ( n21534 , n21531 , n21533 );
buf ( n188812 , n854 );
buf ( n188813 , n874 );
xor ( n21537 , n188812 , n188813 );
buf ( n188815 , n21537 );
buf ( n188816 , n188815 );
not ( n21540 , n188816 );
buf ( n188818 , n18992 );
not ( n21542 , n188818 );
or ( n21543 , n21540 , n21542 );
buf ( n188821 , n186294 );
not ( n21545 , n188821 );
buf ( n188823 , n21545 );
buf ( n188824 , n188823 );
buf ( n188825 , n853 );
buf ( n188826 , n874 );
xor ( n21550 , n188825 , n188826 );
buf ( n188828 , n21550 );
buf ( n188829 , n188828 );
nand ( n21553 , n188824 , n188829 );
buf ( n188831 , n21553 );
buf ( n188832 , n188831 );
nand ( n21556 , n21543 , n188832 );
buf ( n188834 , n21556 );
nand ( n21558 , n21534 , n188834 );
nand ( n21559 , n21527 , n21558 );
buf ( n188837 , n21559 );
nand ( n21561 , n21490 , n188837 );
buf ( n188839 , n21561 );
buf ( n188840 , n188839 );
buf ( n188841 , n188704 );
buf ( n188842 , n21488 );
nand ( n21566 , n188841 , n188842 );
buf ( n188844 , n21566 );
buf ( n188845 , n188844 );
nand ( n21569 , n188840 , n188845 );
buf ( n188847 , n21569 );
buf ( n188848 , n188847 );
and ( n21572 , n21348 , n188848 );
and ( n21573 , n188547 , n188624 );
or ( n21574 , n21572 , n21573 );
buf ( n188852 , n21574 );
not ( n21576 , n188852 );
or ( n21577 , n21257 , n21576 );
nand ( n21578 , n21256 , n21577 );
buf ( n188856 , n21578 );
buf ( n188857 , n21022 );
not ( n21581 , n188857 );
buf ( n188859 , n21581 );
buf ( n188860 , n188859 );
not ( n21584 , n188860 );
and ( n21585 , n20977 , n20986 );
not ( n21586 , n20977 );
and ( n21587 , n21586 , n20907 );
nor ( n21588 , n21585 , n21587 );
buf ( n188866 , n21588 );
not ( n21590 , n188866 );
or ( n21591 , n21584 , n21590 );
buf ( n188869 , n21588 );
buf ( n188870 , n188859 );
or ( n21594 , n188869 , n188870 );
nand ( n21595 , n21591 , n21594 );
buf ( n188873 , n21595 );
buf ( n188874 , n188873 );
buf ( n188875 , n21036 );
not ( n21599 , n188875 );
buf ( n188877 , n188431 );
not ( n21601 , n188877 );
or ( n21602 , n21599 , n21601 );
buf ( n188880 , n21036 );
buf ( n188881 , n188431 );
or ( n21605 , n188880 , n188881 );
nand ( n21606 , n21602 , n21605 );
buf ( n188884 , n21606 );
and ( n21608 , n188884 , n21087 );
not ( n21609 , n188884 );
and ( n21610 , n21609 , n21088 );
or ( n21611 , n21608 , n21610 );
buf ( n188889 , n21611 );
xor ( n21613 , n188874 , n188889 );
xor ( n21614 , n187407 , n187428 );
xor ( n21615 , n21614 , n187491 );
buf ( n188893 , n21615 );
buf ( n188894 , n188893 );
xor ( n21618 , n20273 , n187604 );
xor ( n21619 , n21618 , n187692 );
buf ( n188897 , n21619 );
xor ( n21621 , n188894 , n188897 );
xor ( n21622 , n188056 , n188037 );
buf ( n188900 , n188017 );
buf ( n21624 , n188900 );
buf ( n188902 , n21624 );
xor ( n21626 , n21622 , n188902 );
buf ( n188904 , n21626 );
not ( n21628 , n188904 );
buf ( n188906 , n21628 );
not ( n21630 , n188906 );
buf ( n21631 , n20271 );
not ( n21632 , n21631 );
not ( n21633 , n21632 );
not ( n21634 , n20238 );
not ( n21635 , n21634 );
not ( n21636 , n20252 );
not ( n21637 , n21636 );
or ( n21638 , n21635 , n21637 );
or ( n21639 , n21634 , n21636 );
nand ( n21640 , n21638 , n21639 );
not ( n21641 , n21640 );
or ( n21642 , n21633 , n21641 );
or ( n21643 , n21632 , n21640 );
nand ( n21644 , n21642 , n21643 );
buf ( n188922 , n21644 );
not ( n21646 , n188922 );
buf ( n188924 , n21646 );
not ( n21648 , n188924 );
or ( n21649 , n21630 , n21648 );
not ( n21650 , n21644 );
not ( n21651 , n21626 );
or ( n21652 , n21650 , n21651 );
xor ( n21653 , n20302 , n20321 );
xor ( n21654 , n21653 , n20285 );
nand ( n21655 , n21652 , n21654 );
nand ( n21656 , n21649 , n21655 );
buf ( n188934 , n21656 );
and ( n21658 , n21621 , n188934 );
and ( n21659 , n188894 , n188897 );
or ( n21660 , n21658 , n21659 );
buf ( n188938 , n21660 );
buf ( n188939 , n188938 );
xor ( n21663 , n21613 , n188939 );
buf ( n188941 , n21663 );
buf ( n188942 , n188941 );
xor ( n21666 , n188856 , n188942 );
xor ( n21667 , n188567 , n188584 );
and ( n21668 , n21667 , n188621 );
and ( n21669 , n188567 , n188584 );
or ( n21670 , n21668 , n21669 );
buf ( n188948 , n21670 );
xor ( n21672 , n187434 , n187447 );
xor ( n21673 , n21672 , n187486 );
buf ( n188951 , n21673 );
buf ( n188952 , n188951 );
buf ( n188953 , n188639 );
not ( n21677 , n188953 );
buf ( n188955 , n20811 );
not ( n21679 , n188955 );
or ( n21680 , n21677 , n21679 );
buf ( n188958 , n20993 );
buf ( n188959 , n188571 );
nand ( n21683 , n188958 , n188959 );
buf ( n188961 , n21683 );
buf ( n188962 , n188961 );
nand ( n21686 , n21680 , n188962 );
buf ( n188964 , n21686 );
buf ( n188965 , n188964 );
not ( n21689 , n188965 );
buf ( n188967 , n188664 );
not ( n21691 , n188967 );
buf ( n188969 , n187507 );
not ( n21693 , n188969 );
or ( n21694 , n21691 , n21693 );
buf ( n188972 , n20221 );
buf ( n188973 , n19601 );
nand ( n21697 , n188972 , n188973 );
buf ( n188975 , n21697 );
buf ( n188976 , n188975 );
nand ( n21700 , n21694 , n188976 );
buf ( n188978 , n21700 );
buf ( n188979 , n188978 );
not ( n21703 , n188979 );
or ( n21704 , n21689 , n21703 );
buf ( n188982 , n188964 );
not ( n21706 , n188982 );
buf ( n188984 , n21706 );
buf ( n188985 , n188984 );
not ( n21709 , n188985 );
not ( n21710 , n188978 );
buf ( n188988 , n21710 );
not ( n21712 , n188988 );
or ( n21713 , n21709 , n21712 );
buf ( n188991 , n861 );
buf ( n188992 , n866 );
xor ( n21716 , n188991 , n188992 );
buf ( n188994 , n21716 );
buf ( n188995 , n188994 );
not ( n21719 , n188995 );
buf ( n188997 , n186241 );
not ( n21721 , n188997 );
or ( n21722 , n21719 , n21721 );
buf ( n189000 , n188559 );
buf ( n189001 , n188551 );
nand ( n21725 , n189000 , n189001 );
buf ( n189003 , n21725 );
buf ( n189004 , n189003 );
nand ( n21728 , n21722 , n189004 );
buf ( n189006 , n21728 );
buf ( n189007 , n189006 );
nand ( n21731 , n21713 , n189007 );
buf ( n189009 , n21731 );
buf ( n189010 , n189009 );
nand ( n21734 , n21704 , n189010 );
buf ( n189012 , n21734 );
buf ( n189013 , n189012 );
xor ( n21737 , n188952 , n189013 );
not ( n21738 , n188733 );
not ( n21739 , n20244 );
or ( n21740 , n21738 , n21739 );
buf ( n189018 , n19264 );
buf ( n189019 , n20240 );
nand ( n21743 , n189018 , n189019 );
buf ( n189021 , n21743 );
nand ( n21745 , n21740 , n189021 );
not ( n21746 , n188717 );
not ( n21747 , n20727 );
or ( n21748 , n21746 , n21747 );
buf ( n189026 , n188010 );
buf ( n189027 , n187999 );
nand ( n21751 , n189026 , n189027 );
buf ( n189029 , n21751 );
nand ( n21753 , n21748 , n189029 );
nor ( n21754 , n21745 , n21753 );
buf ( n189032 , n19138 );
not ( n21756 , n189032 );
buf ( n189034 , n21756 );
buf ( n189035 , n189034 );
not ( n21759 , n189035 );
buf ( n189037 , n21759 );
buf ( n189038 , n189037 );
buf ( n189039 , n20269 );
nand ( n21763 , n189038 , n189039 );
buf ( n189041 , n21763 );
nand ( n21765 , n186432 , n188687 );
and ( n21766 , n189041 , n21765 );
or ( n21767 , n21754 , n21766 );
nand ( n21768 , n21745 , n21753 );
nand ( n21769 , n21767 , n21768 );
buf ( n189047 , n21769 );
and ( n21771 , n21737 , n189047 );
and ( n21772 , n188952 , n189013 );
or ( n21773 , n21771 , n21772 );
buf ( n189051 , n21773 );
xor ( n21775 , n188948 , n189051 );
buf ( n189053 , n839 );
buf ( n189054 , n888 );
xor ( n21778 , n189053 , n189054 );
buf ( n189056 , n21778 );
not ( n21780 , n189056 );
not ( n21781 , n20390 );
or ( n21782 , n21780 , n21781 );
buf ( n189060 , n20396 );
buf ( n189061 , n187656 );
nand ( n21785 , n189060 , n189061 );
buf ( n189063 , n21785 );
nand ( n21787 , n21782 , n189063 );
not ( n21788 , n21787 );
not ( n21789 , n21788 );
buf ( n189067 , n835 );
buf ( n189068 , n892 );
xor ( n21792 , n189067 , n189068 );
buf ( n189070 , n21792 );
not ( n21794 , n189070 );
nand ( n21795 , n20197 , n20188 );
not ( n21796 , n21795 );
not ( n21797 , n21796 );
or ( n21798 , n21794 , n21797 );
buf ( n189076 , n187477 );
buf ( n189077 , n187452 );
nand ( n21801 , n189076 , n189077 );
buf ( n189079 , n21801 );
nand ( n21803 , n21798 , n189079 );
not ( n21804 , n21803 );
not ( n21805 , n21804 );
or ( n21806 , n21789 , n21805 );
buf ( n189084 , n863 );
buf ( n189085 , n864 );
xor ( n21809 , n189084 , n189085 );
buf ( n189087 , n21809 );
buf ( n189088 , n189087 );
not ( n21812 , n189088 );
buf ( n189090 , n19031 );
not ( n21814 , n189090 );
or ( n21815 , n21812 , n21814 );
buf ( n189093 , n186340 );
buf ( n189094 , n187609 );
nand ( n21818 , n189093 , n189094 );
buf ( n189096 , n21818 );
buf ( n189097 , n189096 );
nand ( n21821 , n21815 , n189097 );
buf ( n189099 , n21821 );
nand ( n21823 , n21806 , n189099 );
buf ( n189101 , n21823 );
nand ( n21825 , n21787 , n21803 );
buf ( n189103 , n21825 );
nand ( n21827 , n189101 , n189103 );
buf ( n189105 , n21827 );
buf ( n189106 , n189105 );
buf ( n189107 , n847 );
buf ( n189108 , n880 );
xor ( n21832 , n189107 , n189108 );
buf ( n189110 , n21832 );
buf ( n189111 , n189110 );
not ( n21835 , n189111 );
buf ( n189113 , n20675 );
not ( n21837 , n189113 );
or ( n21838 , n21835 , n21837 );
buf ( n189116 , n20358 );
buf ( n189117 , n187629 );
nand ( n21841 , n189116 , n189117 );
buf ( n189119 , n21841 );
buf ( n189120 , n189119 );
nand ( n21844 , n21838 , n189120 );
buf ( n189122 , n21844 );
buf ( n189123 , n189122 );
not ( n21847 , n189123 );
buf ( n189125 , n188793 );
not ( n21849 , n189125 );
and ( n21850 , n20294 , n20295 );
buf ( n189128 , n21850 );
not ( n21852 , n189128 );
or ( n21853 , n21849 , n21852 );
buf ( n189131 , n20558 );
buf ( n189132 , n20300 );
nand ( n21856 , n189131 , n189132 );
buf ( n189134 , n21856 );
buf ( n189135 , n189134 );
nand ( n21859 , n21853 , n189135 );
buf ( n189137 , n21859 );
buf ( n189138 , n189137 );
not ( n21862 , n189138 );
or ( n21863 , n21847 , n21862 );
buf ( n189141 , n189122 );
buf ( n189142 , n189137 );
or ( n21866 , n189141 , n189142 );
buf ( n189144 , n849 );
buf ( n189145 , n878 );
xor ( n21869 , n189144 , n189145 );
buf ( n189147 , n21869 );
buf ( n189148 , n189147 );
not ( n21872 , n189148 );
buf ( n189150 , n186569 );
not ( n21874 , n189150 );
or ( n21875 , n21872 , n21874 );
buf ( n189153 , n186575 );
buf ( n189154 , n187596 );
nand ( n21878 , n189153 , n189154 );
buf ( n189156 , n21878 );
buf ( n189157 , n189156 );
nand ( n21881 , n21875 , n189157 );
buf ( n189159 , n21881 );
buf ( n189160 , n189159 );
nand ( n21884 , n21866 , n189160 );
buf ( n189162 , n21884 );
buf ( n189163 , n189162 );
nand ( n21887 , n21863 , n189163 );
buf ( n189165 , n21887 );
buf ( n189166 , n189165 );
or ( n21890 , n189106 , n189166 );
buf ( n189168 , n188758 );
not ( n21892 , n189168 );
buf ( n189170 , n188751 );
not ( n21894 , n189170 );
or ( n21895 , n21892 , n21894 );
buf ( n189173 , n20902 );
buf ( n189174 , n188022 );
nand ( n21898 , n189173 , n189174 );
buf ( n189176 , n21898 );
buf ( n189177 , n189176 );
nand ( n21901 , n21895 , n189177 );
buf ( n189179 , n21901 );
buf ( n189180 , n189179 );
not ( n21904 , n189180 );
buf ( n189182 , n188781 );
not ( n21906 , n189182 );
buf ( n189184 , n19177 );
not ( n21908 , n189184 );
or ( n21909 , n21906 , n21908 );
buf ( n189187 , n20279 );
buf ( n189188 , n20274 );
nand ( n21912 , n189187 , n189188 );
buf ( n189190 , n21912 );
buf ( n189191 , n189190 );
nand ( n21915 , n21909 , n189191 );
buf ( n189193 , n21915 );
buf ( n189194 , n189193 );
not ( n21918 , n189194 );
or ( n21919 , n21904 , n21918 );
or ( n21920 , n189179 , n189193 );
buf ( n189198 , n188828 );
not ( n21922 , n189198 );
buf ( n189200 , n20582 );
not ( n21924 , n189200 );
or ( n21925 , n21922 , n21924 );
buf ( n189203 , n187865 );
buf ( n189204 , n188043 );
nand ( n21928 , n189203 , n189204 );
buf ( n189206 , n21928 );
buf ( n189207 , n189206 );
nand ( n21931 , n21925 , n189207 );
buf ( n189209 , n21931 );
nand ( n21933 , n21920 , n189209 );
buf ( n189211 , n21933 );
nand ( n21935 , n21919 , n189211 );
buf ( n189213 , n21935 );
buf ( n189214 , n189213 );
nand ( n21938 , n21890 , n189214 );
buf ( n189216 , n21938 );
buf ( n189217 , n189216 );
buf ( n189218 , n189105 );
buf ( n189219 , n189165 );
nand ( n21943 , n189218 , n189219 );
buf ( n189221 , n21943 );
buf ( n189222 , n189221 );
nand ( n21946 , n189217 , n189222 );
buf ( n189224 , n21946 );
xor ( n21948 , n21775 , n189224 );
buf ( n189226 , n21948 );
xor ( n21950 , n188601 , n188618 );
buf ( n189228 , n21950 );
buf ( n189229 , n189228 );
not ( n21953 , n21325 );
not ( n21954 , n895 );
or ( n21955 , n21953 , n21954 );
buf ( n189233 , n895 );
not ( n21957 , n189233 );
buf ( n189235 , n894 );
nand ( n21959 , n21957 , n189235 );
buf ( n189237 , n21959 );
buf ( n189238 , n834 );
buf ( n189239 , n894 );
xor ( n21963 , n189238 , n189239 );
buf ( n189241 , n21963 );
buf ( n189242 , n189241 );
not ( n21966 , n189242 );
buf ( n189244 , n21966 );
or ( n21968 , n189237 , n189244 );
nand ( n21969 , n21955 , n21968 );
buf ( n189247 , n21969 );
buf ( n189248 , n186337 );
buf ( n189249 , n863 );
and ( n21973 , n189248 , n189249 );
buf ( n189251 , n21973 );
buf ( n189252 , n189251 );
xor ( n21976 , n189247 , n189252 );
buf ( n189254 , n836 );
buf ( n189255 , n892 );
xor ( n21979 , n189254 , n189255 );
buf ( n189257 , n21979 );
buf ( n189258 , n189257 );
not ( n21982 , n189258 );
buf ( n189260 , n187469 );
not ( n21984 , n189260 );
or ( n21985 , n21982 , n21984 );
buf ( n189263 , n187477 );
buf ( n189264 , n189070 );
nand ( n21988 , n189263 , n189264 );
buf ( n189266 , n21988 );
buf ( n189267 , n189266 );
nand ( n21991 , n21985 , n189267 );
buf ( n189269 , n21991 );
buf ( n189270 , n189269 );
and ( n21994 , n21976 , n189270 );
and ( n21995 , n189247 , n189252 );
or ( n21996 , n21994 , n21995 );
buf ( n189274 , n21996 );
buf ( n189275 , n189274 );
xor ( n21999 , n189229 , n189275 );
buf ( n189277 , n840 );
buf ( n189278 , n888 );
xor ( n22002 , n189277 , n189278 );
buf ( n189280 , n22002 );
buf ( n189281 , n189280 );
not ( n22005 , n189281 );
buf ( n189283 , n20391 );
not ( n22007 , n189283 );
or ( n22008 , n22005 , n22007 );
buf ( n22009 , n20395 );
buf ( n189287 , n22009 );
buf ( n189288 , n189056 );
nand ( n22012 , n189287 , n189288 );
buf ( n189290 , n22012 );
buf ( n189291 , n189290 );
nand ( n22015 , n22008 , n189291 );
buf ( n189293 , n22015 );
buf ( n189294 , n189293 );
not ( n22018 , n189294 );
and ( n22019 , n848 , n880 );
not ( n22020 , n848 );
and ( n22021 , n22020 , n18856 );
nor ( n22022 , n22019 , n22021 );
buf ( n189300 , n22022 );
not ( n22024 , n189300 );
buf ( n189302 , n18862 );
not ( n22026 , n189302 );
or ( n22027 , n22024 , n22026 );
buf ( n189305 , n20358 );
buf ( n189306 , n189110 );
nand ( n22030 , n189305 , n189306 );
buf ( n189308 , n22030 );
buf ( n189309 , n189308 );
nand ( n22033 , n22027 , n189309 );
buf ( n189311 , n22033 );
buf ( n189312 , n189311 );
not ( n22036 , n189312 );
or ( n22037 , n22018 , n22036 );
buf ( n189315 , n189311 );
not ( n22039 , n189315 );
buf ( n189317 , n22039 );
buf ( n189318 , n189317 );
not ( n22042 , n189318 );
buf ( n189320 , n189293 );
not ( n22044 , n189320 );
buf ( n189322 , n22044 );
buf ( n189323 , n189322 );
not ( n22047 , n189323 );
or ( n22048 , n22042 , n22047 );
buf ( n189326 , n850 );
buf ( n189327 , n878 );
xor ( n22051 , n189326 , n189327 );
buf ( n189329 , n22051 );
buf ( n189330 , n189329 );
not ( n22054 , n189330 );
buf ( n189332 , n186569 );
not ( n22056 , n189332 );
or ( n22057 , n22054 , n22056 );
buf ( n189335 , n186575 );
buf ( n189336 , n189147 );
nand ( n22060 , n189335 , n189336 );
buf ( n189338 , n22060 );
buf ( n189339 , n189338 );
nand ( n22063 , n22057 , n189339 );
buf ( n189341 , n22063 );
buf ( n189342 , n189341 );
nand ( n22066 , n22048 , n189342 );
buf ( n189344 , n22066 );
buf ( n189345 , n189344 );
nand ( n22069 , n22037 , n189345 );
buf ( n189347 , n22069 );
buf ( n189348 , n189347 );
and ( n22072 , n21999 , n189348 );
and ( n22073 , n189229 , n189275 );
or ( n22074 , n22072 , n22073 );
buf ( n189352 , n22074 );
not ( n22076 , n189352 );
xor ( n22077 , n188952 , n189013 );
xor ( n22078 , n22077 , n189047 );
buf ( n189356 , n22078 );
not ( n22080 , n189356 );
not ( n22081 , n22080 );
not ( n22082 , n22081 );
or ( n22083 , n22076 , n22082 );
not ( n22084 , n189352 );
not ( n22085 , n22084 );
not ( n22086 , n22080 );
or ( n22087 , n22085 , n22086 );
not ( n22088 , n189099 );
and ( n22089 , n21803 , n21787 );
not ( n22090 , n21803 );
and ( n22091 , n22090 , n21788 );
nor ( n22092 , n22089 , n22091 );
not ( n22093 , n22092 );
or ( n22094 , n22088 , n22093 );
or ( n22095 , n189099 , n22092 );
nand ( n22096 , n22094 , n22095 );
buf ( n189374 , n22096 );
not ( n22098 , n189374 );
not ( n22099 , n188978 );
not ( n22100 , n188964 );
or ( n22101 , n22099 , n22100 );
nand ( n22102 , n188984 , n21710 );
nand ( n22103 , n22101 , n22102 );
not ( n22104 , n189006 );
and ( n22105 , n22103 , n22104 );
not ( n22106 , n22103 );
and ( n22107 , n22106 , n189006 );
nor ( n22108 , n22105 , n22107 );
not ( n22109 , n22108 );
buf ( n189387 , n22109 );
not ( n22111 , n189387 );
or ( n22112 , n22098 , n22111 );
xor ( n22113 , n189159 , n189137 );
xor ( n22114 , n22113 , n189122 );
buf ( n189392 , n22114 );
nand ( n22116 , n22112 , n189392 );
buf ( n189394 , n22116 );
buf ( n189395 , n189394 );
buf ( n189396 , n22096 );
not ( n22120 , n189396 );
not ( n22121 , n22109 );
buf ( n189399 , n22121 );
nand ( n22123 , n22120 , n189399 );
buf ( n189401 , n22123 );
buf ( n189402 , n189401 );
nand ( n22126 , n189395 , n189402 );
buf ( n189404 , n22126 );
nand ( n22128 , n22087 , n189404 );
nand ( n22129 , n22083 , n22128 );
buf ( n189407 , n22129 );
or ( n22131 , n189226 , n189407 );
xor ( n22132 , n188894 , n188897 );
xor ( n22133 , n22132 , n188934 );
buf ( n189411 , n22133 );
buf ( n189412 , n189411 );
nand ( n22136 , n22131 , n189412 );
buf ( n189414 , n22136 );
buf ( n189415 , n189414 );
buf ( n189416 , n22129 );
buf ( n189417 , n21948 );
nand ( n22141 , n189416 , n189417 );
buf ( n189419 , n22141 );
buf ( n189420 , n189419 );
nand ( n22144 , n189415 , n189420 );
buf ( n189422 , n22144 );
buf ( n189423 , n189422 );
and ( n22147 , n21666 , n189423 );
and ( n22148 , n188856 , n188942 );
or ( n22149 , n22147 , n22148 );
buf ( n189427 , n22149 );
buf ( n189428 , n189427 );
not ( n22152 , n189428 );
buf ( n189430 , n22152 );
buf ( n189431 , n189430 );
not ( n22155 , n189431 );
or ( n22156 , n21225 , n22155 );
xor ( n22157 , n188874 , n188889 );
and ( n22158 , n22157 , n188939 );
and ( n22159 , n188874 , n188889 );
or ( n22160 , n22158 , n22159 );
buf ( n189438 , n22160 );
buf ( n189439 , n189438 );
buf ( n189440 , n860 );
buf ( n189441 , n864 );
and ( n22165 , n189440 , n189441 );
buf ( n189443 , n22165 );
buf ( n189444 , n189443 );
buf ( n189445 , n21062 );
not ( n22169 , n189445 );
buf ( n189447 , n20276 );
not ( n22171 , n189447 );
or ( n22172 , n22169 , n22171 );
buf ( n189450 , n20279 );
xor ( n22174 , n876 , n846 );
buf ( n189452 , n22174 );
nand ( n22176 , n189450 , n189452 );
buf ( n189454 , n22176 );
buf ( n189455 , n189454 );
nand ( n22179 , n22172 , n189455 );
buf ( n189457 , n22179 );
buf ( n189458 , n189457 );
xor ( n22182 , n189444 , n189458 );
not ( n22183 , n21050 );
not ( n22184 , n21046 );
not ( n22185 , n22184 );
or ( n22186 , n22183 , n22185 );
buf ( n189464 , n186575 );
buf ( n189465 , n844 );
buf ( n189466 , n878 );
xor ( n22190 , n189465 , n189466 );
buf ( n189468 , n22190 );
buf ( n189469 , n189468 );
nand ( n22193 , n189464 , n189469 );
buf ( n189471 , n22193 );
nand ( n22195 , n22186 , n189471 );
buf ( n189473 , n22195 );
xor ( n22197 , n22182 , n189473 );
buf ( n189475 , n22197 );
buf ( n189476 , n189475 );
buf ( n189477 , n20197 );
not ( n22201 , n189477 );
buf ( n189479 , n21795 );
not ( n22203 , n189479 );
or ( n22204 , n22201 , n22203 );
buf ( n189482 , n892 );
nand ( n22206 , n22204 , n189482 );
buf ( n189484 , n22206 );
buf ( n189485 , n189484 );
buf ( n189486 , n188162 );
not ( n22210 , n189486 );
buf ( n189488 , n21850 );
not ( n22212 , n189488 );
or ( n22213 , n22210 , n22212 );
buf ( n189491 , n20288 );
buf ( n189492 , n836 );
buf ( n189493 , n886 );
xor ( n22217 , n189492 , n189493 );
buf ( n189495 , n22217 );
buf ( n189496 , n189495 );
nand ( n22220 , n189491 , n189496 );
buf ( n189498 , n22220 );
buf ( n189499 , n189498 );
nand ( n22223 , n22213 , n189499 );
buf ( n189501 , n22223 );
buf ( n189502 , n189501 );
xor ( n22226 , n189485 , n189502 );
buf ( n189504 , n188178 );
not ( n22228 , n189504 );
buf ( n189506 , n188751 );
not ( n22230 , n189506 );
or ( n22231 , n22228 , n22230 );
buf ( n189509 , n20902 );
buf ( n189510 , n832 );
buf ( n189511 , n890 );
xor ( n22235 , n189510 , n189511 );
buf ( n189513 , n22235 );
buf ( n189514 , n189513 );
nand ( n22238 , n189509 , n189514 );
buf ( n189516 , n22238 );
buf ( n189517 , n189516 );
nand ( n22241 , n22231 , n189517 );
buf ( n189519 , n22241 );
buf ( n189520 , n189519 );
xor ( n22244 , n22226 , n189520 );
buf ( n189522 , n22244 );
buf ( n189523 , n189522 );
xor ( n22247 , n189476 , n189523 );
buf ( n22248 , n21119 );
buf ( n189526 , n22248 );
not ( n22250 , n189526 );
buf ( n189528 , n188424 );
not ( n22252 , n189528 );
or ( n22253 , n22250 , n22252 );
buf ( n189531 , n188389 );
nand ( n22255 , n22253 , n189531 );
buf ( n189533 , n22255 );
buf ( n189534 , n189533 );
not ( n22258 , n22248 );
nand ( n22259 , n22258 , n188421 );
buf ( n189537 , n22259 );
nand ( n22261 , n189534 , n189537 );
buf ( n189539 , n22261 );
buf ( n189540 , n189539 );
xor ( n22264 , n22247 , n189540 );
buf ( n189542 , n22264 );
buf ( n189543 , n189542 );
buf ( n189544 , n188383 );
not ( n22268 , n189544 );
buf ( n189546 , n18938 );
buf ( n189547 , n186237 );
nor ( n22271 , n189546 , n189547 );
buf ( n189549 , n22271 );
buf ( n189550 , n189549 );
not ( n22274 , n189550 );
or ( n22275 , n22268 , n22274 );
buf ( n189553 , n186248 );
buf ( n189554 , n856 );
buf ( n189555 , n866 );
xor ( n22279 , n189554 , n189555 );
buf ( n189557 , n22279 );
buf ( n189558 , n189557 );
nand ( n22282 , n189553 , n189558 );
buf ( n189560 , n22282 );
buf ( n189561 , n189560 );
nand ( n22285 , n22275 , n189561 );
buf ( n189563 , n22285 );
buf ( n189564 , n189563 );
not ( n22288 , n20994 );
not ( n22289 , n186194 );
or ( n22290 , n22288 , n22289 );
buf ( n189568 , n20819 );
xor ( n22292 , n868 , n854 );
buf ( n189570 , n22292 );
nand ( n22294 , n189568 , n189570 );
buf ( n189572 , n22294 );
nand ( n22296 , n22290 , n189572 );
buf ( n189574 , n22296 );
xor ( n22298 , n189564 , n189574 );
buf ( n189576 , n21117 );
not ( n22300 , n189576 );
buf ( n189578 , n18862 );
not ( n22302 , n189578 );
or ( n22303 , n22300 , n22302 );
buf ( n22304 , n21116 );
buf ( n189582 , n22304 );
xor ( n22306 , n880 , n842 );
buf ( n189584 , n22306 );
nand ( n22308 , n189582 , n189584 );
buf ( n189586 , n22308 );
buf ( n189587 , n189586 );
nand ( n22311 , n22303 , n189587 );
buf ( n189589 , n22311 );
buf ( n189590 , n189589 );
xor ( n22314 , n22298 , n189590 );
buf ( n189592 , n22314 );
buf ( n189593 , n189592 );
not ( n22317 , n189593 );
not ( n22318 , n188294 );
not ( n22319 , n187507 );
or ( n22320 , n22318 , n22319 );
buf ( n189598 , n19601 );
buf ( n189599 , n840 );
buf ( n189600 , n882 );
xor ( n22324 , n189599 , n189600 );
buf ( n189602 , n22324 );
buf ( n189603 , n189602 );
nand ( n22327 , n189598 , n189603 );
buf ( n189605 , n22327 );
nand ( n22329 , n22320 , n189605 );
not ( n22330 , n188194 );
not ( n22331 , n20382 );
nand ( n22332 , n889 , n890 );
not ( n22333 , n22332 );
not ( n22334 , n22333 );
or ( n22335 , n22331 , n22334 );
nand ( n22336 , n22335 , n20389 );
not ( n22337 , n22336 );
or ( n22338 , n22330 , n22337 );
buf ( n189616 , n20396 );
buf ( n189617 , n834 );
buf ( n189618 , n888 );
xor ( n22342 , n189617 , n189618 );
buf ( n189620 , n22342 );
buf ( n189621 , n189620 );
nand ( n22345 , n189616 , n189621 );
buf ( n189623 , n22345 );
nand ( n22347 , n22338 , n189623 );
not ( n22348 , n22347 );
xor ( n22349 , n22329 , n22348 );
buf ( n189627 , n188281 );
not ( n22351 , n189627 );
buf ( n189629 , n186432 );
not ( n22353 , n189629 );
or ( n22354 , n22351 , n22353 );
buf ( n189632 , n186441 );
xor ( n22356 , n870 , n852 );
buf ( n189634 , n22356 );
nand ( n22358 , n189632 , n189634 );
buf ( n189636 , n22358 );
buf ( n189637 , n189636 );
nand ( n22361 , n22354 , n189637 );
buf ( n189639 , n22361 );
xor ( n22363 , n22349 , n189639 );
buf ( n189641 , n22363 );
not ( n22365 , n189641 );
and ( n22366 , n22317 , n22365 );
buf ( n189644 , n189592 );
buf ( n189645 , n22363 );
and ( n22369 , n189644 , n189645 );
nor ( n22370 , n22366 , n22369 );
buf ( n189648 , n22370 );
buf ( n189649 , n189648 );
not ( n22373 , n20928 );
not ( n22374 , n20769 );
or ( n22375 , n22373 , n22374 );
buf ( n189653 , n18999 );
buf ( n189654 , n848 );
buf ( n189655 , n874 );
xor ( n22379 , n189654 , n189655 );
buf ( n189657 , n22379 );
buf ( n189658 , n189657 );
nand ( n22382 , n189653 , n189658 );
buf ( n189660 , n22382 );
nand ( n22384 , n22375 , n189660 );
buf ( n189662 , n22384 );
not ( n22386 , n189662 );
buf ( n189664 , n21078 );
not ( n22388 , n189664 );
buf ( n189666 , n20463 );
not ( n22390 , n189666 );
or ( n22391 , n22388 , n22390 );
buf ( n189669 , n188010 );
buf ( n189670 , n838 );
buf ( n189671 , n884 );
xor ( n22395 , n189670 , n189671 );
buf ( n189673 , n22395 );
buf ( n189674 , n189673 );
nand ( n22398 , n189669 , n189674 );
buf ( n189676 , n22398 );
buf ( n189677 , n189676 );
nand ( n22401 , n22391 , n189677 );
buf ( n189679 , n22401 );
buf ( n189680 , n189679 );
not ( n22404 , n189680 );
buf ( n189682 , n22404 );
buf ( n189683 , n189682 );
not ( n22407 , n189683 );
or ( n22408 , n22386 , n22407 );
buf ( n189686 , n22384 );
not ( n22410 , n189686 );
buf ( n189688 , n189679 );
nand ( n22412 , n22410 , n189688 );
buf ( n189690 , n22412 );
buf ( n189691 , n189690 );
nand ( n22415 , n22408 , n189691 );
buf ( n189693 , n22415 );
buf ( n189694 , n189693 );
buf ( n189695 , n188224 );
not ( n22419 , n189695 );
buf ( n189697 , n20244 );
not ( n22421 , n189697 );
or ( n22422 , n22419 , n22421 );
buf ( n189700 , n850 );
buf ( n189701 , n872 );
xor ( n22425 , n189700 , n189701 );
buf ( n189703 , n22425 );
buf ( n189704 , n189703 );
buf ( n189705 , n19264 );
nand ( n22429 , n189704 , n189705 );
buf ( n189707 , n22429 );
buf ( n189708 , n189707 );
nand ( n22432 , n22422 , n189708 );
buf ( n189710 , n22432 );
buf ( n189711 , n189710 );
not ( n22435 , n189711 );
buf ( n189713 , n22435 );
buf ( n189714 , n189713 );
and ( n22438 , n189694 , n189714 );
not ( n22439 , n189694 );
buf ( n189717 , n189710 );
and ( n22441 , n22439 , n189717 );
nor ( n22442 , n22438 , n22441 );
buf ( n189720 , n22442 );
buf ( n189721 , n189720 );
and ( n22445 , n189649 , n189721 );
not ( n22446 , n189649 );
buf ( n189724 , n189720 );
not ( n22448 , n189724 );
buf ( n189726 , n22448 );
buf ( n189727 , n189726 );
and ( n22451 , n22446 , n189727 );
nor ( n22452 , n22445 , n22451 );
buf ( n189730 , n22452 );
buf ( n189731 , n189730 );
xor ( n22455 , n189543 , n189731 );
xor ( n22456 , n187907 , n187919 );
and ( n22457 , n22456 , n187980 );
and ( n22458 , n187907 , n187919 );
or ( n22459 , n22457 , n22458 );
buf ( n189737 , n22459 );
buf ( n189738 , n189737 );
buf ( n189739 , n20640 );
buf ( n189740 , n188415 );
not ( n22464 , n189740 );
buf ( n189742 , n19031 );
not ( n22466 , n189742 );
or ( n22467 , n22464 , n22466 );
buf ( n189745 , n186340 );
buf ( n189746 , n858 );
buf ( n189747 , n864 );
xor ( n22471 , n189746 , n189747 );
buf ( n189749 , n22471 );
buf ( n189750 , n189749 );
nand ( n22474 , n189745 , n189750 );
buf ( n189752 , n22474 );
buf ( n189753 , n189752 );
nand ( n22477 , n22467 , n189753 );
buf ( n189755 , n22477 );
buf ( n189756 , n189755 );
xor ( n22480 , n189739 , n189756 );
xor ( n22481 , n188151 , n188168 );
and ( n22482 , n22481 , n188183 );
and ( n22483 , n188151 , n188168 );
or ( n22484 , n22482 , n22483 );
buf ( n189762 , n22484 );
xor ( n22486 , n22480 , n189762 );
buf ( n189764 , n22486 );
buf ( n189765 , n189764 );
xor ( n22489 , n189738 , n189765 );
xor ( n22490 , n187781 , n187826 );
and ( n22491 , n22490 , n187894 );
and ( n22492 , n187781 , n187826 );
or ( n22493 , n22491 , n22492 );
buf ( n189771 , n22493 );
buf ( n189772 , n189771 );
xor ( n22496 , n22489 , n189772 );
buf ( n189774 , n22496 );
buf ( n189775 , n189774 );
xor ( n22499 , n22455 , n189775 );
buf ( n189777 , n22499 );
buf ( n189778 , n189777 );
xor ( n22502 , n189439 , n189778 );
buf ( n189780 , n20419 );
buf ( n189781 , n187703 );
and ( n22505 , n189780 , n189781 );
not ( n22506 , n189780 );
buf ( n189784 , n187495 );
and ( n22508 , n22506 , n189784 );
nor ( n22509 , n22505 , n22508 );
buf ( n189787 , n22509 );
buf ( n189788 , n189787 );
not ( n22512 , n187896 );
buf ( n189790 , n22512 );
and ( n22514 , n189788 , n189790 );
not ( n22515 , n189788 );
buf ( n189793 , n187896 );
and ( n22517 , n22515 , n189793 );
nor ( n22518 , n22514 , n22517 );
buf ( n189796 , n22518 );
buf ( n189797 , n189796 );
not ( n22521 , n189797 );
buf ( n189799 , n22521 );
not ( n22523 , n189799 );
buf ( n189801 , n187982 );
buf ( n189802 , n20843 );
xor ( n22526 , n189801 , n189802 );
buf ( n189804 , n20862 );
xnor ( n22528 , n22526 , n189804 );
buf ( n189806 , n22528 );
buf ( n189807 , n189806 );
not ( n22531 , n189807 );
buf ( n189809 , n22531 );
not ( n22533 , n189809 );
or ( n22534 , n22523 , n22533 );
not ( n22535 , n189796 );
not ( n22536 , n189806 );
or ( n22537 , n22535 , n22536 );
xor ( n22538 , n188948 , n189051 );
and ( n22539 , n22538 , n189224 );
and ( n22540 , n188948 , n189051 );
or ( n22541 , n22539 , n22540 );
nand ( n22542 , n22537 , n22541 );
nand ( n22543 , n22534 , n22542 );
buf ( n189821 , n22543 );
xor ( n22545 , n22502 , n189821 );
buf ( n189823 , n22545 );
buf ( n189824 , n189823 );
nand ( n22548 , n22156 , n189824 );
buf ( n189826 , n22548 );
buf ( n189827 , n189826 );
buf ( n189828 , n188500 );
not ( n22552 , n189828 );
buf ( n189830 , n189427 );
nand ( n22554 , n22552 , n189830 );
buf ( n189832 , n22554 );
buf ( n189833 , n189832 );
nand ( n22557 , n189827 , n189833 );
buf ( n189835 , n22557 );
buf ( n22559 , n189835 );
buf ( n189837 , n189806 );
buf ( n22561 , n189837 );
buf ( n189839 , n22561 );
buf ( n189840 , n189839 );
buf ( n189841 , n189796 );
not ( n22565 , n189841 );
buf ( n189843 , n22541 );
not ( n22567 , n189843 );
and ( n22568 , n22565 , n22567 );
buf ( n189846 , n189796 );
buf ( n189847 , n22541 );
and ( n22571 , n189846 , n189847 );
nor ( n22572 , n22568 , n22571 );
buf ( n189850 , n22572 );
buf ( n189851 , n189850 );
xor ( n22575 , n189840 , n189851 );
buf ( n189853 , n22575 );
buf ( n189854 , n189853 );
xor ( n22578 , n188856 , n188942 );
xor ( n22579 , n22578 , n189423 );
buf ( n189857 , n22579 );
buf ( n189858 , n189857 );
xor ( n22582 , n189854 , n189858 );
xor ( n22583 , n189209 , n189193 );
not ( n22584 , n189179 );
xor ( n22585 , n22583 , n22584 );
buf ( n189863 , n22585 );
not ( n22587 , n189863 );
buf ( n189865 , n22587 );
not ( n22589 , n189865 );
not ( n22590 , n21753 );
not ( n22591 , n21745 );
or ( n22592 , n22590 , n22591 );
or ( n22593 , n21745 , n21753 );
nand ( n22594 , n22592 , n22593 );
not ( n22595 , n21766 );
and ( n22596 , n22594 , n22595 );
not ( n22597 , n22594 );
and ( n22598 , n22597 , n21766 );
nor ( n22599 , n22596 , n22598 );
not ( n22600 , n22599 );
not ( n22601 , n22600 );
or ( n22602 , n22589 , n22601 );
not ( n22603 , n22599 );
not ( n22604 , n22585 );
or ( n22605 , n22603 , n22604 );
xor ( n22606 , n870 , n859 );
buf ( n189884 , n22606 );
not ( n22608 , n189884 );
buf ( n189886 , n20838 );
not ( n22610 , n189886 );
or ( n22611 , n22608 , n22610 );
buf ( n189889 , n19138 );
buf ( n189890 , n21400 );
nand ( n22614 , n189889 , n189890 );
buf ( n189892 , n22614 );
buf ( n189893 , n189892 );
nand ( n22617 , n22611 , n189893 );
buf ( n189895 , n22617 );
not ( n22619 , n189895 );
buf ( n189897 , n847 );
buf ( n189898 , n882 );
xor ( n22622 , n189897 , n189898 );
buf ( n189900 , n22622 );
buf ( n189901 , n189900 );
not ( n22625 , n189901 );
buf ( n189903 , n19613 );
not ( n22627 , n189903 );
or ( n22628 , n22625 , n22627 );
buf ( n189906 , n19942 );
buf ( n189907 , n188654 );
nand ( n22631 , n189906 , n189907 );
buf ( n189909 , n22631 );
buf ( n189910 , n189909 );
nand ( n22634 , n22628 , n189910 );
buf ( n189912 , n22634 );
not ( n22636 , n189912 );
or ( n22637 , n22619 , n22636 );
buf ( n189915 , n189912 );
buf ( n189916 , n189895 );
or ( n22640 , n189915 , n189916 );
buf ( n189918 , n857 );
buf ( n189919 , n872 );
xor ( n22643 , n189918 , n189919 );
buf ( n189921 , n22643 );
buf ( n189922 , n189921 );
not ( n22646 , n189922 );
buf ( n189924 , n20244 );
not ( n22648 , n189924 );
or ( n22649 , n22646 , n22648 );
buf ( n189927 , n19264 );
buf ( n189928 , n188725 );
nand ( n22652 , n189927 , n189928 );
buf ( n189930 , n22652 );
buf ( n189931 , n189930 );
nand ( n22655 , n22649 , n189931 );
buf ( n189933 , n22655 );
buf ( n189934 , n189933 );
nand ( n22658 , n22640 , n189934 );
buf ( n189936 , n22658 );
nand ( n22660 , n22637 , n189936 );
buf ( n189938 , n851 );
buf ( n189939 , n878 );
xor ( n22663 , n189938 , n189939 );
buf ( n189941 , n22663 );
buf ( n189942 , n189941 );
not ( n22666 , n189942 );
buf ( n189944 , n186569 );
not ( n22668 , n189944 );
or ( n22669 , n22666 , n22668 );
buf ( n189947 , n186575 );
buf ( n189948 , n189329 );
nand ( n22672 , n189947 , n189948 );
buf ( n189950 , n22672 );
buf ( n189951 , n189950 );
nand ( n22675 , n22669 , n189951 );
buf ( n189953 , n22675 );
not ( n22677 , n189953 );
buf ( n189955 , n843 );
buf ( n189956 , n886 );
xor ( n22680 , n189955 , n189956 );
buf ( n189958 , n22680 );
nand ( n22682 , n189958 , n20554 );
nand ( n22683 , n20288 , n21523 );
buf ( n189961 , n188771 );
buf ( n189962 , n20279 );
nand ( n22686 , n189961 , n189962 );
buf ( n189964 , n22686 );
buf ( n189965 , n853 );
buf ( n189966 , n876 );
xor ( n22690 , n189965 , n189966 );
buf ( n189968 , n22690 );
nand ( n22692 , n19177 , n189968 );
nand ( n22693 , n22682 , n22683 , n189964 , n22692 );
not ( n22694 , n22693 );
or ( n22695 , n22677 , n22694 );
and ( n22696 , n22692 , n189964 );
not ( n22697 , n22696 );
nand ( n22698 , n22682 , n22683 );
nand ( n22699 , n22697 , n22698 );
nand ( n22700 , n22695 , n22699 );
nor ( n22701 , n22660 , n22700 );
buf ( n189979 , n845 );
buf ( n189980 , n884 );
xor ( n22704 , n189979 , n189980 );
buf ( n189982 , n22704 );
buf ( n189983 , n189982 );
not ( n22707 , n189983 );
buf ( n189985 , n20727 );
not ( n22709 , n189985 );
or ( n22710 , n22707 , n22709 );
buf ( n189988 , n188010 );
buf ( n189989 , n188709 );
nand ( n22713 , n189988 , n189989 );
buf ( n189991 , n22713 );
buf ( n189992 , n189991 );
nand ( n22716 , n22710 , n189992 );
buf ( n189994 , n22716 );
not ( n22718 , n189994 );
buf ( n189996 , n839 );
buf ( n189997 , n890 );
xor ( n22721 , n189996 , n189997 );
buf ( n189999 , n22721 );
buf ( n190000 , n189999 );
not ( n22724 , n190000 );
buf ( n190002 , n188751 );
not ( n22726 , n190002 );
or ( n22727 , n22724 , n22726 );
buf ( n190005 , n20902 );
buf ( n190006 , n188742 );
nand ( n22730 , n190005 , n190006 );
buf ( n190008 , n22730 );
buf ( n190009 , n190008 );
nand ( n22733 , n22727 , n190009 );
buf ( n190011 , n22733 );
not ( n22735 , n190011 );
or ( n22736 , n22718 , n22735 );
buf ( n190014 , n190011 );
buf ( n190015 , n189994 );
or ( n22739 , n190014 , n190015 );
buf ( n190017 , n855 );
buf ( n190018 , n874 );
xor ( n22742 , n190017 , n190018 );
buf ( n190020 , n22742 );
buf ( n190021 , n190020 );
not ( n22745 , n190021 );
buf ( n190023 , n20582 );
not ( n22747 , n190023 );
or ( n22748 , n22745 , n22747 );
buf ( n190026 , n187865 );
buf ( n190027 , n188815 );
nand ( n22751 , n190026 , n190027 );
buf ( n190029 , n22751 );
buf ( n190030 , n190029 );
nand ( n22754 , n22748 , n190030 );
buf ( n190032 , n22754 );
buf ( n190033 , n190032 );
nand ( n22757 , n22739 , n190033 );
buf ( n190035 , n22757 );
nand ( n22759 , n22736 , n190035 );
not ( n22760 , n22759 );
or ( n22761 , n22701 , n22760 );
nand ( n22762 , n22660 , n22700 );
nand ( n22763 , n22761 , n22762 );
nand ( n22764 , n22605 , n22763 );
nand ( n22765 , n22602 , n22764 );
buf ( n190043 , n22765 );
xor ( n22767 , n189213 , n189165 );
xor ( n22768 , n22767 , n189105 );
buf ( n190046 , n22768 );
xor ( n22770 , n190043 , n190046 );
xor ( n22771 , n188924 , n188906 );
xor ( n22772 , n22771 , n21654 );
buf ( n190050 , n22772 );
and ( n22774 , n22770 , n190050 );
and ( n22775 , n190043 , n190046 );
or ( n22776 , n22774 , n22775 );
buf ( n190054 , n22776 );
buf ( n190055 , n190054 );
xor ( n22779 , n188528 , n21227 );
xnor ( n22780 , n22779 , n188852 );
buf ( n190058 , n22780 );
xor ( n22782 , n190055 , n190058 );
xor ( n22783 , n188547 , n188624 );
xor ( n22784 , n22783 , n188848 );
buf ( n190062 , n22784 );
buf ( n190063 , n190062 );
buf ( n190064 , n863 );
buf ( n190065 , n867 );
or ( n22789 , n190064 , n190065 );
buf ( n190067 , n868 );
nand ( n22791 , n22789 , n190067 );
buf ( n190069 , n22791 );
buf ( n190070 , n190069 );
buf ( n190071 , n863 );
buf ( n190072 , n867 );
nand ( n22796 , n190071 , n190072 );
buf ( n190074 , n22796 );
buf ( n190075 , n190074 );
buf ( n190076 , n866 );
and ( n22800 , n190070 , n190075 , n190076 );
buf ( n190078 , n22800 );
buf ( n190079 , n190078 );
buf ( n190080 , n835 );
buf ( n190081 , n894 );
xor ( n22805 , n190080 , n190081 );
buf ( n190083 , n22805 );
buf ( n190084 , n190083 );
not ( n22808 , n190084 );
not ( n22809 , n21329 );
buf ( n190087 , n22809 );
not ( n22811 , n190087 );
or ( n22812 , n22808 , n22811 );
buf ( n190090 , n189241 );
buf ( n190091 , n895 );
nand ( n22815 , n190090 , n190091 );
buf ( n190093 , n22815 );
buf ( n190094 , n190093 );
nand ( n22818 , n22812 , n190094 );
buf ( n190096 , n22818 );
buf ( n190097 , n190096 );
and ( n22821 , n190079 , n190097 );
buf ( n190099 , n22821 );
buf ( n190100 , n190099 );
buf ( n190101 , n862 );
buf ( n190102 , n866 );
xor ( n22826 , n190101 , n190102 );
buf ( n190104 , n22826 );
buf ( n190105 , n190104 );
not ( n22829 , n190105 );
buf ( n190107 , n186241 );
not ( n22831 , n190107 );
or ( n22832 , n22829 , n22831 );
buf ( n190110 , n186254 );
buf ( n190111 , n188994 );
nand ( n22835 , n190110 , n190111 );
buf ( n190113 , n22835 );
buf ( n190114 , n190113 );
nand ( n22838 , n22832 , n190114 );
buf ( n190116 , n22838 );
buf ( n190117 , n190116 );
xor ( n22841 , n190100 , n190117 );
buf ( n190119 , n837 );
buf ( n190120 , n892 );
xor ( n22844 , n190119 , n190120 );
buf ( n190122 , n22844 );
not ( n22846 , n190122 );
not ( n22847 , n20632 );
or ( n22848 , n22846 , n22847 );
buf ( n190126 , n187477 );
buf ( n22850 , n190126 );
buf ( n190128 , n22850 );
buf ( n190129 , n190128 );
buf ( n190130 , n189257 );
nand ( n22854 , n190129 , n190130 );
buf ( n190132 , n22854 );
nand ( n22856 , n22848 , n190132 );
not ( n22857 , n22856 );
not ( n22858 , n21116 );
not ( n22859 , n22022 );
or ( n22860 , n22858 , n22859 );
not ( n22861 , n18860 );
xor ( n22862 , n880 , n849 );
and ( n22863 , n881 , n880 );
not ( n22864 , n881 );
and ( n22865 , n22864 , n18856 );
nor ( n22866 , n22863 , n22865 );
nand ( n22867 , n22861 , n22862 , n22866 );
nand ( n22868 , n22860 , n22867 );
not ( n22869 , n22868 );
or ( n22870 , n22857 , n22869 );
nor ( n22871 , n22856 , n22868 );
buf ( n190149 , n20396 );
buf ( n190150 , n189280 );
nand ( n22874 , n190149 , n190150 );
buf ( n190152 , n22874 );
buf ( n190153 , n841 );
buf ( n190154 , n888 );
xor ( n22878 , n190153 , n190154 );
buf ( n190156 , n22878 );
nand ( n22880 , n190156 , n22336 );
and ( n22881 , n190152 , n22880 );
or ( n22882 , n22871 , n22881 );
nand ( n22883 , n22870 , n22882 );
buf ( n190161 , n22883 );
and ( n22885 , n22841 , n190161 );
and ( n22886 , n190100 , n190117 );
or ( n22887 , n22885 , n22886 );
buf ( n190165 , n22887 );
buf ( n190166 , n190165 );
xor ( n22890 , n189229 , n189275 );
xor ( n22891 , n22890 , n189348 );
buf ( n190169 , n22891 );
buf ( n190170 , n190169 );
xor ( n22894 , n190166 , n190170 );
buf ( n190172 , n21559 );
buf ( n190173 , n188704 );
xor ( n22897 , n190172 , n190173 );
buf ( n190175 , n22897 );
buf ( n190176 , n190175 );
buf ( n190177 , n21488 );
xor ( n22901 , n190176 , n190177 );
buf ( n190179 , n22901 );
buf ( n190180 , n190179 );
and ( n22904 , n22894 , n190180 );
and ( n22905 , n190166 , n190170 );
or ( n22906 , n22904 , n22905 );
buf ( n190184 , n22906 );
buf ( n190185 , n190184 );
xor ( n22909 , n190063 , n190185 );
xor ( n22910 , n21444 , n21460 );
xor ( n22911 , n22910 , n21485 );
xor ( n22912 , n189247 , n189252 );
xor ( n22913 , n22912 , n189270 );
buf ( n190191 , n22913 );
or ( n22915 , n22911 , n190191 );
xor ( n22916 , n188670 , n188648 );
xnor ( n22917 , n22916 , n188693 );
nand ( n22918 , n22915 , n22917 );
buf ( n190196 , n22918 );
buf ( n190197 , n22911 );
buf ( n190198 , n190191 );
nand ( n22922 , n190197 , n190198 );
buf ( n190200 , n22922 );
buf ( n190201 , n190200 );
nand ( n22925 , n190196 , n190201 );
buf ( n190203 , n22925 );
buf ( n190204 , n190203 );
buf ( n190205 , n188834 );
not ( n22929 , n190205 );
buf ( n190207 , n22929 );
not ( n22931 , n188807 );
not ( n22932 , n21532 );
or ( n22933 , n22931 , n22932 );
or ( n22934 , n188807 , n21532 );
nand ( n22935 , n22933 , n22934 );
or ( n22936 , n190207 , n22935 );
nand ( n22937 , n22935 , n190207 );
nand ( n22938 , n22936 , n22937 );
not ( n22939 , n22938 );
buf ( n190217 , n861 );
buf ( n190218 , n868 );
xor ( n22942 , n190217 , n190218 );
buf ( n190220 , n22942 );
buf ( n190221 , n190220 );
not ( n22945 , n190221 );
buf ( n190223 , n186197 );
not ( n22947 , n190223 );
or ( n22948 , n22945 , n22947 );
buf ( n22949 , n20819 );
buf ( n190227 , n22949 );
buf ( n190228 , n188629 );
nand ( n22952 , n190227 , n190228 );
buf ( n190230 , n22952 );
buf ( n190231 , n190230 );
nand ( n22955 , n22948 , n190231 );
buf ( n190233 , n22955 );
buf ( n190234 , n190233 );
not ( n22958 , n190234 );
xor ( n22959 , n190079 , n190097 );
buf ( n190237 , n22959 );
buf ( n190238 , n190237 );
not ( n22962 , n190238 );
or ( n22963 , n22958 , n22962 );
buf ( n190241 , n190220 );
not ( n22965 , n190241 );
buf ( n190243 , n186197 );
not ( n22967 , n190243 );
or ( n22968 , n22965 , n22967 );
buf ( n190246 , n190230 );
nand ( n22970 , n22968 , n190246 );
buf ( n190248 , n22970 );
buf ( n190249 , n190248 );
buf ( n190250 , n190237 );
or ( n22974 , n190249 , n190250 );
buf ( n190252 , n863 );
buf ( n190253 , n866 );
xor ( n22977 , n190252 , n190253 );
buf ( n190255 , n22977 );
not ( n22979 , n190255 );
not ( n22980 , n186241 );
or ( n22981 , n22979 , n22980 );
buf ( n190259 , n186254 );
buf ( n190260 , n190104 );
nand ( n22984 , n190259 , n190260 );
buf ( n190262 , n22984 );
nand ( n22986 , n22981 , n190262 );
buf ( n190264 , n22986 );
nand ( n22988 , n22974 , n190264 );
buf ( n190266 , n22988 );
buf ( n190267 , n190266 );
nand ( n22991 , n22963 , n190267 );
buf ( n190269 , n22991 );
not ( n22993 , n190269 );
not ( n22994 , n22993 );
or ( n22995 , n22939 , n22994 );
buf ( n190273 , n189293 );
not ( n22997 , n190273 );
buf ( n190275 , n189317 );
not ( n22999 , n190275 );
or ( n23000 , n22997 , n22999 );
buf ( n190278 , n189317 );
buf ( n190279 , n189293 );
or ( n23003 , n190278 , n190279 );
nand ( n23004 , n23000 , n23003 );
buf ( n190282 , n23004 );
xor ( n23006 , n189341 , n190282 );
nand ( n23007 , n22995 , n23006 );
buf ( n190285 , n23007 );
not ( n23009 , n22938 );
nand ( n23010 , n190269 , n23009 );
buf ( n190288 , n23010 );
nand ( n23012 , n190285 , n190288 );
buf ( n190290 , n23012 );
buf ( n190291 , n190290 );
xor ( n23015 , n190204 , n190291 );
buf ( n190293 , n22114 );
buf ( n190294 , n22108 );
not ( n23018 , n190294 );
buf ( n190296 , n22096 );
not ( n23020 , n190296 );
or ( n23021 , n23018 , n23020 );
buf ( n190299 , n22108 );
buf ( n190300 , n22096 );
or ( n23024 , n190299 , n190300 );
nand ( n23025 , n23021 , n23024 );
buf ( n190303 , n23025 );
buf ( n190304 , n190303 );
xor ( n23028 , n190293 , n190304 );
buf ( n190306 , n23028 );
buf ( n190307 , n190306 );
and ( n23031 , n23015 , n190307 );
and ( n23032 , n190204 , n190291 );
or ( n23033 , n23031 , n23032 );
buf ( n190311 , n23033 );
buf ( n190312 , n190311 );
and ( n23036 , n22909 , n190312 );
and ( n23037 , n190063 , n190185 );
or ( n23038 , n23036 , n23037 );
buf ( n190316 , n23038 );
buf ( n190317 , n190316 );
and ( n23041 , n22782 , n190317 );
and ( n23042 , n190055 , n190058 );
or ( n23043 , n23041 , n23042 );
buf ( n190321 , n23043 );
buf ( n190322 , n190321 );
xor ( n23046 , n22582 , n190322 );
buf ( n190324 , n23046 );
buf ( n23048 , n190324 );
buf ( n190326 , n862 );
buf ( n190327 , n886 );
xor ( n23051 , n190326 , n190327 );
buf ( n190329 , n23051 );
buf ( n190330 , n190329 );
not ( n23054 , n190330 );
buf ( n190332 , n21850 );
not ( n23056 , n190332 );
buf ( n190334 , n23056 );
buf ( n190335 , n190334 );
not ( n23059 , n190335 );
buf ( n190337 , n23059 );
buf ( n190338 , n190337 );
not ( n23062 , n190338 );
or ( n23063 , n23054 , n23062 );
buf ( n190341 , n20558 );
buf ( n190342 , n861 );
buf ( n190343 , n886 );
xor ( n23067 , n190342 , n190343 );
buf ( n190345 , n23067 );
buf ( n190346 , n190345 );
nand ( n23070 , n190341 , n190346 );
buf ( n190348 , n23070 );
buf ( n190349 , n190348 );
nand ( n23073 , n23063 , n190349 );
buf ( n190351 , n23073 );
buf ( n190352 , n854 );
buf ( n190353 , n894 );
xor ( n23077 , n190352 , n190353 );
buf ( n190355 , n23077 );
buf ( n190356 , n190355 );
not ( n23080 , n190356 );
buf ( n190358 , n22809 );
not ( n23082 , n190358 );
or ( n23083 , n23080 , n23082 );
buf ( n190361 , n853 );
buf ( n190362 , n894 );
xor ( n23086 , n190361 , n190362 );
buf ( n190364 , n23086 );
buf ( n190365 , n190364 );
buf ( n190366 , n895 );
nand ( n23090 , n190365 , n190366 );
buf ( n190368 , n23090 );
buf ( n190369 , n190368 );
nand ( n23093 , n23083 , n190369 );
buf ( n190371 , n23093 );
xor ( n23095 , n190351 , n190371 );
buf ( n190373 , n858 );
buf ( n190374 , n890 );
xor ( n23098 , n190373 , n190374 );
buf ( n190376 , n23098 );
buf ( n190377 , n190376 );
not ( n23101 , n190377 );
buf ( n190379 , n188751 );
not ( n23103 , n190379 );
or ( n23104 , n23101 , n23103 );
buf ( n190382 , n20902 );
buf ( n190383 , n857 );
buf ( n190384 , n890 );
xor ( n23108 , n190383 , n190384 );
buf ( n190386 , n23108 );
buf ( n190387 , n190386 );
nand ( n23111 , n190382 , n190387 );
buf ( n190389 , n23111 );
buf ( n190390 , n190389 );
nand ( n23114 , n23104 , n190390 );
buf ( n190392 , n23114 );
xor ( n23116 , n23095 , n190392 );
buf ( n190394 , n23116 );
buf ( n190395 , n859 );
buf ( n190396 , n890 );
xor ( n23120 , n190395 , n190396 );
buf ( n190398 , n23120 );
buf ( n190399 , n190398 );
not ( n23123 , n190399 );
buf ( n190401 , n188751 );
not ( n23125 , n190401 );
or ( n23126 , n23123 , n23125 );
buf ( n23127 , n20902 );
buf ( n190405 , n23127 );
buf ( n190406 , n190376 );
nand ( n23130 , n190405 , n190406 );
buf ( n190408 , n23130 );
buf ( n190409 , n190408 );
nand ( n23133 , n23126 , n190409 );
buf ( n190411 , n23133 );
buf ( n190412 , n190411 );
buf ( n190413 , n20558 );
buf ( n190414 , n863 );
nand ( n23138 , n190413 , n190414 );
buf ( n190416 , n23138 );
buf ( n190417 , n190416 );
not ( n23141 , n190417 );
buf ( n190419 , n23141 );
buf ( n190420 , n190419 );
not ( n23144 , n190420 );
not ( n23145 , n189237 );
buf ( n190423 , n856 );
buf ( n190424 , n894 );
xor ( n23148 , n190423 , n190424 );
buf ( n190426 , n23148 );
buf ( n190427 , n190426 );
not ( n23151 , n190427 );
buf ( n190429 , n23151 );
not ( n23153 , n190429 );
and ( n23154 , n23145 , n23153 );
xor ( n23155 , n894 , n855 );
and ( n23156 , n23155 , n895 );
nor ( n23157 , n23154 , n23156 );
buf ( n190435 , n23157 );
not ( n23159 , n190435 );
buf ( n190437 , n23159 );
buf ( n190438 , n190437 );
not ( n23162 , n190438 );
or ( n23163 , n23144 , n23162 );
buf ( n190441 , n190416 );
not ( n23165 , n190441 );
buf ( n190443 , n23157 );
not ( n23167 , n190443 );
or ( n23168 , n23165 , n23167 );
buf ( n190446 , n862 );
buf ( n190447 , n888 );
xor ( n23171 , n190446 , n190447 );
buf ( n190449 , n23171 );
buf ( n190450 , n190449 );
not ( n23174 , n190450 );
buf ( n190452 , n22336 );
buf ( n23176 , n190452 );
buf ( n190454 , n23176 );
buf ( n190455 , n190454 );
not ( n23179 , n190455 );
or ( n23180 , n23174 , n23179 );
buf ( n190458 , n20396 );
buf ( n190459 , n861 );
buf ( n190460 , n888 );
xor ( n23184 , n190459 , n190460 );
buf ( n190462 , n23184 );
buf ( n190463 , n190462 );
nand ( n23187 , n190458 , n190463 );
buf ( n190465 , n23187 );
buf ( n190466 , n190465 );
nand ( n23190 , n23180 , n190466 );
buf ( n190468 , n23190 );
buf ( n190469 , n190468 );
nand ( n23193 , n23168 , n190469 );
buf ( n190471 , n23193 );
buf ( n190472 , n190471 );
nand ( n23196 , n23163 , n190472 );
buf ( n190474 , n23196 );
buf ( n190475 , n190474 );
xor ( n23199 , n190412 , n190475 );
buf ( n190477 , n857 );
buf ( n190478 , n892 );
xor ( n23202 , n190477 , n190478 );
buf ( n190480 , n23202 );
buf ( n190481 , n190480 );
not ( n23205 , n190481 );
buf ( n190483 , n187469 );
buf ( n23207 , n190483 );
buf ( n190485 , n23207 );
buf ( n190486 , n190485 );
not ( n23210 , n190486 );
or ( n23211 , n23205 , n23210 );
buf ( n190489 , n20197 );
not ( n23213 , n190489 );
buf ( n190491 , n23213 );
buf ( n190492 , n190491 );
buf ( n190493 , n856 );
buf ( n190494 , n892 );
xor ( n23218 , n190493 , n190494 );
buf ( n190496 , n23218 );
buf ( n190497 , n190496 );
nand ( n23221 , n190492 , n190497 );
buf ( n190499 , n23221 );
buf ( n190500 , n190499 );
nand ( n23224 , n23211 , n190500 );
buf ( n190502 , n23224 );
buf ( n190503 , n190502 );
not ( n23227 , n190503 );
buf ( n190505 , n863 );
buf ( n190506 , n887 );
or ( n23230 , n190505 , n190506 );
buf ( n190508 , n888 );
nand ( n23232 , n23230 , n190508 );
buf ( n190510 , n23232 );
buf ( n190511 , n190510 );
buf ( n190512 , n863 );
buf ( n190513 , n887 );
nand ( n23237 , n190512 , n190513 );
buf ( n190515 , n23237 );
buf ( n190516 , n190515 );
buf ( n190517 , n886 );
nand ( n23241 , n190511 , n190516 , n190517 );
buf ( n190519 , n23241 );
buf ( n190520 , n190519 );
not ( n23244 , n190520 );
or ( n23245 , n23227 , n23244 );
buf ( n190523 , n190519 );
buf ( n190524 , n190502 );
or ( n23248 , n190523 , n190524 );
nand ( n23249 , n23245 , n23248 );
buf ( n190527 , n23249 );
buf ( n190528 , n190527 );
and ( n23252 , n23199 , n190528 );
and ( n23253 , n190412 , n190475 );
or ( n23254 , n23252 , n23253 );
buf ( n190532 , n23254 );
buf ( n190533 , n190532 );
xor ( n23257 , n190394 , n190533 );
buf ( n190535 , n190502 );
not ( n23259 , n190535 );
buf ( n190537 , n190519 );
nor ( n23261 , n23259 , n190537 );
buf ( n190539 , n23261 );
buf ( n190540 , n190539 );
buf ( n190541 , n188010 );
buf ( n23265 , n190541 );
buf ( n190543 , n23265 );
buf ( n190544 , n190543 );
not ( n23268 , n190544 );
buf ( n190546 , n863 );
not ( n23270 , n190546 );
buf ( n190548 , n23270 );
buf ( n190549 , n190548 );
nor ( n23273 , n23268 , n190549 );
buf ( n190551 , n23273 );
buf ( n190552 , n190551 );
buf ( n190553 , n860 );
buf ( n190554 , n888 );
xor ( n23278 , n190553 , n190554 );
buf ( n190556 , n23278 );
buf ( n190557 , n190556 );
not ( n23281 , n190557 );
buf ( n190559 , n190454 );
not ( n23283 , n190559 );
or ( n23284 , n23281 , n23283 );
buf ( n190562 , n20396 );
buf ( n190563 , n859 );
buf ( n190564 , n888 );
xor ( n23288 , n190563 , n190564 );
buf ( n190566 , n23288 );
buf ( n190567 , n190566 );
nand ( n23291 , n190562 , n190567 );
buf ( n190569 , n23291 );
buf ( n190570 , n190569 );
nand ( n23294 , n23284 , n190570 );
buf ( n190572 , n23294 );
buf ( n190573 , n190572 );
xor ( n23297 , n190552 , n190573 );
buf ( n190575 , n190496 );
not ( n23299 , n190575 );
buf ( n190577 , n190485 );
not ( n23301 , n190577 );
or ( n23302 , n23299 , n23301 );
buf ( n190580 , n190491 );
buf ( n190581 , n855 );
buf ( n190582 , n892 );
xor ( n23306 , n190581 , n190582 );
buf ( n190584 , n23306 );
buf ( n190585 , n190584 );
nand ( n23309 , n190580 , n190585 );
buf ( n190587 , n23309 );
buf ( n190588 , n190587 );
nand ( n23312 , n23302 , n190588 );
buf ( n190590 , n23312 );
buf ( n190591 , n190590 );
xor ( n23315 , n23297 , n190591 );
buf ( n190593 , n23315 );
buf ( n190594 , n190593 );
xor ( n23318 , n190540 , n190594 );
buf ( n190596 , n23155 );
not ( n23320 , n190596 );
buf ( n23321 , n20165 );
buf ( n190599 , n23321 );
not ( n23323 , n190599 );
or ( n23324 , n23320 , n23323 );
buf ( n190602 , n190355 );
buf ( n190603 , n895 );
nand ( n23327 , n190602 , n190603 );
buf ( n190605 , n23327 );
buf ( n190606 , n190605 );
nand ( n23330 , n23324 , n190606 );
buf ( n190608 , n23330 );
buf ( n190609 , n190608 );
buf ( n190610 , n190462 );
not ( n23334 , n190610 );
buf ( n190612 , n190454 );
not ( n23336 , n190612 );
or ( n23337 , n23334 , n23336 );
buf ( n190615 , n20396 );
buf ( n190616 , n190556 );
nand ( n23340 , n190615 , n190616 );
buf ( n190618 , n23340 );
buf ( n190619 , n190618 );
nand ( n23343 , n23337 , n190619 );
buf ( n190621 , n23343 );
buf ( n190622 , n190621 );
xor ( n23346 , n190609 , n190622 );
xor ( n23347 , n886 , n863 );
buf ( n190625 , n23347 );
not ( n23349 , n190625 );
buf ( n190627 , n190337 );
not ( n23351 , n190627 );
or ( n23352 , n23349 , n23351 );
buf ( n23353 , n20293 );
buf ( n190631 , n23353 );
buf ( n190632 , n190329 );
nand ( n23356 , n190631 , n190632 );
buf ( n190634 , n23356 );
buf ( n190635 , n190634 );
nand ( n23359 , n23352 , n190635 );
buf ( n190637 , n23359 );
buf ( n190638 , n190637 );
and ( n23362 , n23346 , n190638 );
and ( n23363 , n190609 , n190622 );
or ( n23364 , n23362 , n23363 );
buf ( n190642 , n23364 );
buf ( n190643 , n190642 );
xor ( n23367 , n23318 , n190643 );
buf ( n190645 , n23367 );
buf ( n190646 , n190645 );
xor ( n23370 , n23257 , n190646 );
buf ( n190648 , n23370 );
buf ( n23372 , n190648 );
buf ( n190650 , n859 );
buf ( n190651 , n864 );
and ( n23375 , n190650 , n190651 );
buf ( n190653 , n23375 );
buf ( n190654 , n190653 );
buf ( n190655 , n189749 );
not ( n23379 , n190655 );
buf ( n190657 , n20335 );
not ( n23381 , n190657 );
or ( n23382 , n23379 , n23381 );
buf ( n190660 , n186340 );
buf ( n190661 , n857 );
buf ( n190662 , n864 );
xor ( n23386 , n190661 , n190662 );
buf ( n190664 , n23386 );
buf ( n190665 , n190664 );
nand ( n23389 , n190660 , n190665 );
buf ( n190667 , n23389 );
buf ( n190668 , n190667 );
nand ( n23392 , n23382 , n190668 );
buf ( n190670 , n23392 );
buf ( n190671 , n190670 );
xor ( n23395 , n190654 , n190671 );
buf ( n190673 , n189513 );
not ( n23397 , n190673 );
buf ( n190675 , n20437 );
not ( n23399 , n190675 );
or ( n23400 , n23397 , n23399 );
buf ( n190678 , n20902 );
buf ( n190679 , n890 );
nand ( n23403 , n190678 , n190679 );
buf ( n190681 , n23403 );
buf ( n190682 , n190681 );
nand ( n23406 , n23400 , n190682 );
buf ( n190684 , n23406 );
buf ( n190685 , n190684 );
not ( n23409 , n190685 );
buf ( n190687 , n23409 );
buf ( n190688 , n190687 );
xor ( n23412 , n23395 , n190688 );
buf ( n190690 , n23412 );
buf ( n190691 , n190690 );
xor ( n23415 , n189739 , n189756 );
and ( n23416 , n23415 , n189762 );
and ( n23417 , n189739 , n189756 );
or ( n23418 , n23416 , n23417 );
buf ( n190696 , n23418 );
buf ( n190697 , n190696 );
xor ( n23421 , n190691 , n190697 );
not ( n23422 , n21186 );
not ( n23423 , n21197 );
or ( n23424 , n23422 , n23423 );
not ( n23425 , n188468 );
not ( n23426 , n21198 );
or ( n23427 , n23425 , n23426 );
nand ( n23428 , n23427 , n188457 );
nand ( n23429 , n23424 , n23428 );
buf ( n190707 , n23429 );
and ( n23431 , n23421 , n190707 );
and ( n23432 , n190691 , n190697 );
or ( n23433 , n23431 , n23432 );
buf ( n190711 , n23433 );
xor ( n23435 , n189564 , n189574 );
and ( n23436 , n23435 , n189590 );
and ( n23437 , n189564 , n189574 );
or ( n23438 , n23436 , n23437 );
buf ( n190716 , n23438 );
not ( n23440 , n22329 );
not ( n23441 , n22347 );
or ( n23442 , n23440 , n23441 );
not ( n23443 , n22329 );
not ( n23444 , n23443 );
not ( n23445 , n22348 );
or ( n23446 , n23444 , n23445 );
nand ( n23447 , n23446 , n189639 );
nand ( n23448 , n23442 , n23447 );
or ( n23449 , n190716 , n23448 );
buf ( n190727 , n189673 );
not ( n23451 , n190727 );
buf ( n190729 , n20727 );
not ( n23453 , n190729 );
or ( n23454 , n23451 , n23453 );
buf ( n190732 , n190543 );
buf ( n190733 , n837 );
buf ( n190734 , n884 );
xor ( n23458 , n190733 , n190734 );
buf ( n190736 , n23458 );
buf ( n190737 , n190736 );
nand ( n23461 , n190732 , n190737 );
buf ( n190739 , n23461 );
buf ( n190740 , n190739 );
nand ( n23464 , n23454 , n190740 );
buf ( n190742 , n23464 );
buf ( n190743 , n190742 );
buf ( n190744 , n189620 );
not ( n23468 , n190744 );
buf ( n190746 , n20391 );
not ( n23470 , n190746 );
or ( n23471 , n23468 , n23470 );
buf ( n190749 , n833 );
buf ( n190750 , n888 );
xor ( n23474 , n190749 , n190750 );
buf ( n190752 , n23474 );
buf ( n190753 , n190752 );
buf ( n190754 , n20396 );
nand ( n23478 , n190753 , n190754 );
buf ( n190756 , n23478 );
buf ( n190757 , n190756 );
nand ( n23481 , n23471 , n190757 );
buf ( n190759 , n23481 );
buf ( n190760 , n190759 );
buf ( n190761 , n22174 );
not ( n23485 , n190761 );
buf ( n190763 , n20276 );
not ( n23487 , n190763 );
or ( n23488 , n23485 , n23487 );
and ( n23489 , n845 , n876 );
not ( n23490 , n845 );
and ( n23491 , n23490 , n19089 );
nor ( n23492 , n23489 , n23491 );
nand ( n23493 , n20279 , n23492 );
buf ( n190771 , n23493 );
nand ( n23495 , n23488 , n190771 );
buf ( n190773 , n23495 );
buf ( n190774 , n190773 );
and ( n23498 , n190760 , n190774 );
not ( n23499 , n190760 );
buf ( n190777 , n190773 );
not ( n23501 , n190777 );
buf ( n190779 , n23501 );
buf ( n190780 , n190779 );
and ( n23504 , n23499 , n190780 );
nor ( n23505 , n23498 , n23504 );
buf ( n190783 , n23505 );
buf ( n190784 , n190783 );
xor ( n23508 , n190743 , n190784 );
buf ( n190786 , n23508 );
nand ( n23510 , n23449 , n190786 );
buf ( n190788 , n190716 );
buf ( n190789 , n23448 );
nand ( n23513 , n190788 , n190789 );
buf ( n190791 , n23513 );
nand ( n23515 , n23510 , n190791 );
buf ( n190793 , n190684 );
buf ( n190794 , n190773 );
not ( n23518 , n190794 );
buf ( n190796 , n190759 );
not ( n23520 , n190796 );
or ( n23521 , n23518 , n23520 );
buf ( n190799 , n190759 );
buf ( n190800 , n190773 );
or ( n23524 , n190799 , n190800 );
buf ( n190802 , n190742 );
nand ( n23526 , n23524 , n190802 );
buf ( n190804 , n23526 );
buf ( n190805 , n190804 );
nand ( n23529 , n23521 , n190805 );
buf ( n190807 , n23529 );
buf ( n190808 , n190807 );
xor ( n23532 , n190793 , n190808 );
not ( n23533 , n20800 );
xor ( n23534 , n882 , n839 );
not ( n23535 , n23534 );
or ( n23536 , n23533 , n23535 );
nand ( n23537 , n189602 , n19602 , n19609 );
nand ( n23538 , n23536 , n23537 );
buf ( n190816 , n23538 );
not ( n23540 , n189657 );
not ( n23541 , n20769 );
or ( n23542 , n23540 , n23541 );
buf ( n190820 , n187865 );
buf ( n190821 , n847 );
buf ( n190822 , n874 );
xor ( n23546 , n190821 , n190822 );
buf ( n190824 , n23546 );
buf ( n190825 , n190824 );
nand ( n23549 , n190820 , n190825 );
buf ( n190827 , n23549 );
nand ( n23551 , n23542 , n190827 );
buf ( n190829 , n23551 );
xor ( n23553 , n190816 , n190829 );
buf ( n190831 , n189703 );
not ( n23555 , n190831 );
buf ( n190833 , n19260 );
not ( n23557 , n190833 );
or ( n23558 , n23555 , n23557 );
buf ( n190836 , n19265 );
buf ( n190837 , n849 );
buf ( n190838 , n872 );
xor ( n23562 , n190837 , n190838 );
buf ( n190840 , n23562 );
buf ( n190841 , n190840 );
nand ( n23565 , n190836 , n190841 );
buf ( n190843 , n23565 );
buf ( n190844 , n190843 );
nand ( n23568 , n23558 , n190844 );
buf ( n190846 , n23568 );
buf ( n190847 , n190846 );
and ( n23571 , n23553 , n190847 );
and ( n23572 , n190816 , n190829 );
or ( n23573 , n23571 , n23572 );
buf ( n190851 , n23573 );
buf ( n190852 , n190851 );
xor ( n23576 , n23532 , n190852 );
buf ( n190854 , n23576 );
xor ( n23578 , n23515 , n190854 );
not ( n23579 , n189557 );
not ( n23580 , n189549 );
or ( n23581 , n23579 , n23580 );
buf ( n190859 , n186248 );
xor ( n23583 , n866 , n855 );
buf ( n190861 , n23583 );
nand ( n23585 , n190859 , n190861 );
buf ( n190863 , n23585 );
nand ( n23587 , n23581 , n190863 );
not ( n23588 , n22292 );
not ( n23589 , n186194 );
or ( n23590 , n23588 , n23589 );
buf ( n190868 , n20819 );
xor ( n23592 , n868 , n853 );
buf ( n190870 , n23592 );
nand ( n23594 , n190868 , n190870 );
buf ( n190872 , n23594 );
nand ( n23596 , n23590 , n190872 );
xor ( n23597 , n23587 , n23596 );
not ( n23598 , n189468 );
buf ( n190876 , n21043 );
buf ( n190877 , n186565 );
nor ( n23601 , n190876 , n190877 );
buf ( n190879 , n23601 );
not ( n23603 , n190879 );
or ( n23604 , n23598 , n23603 );
buf ( n190882 , n843 );
buf ( n190883 , n878 );
xor ( n23607 , n190882 , n190883 );
buf ( n190885 , n23607 );
nand ( n23609 , n190885 , n186575 );
nand ( n23610 , n23604 , n23609 );
and ( n23611 , n23597 , n23610 );
and ( n23612 , n23587 , n23596 );
or ( n23613 , n23611 , n23612 );
not ( n23614 , n23613 );
buf ( n190892 , n22306 );
not ( n23616 , n190892 );
buf ( n190894 , n20675 );
not ( n23618 , n190894 );
or ( n23619 , n23616 , n23618 );
xor ( n23620 , n880 , n841 );
nand ( n23621 , n21116 , n23620 );
buf ( n190899 , n23621 );
nand ( n23623 , n23619 , n190899 );
buf ( n190901 , n23623 );
buf ( n190902 , n190901 );
buf ( n190903 , n22356 );
not ( n23627 , n190903 );
buf ( n190905 , n186429 );
not ( n23629 , n190905 );
or ( n23630 , n23627 , n23629 );
xor ( n23631 , n870 , n851 );
nand ( n23632 , n23631 , n20259 );
buf ( n190910 , n23632 );
nand ( n23634 , n23630 , n190910 );
buf ( n190912 , n23634 );
buf ( n190913 , n190912 );
xor ( n23637 , n190902 , n190913 );
buf ( n190915 , n189495 );
not ( n23639 , n190915 );
buf ( n190917 , n20554 );
not ( n23641 , n190917 );
or ( n23642 , n23639 , n23641 );
buf ( n190920 , n20558 );
xor ( n23644 , n886 , n835 );
buf ( n190922 , n23644 );
nand ( n23646 , n190920 , n190922 );
buf ( n190924 , n23646 );
buf ( n190925 , n190924 );
nand ( n23649 , n23642 , n190925 );
buf ( n190927 , n23649 );
buf ( n190928 , n190927 );
and ( n23652 , n23637 , n190928 );
and ( n23653 , n190902 , n190913 );
or ( n23654 , n23652 , n23653 );
buf ( n190932 , n23654 );
not ( n23656 , n190932 );
not ( n23657 , n23656 );
or ( n23658 , n23614 , n23657 );
not ( n23659 , n23613 );
nand ( n23660 , n190932 , n23659 );
nand ( n23661 , n23658 , n23660 );
buf ( n190939 , n190824 );
not ( n23663 , n190939 );
buf ( n190941 , n20582 );
not ( n23665 , n190941 );
or ( n23666 , n23663 , n23665 );
buf ( n190944 , n187865 );
buf ( n190945 , n846 );
buf ( n190946 , n874 );
xor ( n23670 , n190945 , n190946 );
buf ( n190948 , n23670 );
buf ( n190949 , n190948 );
nand ( n23673 , n190944 , n190949 );
buf ( n190951 , n23673 );
buf ( n190952 , n190951 );
nand ( n23676 , n23666 , n190952 );
buf ( n190954 , n23676 );
buf ( n190955 , n23534 );
not ( n23679 , n190955 );
buf ( n190957 , n19613 );
not ( n23681 , n190957 );
or ( n23682 , n23679 , n23681 );
buf ( n190960 , n19942 );
buf ( n190961 , n838 );
buf ( n190962 , n882 );
xor ( n23686 , n190961 , n190962 );
buf ( n190964 , n23686 );
buf ( n190965 , n190964 );
nand ( n23689 , n190960 , n190965 );
buf ( n190967 , n23689 );
buf ( n190968 , n190967 );
nand ( n23692 , n23682 , n190968 );
buf ( n190970 , n23692 );
not ( n23694 , n190970 );
and ( n23695 , n190954 , n23694 );
not ( n23696 , n190954 );
and ( n23697 , n23696 , n190970 );
nor ( n23698 , n23695 , n23697 );
buf ( n190976 , n19103 );
buf ( n190977 , n844 );
buf ( n190978 , n876 );
xor ( n23702 , n190977 , n190978 );
buf ( n190980 , n23702 );
buf ( n190981 , n190980 );
nand ( n23705 , n190976 , n190981 );
buf ( n190983 , n23705 );
nand ( n23707 , n23492 , n19098 );
nand ( n23708 , n190983 , n23707 );
not ( n23709 , n23708 );
xor ( n23710 , n23698 , n23709 );
and ( n23711 , n23661 , n23710 );
not ( n23712 , n23661 );
not ( n23713 , n23710 );
and ( n23714 , n23712 , n23713 );
nor ( n23715 , n23711 , n23714 );
xor ( n23716 , n23578 , n23715 );
xor ( n23717 , n190711 , n23716 );
xor ( n23718 , n189444 , n189458 );
and ( n23719 , n23718 , n189473 );
and ( n23720 , n189444 , n189458 );
or ( n23721 , n23719 , n23720 );
buf ( n190999 , n23721 );
buf ( n191000 , n190999 );
xor ( n23724 , n189485 , n189502 );
and ( n23725 , n23724 , n189520 );
and ( n23726 , n189485 , n189502 );
or ( n23727 , n23725 , n23726 );
buf ( n191005 , n23727 );
buf ( n191006 , n191005 );
xor ( n23730 , n191000 , n191006 );
buf ( n191008 , n189682 );
not ( n23732 , n191008 );
buf ( n191010 , n189713 );
not ( n23734 , n191010 );
or ( n23735 , n23732 , n23734 );
buf ( n191013 , n22384 );
nand ( n23737 , n23735 , n191013 );
buf ( n191015 , n23737 );
buf ( n191016 , n191015 );
buf ( n191017 , n189710 );
buf ( n191018 , n189679 );
nand ( n23742 , n191017 , n191018 );
buf ( n191020 , n23742 );
buf ( n191021 , n191020 );
nand ( n23745 , n191016 , n191021 );
buf ( n191023 , n23745 );
buf ( n191024 , n191023 );
xor ( n23748 , n23730 , n191024 );
buf ( n191026 , n23748 );
buf ( n191027 , n191026 );
xor ( n23751 , n189476 , n189523 );
and ( n23752 , n23751 , n189540 );
and ( n23753 , n189476 , n189523 );
or ( n23754 , n23752 , n23753 );
buf ( n191032 , n23754 );
buf ( n191033 , n191032 );
xor ( n23757 , n191027 , n191033 );
xor ( n23758 , n23448 , n190716 );
buf ( n191036 , n23758 );
buf ( n191037 , n190786 );
and ( n23761 , n191036 , n191037 );
not ( n23762 , n191036 );
buf ( n191040 , n190786 );
not ( n23764 , n191040 );
buf ( n191042 , n23764 );
buf ( n191043 , n191042 );
and ( n23767 , n23762 , n191043 );
nor ( n23768 , n23761 , n23767 );
buf ( n191046 , n23768 );
buf ( n191047 , n191046 );
and ( n23771 , n23757 , n191047 );
and ( n23772 , n191027 , n191033 );
or ( n23773 , n23771 , n23772 );
buf ( n191051 , n23773 );
xor ( n23775 , n23717 , n191051 );
not ( n23776 , n23775 );
not ( n23777 , n23776 );
buf ( n191055 , n189720 );
not ( n23779 , n191055 );
buf ( n191057 , n22363 );
not ( n23781 , n191057 );
or ( n23782 , n23779 , n23781 );
buf ( n191060 , n189592 );
nand ( n23784 , n23782 , n191060 );
buf ( n191062 , n23784 );
buf ( n191063 , n191062 );
buf ( n191064 , n22363 );
not ( n23788 , n191064 );
buf ( n191066 , n189726 );
nand ( n23790 , n23788 , n191066 );
buf ( n191068 , n23790 );
buf ( n191069 , n191068 );
nand ( n23793 , n191063 , n191069 );
buf ( n191071 , n23793 );
buf ( n191072 , n191071 );
xor ( n23796 , n23587 , n23596 );
xor ( n23797 , n23796 , n23610 );
buf ( n191075 , n23797 );
xor ( n23799 , n190816 , n190829 );
xor ( n23800 , n23799 , n190847 );
buf ( n191078 , n23800 );
buf ( n191079 , n191078 );
xor ( n23803 , n191075 , n191079 );
xor ( n23804 , n190902 , n190913 );
xor ( n23805 , n23804 , n190928 );
buf ( n191083 , n23805 );
buf ( n191084 , n191083 );
xor ( n23808 , n23803 , n191084 );
buf ( n191086 , n23808 );
buf ( n191087 , n191086 );
xor ( n23811 , n191072 , n191087 );
xor ( n23812 , n189738 , n189765 );
and ( n23813 , n23812 , n189772 );
and ( n23814 , n189738 , n189765 );
or ( n23815 , n23813 , n23814 );
buf ( n191093 , n23815 );
buf ( n191094 , n191093 );
and ( n23818 , n23811 , n191094 );
and ( n23819 , n191072 , n191087 );
or ( n23820 , n23818 , n23819 );
buf ( n191098 , n23820 );
xor ( n23822 , n191075 , n191079 );
and ( n23823 , n23822 , n191084 );
and ( n23824 , n191075 , n191079 );
or ( n23825 , n23823 , n23824 );
buf ( n191103 , n23825 );
buf ( n191104 , n191103 );
buf ( n191105 , n858 );
buf ( n191106 , n864 );
and ( n23830 , n191105 , n191106 );
buf ( n191108 , n23830 );
buf ( n191109 , n191108 );
buf ( n191110 , n190664 );
not ( n23834 , n191110 );
buf ( n191112 , n20335 );
not ( n23836 , n191112 );
or ( n23837 , n23834 , n23836 );
buf ( n191115 , n186337 );
buf ( n191116 , n856 );
buf ( n191117 , n864 );
xor ( n23841 , n191116 , n191117 );
buf ( n191119 , n23841 );
buf ( n191120 , n191119 );
nand ( n23844 , n191115 , n191120 );
buf ( n191122 , n23844 );
buf ( n191123 , n191122 );
nand ( n23847 , n23837 , n191123 );
buf ( n191125 , n23847 );
buf ( n191126 , n191125 );
xor ( n23850 , n191109 , n191126 );
buf ( n191128 , n190885 );
not ( n23852 , n191128 );
buf ( n191130 , n186569 );
not ( n23854 , n191130 );
or ( n23855 , n23852 , n23854 );
buf ( n191133 , n186575 );
buf ( n191134 , n842 );
buf ( n191135 , n878 );
xor ( n23859 , n191134 , n191135 );
buf ( n191137 , n23859 );
buf ( n191138 , n191137 );
nand ( n23862 , n191133 , n191138 );
buf ( n191140 , n23862 );
buf ( n191141 , n191140 );
nand ( n23865 , n23855 , n191141 );
buf ( n191143 , n23865 );
buf ( n191144 , n191143 );
xor ( n23868 , n23850 , n191144 );
buf ( n191146 , n23868 );
buf ( n191147 , n20437 );
not ( n23871 , n191147 );
buf ( n191149 , n23871 );
not ( n23873 , n20902 );
nand ( n23874 , n191149 , n23873 );
nand ( n23875 , n23874 , n890 );
nand ( n23876 , n22336 , n190752 );
buf ( n191154 , n20396 );
buf ( n191155 , n832 );
buf ( n191156 , n888 );
xor ( n23880 , n191155 , n191156 );
buf ( n191158 , n23880 );
buf ( n191159 , n191158 );
nand ( n23883 , n191154 , n191159 );
buf ( n191161 , n23883 );
nand ( n23885 , n23876 , n191161 );
not ( n23886 , n23885 );
and ( n23887 , n23875 , n23886 );
not ( n23888 , n23875 );
and ( n23889 , n23888 , n23885 );
nor ( n23890 , n23887 , n23889 );
not ( n23891 , n190736 );
not ( n23892 , n20727 );
or ( n23893 , n23891 , n23892 );
buf ( n191171 , n188010 );
buf ( n191172 , n836 );
buf ( n191173 , n884 );
xor ( n23897 , n191172 , n191173 );
buf ( n191175 , n23897 );
buf ( n191176 , n191175 );
nand ( n23900 , n191171 , n191176 );
buf ( n191178 , n23900 );
nand ( n23902 , n23893 , n191178 );
xnor ( n23903 , n23890 , n23902 );
xor ( n23904 , n191146 , n23903 );
buf ( n191182 , n23583 );
not ( n23906 , n191182 );
buf ( n191184 , n186241 );
not ( n23908 , n191184 );
or ( n23909 , n23906 , n23908 );
buf ( n191187 , n188559 );
buf ( n191188 , n854 );
buf ( n191189 , n866 );
xor ( n23913 , n191188 , n191189 );
buf ( n191191 , n23913 );
buf ( n191192 , n191191 );
nand ( n23916 , n191187 , n191192 );
buf ( n191194 , n23916 );
buf ( n191195 , n191194 );
nand ( n23919 , n23909 , n191195 );
buf ( n191197 , n23919 );
buf ( n191198 , n23592 );
not ( n23922 , n191198 );
buf ( n191200 , n18891 );
buf ( n191201 , n186191 );
and ( n23925 , n191200 , n191201 );
buf ( n191203 , n23925 );
buf ( n191204 , n191203 );
not ( n23928 , n191204 );
or ( n23929 , n23922 , n23928 );
buf ( n191207 , n18907 );
buf ( n191208 , n852 );
buf ( n191209 , n868 );
xor ( n23933 , n191208 , n191209 );
buf ( n191211 , n23933 );
buf ( n191212 , n191211 );
nand ( n23936 , n191207 , n191212 );
buf ( n191214 , n23936 );
buf ( n191215 , n191214 );
nand ( n23939 , n23929 , n191215 );
buf ( n191217 , n23939 );
xor ( n23941 , n191197 , n191217 );
buf ( n191219 , n23941 );
buf ( n191220 , n23620 );
not ( n23944 , n191220 );
buf ( n191222 , n186924 );
not ( n23946 , n191222 );
or ( n23947 , n23944 , n23946 );
buf ( n191225 , n20358 );
buf ( n23949 , n191225 );
buf ( n191227 , n23949 );
buf ( n191228 , n191227 );
buf ( n191229 , n840 );
buf ( n191230 , n880 );
xor ( n23954 , n191229 , n191230 );
buf ( n191232 , n23954 );
buf ( n191233 , n191232 );
nand ( n23957 , n191228 , n191233 );
buf ( n191235 , n23957 );
buf ( n191236 , n191235 );
nand ( n23960 , n23947 , n191236 );
buf ( n191238 , n23960 );
buf ( n191239 , n191238 );
xor ( n23963 , n191219 , n191239 );
buf ( n191241 , n23963 );
xor ( n23965 , n23904 , n191241 );
buf ( n191243 , n23965 );
xor ( n23967 , n191104 , n191243 );
xor ( n23968 , n190654 , n190671 );
and ( n23969 , n23968 , n190688 );
and ( n23970 , n190654 , n190671 );
or ( n23971 , n23969 , n23970 );
buf ( n191249 , n23971 );
buf ( n191250 , n191249 );
buf ( n191251 , n23631 );
not ( n23975 , n191251 );
buf ( n191253 , n186432 );
not ( n23977 , n191253 );
or ( n23978 , n23975 , n23977 );
buf ( n191256 , n186441 );
buf ( n191257 , n850 );
buf ( n191258 , n870 );
xor ( n23982 , n191257 , n191258 );
buf ( n191260 , n23982 );
buf ( n191261 , n191260 );
nand ( n23985 , n191256 , n191261 );
buf ( n191263 , n23985 );
buf ( n191264 , n191263 );
nand ( n23988 , n23978 , n191264 );
buf ( n191266 , n23988 );
buf ( n191267 , n190840 );
not ( n23991 , n191267 );
buf ( n191269 , n20244 );
not ( n23993 , n191269 );
or ( n23994 , n23991 , n23993 );
buf ( n191272 , n19264 );
buf ( n191273 , n848 );
buf ( n191274 , n872 );
xor ( n23998 , n191273 , n191274 );
buf ( n191276 , n23998 );
buf ( n191277 , n191276 );
nand ( n24001 , n191272 , n191277 );
buf ( n191279 , n24001 );
buf ( n191280 , n191279 );
nand ( n24004 , n23994 , n191280 );
buf ( n191282 , n24004 );
xor ( n24006 , n191266 , n191282 );
buf ( n191284 , n23644 );
not ( n24008 , n191284 );
buf ( n191286 , n20554 );
not ( n24010 , n191286 );
or ( n24011 , n24008 , n24010 );
buf ( n191289 , n20558 );
buf ( n191290 , n834 );
buf ( n191291 , n886 );
xor ( n24015 , n191290 , n191291 );
buf ( n191293 , n24015 );
buf ( n191294 , n191293 );
nand ( n24018 , n191289 , n191294 );
buf ( n191296 , n24018 );
buf ( n191297 , n191296 );
nand ( n24021 , n24011 , n191297 );
buf ( n191299 , n24021 );
xor ( n24023 , n24006 , n191299 );
buf ( n191301 , n24023 );
xor ( n24025 , n191250 , n191301 );
xor ( n24026 , n191000 , n191006 );
and ( n24027 , n24026 , n191024 );
and ( n24028 , n191000 , n191006 );
or ( n24029 , n24027 , n24028 );
buf ( n191307 , n24029 );
buf ( n191308 , n191307 );
xor ( n24032 , n24025 , n191308 );
buf ( n191310 , n24032 );
buf ( n191311 , n191310 );
xor ( n24035 , n23967 , n191311 );
buf ( n191313 , n24035 );
xor ( n24037 , n191098 , n191313 );
xor ( n24038 , n190691 , n190697 );
xor ( n24039 , n24038 , n190707 );
buf ( n191317 , n24039 );
buf ( n191318 , n191317 );
not ( n24042 , n188485 );
not ( n24043 , n21159 );
or ( n24044 , n24042 , n24043 );
not ( n24045 , n21160 );
not ( n24046 , n21202 );
or ( n24047 , n24045 , n24046 );
nand ( n24048 , n24047 , n188305 );
nand ( n24049 , n24044 , n24048 );
buf ( n191327 , n24049 );
xor ( n24051 , n191318 , n191327 );
xor ( n24052 , n191027 , n191033 );
xor ( n24053 , n24052 , n191047 );
buf ( n191331 , n24053 );
buf ( n191332 , n191331 );
and ( n24056 , n24051 , n191332 );
and ( n24057 , n191318 , n191327 );
or ( n24058 , n24056 , n24057 );
buf ( n191336 , n24058 );
xor ( n24060 , n24037 , n191336 );
not ( n24061 , n24060 );
not ( n24062 , n24061 );
or ( n24063 , n23777 , n24062 );
xor ( n24064 , n191072 , n191087 );
xor ( n24065 , n24064 , n191094 );
buf ( n191343 , n24065 );
not ( n24067 , n191343 );
xor ( n24068 , n189543 , n189731 );
and ( n24069 , n24068 , n189775 );
and ( n24070 , n189543 , n189731 );
or ( n24071 , n24069 , n24070 );
buf ( n191349 , n24071 );
not ( n24073 , n191349 );
or ( n24074 , n24067 , n24073 );
not ( n24075 , n191349 );
not ( n24076 , n24075 );
not ( n24077 , n191343 );
not ( n24078 , n24077 );
or ( n24079 , n24076 , n24078 );
buf ( n191357 , n188143 );
buf ( n191358 , n187902 );
or ( n24082 , n191357 , n191358 );
buf ( n191360 , n21210 );
nand ( n24084 , n24082 , n191360 );
buf ( n191362 , n24084 );
buf ( n191363 , n191362 );
buf ( n191364 , n188143 );
buf ( n191365 , n187495 );
not ( n24089 , n191365 );
buf ( n191367 , n20420 );
not ( n24091 , n191367 );
or ( n24092 , n24089 , n24091 );
buf ( n191370 , n187899 );
nand ( n24094 , n24092 , n191370 );
buf ( n191372 , n24094 );
buf ( n191373 , n191372 );
nand ( n24097 , n191364 , n191373 );
buf ( n191375 , n24097 );
buf ( n191376 , n191375 );
nand ( n24100 , n191363 , n191376 );
buf ( n191378 , n24100 );
nand ( n24102 , n24079 , n191378 );
nand ( n24103 , n24074 , n24102 );
buf ( n24104 , n24103 );
nand ( n24105 , n24063 , n24104 );
nand ( n24106 , n24060 , n23775 );
nand ( n24107 , n24105 , n24106 );
buf ( n24108 , n24107 );
buf ( n191386 , n22763 );
not ( n24110 , n191386 );
not ( n24111 , n22600 );
not ( n24112 , n189865 );
or ( n24113 , n24111 , n24112 );
or ( n24114 , n189865 , n22600 );
nand ( n24115 , n24113 , n24114 );
buf ( n191393 , n24115 );
not ( n24117 , n191393 );
or ( n24118 , n24110 , n24117 );
buf ( n191396 , n24115 );
buf ( n191397 , n22763 );
or ( n24121 , n191396 , n191397 );
nand ( n24122 , n24118 , n24121 );
buf ( n191400 , n24122 );
buf ( n191401 , n191400 );
xor ( n24125 , n190100 , n190117 );
xor ( n24126 , n24125 , n190161 );
buf ( n191404 , n24126 );
buf ( n191405 , n191404 );
buf ( n191406 , n842 );
buf ( n191407 , n888 );
xor ( n24131 , n191406 , n191407 );
buf ( n191409 , n24131 );
buf ( n191410 , n191409 );
not ( n24134 , n191410 );
buf ( n191412 , n190454 );
not ( n24136 , n191412 );
or ( n24137 , n24134 , n24136 );
buf ( n191415 , n20396 );
buf ( n191416 , n190156 );
nand ( n24140 , n191415 , n191416 );
buf ( n191418 , n24140 );
buf ( n191419 , n191418 );
nand ( n24143 , n24137 , n191419 );
buf ( n191421 , n24143 );
not ( n24145 , n191421 );
buf ( n191423 , n188559 );
buf ( n191424 , n863 );
and ( n24148 , n191423 , n191424 );
buf ( n191426 , n24148 );
not ( n24150 , n191426 );
or ( n24151 , n24145 , n24150 );
buf ( n191429 , n191421 );
buf ( n191430 , n191426 );
nor ( n24154 , n191429 , n191430 );
buf ( n191432 , n24154 );
buf ( n191433 , n838 );
buf ( n191434 , n892 );
xor ( n24158 , n191433 , n191434 );
buf ( n191436 , n24158 );
buf ( n191437 , n191436 );
not ( n24161 , n191437 );
buf ( n191439 , n190485 );
not ( n24163 , n191439 );
or ( n24164 , n24161 , n24163 );
buf ( n191442 , n190491 );
buf ( n191443 , n190122 );
nand ( n24167 , n191442 , n191443 );
buf ( n191445 , n24167 );
buf ( n191446 , n191445 );
nand ( n24170 , n24164 , n191446 );
buf ( n191448 , n24170 );
buf ( n191449 , n191448 );
not ( n24173 , n191449 );
buf ( n191451 , n24173 );
or ( n24175 , n191432 , n191451 );
nand ( n24176 , n24151 , n24175 );
not ( n24177 , n24176 );
buf ( n191455 , n24177 );
not ( n24179 , n191455 );
buf ( n191457 , n850 );
buf ( n191458 , n880 );
xor ( n24182 , n191457 , n191458 );
buf ( n191460 , n24182 );
buf ( n191461 , n191460 );
not ( n24185 , n191461 );
buf ( n191463 , n18862 );
not ( n24187 , n191463 );
or ( n24188 , n24185 , n24187 );
nand ( n24189 , n22304 , n22862 );
buf ( n191467 , n24189 );
nand ( n24191 , n24188 , n191467 );
buf ( n191469 , n24191 );
buf ( n191470 , n191469 );
buf ( n191471 , n852 );
buf ( n191472 , n878 );
xor ( n24196 , n191471 , n191472 );
buf ( n191474 , n24196 );
buf ( n191475 , n191474 );
not ( n24199 , n191475 );
buf ( n191477 , n186569 );
not ( n24201 , n191477 );
or ( n24202 , n24199 , n24201 );
buf ( n191480 , n186575 );
buf ( n191481 , n189941 );
nand ( n24205 , n191480 , n191481 );
buf ( n191483 , n24205 );
buf ( n191484 , n191483 );
nand ( n24208 , n24202 , n191484 );
buf ( n191486 , n24208 );
buf ( n191487 , n191486 );
xor ( n24211 , n191470 , n191487 );
buf ( n191489 , n844 );
buf ( n191490 , n886 );
xor ( n24214 , n191489 , n191490 );
buf ( n191492 , n24214 );
buf ( n191493 , n191492 );
not ( n24217 , n191493 );
buf ( n191495 , n20554 );
not ( n24219 , n191495 );
or ( n24220 , n24217 , n24219 );
buf ( n191498 , n20558 );
buf ( n191499 , n189958 );
nand ( n24223 , n191498 , n191499 );
buf ( n191501 , n24223 );
buf ( n191502 , n191501 );
nand ( n24226 , n24220 , n191502 );
buf ( n191504 , n24226 );
buf ( n191505 , n191504 );
and ( n24229 , n24211 , n191505 );
and ( n24230 , n191470 , n191487 );
or ( n24231 , n24229 , n24230 );
buf ( n191509 , n24231 );
buf ( n191510 , n191509 );
not ( n24234 , n191510 );
buf ( n191512 , n24234 );
buf ( n191513 , n191512 );
not ( n24237 , n191513 );
or ( n24238 , n24179 , n24237 );
buf ( n191516 , n836 );
buf ( n191517 , n894 );
xor ( n24241 , n191516 , n191517 );
buf ( n191519 , n24241 );
buf ( n191520 , n191519 );
not ( n24244 , n191520 );
buf ( n191522 , n22809 );
not ( n24246 , n191522 );
or ( n24247 , n24244 , n24246 );
buf ( n191525 , n190083 );
buf ( n191526 , n895 );
nand ( n24250 , n191525 , n191526 );
buf ( n191528 , n24250 );
buf ( n191529 , n191528 );
nand ( n24253 , n24247 , n191529 );
buf ( n191531 , n24253 );
not ( n24255 , n191531 );
buf ( n191533 , n854 );
buf ( n191534 , n876 );
xor ( n24258 , n191533 , n191534 );
buf ( n191536 , n24258 );
not ( n24260 , n191536 );
not ( n24261 , n19177 );
or ( n24262 , n24260 , n24261 );
buf ( n191540 , n20279 );
buf ( n191541 , n189968 );
nand ( n24265 , n191540 , n191541 );
buf ( n191543 , n24265 );
nand ( n24267 , n24262 , n191543 );
not ( n24268 , n24267 );
or ( n24269 , n24255 , n24268 );
buf ( n191547 , n24267 );
buf ( n191548 , n191531 );
nor ( n24272 , n191547 , n191548 );
buf ( n191550 , n24272 );
buf ( n191551 , n20582 );
buf ( n191552 , n856 );
buf ( n191553 , n874 );
xor ( n24277 , n191552 , n191553 );
buf ( n191555 , n24277 );
buf ( n191556 , n191555 );
and ( n24280 , n191551 , n191556 );
buf ( n191558 , n187865 );
buf ( n191559 , n190020 );
and ( n24283 , n191558 , n191559 );
nor ( n24284 , n24280 , n24283 );
buf ( n191562 , n24284 );
or ( n24286 , n191550 , n191562 );
nand ( n24287 , n24269 , n24286 );
buf ( n24288 , n24287 );
buf ( n191566 , n24288 );
nand ( n24290 , n24238 , n191566 );
buf ( n191568 , n24290 );
buf ( n191569 , n191568 );
buf ( n191570 , n191509 );
buf ( n191571 , n24176 );
nand ( n24295 , n191570 , n191571 );
buf ( n191573 , n24295 );
buf ( n191574 , n191573 );
nand ( n24298 , n191569 , n191574 );
buf ( n191576 , n24298 );
buf ( n191577 , n191576 );
xor ( n24301 , n191405 , n191577 );
not ( n24302 , n189895 );
not ( n24303 , n189933 );
not ( n24304 , n24303 );
or ( n24305 , n24302 , n24304 );
not ( n24306 , n189895 );
nand ( n24307 , n24306 , n189933 );
nand ( n24308 , n24305 , n24307 );
and ( n24309 , n24308 , n189912 );
not ( n24310 , n24308 );
not ( n24311 , n189912 );
and ( n24312 , n24310 , n24311 );
nor ( n24313 , n24309 , n24312 );
not ( n24314 , n22697 );
not ( n24315 , n22698 );
not ( n24316 , n24315 );
or ( n24317 , n24314 , n24316 );
nand ( n24318 , n22698 , n22696 );
nand ( n24319 , n24317 , n24318 );
buf ( n191597 , n24319 );
buf ( n191598 , n189953 );
xor ( n24322 , n191597 , n191598 );
buf ( n191600 , n24322 );
xor ( n24324 , n24313 , n191600 );
buf ( n191602 , n190011 );
buf ( n191603 , n190032 );
xor ( n24327 , n191602 , n191603 );
buf ( n191605 , n24327 );
buf ( n191606 , n191605 );
buf ( n191607 , n189994 );
xor ( n24331 , n191606 , n191607 );
buf ( n191609 , n24331 );
and ( n24333 , n24324 , n191609 );
and ( n24334 , n24313 , n191600 );
or ( n24335 , n24333 , n24334 );
buf ( n191613 , n24335 );
and ( n24337 , n24301 , n191613 );
and ( n24338 , n191405 , n191577 );
or ( n24339 , n24337 , n24338 );
buf ( n191617 , n24339 );
buf ( n191618 , n191617 );
xor ( n24342 , n191401 , n191618 );
not ( n24343 , n22700 );
not ( n24344 , n22759 );
and ( n24345 , n24343 , n24344 );
and ( n24346 , n22700 , n22759 );
nor ( n24347 , n24345 , n24346 );
and ( n24348 , n24347 , n22660 );
not ( n24349 , n24347 );
buf ( n191627 , n22660 );
not ( n24351 , n191627 );
buf ( n191629 , n24351 );
and ( n24353 , n24349 , n191629 );
nor ( n24354 , n24348 , n24353 );
buf ( n191632 , n24354 );
buf ( n191633 , n848 );
buf ( n191634 , n882 );
xor ( n24358 , n191633 , n191634 );
buf ( n191636 , n24358 );
not ( n24360 , n191636 );
not ( n24361 , n19613 );
or ( n24362 , n24360 , n24361 );
buf ( n191640 , n20800 );
buf ( n191641 , n189900 );
nand ( n24365 , n191640 , n191641 );
buf ( n191643 , n24365 );
nand ( n24367 , n24362 , n191643 );
not ( n24368 , n24367 );
buf ( n191646 , n862 );
buf ( n191647 , n868 );
xor ( n24371 , n191646 , n191647 );
buf ( n191649 , n24371 );
buf ( n191650 , n191649 );
not ( n24374 , n191650 );
buf ( n191652 , n191203 );
not ( n24376 , n191652 );
or ( n24377 , n24374 , n24376 );
buf ( n191655 , n18907 );
buf ( n191656 , n190220 );
nand ( n24380 , n191655 , n191656 );
buf ( n191658 , n24380 );
buf ( n191659 , n191658 );
nand ( n24383 , n24377 , n191659 );
buf ( n191661 , n24383 );
not ( n24385 , n191661 );
or ( n24386 , n24368 , n24385 );
or ( n24387 , n191661 , n24367 );
buf ( n191665 , n840 );
buf ( n191666 , n890 );
xor ( n24390 , n191665 , n191666 );
buf ( n191668 , n24390 );
buf ( n191669 , n191668 );
not ( n24393 , n191669 );
buf ( n191671 , n188751 );
not ( n24395 , n191671 );
or ( n24396 , n24393 , n24395 );
buf ( n191674 , n20902 );
buf ( n191675 , n189999 );
nand ( n24399 , n191674 , n191675 );
buf ( n191677 , n24399 );
buf ( n191678 , n191677 );
nand ( n24402 , n24396 , n191678 );
buf ( n191680 , n24402 );
nand ( n24404 , n24387 , n191680 );
nand ( n24405 , n24386 , n24404 );
buf ( n191683 , n858 );
buf ( n191684 , n872 );
xor ( n24408 , n191683 , n191684 );
buf ( n191686 , n24408 );
buf ( n191687 , n191686 );
not ( n24411 , n191687 );
buf ( n191689 , n20244 );
not ( n24413 , n191689 );
or ( n24414 , n24411 , n24413 );
buf ( n191692 , n189921 );
buf ( n191693 , n19264 );
nand ( n24417 , n191692 , n191693 );
buf ( n191695 , n24417 );
buf ( n191696 , n191695 );
nand ( n24420 , n24414 , n191696 );
buf ( n191698 , n24420 );
buf ( n191699 , n191698 );
not ( n24423 , n191699 );
buf ( n191701 , n846 );
buf ( n191702 , n884 );
xor ( n24426 , n191701 , n191702 );
buf ( n191704 , n24426 );
buf ( n191705 , n191704 );
not ( n24429 , n191705 );
buf ( n191707 , n20727 );
not ( n24431 , n191707 );
or ( n24432 , n24429 , n24431 );
buf ( n191710 , n188010 );
buf ( n191711 , n189982 );
nand ( n24435 , n191710 , n191711 );
buf ( n191713 , n24435 );
buf ( n191714 , n191713 );
nand ( n24438 , n24432 , n191714 );
buf ( n191716 , n24438 );
buf ( n191717 , n191716 );
not ( n24441 , n191717 );
or ( n24442 , n24423 , n24441 );
or ( n24443 , n191716 , n191698 );
buf ( n191721 , n860 );
buf ( n191722 , n870 );
xor ( n24446 , n191721 , n191722 );
buf ( n191724 , n24446 );
not ( n24448 , n191724 );
not ( n24449 , n186432 );
or ( n24450 , n24448 , n24449 );
buf ( n191728 , n22606 );
buf ( n191729 , n189037 );
nand ( n24453 , n191728 , n191729 );
buf ( n191731 , n24453 );
nand ( n24455 , n24450 , n191731 );
nand ( n24456 , n24443 , n24455 );
buf ( n191734 , n24456 );
nand ( n24458 , n24442 , n191734 );
buf ( n191736 , n24458 );
or ( n24460 , n24405 , n191736 );
not ( n24461 , n24460 );
xor ( n24462 , n22868 , n22881 );
xnor ( n24463 , n24462 , n22856 );
not ( n24464 , n24463 );
or ( n24465 , n24461 , n24464 );
nand ( n24466 , n191736 , n24405 );
nand ( n24467 , n24465 , n24466 );
buf ( n191745 , n24467 );
xor ( n24469 , n191632 , n191745 );
xor ( n24470 , n190269 , n23009 );
xor ( n24471 , n24470 , n23006 );
buf ( n191749 , n24471 );
and ( n24473 , n24469 , n191749 );
and ( n24474 , n191632 , n191745 );
or ( n24475 , n24473 , n24474 );
buf ( n191753 , n24475 );
buf ( n191754 , n191753 );
and ( n24478 , n24342 , n191754 );
and ( n24479 , n191401 , n191618 );
or ( n24480 , n24478 , n24479 );
buf ( n191758 , n24480 );
buf ( n191759 , n191758 );
xor ( n24483 , n190166 , n190170 );
xor ( n24484 , n24483 , n190180 );
buf ( n191762 , n24484 );
buf ( n191763 , n191762 );
xor ( n24487 , n190204 , n190291 );
xor ( n24488 , n24487 , n190307 );
buf ( n191766 , n24488 );
buf ( n191767 , n191766 );
xor ( n24491 , n191763 , n191767 );
xor ( n24492 , n22911 , n22917 );
xor ( n24493 , n24492 , n190191 );
buf ( n191771 , n24493 );
xor ( n24495 , n22986 , n190233 );
xor ( n24496 , n24495 , n190237 );
buf ( n191774 , n24496 );
buf ( n191775 , n839 );
buf ( n191776 , n892 );
xor ( n24500 , n191775 , n191776 );
buf ( n191778 , n24500 );
not ( n24502 , n191778 );
not ( n24503 , n20632 );
or ( n24504 , n24502 , n24503 );
buf ( n191782 , n190491 );
buf ( n191783 , n191436 );
nand ( n24507 , n191782 , n191783 );
buf ( n191785 , n24507 );
nand ( n24509 , n24504 , n191785 );
buf ( n191787 , n24509 );
buf ( n191788 , n863 );
buf ( n191789 , n869 );
or ( n24513 , n191788 , n191789 );
buf ( n191791 , n870 );
nand ( n24515 , n24513 , n191791 );
buf ( n191793 , n24515 );
buf ( n191794 , n863 );
buf ( n191795 , n869 );
nand ( n24519 , n191794 , n191795 );
buf ( n191797 , n24519 );
and ( n24521 , n191793 , n191797 , n868 );
buf ( n191799 , n24521 );
and ( n24523 , n191787 , n191799 );
buf ( n191801 , n24523 );
not ( n24525 , n191460 );
not ( n24526 , n20358 );
or ( n24527 , n24525 , n24526 );
not ( n24528 , n18859 );
buf ( n191806 , n851 );
buf ( n191807 , n880 );
xor ( n24531 , n191806 , n191807 );
buf ( n191809 , n24531 );
nand ( n24533 , n24528 , n191809 , n22861 );
nand ( n24534 , n24527 , n24533 );
buf ( n191812 , n24534 );
not ( n24536 , n191812 );
buf ( n191814 , n24536 );
not ( n24538 , n191814 );
buf ( n191816 , n843 );
buf ( n191817 , n888 );
xor ( n24541 , n191816 , n191817 );
buf ( n191819 , n24541 );
buf ( n191820 , n191819 );
not ( n24544 , n191820 );
buf ( n191822 , n20390 );
not ( n24546 , n191822 );
or ( n24547 , n24544 , n24546 );
buf ( n191825 , n20396 );
buf ( n191826 , n191409 );
nand ( n24550 , n191825 , n191826 );
buf ( n191828 , n24550 );
buf ( n191829 , n191828 );
nand ( n24553 , n24547 , n191829 );
buf ( n191831 , n24553 );
buf ( n191832 , n191831 );
not ( n24556 , n191832 );
buf ( n191834 , n24556 );
not ( n24558 , n191834 );
or ( n24559 , n24538 , n24558 );
buf ( n191837 , n853 );
buf ( n191838 , n878 );
xor ( n24562 , n191837 , n191838 );
buf ( n191840 , n24562 );
buf ( n191841 , n191840 );
not ( n24565 , n191841 );
buf ( n191843 , n186569 );
not ( n24567 , n191843 );
or ( n24568 , n24565 , n24567 );
buf ( n191846 , n186575 );
buf ( n191847 , n191474 );
nand ( n24571 , n191846 , n191847 );
buf ( n191849 , n24571 );
buf ( n191850 , n191849 );
nand ( n24574 , n24568 , n191850 );
buf ( n191852 , n24574 );
nand ( n24576 , n24559 , n191852 );
buf ( n191854 , n191831 );
buf ( n191855 , n24534 );
nand ( n24579 , n191854 , n191855 );
buf ( n191857 , n24579 );
nand ( n24581 , n24576 , n191857 );
xor ( n24582 , n191801 , n24581 );
buf ( n191860 , n845 );
buf ( n191861 , n886 );
xor ( n24585 , n191860 , n191861 );
buf ( n191863 , n24585 );
buf ( n191864 , n191863 );
not ( n24588 , n191864 );
buf ( n191866 , n20554 );
not ( n24590 , n191866 );
or ( n24591 , n24588 , n24590 );
buf ( n191869 , n20558 );
buf ( n191870 , n191492 );
nand ( n24594 , n191869 , n191870 );
buf ( n191872 , n24594 );
buf ( n191873 , n191872 );
nand ( n24597 , n24591 , n191873 );
buf ( n191875 , n24597 );
not ( n24599 , n191875 );
buf ( n191877 , n855 );
buf ( n191878 , n876 );
xor ( n24602 , n191877 , n191878 );
buf ( n191880 , n24602 );
buf ( n191881 , n191880 );
not ( n24605 , n191881 );
buf ( n191883 , n19098 );
not ( n24607 , n191883 );
or ( n24608 , n24605 , n24607 );
buf ( n191886 , n19103 );
buf ( n191887 , n191536 );
nand ( n24611 , n191886 , n191887 );
buf ( n191889 , n24611 );
buf ( n191890 , n191889 );
nand ( n24614 , n24608 , n191890 );
buf ( n191892 , n24614 );
not ( n24616 , n191892 );
or ( n24617 , n24599 , n24616 );
buf ( n191895 , n191875 );
buf ( n191896 , n191892 );
nor ( n24620 , n191895 , n191896 );
buf ( n191898 , n24620 );
buf ( n191899 , n186287 );
buf ( n191900 , n857 );
buf ( n191901 , n874 );
xor ( n24625 , n191900 , n191901 );
buf ( n191903 , n24625 );
buf ( n191904 , n191903 );
and ( n24628 , n191899 , n191904 );
buf ( n191906 , n187865 );
buf ( n191907 , n191555 );
and ( n24631 , n191906 , n191907 );
nor ( n24632 , n24628 , n24631 );
buf ( n191910 , n24632 );
or ( n24634 , n191898 , n191910 );
nand ( n24635 , n24617 , n24634 );
and ( n24636 , n24582 , n24635 );
and ( n24637 , n191801 , n24581 );
or ( n24638 , n24636 , n24637 );
buf ( n191916 , n24638 );
xor ( n24640 , n191774 , n191916 );
buf ( n191918 , n186254 );
buf ( n191919 , n863 );
nand ( n24643 , n191918 , n191919 );
buf ( n191921 , n24643 );
buf ( n191922 , n191921 );
buf ( n191923 , n191448 );
xor ( n24647 , n191922 , n191923 );
buf ( n191925 , n191421 );
xor ( n24649 , n24647 , n191925 );
buf ( n191927 , n24649 );
buf ( n191928 , n191927 );
not ( n24652 , n191928 );
not ( n24653 , n191661 );
not ( n24654 , n24367 );
not ( n24655 , n191680 );
and ( n24656 , n24654 , n24655 );
and ( n24657 , n24367 , n191680 );
nor ( n24658 , n24656 , n24657 );
not ( n24659 , n24658 );
or ( n24660 , n24653 , n24659 );
or ( n24661 , n191661 , n24658 );
nand ( n24662 , n24660 , n24661 );
buf ( n191940 , n24662 );
not ( n24664 , n191940 );
or ( n24665 , n24652 , n24664 );
buf ( n191943 , n191531 );
buf ( n191944 , n24267 );
xor ( n24668 , n191943 , n191944 );
buf ( n191946 , n191562 );
xnor ( n24670 , n24668 , n191946 );
buf ( n191948 , n24670 );
buf ( n191949 , n191948 );
nand ( n24673 , n24665 , n191949 );
buf ( n191951 , n24673 );
buf ( n191952 , n191951 );
buf ( n191953 , n24662 );
not ( n24677 , n191953 );
buf ( n191955 , n191927 );
not ( n24679 , n191955 );
buf ( n191957 , n24679 );
buf ( n191958 , n191957 );
nand ( n24682 , n24677 , n191958 );
buf ( n191960 , n24682 );
buf ( n191961 , n191960 );
nand ( n24685 , n191952 , n191961 );
buf ( n191963 , n24685 );
buf ( n191964 , n191963 );
and ( n24688 , n24640 , n191964 );
and ( n24689 , n191774 , n191916 );
or ( n24690 , n24688 , n24689 );
buf ( n191968 , n24690 );
buf ( n191969 , n191968 );
xor ( n24693 , n191771 , n191969 );
not ( n24694 , n24288 );
not ( n24695 , n24177 );
or ( n24696 , n24694 , n24695 );
buf ( n191974 , n24287 );
not ( n24698 , n191974 );
buf ( n191976 , n24176 );
nand ( n24700 , n24698 , n191976 );
buf ( n191978 , n24700 );
nand ( n24702 , n24696 , n191978 );
and ( n24703 , n24702 , n191512 );
not ( n24704 , n24702 );
and ( n24705 , n24704 , n191509 );
nor ( n24706 , n24703 , n24705 );
buf ( n191984 , n24706 );
not ( n24708 , n191984 );
buf ( n191986 , n191736 );
buf ( n191987 , n24405 );
xor ( n24711 , n191986 , n191987 );
buf ( n191989 , n24463 );
xnor ( n24713 , n24711 , n191989 );
buf ( n191991 , n24713 );
buf ( n191992 , n191991 );
not ( n24716 , n191992 );
or ( n24717 , n24708 , n24716 );
buf ( n191995 , n837 );
buf ( n191996 , n894 );
xor ( n24720 , n191995 , n191996 );
buf ( n191998 , n24720 );
buf ( n191999 , n191998 );
not ( n24723 , n191999 );
buf ( n192001 , n21330 );
not ( n24725 , n192001 );
or ( n24726 , n24723 , n24725 );
buf ( n192004 , n191519 );
buf ( n192005 , n895 );
nand ( n24729 , n192004 , n192005 );
buf ( n192007 , n24729 );
buf ( n192008 , n192007 );
nand ( n24732 , n24726 , n192008 );
buf ( n192010 , n24732 );
buf ( n192011 , n192010 );
buf ( n192012 , n847 );
buf ( n192013 , n884 );
xor ( n24737 , n192012 , n192013 );
buf ( n192015 , n24737 );
buf ( n192016 , n192015 );
not ( n24740 , n192016 );
buf ( n192018 , n20727 );
not ( n24742 , n192018 );
or ( n24743 , n24740 , n24742 );
buf ( n192021 , n188010 );
buf ( n192022 , n191704 );
nand ( n24746 , n192021 , n192022 );
buf ( n192024 , n24746 );
buf ( n192025 , n192024 );
nand ( n24749 , n24743 , n192025 );
buf ( n192027 , n24749 );
buf ( n192028 , n192027 );
xor ( n24752 , n192011 , n192028 );
xor ( n24753 , n872 , n859 );
buf ( n192031 , n24753 );
not ( n24755 , n192031 );
buf ( n192033 , n19260 );
not ( n24757 , n192033 );
or ( n24758 , n24755 , n24757 );
buf ( n192036 , n19264 );
buf ( n192037 , n191686 );
nand ( n24761 , n192036 , n192037 );
buf ( n192039 , n24761 );
buf ( n192040 , n192039 );
nand ( n24764 , n24758 , n192040 );
buf ( n192042 , n24764 );
buf ( n192043 , n192042 );
and ( n24767 , n24752 , n192043 );
and ( n24768 , n192011 , n192028 );
or ( n24769 , n24767 , n24768 );
buf ( n192047 , n24769 );
buf ( n192048 , n192047 );
buf ( n192049 , n841 );
buf ( n192050 , n890 );
xor ( n24774 , n192049 , n192050 );
buf ( n192052 , n24774 );
buf ( n192053 , n192052 );
not ( n24777 , n192053 );
buf ( n192055 , n188751 );
not ( n24779 , n192055 );
or ( n24780 , n24777 , n24779 );
buf ( n192058 , n20902 );
buf ( n192059 , n191668 );
nand ( n24783 , n192058 , n192059 );
buf ( n192061 , n24783 );
buf ( n192062 , n192061 );
nand ( n24786 , n24780 , n192062 );
buf ( n192064 , n24786 );
buf ( n192065 , n192064 );
not ( n24789 , n192065 );
buf ( n192067 , n863 );
buf ( n192068 , n868 );
xor ( n24792 , n192067 , n192068 );
buf ( n192070 , n24792 );
buf ( n192071 , n192070 );
not ( n24795 , n192071 );
buf ( n192073 , n191203 );
not ( n24797 , n192073 );
or ( n24798 , n24795 , n24797 );
buf ( n192076 , n22949 );
buf ( n192077 , n191649 );
nand ( n24801 , n192076 , n192077 );
buf ( n192079 , n24801 );
buf ( n192080 , n192079 );
nand ( n24804 , n24798 , n192080 );
buf ( n192082 , n24804 );
buf ( n192083 , n192082 );
not ( n24807 , n192083 );
or ( n24808 , n24789 , n24807 );
buf ( n192086 , n192064 );
buf ( n192087 , n192082 );
or ( n24811 , n192086 , n192087 );
buf ( n192089 , n861 );
buf ( n192090 , n870 );
xor ( n24814 , n192089 , n192090 );
buf ( n192092 , n24814 );
buf ( n192093 , n192092 );
not ( n24817 , n192093 );
buf ( n192095 , n186432 );
not ( n24819 , n192095 );
or ( n24820 , n24817 , n24819 );
buf ( n192098 , n189037 );
buf ( n192099 , n191724 );
nand ( n24823 , n192098 , n192099 );
buf ( n192101 , n24823 );
buf ( n192102 , n192101 );
nand ( n24826 , n24820 , n192102 );
buf ( n192104 , n24826 );
buf ( n192105 , n192104 );
nand ( n24829 , n24811 , n192105 );
buf ( n192107 , n24829 );
buf ( n192108 , n192107 );
nand ( n24832 , n24808 , n192108 );
buf ( n192110 , n24832 );
buf ( n192111 , n192110 );
xor ( n24835 , n192048 , n192111 );
xor ( n24836 , n191470 , n191487 );
xor ( n24837 , n24836 , n191505 );
buf ( n192115 , n24837 );
buf ( n192116 , n192115 );
and ( n24840 , n24835 , n192116 );
and ( n24841 , n192048 , n192111 );
or ( n24842 , n24840 , n24841 );
buf ( n192120 , n24842 );
buf ( n192121 , n192120 );
nand ( n24845 , n24717 , n192121 );
buf ( n192123 , n24845 );
buf ( n192124 , n192123 );
buf ( n192125 , n24706 );
not ( n24849 , n192125 );
buf ( n192127 , n191991 );
not ( n24851 , n192127 );
buf ( n192129 , n24851 );
buf ( n192130 , n192129 );
nand ( n24854 , n24849 , n192130 );
buf ( n192132 , n24854 );
buf ( n192133 , n192132 );
nand ( n24857 , n192124 , n192133 );
buf ( n192135 , n24857 );
buf ( n192136 , n192135 );
and ( n24860 , n24693 , n192136 );
and ( n24861 , n191771 , n191969 );
or ( n24862 , n24860 , n24861 );
buf ( n192140 , n24862 );
buf ( n192141 , n192140 );
and ( n24865 , n24491 , n192141 );
and ( n24866 , n191763 , n191767 );
or ( n24867 , n24865 , n24866 );
buf ( n192145 , n24867 );
buf ( n192146 , n192145 );
xor ( n24870 , n191759 , n192146 );
xor ( n24871 , n189352 , n22081 );
xor ( n24872 , n24871 , n189404 );
buf ( n192150 , n24872 );
xor ( n24874 , n190043 , n190046 );
xor ( n24875 , n24874 , n190050 );
buf ( n192153 , n24875 );
buf ( n192154 , n192153 );
xor ( n24878 , n192150 , n192154 );
xor ( n24879 , n190063 , n190185 );
xor ( n24880 , n24879 , n190312 );
buf ( n192158 , n24880 );
buf ( n192159 , n192158 );
xor ( n24883 , n24878 , n192159 );
buf ( n192161 , n24883 );
buf ( n192162 , n192161 );
xor ( n24886 , n24870 , n192162 );
buf ( n192164 , n24886 );
buf ( n24888 , n192164 );
buf ( n192166 , n851 );
buf ( n192167 , n866 );
xor ( n24891 , n192166 , n192167 );
buf ( n192169 , n24891 );
buf ( n192170 , n192169 );
not ( n24894 , n192170 );
buf ( n192172 , n186241 );
not ( n24896 , n192172 );
or ( n24897 , n24894 , n24896 );
buf ( n192175 , n188559 );
buf ( n192176 , n850 );
buf ( n192177 , n866 );
xor ( n24901 , n192176 , n192177 );
buf ( n192179 , n24901 );
buf ( n192180 , n192179 );
nand ( n24904 , n192175 , n192180 );
buf ( n192182 , n24904 );
buf ( n192183 , n192182 );
nand ( n24907 , n24897 , n192183 );
buf ( n192185 , n24907 );
buf ( n192186 , n849 );
buf ( n192187 , n868 );
xor ( n24911 , n192186 , n192187 );
buf ( n192189 , n24911 );
buf ( n192190 , n192189 );
not ( n24914 , n192190 );
buf ( n192192 , n186197 );
not ( n24916 , n192192 );
or ( n24917 , n24914 , n24916 );
buf ( n192195 , n22949 );
buf ( n192196 , n848 );
buf ( n192197 , n868 );
xor ( n24921 , n192196 , n192197 );
buf ( n192199 , n24921 );
buf ( n192200 , n192199 );
nand ( n24924 , n192195 , n192200 );
buf ( n192202 , n24924 );
buf ( n192203 , n192202 );
nand ( n24927 , n24917 , n192203 );
buf ( n192205 , n24927 );
xor ( n24929 , n192185 , n192205 );
buf ( n192207 , n835 );
buf ( n192208 , n882 );
xor ( n24932 , n192207 , n192208 );
buf ( n192210 , n24932 );
buf ( n192211 , n192210 );
not ( n24935 , n192211 );
buf ( n192213 , n19613 );
not ( n24937 , n192213 );
or ( n24938 , n24935 , n24937 );
buf ( n192216 , n19942 );
buf ( n192217 , n834 );
buf ( n192218 , n882 );
xor ( n24942 , n192217 , n192218 );
buf ( n192220 , n24942 );
buf ( n192221 , n192220 );
nand ( n24945 , n192216 , n192221 );
buf ( n192223 , n24945 );
buf ( n192224 , n192223 );
nand ( n24948 , n24938 , n192224 );
buf ( n192226 , n24948 );
not ( n24950 , n192226 );
and ( n24951 , n24929 , n24950 );
not ( n24952 , n24929 );
and ( n24953 , n24952 , n192226 );
nor ( n24954 , n24951 , n24953 );
buf ( n192232 , n847 );
buf ( n192233 , n870 );
xor ( n24957 , n192232 , n192233 );
buf ( n192235 , n24957 );
buf ( n192236 , n192235 );
not ( n24960 , n192236 );
buf ( n192238 , n186432 );
not ( n24962 , n192238 );
or ( n24963 , n24960 , n24962 );
buf ( n192241 , n186441 );
buf ( n192242 , n846 );
buf ( n192243 , n870 );
xor ( n24967 , n192242 , n192243 );
buf ( n192245 , n24967 );
buf ( n192246 , n192245 );
nand ( n24970 , n192241 , n192246 );
buf ( n192248 , n24970 );
buf ( n192249 , n192248 );
nand ( n24973 , n24963 , n192249 );
buf ( n192251 , n24973 );
buf ( n192252 , n192251 );
buf ( n192253 , n845 );
buf ( n192254 , n872 );
xor ( n24978 , n192253 , n192254 );
buf ( n192256 , n24978 );
buf ( n192257 , n192256 );
not ( n24981 , n192257 );
buf ( n192259 , n19260 );
not ( n24983 , n192259 );
or ( n24984 , n24981 , n24983 );
buf ( n192262 , n19265 );
buf ( n192263 , n844 );
buf ( n192264 , n872 );
xor ( n24988 , n192263 , n192264 );
buf ( n192266 , n24988 );
buf ( n192267 , n192266 );
nand ( n24991 , n192262 , n192267 );
buf ( n192269 , n24991 );
buf ( n192270 , n192269 );
nand ( n24994 , n24984 , n192270 );
buf ( n192272 , n24994 );
buf ( n192273 , n192272 );
xor ( n24997 , n192252 , n192273 );
buf ( n192275 , n839 );
buf ( n192276 , n878 );
xor ( n25000 , n192275 , n192276 );
buf ( n192278 , n25000 );
buf ( n192279 , n192278 );
not ( n25003 , n192279 );
buf ( n192281 , n186569 );
not ( n25005 , n192281 );
or ( n25006 , n25003 , n25005 );
buf ( n192284 , n186575 );
buf ( n192285 , n838 );
buf ( n192286 , n878 );
xor ( n25010 , n192285 , n192286 );
buf ( n192288 , n25010 );
buf ( n192289 , n192288 );
nand ( n25013 , n192284 , n192289 );
buf ( n192291 , n25013 );
buf ( n192292 , n192291 );
nand ( n25016 , n25006 , n192292 );
buf ( n192294 , n25016 );
buf ( n192295 , n192294 );
xor ( n25019 , n24997 , n192295 );
buf ( n192297 , n25019 );
not ( n25021 , n192297 );
xor ( n25022 , n24954 , n25021 );
not ( n25023 , n20558 );
not ( n25024 , n25023 );
buf ( n192302 , n20554 );
not ( n25026 , n192302 );
buf ( n192304 , n25026 );
not ( n25028 , n192304 );
or ( n25029 , n25024 , n25028 );
nand ( n25030 , n25029 , n886 );
buf ( n192308 , n837 );
buf ( n192309 , n880 );
xor ( n25033 , n192308 , n192309 );
buf ( n192311 , n25033 );
not ( n25035 , n192311 );
not ( n25036 , n18862 );
or ( n25037 , n25035 , n25036 );
buf ( n192315 , n22304 );
buf ( n192316 , n836 );
buf ( n192317 , n880 );
xor ( n25041 , n192316 , n192317 );
buf ( n192319 , n25041 );
buf ( n192320 , n192319 );
nand ( n25044 , n192315 , n192320 );
buf ( n192322 , n25044 );
nand ( n25046 , n25037 , n192322 );
xor ( n25047 , n25030 , n25046 );
buf ( n192325 , n833 );
buf ( n192326 , n884 );
xor ( n25050 , n192325 , n192326 );
buf ( n192328 , n25050 );
not ( n25052 , n192328 );
buf ( n192330 , n20727 );
buf ( n25054 , n192330 );
buf ( n192332 , n25054 );
not ( n25056 , n192332 );
or ( n25057 , n25052 , n25056 );
buf ( n192335 , n190543 );
buf ( n192336 , n832 );
buf ( n192337 , n884 );
xor ( n25061 , n192336 , n192337 );
buf ( n192339 , n25061 );
buf ( n192340 , n192339 );
nand ( n25064 , n192335 , n192340 );
buf ( n192342 , n25064 );
nand ( n25066 , n25057 , n192342 );
xor ( n25067 , n25047 , n25066 );
xor ( n25068 , n25022 , n25067 );
buf ( n192346 , n854 );
buf ( n192347 , n864 );
and ( n25071 , n192346 , n192347 );
buf ( n192349 , n25071 );
buf ( n192350 , n192349 );
buf ( n192351 , n853 );
buf ( n192352 , n864 );
xor ( n25076 , n192351 , n192352 );
buf ( n192354 , n25076 );
buf ( n192355 , n192354 );
not ( n25079 , n192355 );
buf ( n192357 , n19031 );
not ( n25081 , n192357 );
or ( n25082 , n25079 , n25081 );
buf ( n192360 , n186340 );
buf ( n192361 , n852 );
buf ( n192362 , n864 );
xor ( n25086 , n192361 , n192362 );
buf ( n192364 , n25086 );
buf ( n192365 , n192364 );
nand ( n25089 , n192360 , n192365 );
buf ( n192367 , n25089 );
buf ( n192368 , n192367 );
nand ( n25092 , n25082 , n192368 );
buf ( n192370 , n25092 );
buf ( n192371 , n192370 );
xor ( n25095 , n192350 , n192371 );
buf ( n192373 , n841 );
buf ( n192374 , n876 );
xor ( n25098 , n192373 , n192374 );
buf ( n192376 , n25098 );
buf ( n192377 , n192376 );
not ( n25101 , n192377 );
buf ( n192379 , n19098 );
not ( n25103 , n192379 );
or ( n25104 , n25101 , n25103 );
buf ( n192382 , n20279 );
buf ( n192383 , n840 );
buf ( n192384 , n876 );
xor ( n25108 , n192383 , n192384 );
buf ( n192386 , n25108 );
buf ( n192387 , n192386 );
nand ( n25111 , n192382 , n192387 );
buf ( n192389 , n25111 );
buf ( n192390 , n192389 );
nand ( n25114 , n25104 , n192390 );
buf ( n192392 , n25114 );
buf ( n192393 , n192392 );
xor ( n25117 , n25095 , n192393 );
buf ( n192395 , n25117 );
buf ( n192396 , n192395 );
xor ( n25120 , n874 , n843 );
buf ( n192398 , n25120 );
not ( n25122 , n192398 );
buf ( n192400 , n20582 );
not ( n25124 , n192400 );
or ( n25125 , n25122 , n25124 );
buf ( n192403 , n186297 );
buf ( n192404 , n842 );
buf ( n192405 , n874 );
xor ( n25129 , n192404 , n192405 );
buf ( n192407 , n25129 );
buf ( n192408 , n192407 );
nand ( n25132 , n192403 , n192408 );
buf ( n192410 , n25132 );
buf ( n192411 , n192410 );
nand ( n25135 , n25125 , n192411 );
buf ( n192413 , n25135 );
buf ( n192414 , n192413 );
buf ( n192415 , n834 );
buf ( n192416 , n884 );
xor ( n25140 , n192415 , n192416 );
buf ( n192418 , n25140 );
buf ( n192419 , n192418 );
not ( n25143 , n192419 );
buf ( n192421 , n192332 );
not ( n25145 , n192421 );
or ( n25146 , n25143 , n25145 );
buf ( n192424 , n190543 );
buf ( n192425 , n192328 );
nand ( n25149 , n192424 , n192425 );
buf ( n192427 , n25149 );
buf ( n192428 , n192427 );
nand ( n25152 , n25146 , n192428 );
buf ( n192430 , n25152 );
buf ( n192431 , n192430 );
xor ( n25155 , n192414 , n192431 );
buf ( n192433 , n850 );
buf ( n192434 , n868 );
xor ( n25158 , n192433 , n192434 );
buf ( n192436 , n25158 );
buf ( n192437 , n192436 );
not ( n25161 , n192437 );
buf ( n192439 , n191203 );
not ( n25163 , n192439 );
or ( n25164 , n25161 , n25163 );
buf ( n192442 , n22949 );
buf ( n192443 , n192189 );
nand ( n25167 , n192442 , n192443 );
buf ( n192445 , n25167 );
buf ( n192446 , n192445 );
nand ( n25170 , n25164 , n192446 );
buf ( n192448 , n25170 );
not ( n25172 , n192448 );
buf ( n192450 , n852 );
buf ( n192451 , n866 );
xor ( n25175 , n192450 , n192451 );
buf ( n192453 , n25175 );
buf ( n192454 , n192453 );
not ( n25178 , n192454 );
buf ( n192456 , n186241 );
not ( n25180 , n192456 );
or ( n25181 , n25178 , n25180 );
buf ( n192459 , n186248 );
buf ( n192460 , n192169 );
nand ( n25184 , n192459 , n192460 );
buf ( n192462 , n25184 );
buf ( n192463 , n192462 );
nand ( n25187 , n25181 , n192463 );
buf ( n192465 , n25187 );
not ( n25189 , n192465 );
or ( n25190 , n25172 , n25189 );
buf ( n192468 , n192448 );
buf ( n192469 , n192465 );
nor ( n25193 , n192468 , n192469 );
buf ( n192471 , n25193 );
buf ( n192472 , n840 );
buf ( n192473 , n878 );
xor ( n25197 , n192472 , n192473 );
buf ( n192475 , n25197 );
buf ( n192476 , n192475 );
not ( n25200 , n192476 );
buf ( n192478 , n186569 );
not ( n25202 , n192478 );
or ( n25203 , n25200 , n25202 );
buf ( n192481 , n186575 );
buf ( n192482 , n192278 );
nand ( n25206 , n192481 , n192482 );
buf ( n192484 , n25206 );
buf ( n192485 , n192484 );
nand ( n25209 , n25203 , n192485 );
buf ( n192487 , n25209 );
buf ( n192488 , n192487 );
not ( n25212 , n192488 );
buf ( n192490 , n25212 );
or ( n25214 , n192471 , n192490 );
nand ( n25215 , n25190 , n25214 );
buf ( n192493 , n25215 );
xor ( n25217 , n25155 , n192493 );
buf ( n192495 , n25217 );
buf ( n192496 , n192495 );
xor ( n25220 , n192396 , n192496 );
buf ( n192498 , n192418 );
not ( n25222 , n192498 );
buf ( n192500 , n192332 );
not ( n25224 , n192500 );
or ( n25225 , n25222 , n25224 );
buf ( n192503 , n192427 );
nand ( n25227 , n25225 , n192503 );
buf ( n192505 , n25227 );
buf ( n192506 , n192505 );
not ( n25230 , n192506 );
buf ( n192508 , n25230 );
buf ( n192509 , n192508 );
buf ( n192510 , n851 );
buf ( n192511 , n868 );
xor ( n25235 , n192510 , n192511 );
buf ( n192513 , n25235 );
buf ( n192514 , n192513 );
not ( n25238 , n192514 );
buf ( n192516 , n191203 );
not ( n25240 , n192516 );
or ( n25241 , n25238 , n25240 );
buf ( n192519 , n18907 );
buf ( n192520 , n192436 );
nand ( n25244 , n192519 , n192520 );
buf ( n192522 , n25244 );
buf ( n192523 , n192522 );
nand ( n25247 , n25241 , n192523 );
buf ( n192525 , n25247 );
buf ( n192526 , n192525 );
not ( n25250 , n192526 );
buf ( n192528 , n849 );
buf ( n192529 , n870 );
xor ( n25253 , n192528 , n192529 );
buf ( n192531 , n25253 );
buf ( n192532 , n192531 );
not ( n25256 , n192532 );
buf ( n192534 , n20838 );
not ( n25258 , n192534 );
or ( n25259 , n25256 , n25258 );
buf ( n192537 , n186441 );
buf ( n192538 , n848 );
buf ( n192539 , n870 );
xor ( n25263 , n192538 , n192539 );
buf ( n192541 , n25263 );
buf ( n192542 , n192541 );
nand ( n25266 , n192537 , n192542 );
buf ( n192544 , n25266 );
buf ( n192545 , n192544 );
nand ( n25269 , n25259 , n192545 );
buf ( n192547 , n25269 );
buf ( n192548 , n192547 );
not ( n25272 , n192548 );
or ( n25273 , n25250 , n25272 );
buf ( n192551 , n192547 );
not ( n25275 , n192551 );
buf ( n192553 , n25275 );
buf ( n192554 , n192553 );
not ( n25278 , n192554 );
buf ( n192556 , n192525 );
not ( n25280 , n192556 );
buf ( n192558 , n25280 );
buf ( n192559 , n192558 );
not ( n25283 , n192559 );
or ( n25284 , n25278 , n25283 );
buf ( n192562 , n835 );
buf ( n192563 , n884 );
xor ( n25287 , n192562 , n192563 );
buf ( n192565 , n25287 );
buf ( n192566 , n192565 );
not ( n25290 , n192566 );
buf ( n192568 , n192332 );
not ( n25292 , n192568 );
or ( n25293 , n25290 , n25292 );
buf ( n192571 , n188010 );
buf ( n25295 , n192571 );
buf ( n192573 , n25295 );
buf ( n192574 , n192573 );
buf ( n192575 , n192418 );
nand ( n25299 , n192574 , n192575 );
buf ( n192577 , n25299 );
buf ( n192578 , n192577 );
nand ( n25302 , n25293 , n192578 );
buf ( n192580 , n25302 );
buf ( n192581 , n192580 );
nand ( n25305 , n25284 , n192581 );
buf ( n192583 , n25305 );
buf ( n192584 , n192583 );
nand ( n25308 , n25273 , n192584 );
buf ( n192586 , n25308 );
buf ( n192587 , n192586 );
xor ( n25311 , n192509 , n192587 );
buf ( n192589 , n847 );
buf ( n192590 , n872 );
xor ( n25314 , n192589 , n192590 );
buf ( n192592 , n25314 );
buf ( n192593 , n192592 );
not ( n25317 , n192593 );
not ( n25318 , n20243 );
buf ( n192596 , n25318 );
not ( n25320 , n192596 );
or ( n25321 , n25317 , n25320 );
buf ( n192599 , n19264 );
buf ( n192600 , n846 );
buf ( n192601 , n872 );
xor ( n25325 , n192600 , n192601 );
buf ( n192603 , n25325 );
buf ( n192604 , n192603 );
nand ( n25328 , n192599 , n192604 );
buf ( n192606 , n25328 );
buf ( n192607 , n192606 );
nand ( n25331 , n25321 , n192607 );
buf ( n192609 , n25331 );
buf ( n192610 , n192609 );
buf ( n192611 , n845 );
buf ( n192612 , n874 );
xor ( n25336 , n192611 , n192612 );
buf ( n192614 , n25336 );
buf ( n192615 , n192614 );
not ( n25339 , n192615 );
buf ( n192617 , n18992 );
not ( n25341 , n192617 );
or ( n25342 , n25339 , n25341 );
buf ( n192620 , n188823 );
xor ( n25344 , n874 , n844 );
buf ( n192622 , n25344 );
nand ( n25346 , n192620 , n192622 );
buf ( n192624 , n25346 );
buf ( n192625 , n192624 );
nand ( n25349 , n25342 , n192625 );
buf ( n192627 , n25349 );
buf ( n192628 , n192627 );
xor ( n25352 , n192610 , n192628 );
buf ( n192630 , n839 );
buf ( n192631 , n880 );
xor ( n25355 , n192630 , n192631 );
buf ( n192633 , n25355 );
buf ( n192634 , n192633 );
not ( n25358 , n192634 );
buf ( n192636 , n18862 );
not ( n25360 , n192636 );
or ( n25361 , n25358 , n25360 );
buf ( n192639 , n191227 );
buf ( n192640 , n838 );
buf ( n192641 , n880 );
xor ( n25365 , n192640 , n192641 );
buf ( n192643 , n25365 );
buf ( n192644 , n192643 );
nand ( n25368 , n192639 , n192644 );
buf ( n192646 , n25368 );
buf ( n192647 , n192646 );
nand ( n25371 , n25361 , n192647 );
buf ( n192649 , n25371 );
buf ( n192650 , n192649 );
and ( n25374 , n25352 , n192650 );
and ( n25375 , n192610 , n192628 );
or ( n25376 , n25374 , n25375 );
buf ( n192654 , n25376 );
buf ( n192655 , n192654 );
and ( n25379 , n25311 , n192655 );
and ( n25380 , n192509 , n192587 );
or ( n25381 , n25379 , n25380 );
buf ( n192659 , n25381 );
buf ( n192660 , n192659 );
xor ( n25384 , n25220 , n192660 );
buf ( n192662 , n25384 );
xor ( n25386 , n25068 , n192662 );
buf ( n192664 , n856 );
buf ( n192665 , n864 );
and ( n25389 , n192664 , n192665 );
buf ( n192667 , n25389 );
buf ( n192668 , n192667 );
buf ( n192669 , n843 );
buf ( n192670 , n876 );
xor ( n25394 , n192669 , n192670 );
buf ( n192672 , n25394 );
buf ( n192673 , n192672 );
not ( n25397 , n192673 );
buf ( n192675 , n19177 );
not ( n25399 , n192675 );
or ( n25400 , n25397 , n25399 );
buf ( n192678 , n19103 );
buf ( n192679 , n842 );
buf ( n192680 , n876 );
xor ( n25404 , n192679 , n192680 );
buf ( n192682 , n25404 );
buf ( n192683 , n192682 );
nand ( n25407 , n192678 , n192683 );
buf ( n192685 , n25407 );
buf ( n192686 , n192685 );
nand ( n25410 , n25400 , n192686 );
buf ( n192688 , n25410 );
buf ( n192689 , n192688 );
xor ( n25413 , n192668 , n192689 );
buf ( n192691 , n191293 );
not ( n25415 , n192691 );
buf ( n192693 , n20554 );
not ( n25417 , n192693 );
or ( n25418 , n25415 , n25417 );
buf ( n192696 , n20558 );
buf ( n192697 , n833 );
buf ( n192698 , n886 );
xor ( n25422 , n192697 , n192698 );
buf ( n192700 , n25422 );
buf ( n192701 , n192700 );
nand ( n25425 , n192696 , n192701 );
buf ( n192703 , n25425 );
buf ( n192704 , n192703 );
nand ( n25428 , n25418 , n192704 );
buf ( n192706 , n25428 );
buf ( n192707 , n192706 );
and ( n25431 , n25413 , n192707 );
and ( n25432 , n192668 , n192689 );
or ( n25433 , n25431 , n25432 );
buf ( n192711 , n25433 );
buf ( n192712 , n192711 );
buf ( n192713 , n191232 );
not ( n25437 , n192713 );
buf ( n192715 , n20675 );
not ( n25439 , n192715 );
or ( n25440 , n25437 , n25439 );
buf ( n192718 , n20358 );
buf ( n192719 , n192633 );
nand ( n25443 , n192718 , n192719 );
buf ( n192721 , n25443 );
buf ( n192722 , n192721 );
nand ( n25446 , n25440 , n192722 );
buf ( n192724 , n25446 );
buf ( n192725 , n192724 );
buf ( n192726 , n191211 );
not ( n25450 , n192726 );
buf ( n192728 , n191203 );
not ( n25452 , n192728 );
or ( n25453 , n25450 , n25452 );
buf ( n192731 , n18907 );
buf ( n192732 , n192513 );
nand ( n25456 , n192731 , n192732 );
buf ( n192734 , n25456 );
buf ( n192735 , n192734 );
nand ( n25459 , n25453 , n192735 );
buf ( n192737 , n25459 );
buf ( n192738 , n192737 );
or ( n25462 , n192725 , n192738 );
buf ( n192740 , n191260 );
not ( n25464 , n192740 );
buf ( n192742 , n186432 );
not ( n25466 , n192742 );
or ( n25467 , n25464 , n25466 );
buf ( n192745 , n189037 );
buf ( n192746 , n192531 );
nand ( n25470 , n192745 , n192746 );
buf ( n192748 , n25470 );
buf ( n192749 , n192748 );
nand ( n25473 , n25467 , n192749 );
buf ( n192751 , n25473 );
buf ( n192752 , n192751 );
nand ( n25476 , n25462 , n192752 );
buf ( n192754 , n25476 );
buf ( n192755 , n192754 );
buf ( n192756 , n192737 );
buf ( n192757 , n192724 );
nand ( n25481 , n192756 , n192757 );
buf ( n192759 , n25481 );
buf ( n192760 , n192759 );
nand ( n25484 , n192755 , n192760 );
buf ( n192762 , n25484 );
buf ( n192763 , n192762 );
buf ( n192764 , n25318 );
buf ( n192765 , n191276 );
and ( n25489 , n192764 , n192765 );
buf ( n192767 , n19264 );
buf ( n192768 , n192592 );
and ( n25492 , n192767 , n192768 );
nor ( n25493 , n25489 , n25492 );
buf ( n192771 , n25493 );
buf ( n192772 , n192771 );
not ( n25496 , n192772 );
buf ( n192774 , n25496 );
buf ( n192775 , n192774 );
not ( n25499 , n192775 );
buf ( n192777 , n190964 );
not ( n25501 , n192777 );
buf ( n192779 , n19613 );
not ( n25503 , n192779 );
or ( n25504 , n25501 , n25503 );
buf ( n192782 , n837 );
buf ( n192783 , n882 );
xor ( n25507 , n192782 , n192783 );
buf ( n192785 , n25507 );
buf ( n192786 , n192785 );
buf ( n192787 , n19942 );
nand ( n25511 , n192786 , n192787 );
buf ( n192789 , n25511 );
buf ( n192790 , n192789 );
nand ( n25514 , n25504 , n192790 );
buf ( n192792 , n25514 );
buf ( n192793 , n192792 );
not ( n25517 , n192793 );
or ( n25518 , n25499 , n25517 );
not ( n25519 , n192792 );
buf ( n192797 , n25519 );
not ( n25521 , n192797 );
buf ( n192799 , n192771 );
not ( n25523 , n192799 );
or ( n25524 , n25521 , n25523 );
buf ( n192802 , n190948 );
not ( n25526 , n192802 );
buf ( n192804 , n18992 );
not ( n25528 , n192804 );
or ( n25529 , n25526 , n25528 );
buf ( n192807 , n187865 );
buf ( n192808 , n192614 );
nand ( n25532 , n192807 , n192808 );
buf ( n192810 , n25532 );
buf ( n192811 , n192810 );
nand ( n25535 , n25529 , n192811 );
buf ( n192813 , n25535 );
buf ( n192814 , n192813 );
nand ( n25538 , n25524 , n192814 );
buf ( n192816 , n25538 );
buf ( n192817 , n192816 );
nand ( n25541 , n25518 , n192817 );
buf ( n192819 , n25541 );
buf ( n192820 , n192819 );
xor ( n25544 , n192763 , n192820 );
not ( n25545 , n20396 );
not ( n25546 , n888 );
or ( n25547 , n25545 , n25546 );
nand ( n25548 , n191158 , n22336 );
nand ( n25549 , n25547 , n25548 );
buf ( n192827 , n25549 );
not ( n25551 , n192827 );
buf ( n192829 , n25551 );
buf ( n192830 , n192829 );
not ( n25554 , n192830 );
buf ( n192832 , n191191 );
not ( n25556 , n192832 );
buf ( n192834 , n186241 );
not ( n25558 , n192834 );
or ( n25559 , n25556 , n25558 );
buf ( n192837 , n188559 );
buf ( n192838 , n853 );
buf ( n192839 , n866 );
xor ( n25563 , n192838 , n192839 );
buf ( n192841 , n25563 );
buf ( n192842 , n192841 );
nand ( n25566 , n192837 , n192842 );
buf ( n192844 , n25566 );
buf ( n192845 , n192844 );
nand ( n25569 , n25559 , n192845 );
buf ( n192847 , n25569 );
buf ( n192848 , n192847 );
not ( n25572 , n192848 );
buf ( n192850 , n25572 );
buf ( n192851 , n192850 );
not ( n25575 , n192851 );
or ( n25576 , n25554 , n25575 );
buf ( n192854 , n191137 );
not ( n25578 , n192854 );
buf ( n192856 , n186789 );
not ( n25580 , n192856 );
or ( n25581 , n25578 , n25580 );
buf ( n192859 , n186575 );
buf ( n192860 , n841 );
buf ( n192861 , n878 );
xor ( n25585 , n192860 , n192861 );
buf ( n192863 , n25585 );
buf ( n192864 , n192863 );
nand ( n25588 , n192859 , n192864 );
buf ( n192866 , n25588 );
buf ( n192867 , n192866 );
nand ( n25591 , n25581 , n192867 );
buf ( n192869 , n25591 );
buf ( n192870 , n192869 );
nand ( n25594 , n25576 , n192870 );
buf ( n192872 , n25594 );
buf ( n192873 , n192872 );
buf ( n192874 , n25549 );
buf ( n192875 , n192847 );
nand ( n25599 , n192874 , n192875 );
buf ( n192877 , n25599 );
buf ( n192878 , n192877 );
nand ( n25602 , n192873 , n192878 );
buf ( n192880 , n25602 );
buf ( n192881 , n192880 );
and ( n25605 , n25544 , n192881 );
and ( n25606 , n192763 , n192820 );
or ( n25607 , n25605 , n25606 );
buf ( n192885 , n25607 );
buf ( n192886 , n192885 );
xor ( n25610 , n192712 , n192886 );
xor ( n25611 , n192509 , n192587 );
xor ( n25612 , n25611 , n192655 );
buf ( n192890 , n25612 );
buf ( n192891 , n192890 );
and ( n25615 , n25610 , n192891 );
and ( n25616 , n192712 , n192886 );
or ( n25617 , n25615 , n25616 );
buf ( n192895 , n25617 );
xor ( n25619 , n25386 , n192895 );
buf ( n192897 , n25619 );
buf ( n192898 , n192863 );
not ( n25622 , n192898 );
buf ( n192900 , n186569 );
not ( n25624 , n192900 );
or ( n25625 , n25622 , n25624 );
buf ( n192903 , n186575 );
buf ( n192904 , n192475 );
nand ( n25628 , n192903 , n192904 );
buf ( n192906 , n25628 );
buf ( n192907 , n192906 );
nand ( n25631 , n25625 , n192907 );
buf ( n192909 , n25631 );
buf ( n192910 , n192909 );
not ( n25634 , n192910 );
buf ( n192912 , n192841 );
not ( n25636 , n192912 );
buf ( n192914 , n186241 );
not ( n25638 , n192914 );
or ( n25639 , n25636 , n25638 );
buf ( n192917 , n188559 );
buf ( n192918 , n192453 );
nand ( n25642 , n192917 , n192918 );
buf ( n192920 , n25642 );
buf ( n192921 , n192920 );
nand ( n25645 , n25639 , n192921 );
buf ( n192923 , n25645 );
buf ( n192924 , n192923 );
not ( n25648 , n192924 );
buf ( n192926 , n25648 );
buf ( n192927 , n192926 );
not ( n25651 , n192927 );
or ( n25652 , n25634 , n25651 );
buf ( n192930 , n192909 );
not ( n25654 , n192930 );
buf ( n192932 , n192923 );
nand ( n25656 , n25654 , n192932 );
buf ( n192934 , n25656 );
buf ( n192935 , n192934 );
nand ( n25659 , n25652 , n192935 );
buf ( n192937 , n25659 );
buf ( n192938 , n192937 );
buf ( n192939 , n855 );
buf ( n192940 , n864 );
xor ( n25664 , n192939 , n192940 );
buf ( n192942 , n25664 );
buf ( n192943 , n192942 );
not ( n25667 , n192943 );
buf ( n192945 , n19031 );
not ( n25669 , n192945 );
or ( n25670 , n25667 , n25669 );
buf ( n192948 , n186340 );
buf ( n192949 , n854 );
buf ( n192950 , n864 );
xor ( n25674 , n192949 , n192950 );
buf ( n192952 , n25674 );
buf ( n192953 , n192952 );
nand ( n25677 , n192948 , n192953 );
buf ( n192955 , n25677 );
buf ( n192956 , n192955 );
nand ( n25680 , n25670 , n192956 );
buf ( n192958 , n25680 );
buf ( n192959 , n192958 );
not ( n25683 , n192959 );
buf ( n192961 , n25683 );
buf ( n192962 , n192961 );
and ( n25686 , n192938 , n192962 );
not ( n25687 , n192938 );
buf ( n192965 , n192958 );
and ( n25689 , n25687 , n192965 );
nor ( n25690 , n25686 , n25689 );
buf ( n192968 , n25690 );
buf ( n192969 , n192968 );
not ( n25693 , n192969 );
buf ( n192971 , n25693 );
not ( n25695 , n192971 );
xor ( n25696 , n192668 , n192689 );
xor ( n25697 , n25696 , n192707 );
buf ( n192975 , n25697 );
not ( n25699 , n192975 );
or ( n25700 , n25695 , n25699 );
buf ( n192978 , n192971 );
buf ( n192979 , n192975 );
or ( n25703 , n192978 , n192979 );
xor ( n25704 , n192547 , n192558 );
xnor ( n25705 , n25704 , n192580 );
buf ( n192983 , n25705 );
nand ( n25707 , n25703 , n192983 );
buf ( n192985 , n25707 );
nand ( n25709 , n25700 , n192985 );
buf ( n192987 , n25709 );
buf ( n192988 , n857 );
buf ( n192989 , n864 );
and ( n25713 , n192988 , n192989 );
buf ( n192991 , n25713 );
buf ( n192992 , n192991 );
buf ( n192993 , n191119 );
not ( n25717 , n192993 );
buf ( n192995 , n19031 );
not ( n25719 , n192995 );
or ( n25720 , n25717 , n25719 );
buf ( n192998 , n186340 );
buf ( n192999 , n192942 );
nand ( n25723 , n192998 , n192999 );
buf ( n193001 , n25723 );
buf ( n193002 , n193001 );
nand ( n25726 , n25720 , n193002 );
buf ( n193004 , n25726 );
buf ( n193005 , n193004 );
xor ( n25729 , n192992 , n193005 );
buf ( n193007 , n191175 );
not ( n25731 , n193007 );
buf ( n193009 , n192332 );
not ( n25733 , n193009 );
or ( n25734 , n25731 , n25733 );
buf ( n193012 , n192573 );
buf ( n193013 , n192565 );
nand ( n25737 , n193012 , n193013 );
buf ( n193015 , n25737 );
buf ( n193016 , n193015 );
nand ( n25740 , n25734 , n193016 );
buf ( n193018 , n25740 );
buf ( n193019 , n193018 );
and ( n25743 , n25729 , n193019 );
and ( n25744 , n192992 , n193005 );
or ( n25745 , n25743 , n25744 );
buf ( n193023 , n25745 );
buf ( n193024 , n193023 );
xor ( n25748 , n192610 , n192628 );
xor ( n25749 , n25748 , n192650 );
buf ( n193027 , n25749 );
buf ( n193028 , n193027 );
xor ( n25752 , n193024 , n193028 );
not ( n25753 , n20391 );
not ( n25754 , n25753 );
buf ( n193032 , n20396 );
not ( n25756 , n193032 );
buf ( n193034 , n25756 );
not ( n25758 , n193034 );
or ( n25759 , n25754 , n25758 );
nand ( n25760 , n25759 , n888 );
buf ( n193038 , n25760 );
buf ( n193039 , n192700 );
not ( n25763 , n193039 );
buf ( n193041 , n20554 );
not ( n25765 , n193041 );
or ( n25766 , n25763 , n25765 );
buf ( n193044 , n20558 );
buf ( n193045 , n832 );
buf ( n193046 , n886 );
xor ( n25770 , n193045 , n193046 );
buf ( n193048 , n25770 );
buf ( n193049 , n193048 );
nand ( n25773 , n193044 , n193049 );
buf ( n193051 , n25773 );
buf ( n193052 , n193051 );
nand ( n25776 , n25766 , n193052 );
buf ( n193054 , n25776 );
buf ( n193055 , n193054 );
xor ( n25779 , n193038 , n193055 );
buf ( n193057 , n192785 );
not ( n25781 , n193057 );
buf ( n193059 , n19613 );
not ( n25783 , n193059 );
or ( n25784 , n25781 , n25783 );
buf ( n193062 , n19943 );
buf ( n193063 , n836 );
buf ( n193064 , n882 );
xor ( n25788 , n193063 , n193064 );
buf ( n193066 , n25788 );
buf ( n193067 , n193066 );
nand ( n25791 , n193062 , n193067 );
buf ( n193069 , n25791 );
buf ( n193070 , n193069 );
nand ( n25794 , n25784 , n193070 );
buf ( n193072 , n25794 );
buf ( n193073 , n193072 );
xor ( n25797 , n25779 , n193073 );
buf ( n193075 , n25797 );
buf ( n193076 , n193075 );
and ( n25800 , n25752 , n193076 );
and ( n25801 , n193024 , n193028 );
or ( n25802 , n25800 , n25801 );
buf ( n193080 , n25802 );
buf ( n193081 , n193080 );
xor ( n25805 , n192987 , n193081 );
buf ( n193083 , n192926 );
not ( n25807 , n193083 );
buf ( n193085 , n192961 );
not ( n25809 , n193085 );
or ( n25810 , n25807 , n25809 );
buf ( n193088 , n192909 );
nand ( n25812 , n25810 , n193088 );
buf ( n193090 , n25812 );
buf ( n193091 , n193090 );
buf ( n193092 , n192958 );
buf ( n193093 , n192923 );
nand ( n25817 , n193092 , n193093 );
buf ( n193095 , n25817 );
buf ( n193096 , n193095 );
nand ( n25820 , n193091 , n193096 );
buf ( n193098 , n25820 );
buf ( n193099 , n193098 );
buf ( n193100 , n855 );
buf ( n193101 , n864 );
and ( n25825 , n193100 , n193101 );
buf ( n193103 , n25825 );
buf ( n193104 , n193103 );
buf ( n193105 , n25344 );
not ( n25829 , n193105 );
buf ( n193107 , n20582 );
not ( n25831 , n193107 );
or ( n25832 , n25829 , n25831 );
buf ( n193110 , n188823 );
buf ( n193111 , n25120 );
nand ( n25835 , n193110 , n193111 );
buf ( n193113 , n25835 );
buf ( n193114 , n193113 );
nand ( n25838 , n25832 , n193114 );
buf ( n193116 , n25838 );
buf ( n193117 , n193116 );
xor ( n25841 , n193104 , n193117 );
buf ( n193119 , n193066 );
not ( n25843 , n193119 );
buf ( n193121 , n19613 );
not ( n25845 , n193121 );
or ( n25846 , n25843 , n25845 );
buf ( n193124 , n19943 );
buf ( n193125 , n192210 );
nand ( n25849 , n193124 , n193125 );
buf ( n193127 , n25849 );
buf ( n193128 , n193127 );
nand ( n25852 , n25846 , n193128 );
buf ( n193130 , n25852 );
buf ( n193131 , n193130 );
xor ( n25855 , n25841 , n193131 );
buf ( n193133 , n25855 );
buf ( n193134 , n193133 );
xor ( n25858 , n193099 , n193134 );
xor ( n25859 , n193038 , n193055 );
and ( n25860 , n25859 , n193073 );
and ( n25861 , n193038 , n193055 );
or ( n25862 , n25860 , n25861 );
buf ( n193140 , n25862 );
buf ( n193141 , n193140 );
xor ( n25865 , n25858 , n193141 );
buf ( n193143 , n25865 );
buf ( n193144 , n193143 );
xor ( n25868 , n25805 , n193144 );
buf ( n193146 , n25868 );
buf ( n193147 , n193146 );
xor ( n25871 , n193024 , n193028 );
xor ( n25872 , n25871 , n193076 );
buf ( n193150 , n25872 );
buf ( n193151 , n193150 );
xor ( n25875 , n191109 , n191126 );
and ( n25876 , n25875 , n191144 );
and ( n25877 , n191109 , n191126 );
or ( n25878 , n25876 , n25877 );
buf ( n193156 , n25878 );
buf ( n193157 , n193156 );
xor ( n25881 , n192992 , n193005 );
xor ( n25882 , n25881 , n193019 );
buf ( n193160 , n25882 );
buf ( n193161 , n193160 );
xor ( n25885 , n193157 , n193161 );
and ( n25886 , n192813 , n25519 );
not ( n25887 , n192813 );
and ( n25888 , n25887 , n192792 );
or ( n25889 , n25886 , n25888 );
and ( n25890 , n25889 , n192774 );
not ( n25891 , n25889 );
and ( n25892 , n25891 , n192771 );
nor ( n25893 , n25890 , n25892 );
buf ( n193171 , n25893 );
and ( n25895 , n25885 , n193171 );
and ( n25896 , n193157 , n193161 );
or ( n25897 , n25895 , n25896 );
buf ( n193175 , n25897 );
buf ( n193176 , n193175 );
xor ( n25900 , n193151 , n193176 );
xor ( n25901 , n192968 , n25705 );
not ( n25902 , n192975 );
xor ( n25903 , n25901 , n25902 );
buf ( n193181 , n25903 );
and ( n25905 , n25900 , n193181 );
and ( n25906 , n193151 , n193176 );
or ( n25907 , n25905 , n25906 );
buf ( n193185 , n25907 );
buf ( n193186 , n193185 );
xor ( n25910 , n193147 , n193186 );
xnor ( n25911 , n192737 , n192724 );
buf ( n193189 , n25911 );
buf ( n193190 , n192751 );
buf ( n25914 , n193190 );
buf ( n193192 , n25914 );
buf ( n193193 , n193192 );
not ( n25917 , n193193 );
buf ( n193195 , n25917 );
buf ( n193196 , n193195 );
and ( n25920 , n193189 , n193196 );
not ( n25921 , n193189 );
buf ( n193199 , n193192 );
and ( n25923 , n25921 , n193199 );
nor ( n25924 , n25920 , n25923 );
buf ( n193202 , n25924 );
buf ( n193203 , n193202 );
xnor ( n25927 , n192850 , n25549 );
xor ( n25928 , n192869 , n25927 );
buf ( n193206 , n25928 );
xor ( n25930 , n193203 , n193206 );
buf ( n193208 , n190980 );
not ( n25932 , n193208 );
buf ( n193210 , n19177 );
not ( n25934 , n193210 );
or ( n25935 , n25932 , n25934 );
buf ( n193213 , n19103 );
buf ( n193214 , n192672 );
nand ( n25938 , n193213 , n193214 );
buf ( n193216 , n25938 );
buf ( n193217 , n193216 );
nand ( n25941 , n25935 , n193217 );
buf ( n193219 , n25941 );
buf ( n193220 , n193219 );
buf ( n193221 , n192706 );
not ( n25945 , n193221 );
buf ( n193223 , n25945 );
buf ( n193224 , n193223 );
xor ( n25948 , n193220 , n193224 );
buf ( n193226 , n191197 );
buf ( n193227 , n191217 );
or ( n25951 , n193226 , n193227 );
buf ( n193229 , n191238 );
nand ( n25953 , n25951 , n193229 );
buf ( n193231 , n25953 );
buf ( n193232 , n193231 );
buf ( n193233 , n191197 );
buf ( n193234 , n191217 );
nand ( n25958 , n193233 , n193234 );
buf ( n193236 , n25958 );
buf ( n193237 , n193236 );
nand ( n25961 , n193232 , n193237 );
buf ( n193239 , n25961 );
buf ( n193240 , n193239 );
xor ( n25964 , n25948 , n193240 );
buf ( n193242 , n25964 );
buf ( n193243 , n193242 );
and ( n25967 , n25930 , n193243 );
and ( n25968 , n193203 , n193206 );
or ( n25969 , n25967 , n25968 );
buf ( n193247 , n25969 );
buf ( n193248 , n193247 );
xor ( n25972 , n190793 , n190808 );
and ( n25973 , n25972 , n190852 );
and ( n25974 , n190793 , n190808 );
or ( n25975 , n25973 , n25974 );
buf ( n193253 , n25975 );
buf ( n193254 , n193253 );
not ( n25978 , n23613 );
not ( n25979 , n190932 );
or ( n25980 , n25978 , n25979 );
not ( n25981 , n23659 );
not ( n25982 , n23656 );
or ( n25983 , n25981 , n25982 );
nand ( n25984 , n25983 , n23710 );
nand ( n25985 , n25980 , n25984 );
buf ( n193263 , n25985 );
xor ( n25987 , n193254 , n193263 );
not ( n25988 , n23875 );
not ( n25989 , n23885 );
or ( n25990 , n25988 , n25989 );
not ( n25991 , n23874 );
and ( n25992 , n23876 , n191161 , n890 );
not ( n25993 , n25992 );
or ( n25994 , n25991 , n25993 );
nand ( n25995 , n25994 , n23902 );
nand ( n25996 , n25990 , n25995 );
buf ( n193274 , n25996 );
or ( n25998 , n191299 , n191282 );
nand ( n25999 , n25998 , n191266 );
buf ( n193277 , n191299 );
buf ( n193278 , n191282 );
nand ( n26002 , n193277 , n193278 );
buf ( n193280 , n26002 );
nand ( n26004 , n25999 , n193280 );
buf ( n193282 , n26004 );
xor ( n26006 , n193274 , n193282 );
not ( n26007 , n190954 );
nand ( n26008 , n26007 , n23694 );
nand ( n26009 , n23708 , n26008 );
not ( n26010 , n23694 );
nand ( n26011 , n26010 , n190954 );
nand ( n26012 , n26009 , n26011 );
buf ( n193290 , n26012 );
xor ( n26014 , n26006 , n193290 );
buf ( n193292 , n26014 );
buf ( n193293 , n193292 );
and ( n26017 , n25987 , n193293 );
and ( n26018 , n193254 , n193263 );
or ( n26019 , n26017 , n26018 );
buf ( n193297 , n26019 );
buf ( n193298 , n193297 );
xor ( n26022 , n193248 , n193298 );
xor ( n26023 , n193220 , n193224 );
and ( n26024 , n26023 , n193240 );
and ( n26025 , n193220 , n193224 );
or ( n26026 , n26024 , n26025 );
buf ( n193304 , n26026 );
buf ( n193305 , n193304 );
xor ( n26029 , n193274 , n193282 );
and ( n26030 , n26029 , n193290 );
and ( n26031 , n193274 , n193282 );
or ( n26032 , n26030 , n26031 );
buf ( n193310 , n26032 );
buf ( n193311 , n193310 );
xor ( n26035 , n193305 , n193311 );
xor ( n26036 , n192763 , n192820 );
xor ( n26037 , n26036 , n192881 );
buf ( n193315 , n26037 );
buf ( n193316 , n193315 );
xor ( n26040 , n26035 , n193316 );
buf ( n193318 , n26040 );
buf ( n193319 , n193318 );
and ( n26043 , n26022 , n193319 );
and ( n26044 , n193248 , n193298 );
or ( n26045 , n26043 , n26044 );
buf ( n193323 , n26045 );
buf ( n193324 , n193323 );
and ( n26048 , n25910 , n193324 );
and ( n26049 , n193147 , n193186 );
or ( n26050 , n26048 , n26049 );
buf ( n193328 , n26050 );
buf ( n193329 , n193328 );
xor ( n26053 , n192897 , n193329 );
xor ( n26054 , n192987 , n193081 );
and ( n26055 , n26054 , n193144 );
and ( n26056 , n192987 , n193081 );
or ( n26057 , n26055 , n26056 );
buf ( n193335 , n26057 );
buf ( n193336 , n193335 );
xor ( n26060 , n193099 , n193134 );
and ( n26061 , n26060 , n193141 );
and ( n26062 , n193099 , n193134 );
or ( n26063 , n26061 , n26062 );
buf ( n193341 , n26063 );
buf ( n193342 , n193341 );
buf ( n193343 , n192682 );
not ( n26067 , n193343 );
buf ( n193345 , n19177 );
not ( n26069 , n193345 );
or ( n26070 , n26067 , n26069 );
buf ( n193348 , n20279 );
buf ( n193349 , n192376 );
nand ( n26073 , n193348 , n193349 );
buf ( n193351 , n26073 );
buf ( n193352 , n193351 );
nand ( n26076 , n26070 , n193352 );
buf ( n193354 , n26076 );
buf ( n193355 , n192952 );
not ( n26079 , n193355 );
buf ( n193357 , n20335 );
not ( n26081 , n193357 );
or ( n26082 , n26079 , n26081 );
buf ( n193360 , n186337 );
buf ( n193361 , n192354 );
nand ( n26085 , n193360 , n193361 );
buf ( n193363 , n26085 );
buf ( n193364 , n193363 );
nand ( n26088 , n26082 , n193364 );
buf ( n193366 , n26088 );
or ( n26090 , n193354 , n193366 );
buf ( n193368 , n193048 );
not ( n26092 , n193368 );
buf ( n193370 , n20554 );
not ( n26094 , n193370 );
or ( n26095 , n26092 , n26094 );
buf ( n193373 , n20558 );
buf ( n193374 , n886 );
nand ( n26098 , n193373 , n193374 );
buf ( n193376 , n26098 );
buf ( n193377 , n193376 );
nand ( n26101 , n26095 , n193377 );
buf ( n193379 , n26101 );
nand ( n26103 , n26090 , n193379 );
buf ( n193381 , n192682 );
not ( n26105 , n193381 );
buf ( n193383 , n19098 );
not ( n26107 , n193383 );
or ( n26108 , n26105 , n26107 );
buf ( n193386 , n193351 );
nand ( n26110 , n26108 , n193386 );
buf ( n193388 , n26110 );
buf ( n193389 , n193388 );
buf ( n193390 , n193366 );
nand ( n26114 , n193389 , n193390 );
buf ( n193392 , n26114 );
nand ( n26116 , n26103 , n193392 );
buf ( n193394 , n26116 );
xor ( n26118 , n193104 , n193117 );
and ( n26119 , n26118 , n193131 );
and ( n26120 , n193104 , n193117 );
or ( n26121 , n26119 , n26120 );
buf ( n193399 , n26121 );
buf ( n193400 , n193399 );
xor ( n26124 , n193394 , n193400 );
buf ( n193402 , n192643 );
not ( n26126 , n193402 );
buf ( n193404 , n186924 );
not ( n26128 , n193404 );
or ( n26129 , n26126 , n26128 );
buf ( n193407 , n18875 );
buf ( n193408 , n192311 );
nand ( n26132 , n193407 , n193408 );
buf ( n193410 , n26132 );
buf ( n193411 , n193410 );
nand ( n26135 , n26129 , n193411 );
buf ( n193413 , n26135 );
buf ( n193414 , n192603 );
not ( n26138 , n193414 );
buf ( n193416 , n19260 );
not ( n26140 , n193416 );
or ( n26141 , n26138 , n26140 );
buf ( n193419 , n19265 );
buf ( n193420 , n192256 );
nand ( n26144 , n193419 , n193420 );
buf ( n193422 , n26144 );
buf ( n193423 , n193422 );
nand ( n26147 , n26141 , n193423 );
buf ( n193425 , n26147 );
xor ( n26149 , n193413 , n193425 );
buf ( n193427 , n192541 );
not ( n26151 , n193427 );
buf ( n193429 , n186435 );
not ( n26153 , n193429 );
or ( n26154 , n26151 , n26153 );
buf ( n193432 , n186444 );
buf ( n193433 , n192235 );
nand ( n26157 , n193432 , n193433 );
buf ( n193435 , n26157 );
buf ( n193436 , n193435 );
nand ( n26160 , n26154 , n193436 );
buf ( n193438 , n26160 );
and ( n26162 , n26149 , n193438 );
and ( n26163 , n193413 , n193425 );
or ( n26164 , n26162 , n26163 );
buf ( n193442 , n26164 );
xor ( n26166 , n26124 , n193442 );
buf ( n193444 , n26166 );
buf ( n193445 , n193444 );
xor ( n26169 , n193342 , n193445 );
xor ( n26170 , n193379 , n193388 );
buf ( n193448 , n26170 );
buf ( n193449 , n193366 );
xor ( n26173 , n193448 , n193449 );
buf ( n193451 , n26173 );
buf ( n193452 , n193451 );
xor ( n26176 , n192465 , n192448 );
and ( n26177 , n26176 , n192487 );
not ( n26178 , n26176 );
and ( n26179 , n26178 , n192490 );
nor ( n26180 , n26177 , n26179 );
buf ( n193458 , n26180 );
xor ( n26182 , n193452 , n193458 );
xor ( n26183 , n193413 , n193425 );
xor ( n26184 , n26183 , n193438 );
buf ( n193462 , n26184 );
and ( n26186 , n26182 , n193462 );
and ( n26187 , n193452 , n193458 );
or ( n26188 , n26186 , n26187 );
buf ( n193466 , n26188 );
buf ( n193467 , n193466 );
xor ( n26191 , n26169 , n193467 );
buf ( n193469 , n26191 );
buf ( n193470 , n193469 );
xor ( n26194 , n193336 , n193470 );
xor ( n26195 , n193452 , n193458 );
xor ( n26196 , n26195 , n193462 );
buf ( n193474 , n26196 );
xor ( n26198 , n192712 , n192886 );
xor ( n26199 , n26198 , n192891 );
buf ( n193477 , n26199 );
nand ( n26201 , n193474 , n193477 );
xor ( n26202 , n193305 , n193311 );
and ( n26203 , n26202 , n193316 );
and ( n26204 , n193305 , n193311 );
or ( n26205 , n26203 , n26204 );
buf ( n193483 , n26205 );
nand ( n26207 , n193474 , n193483 );
nand ( n26208 , n193477 , n193483 );
nand ( n26209 , n26201 , n26207 , n26208 );
buf ( n193487 , n26209 );
xor ( n26211 , n26194 , n193487 );
buf ( n193489 , n26211 );
buf ( n193490 , n193489 );
xor ( n26214 , n26053 , n193490 );
buf ( n193492 , n26214 );
buf ( n26216 , n193492 );
xor ( n26217 , n186765 , n186783 );
and ( n26218 , n26217 , n186803 );
and ( n26219 , n186765 , n186783 );
or ( n26220 , n26218 , n26219 );
buf ( n193498 , n26220 );
buf ( n193499 , n193498 );
xor ( n26223 , n186609 , n186657 );
and ( n26224 , n26223 , n186705 );
and ( n26225 , n186609 , n186657 );
or ( n26226 , n26224 , n26225 );
buf ( n193504 , n26226 );
buf ( n193505 , n193504 );
xor ( n26229 , n193499 , n193505 );
buf ( n193507 , n186799 );
xor ( n26231 , n186716 , n186730 );
and ( n26232 , n26231 , n186745 );
and ( n26233 , n186716 , n186730 );
or ( n26234 , n26232 , n26233 );
buf ( n193512 , n26234 );
buf ( n193513 , n193512 );
xor ( n26237 , n193507 , n193513 );
xor ( n26238 , n186821 , n186835 );
and ( n26239 , n26238 , n186850 );
and ( n26240 , n186821 , n186835 );
or ( n26241 , n26239 , n26240 );
buf ( n193519 , n26241 );
buf ( n193520 , n193519 );
xor ( n26244 , n26237 , n193520 );
buf ( n193522 , n26244 );
buf ( n193523 , n193522 );
xor ( n26247 , n26229 , n193523 );
buf ( n193525 , n26247 );
buf ( n193526 , n193525 );
xor ( n26250 , n186748 , n186806 );
and ( n26251 , n26250 , n186853 );
and ( n26252 , n186748 , n186806 );
or ( n26253 , n26251 , n26252 );
buf ( n193531 , n26253 );
buf ( n193532 , n193531 );
buf ( n193533 , n846 );
buf ( n193534 , n864 );
and ( n26258 , n193533 , n193534 );
buf ( n193536 , n26258 );
buf ( n193537 , n193536 );
buf ( n193538 , n19446 );
not ( n26262 , n193538 );
buf ( n193540 , n186640 );
not ( n26264 , n193540 );
or ( n26265 , n26262 , n26264 );
buf ( n193543 , n186340 );
buf ( n193544 , n864 );
buf ( n193545 , n844 );
xor ( n26269 , n193544 , n193545 );
buf ( n193547 , n26269 );
buf ( n193548 , n193547 );
nand ( n26272 , n193543 , n193548 );
buf ( n193550 , n26272 );
buf ( n193551 , n193550 );
nand ( n26275 , n26265 , n193551 );
buf ( n193553 , n26275 );
buf ( n193554 , n193553 );
xor ( n26278 , n193537 , n193554 );
buf ( n193556 , n19537 );
not ( n26280 , n193556 );
buf ( n193558 , n186435 );
not ( n26282 , n193558 );
or ( n26283 , n26280 , n26282 );
buf ( n193561 , n186444 );
buf ( n193562 , n838 );
buf ( n193563 , n870 );
xor ( n26287 , n193562 , n193563 );
buf ( n193565 , n26287 );
buf ( n193566 , n193565 );
nand ( n26290 , n193561 , n193566 );
buf ( n193568 , n26290 );
buf ( n193569 , n193568 );
nand ( n26293 , n26283 , n193569 );
buf ( n193571 , n26293 );
buf ( n193572 , n193571 );
xor ( n26296 , n26278 , n193572 );
buf ( n193574 , n26296 );
buf ( n193575 , n193574 );
buf ( n193576 , n186758 );
not ( n26300 , n193576 );
buf ( n193578 , n186241 );
not ( n26302 , n193578 );
or ( n26303 , n26300 , n26302 );
buf ( n193581 , n186254 );
buf ( n193582 , n842 );
buf ( n193583 , n866 );
xor ( n26307 , n193582 , n193583 );
buf ( n193585 , n26307 );
buf ( n193586 , n193585 );
nand ( n26310 , n193581 , n193586 );
buf ( n193588 , n26310 );
buf ( n193589 , n193588 );
nand ( n26313 , n26303 , n193589 );
buf ( n193591 , n26313 );
buf ( n193592 , n193591 );
buf ( n193593 , n19551 );
not ( n26317 , n193593 );
buf ( n193595 , n186287 );
not ( n26319 , n193595 );
or ( n26320 , n26317 , n26319 );
buf ( n193598 , n186297 );
buf ( n193599 , n834 );
buf ( n193600 , n874 );
xor ( n26324 , n193599 , n193600 );
buf ( n193602 , n26324 );
buf ( n193603 , n193602 );
nand ( n26327 , n193598 , n193603 );
buf ( n193605 , n26327 );
buf ( n193606 , n193605 );
nand ( n26330 , n26320 , n193606 );
buf ( n193608 , n26330 );
buf ( n193609 , n193608 );
xor ( n26333 , n193592 , n193609 );
buf ( n193611 , n186776 );
not ( n26335 , n193611 );
buf ( n193613 , n186197 );
not ( n26337 , n193613 );
or ( n26338 , n26335 , n26337 );
buf ( n193616 , n186208 );
buf ( n193617 , n840 );
buf ( n193618 , n868 );
xor ( n26342 , n193617 , n193618 );
buf ( n193620 , n26342 );
buf ( n193621 , n193620 );
nand ( n26345 , n193616 , n193621 );
buf ( n193623 , n26345 );
buf ( n193624 , n193623 );
nand ( n26348 , n26338 , n193624 );
buf ( n193626 , n26348 );
buf ( n193627 , n193626 );
xor ( n26351 , n26333 , n193627 );
buf ( n193629 , n26351 );
buf ( n193630 , n193629 );
xor ( n26354 , n193575 , n193630 );
buf ( n193632 , n19461 );
not ( n26356 , n193632 );
buf ( n193634 , n19260 );
not ( n26358 , n193634 );
or ( n26359 , n26356 , n26358 );
buf ( n193637 , n19265 );
xor ( n26361 , n872 , n836 );
buf ( n193639 , n26361 );
nand ( n26363 , n193637 , n193639 );
buf ( n193641 , n26363 );
buf ( n193642 , n193641 );
nand ( n26366 , n26359 , n193642 );
buf ( n193644 , n26366 );
buf ( n193645 , n19566 );
not ( n26369 , n193645 );
buf ( n193647 , n19177 );
not ( n26371 , n193647 );
or ( n26372 , n26369 , n26371 );
buf ( n193650 , n186395 );
xor ( n26374 , n876 , n832 );
buf ( n193652 , n26374 );
nand ( n26376 , n193650 , n193652 );
buf ( n193654 , n26376 );
buf ( n193655 , n193654 );
nand ( n26379 , n26372 , n193655 );
buf ( n193657 , n26379 );
xor ( n26381 , n193644 , n193657 );
buf ( n193659 , n186789 );
buf ( n193660 , n186575 );
or ( n26384 , n193659 , n193660 );
buf ( n193662 , n878 );
nand ( n26386 , n26384 , n193662 );
buf ( n193664 , n26386 );
xor ( n26388 , n26381 , n193664 );
buf ( n193666 , n26388 );
xor ( n26390 , n26354 , n193666 );
buf ( n193668 , n26390 );
buf ( n193669 , n193668 );
xor ( n26393 , n193532 , n193669 );
xor ( n26394 , n186366 , n186593 );
and ( n26395 , n26394 , n186708 );
and ( n26396 , n186366 , n186593 );
or ( n26397 , n26395 , n26396 );
buf ( n193675 , n26397 );
buf ( n193676 , n193675 );
xor ( n26400 , n26393 , n193676 );
buf ( n193678 , n26400 );
buf ( n193679 , n193678 );
xor ( n26403 , n193526 , n193679 );
xor ( n26404 , n186856 , n186874 );
and ( n26405 , n26404 , n187087 );
and ( n26406 , n186856 , n186874 );
or ( n26407 , n26405 , n26406 );
buf ( n193685 , n26407 );
buf ( n193686 , n193685 );
xor ( n26410 , n26403 , n193686 );
buf ( n193688 , n26410 );
buf ( n26412 , n193688 );
xor ( n26413 , n192897 , n193329 );
and ( n26414 , n26413 , n193490 );
and ( n26415 , n192897 , n193329 );
or ( n26416 , n26414 , n26415 );
buf ( n193694 , n26416 );
buf ( n26418 , n193694 );
buf ( n193696 , n856 );
buf ( n193697 , n886 );
xor ( n26421 , n193696 , n193697 );
buf ( n193699 , n26421 );
not ( n26423 , n193699 );
not ( n26424 , n20554 );
or ( n26425 , n26423 , n26424 );
buf ( n193703 , n855 );
buf ( n193704 , n886 );
xor ( n26428 , n193703 , n193704 );
buf ( n193706 , n26428 );
nand ( n26430 , n20558 , n193706 );
nand ( n26431 , n26425 , n26430 );
buf ( n193709 , n862 );
buf ( n193710 , n880 );
xor ( n26434 , n193709 , n193710 );
buf ( n193712 , n26434 );
buf ( n193713 , n193712 );
not ( n26437 , n193713 );
buf ( n193715 , n186924 );
not ( n26439 , n193715 );
or ( n26440 , n26437 , n26439 );
buf ( n193718 , n18875 );
buf ( n193719 , n861 );
buf ( n193720 , n880 );
xor ( n26444 , n193719 , n193720 );
buf ( n193722 , n26444 );
buf ( n193723 , n193722 );
nand ( n26447 , n193718 , n193723 );
buf ( n193725 , n26447 );
buf ( n193726 , n193725 );
nand ( n26450 , n26440 , n193726 );
buf ( n193728 , n26450 );
xor ( n26452 , n26431 , n193728 );
buf ( n193730 , n854 );
buf ( n193731 , n888 );
xor ( n26455 , n193730 , n193731 );
buf ( n193733 , n26455 );
buf ( n193734 , n193733 );
not ( n26458 , n193734 );
buf ( n193736 , n20391 );
not ( n26460 , n193736 );
or ( n26461 , n26458 , n26460 );
buf ( n193739 , n20396 );
buf ( n193740 , n853 );
buf ( n193741 , n888 );
xor ( n26465 , n193740 , n193741 );
buf ( n193743 , n26465 );
buf ( n193744 , n193743 );
nand ( n26468 , n193739 , n193744 );
buf ( n193746 , n26468 );
buf ( n193747 , n193746 );
nand ( n26471 , n26461 , n193747 );
buf ( n193749 , n26471 );
xor ( n26473 , n26452 , n193749 );
buf ( n193751 , n850 );
buf ( n193752 , n892 );
xor ( n26476 , n193751 , n193752 );
buf ( n193754 , n26476 );
buf ( n193755 , n193754 );
not ( n26479 , n193755 );
buf ( n193757 , n190485 );
not ( n26481 , n193757 );
or ( n26482 , n26479 , n26481 );
buf ( n193760 , n190128 );
buf ( n193761 , n849 );
buf ( n193762 , n892 );
xor ( n26486 , n193761 , n193762 );
buf ( n193764 , n26486 );
buf ( n193765 , n193764 );
nand ( n26489 , n193760 , n193765 );
buf ( n193767 , n26489 );
buf ( n193768 , n193767 );
nand ( n26492 , n26482 , n193768 );
buf ( n193770 , n26492 );
not ( n26494 , n21330 );
buf ( n193772 , n848 );
buf ( n193773 , n894 );
xor ( n26497 , n193772 , n193773 );
buf ( n193775 , n26497 );
not ( n26499 , n193775 );
or ( n26500 , n26494 , n26499 );
buf ( n193778 , n847 );
buf ( n193779 , n894 );
xor ( n26503 , n193778 , n193779 );
buf ( n193781 , n26503 );
buf ( n193782 , n193781 );
buf ( n193783 , n895 );
nand ( n26507 , n193782 , n193783 );
buf ( n193785 , n26507 );
nand ( n26509 , n26500 , n193785 );
not ( n26510 , n26509 );
nand ( n26511 , n863 , n186575 );
and ( n26512 , n26510 , n26511 );
not ( n26513 , n26510 );
nand ( n26514 , n186575 , n863 );
not ( n26515 , n26514 );
and ( n26516 , n26513 , n26515 );
nor ( n26517 , n26512 , n26516 );
xor ( n26518 , n193770 , n26517 );
buf ( n26519 , n26518 );
buf ( n193797 , n852 );
buf ( n193798 , n890 );
xor ( n26522 , n193797 , n193798 );
buf ( n193800 , n26522 );
buf ( n193801 , n193800 );
not ( n26525 , n193801 );
buf ( n193803 , n188751 );
not ( n26527 , n193803 );
or ( n26528 , n26525 , n26527 );
buf ( n193806 , n20902 );
buf ( n193807 , n851 );
buf ( n193808 , n890 );
xor ( n26532 , n193807 , n193808 );
buf ( n193810 , n26532 );
buf ( n193811 , n193810 );
nand ( n26535 , n193806 , n193811 );
buf ( n193813 , n26535 );
buf ( n193814 , n193813 );
nand ( n26538 , n26528 , n193814 );
buf ( n193816 , n26538 );
buf ( n193817 , n858 );
buf ( n193818 , n884 );
xor ( n26542 , n193817 , n193818 );
buf ( n193820 , n26542 );
buf ( n193821 , n193820 );
not ( n26545 , n193821 );
buf ( n193823 , n192332 );
not ( n26547 , n193823 );
or ( n26548 , n26545 , n26547 );
buf ( n193826 , n190543 );
buf ( n193827 , n857 );
buf ( n193828 , n884 );
xor ( n26552 , n193827 , n193828 );
buf ( n193830 , n26552 );
buf ( n193831 , n193830 );
nand ( n26555 , n193826 , n193831 );
buf ( n193833 , n26555 );
buf ( n193834 , n193833 );
nand ( n26558 , n26548 , n193834 );
buf ( n193836 , n26558 );
xor ( n26560 , n193816 , n193836 );
buf ( n193838 , n860 );
buf ( n193839 , n882 );
xor ( n26563 , n193838 , n193839 );
buf ( n193841 , n26563 );
buf ( n193842 , n193841 );
not ( n26566 , n193842 );
buf ( n26567 , n19613 );
buf ( n193845 , n26567 );
not ( n26569 , n193845 );
or ( n26570 , n26566 , n26569 );
not ( n26571 , n19602 );
buf ( n193849 , n26571 );
buf ( n193850 , n859 );
buf ( n193851 , n882 );
xor ( n26575 , n193850 , n193851 );
buf ( n193853 , n26575 );
buf ( n193854 , n193853 );
nand ( n26578 , n193849 , n193854 );
buf ( n193856 , n26578 );
buf ( n193857 , n193856 );
nand ( n26581 , n26570 , n193857 );
buf ( n193859 , n26581 );
xor ( n26583 , n26560 , n193859 );
nand ( n26584 , n26473 , n26519 , n26583 );
not ( n26585 , n26519 );
not ( n26586 , n26583 );
nand ( n26587 , n26585 , n26586 );
not ( n26588 , n26587 );
nand ( n26589 , n26588 , n26473 );
not ( n26590 , n26473 );
not ( n26591 , n26583 );
nor ( n26592 , n26591 , n26519 );
nand ( n26593 , n26590 , n26592 );
nand ( n26594 , n26590 , n26519 , n26586 );
nand ( n26595 , n26584 , n26589 , n26593 , n26594 );
buf ( n193873 , n26595 );
buf ( n193874 , n851 );
buf ( n193875 , n894 );
xor ( n26599 , n193874 , n193875 );
buf ( n193877 , n26599 );
buf ( n193878 , n193877 );
not ( n26602 , n193878 );
buf ( n193880 , n23321 );
not ( n26604 , n193880 );
or ( n26605 , n26602 , n26604 );
buf ( n193883 , n850 );
buf ( n193884 , n894 );
xor ( n26608 , n193883 , n193884 );
buf ( n193886 , n26608 );
buf ( n193887 , n193886 );
buf ( n193888 , n895 );
nand ( n26612 , n193887 , n193888 );
buf ( n193890 , n26612 );
buf ( n193891 , n193890 );
nand ( n26615 , n26605 , n193891 );
buf ( n193893 , n26615 );
buf ( n193894 , n193893 );
buf ( n193895 , n863 );
buf ( n193896 , n883 );
or ( n26620 , n193895 , n193896 );
buf ( n193898 , n884 );
nand ( n26622 , n26620 , n193898 );
buf ( n193900 , n26622 );
buf ( n193901 , n863 );
buf ( n193902 , n883 );
nand ( n26626 , n193901 , n193902 );
buf ( n193904 , n26626 );
and ( n26628 , n193900 , n193904 , n882 );
buf ( n193906 , n26628 );
and ( n26630 , n193894 , n193906 );
buf ( n193908 , n26630 );
buf ( n193909 , n193908 );
xor ( n26633 , n882 , n862 );
buf ( n193911 , n26633 );
not ( n26635 , n193911 );
buf ( n193913 , n19613 );
not ( n26637 , n193913 );
or ( n26638 , n26635 , n26637 );
buf ( n193916 , n19943 );
buf ( n193917 , n861 );
buf ( n193918 , n882 );
xor ( n26642 , n193917 , n193918 );
buf ( n193920 , n26642 );
buf ( n193921 , n193920 );
nand ( n26645 , n193916 , n193921 );
buf ( n193923 , n26645 );
buf ( n193924 , n193923 );
nand ( n26648 , n26638 , n193924 );
buf ( n193926 , n26648 );
buf ( n193927 , n193926 );
xor ( n26651 , n193909 , n193927 );
xor ( n26652 , n884 , n860 );
buf ( n193930 , n26652 );
not ( n26654 , n193930 );
buf ( n193932 , n192332 );
not ( n26656 , n193932 );
or ( n26657 , n26654 , n26656 );
buf ( n193935 , n192573 );
buf ( n193936 , n859 );
buf ( n193937 , n884 );
xor ( n26661 , n193936 , n193937 );
buf ( n193939 , n26661 );
buf ( n193940 , n193939 );
nand ( n26664 , n193935 , n193940 );
buf ( n193942 , n26664 );
buf ( n193943 , n193942 );
nand ( n26667 , n26657 , n193943 );
buf ( n193945 , n26667 );
buf ( n193946 , n193945 );
and ( n26670 , n26651 , n193946 );
and ( n26671 , n193909 , n193927 );
or ( n26672 , n26670 , n26671 );
buf ( n193950 , n26672 );
buf ( n193951 , n193950 );
buf ( n193952 , n193920 );
not ( n26676 , n193952 );
buf ( n193954 , n26567 );
not ( n26678 , n193954 );
or ( n26679 , n26676 , n26678 );
buf ( n193957 , n19943 );
buf ( n193958 , n193841 );
nand ( n26682 , n193957 , n193958 );
buf ( n193960 , n26682 );
buf ( n193961 , n193960 );
nand ( n26685 , n26679 , n193961 );
buf ( n193963 , n26685 );
buf ( n193964 , n193963 );
buf ( n193965 , n863 );
buf ( n193966 , n881 );
or ( n26690 , n193965 , n193966 );
buf ( n193968 , n882 );
nand ( n26692 , n26690 , n193968 );
buf ( n193970 , n26692 );
buf ( n193971 , n193970 );
buf ( n193972 , n863 );
buf ( n193973 , n881 );
nand ( n26697 , n193972 , n193973 );
buf ( n193975 , n26697 );
buf ( n193976 , n193975 );
buf ( n193977 , n880 );
and ( n26701 , n193971 , n193976 , n193977 );
buf ( n193979 , n26701 );
buf ( n193980 , n193979 );
buf ( n193981 , n849 );
buf ( n193982 , n894 );
xor ( n26706 , n193981 , n193982 );
buf ( n193984 , n26706 );
buf ( n193985 , n193984 );
not ( n26709 , n193985 );
buf ( n193987 , n21330 );
not ( n26711 , n193987 );
or ( n26712 , n26709 , n26711 );
buf ( n193990 , n193775 );
buf ( n193991 , n895 );
nand ( n26715 , n193990 , n193991 );
buf ( n193993 , n26715 );
buf ( n193994 , n193993 );
nand ( n26718 , n26712 , n193994 );
buf ( n193996 , n26718 );
buf ( n193997 , n193996 );
xor ( n26721 , n193980 , n193997 );
buf ( n193999 , n26721 );
buf ( n194000 , n193999 );
xor ( n26724 , n193964 , n194000 );
buf ( n194002 , n20358 );
buf ( n194003 , n863 );
and ( n26727 , n194002 , n194003 );
buf ( n194005 , n26727 );
buf ( n194006 , n194005 );
buf ( n194007 , n193886 );
not ( n26731 , n194007 );
buf ( n194009 , n21330 );
not ( n26733 , n194009 );
or ( n26734 , n26731 , n26733 );
buf ( n194012 , n193984 );
buf ( n194013 , n895 );
nand ( n26737 , n194012 , n194013 );
buf ( n194015 , n26737 );
buf ( n194016 , n194015 );
nand ( n26740 , n26734 , n194016 );
buf ( n194018 , n26740 );
buf ( n194019 , n194018 );
xor ( n26743 , n194006 , n194019 );
buf ( n194021 , n852 );
buf ( n194022 , n892 );
xor ( n26746 , n194021 , n194022 );
buf ( n194024 , n26746 );
buf ( n194025 , n194024 );
not ( n26749 , n194025 );
buf ( n194027 , n190485 );
not ( n26751 , n194027 );
or ( n26752 , n26749 , n26751 );
buf ( n194030 , n190128 );
buf ( n194031 , n851 );
buf ( n194032 , n892 );
xor ( n26756 , n194031 , n194032 );
buf ( n194034 , n26756 );
buf ( n194035 , n194034 );
nand ( n26759 , n194030 , n194035 );
buf ( n194037 , n26759 );
buf ( n194038 , n194037 );
nand ( n26762 , n26752 , n194038 );
buf ( n194040 , n26762 );
buf ( n194041 , n194040 );
and ( n26765 , n26743 , n194041 );
and ( n26766 , n194006 , n194019 );
or ( n26767 , n26765 , n26766 );
buf ( n194045 , n26767 );
buf ( n194046 , n194045 );
xor ( n26770 , n26724 , n194046 );
buf ( n194048 , n26770 );
buf ( n194049 , n194048 );
xor ( n26773 , n193951 , n194049 );
xor ( n26774 , n194006 , n194019 );
xor ( n26775 , n26774 , n194041 );
buf ( n194053 , n26775 );
buf ( n194054 , n194053 );
buf ( n194055 , n857 );
buf ( n194056 , n888 );
xor ( n26780 , n194055 , n194056 );
buf ( n194058 , n26780 );
buf ( n194059 , n194058 );
not ( n26783 , n194059 );
buf ( n194061 , n20391 );
not ( n26785 , n194061 );
or ( n26786 , n26783 , n26785 );
buf ( n194064 , n20396 );
buf ( n194065 , n856 );
buf ( n194066 , n888 );
xor ( n26790 , n194065 , n194066 );
buf ( n194068 , n26790 );
buf ( n194069 , n194068 );
nand ( n26793 , n194064 , n194069 );
buf ( n194071 , n26793 );
buf ( n194072 , n194071 );
nand ( n26796 , n26786 , n194072 );
buf ( n194074 , n26796 );
buf ( n194075 , n194074 );
not ( n26799 , n194075 );
buf ( n194077 , n859 );
buf ( n194078 , n886 );
xor ( n26802 , n194077 , n194078 );
buf ( n194080 , n26802 );
buf ( n194081 , n194080 );
not ( n26805 , n194081 );
buf ( n194083 , n20554 );
not ( n26807 , n194083 );
or ( n26808 , n26805 , n26807 );
buf ( n194086 , n20558 );
buf ( n194087 , n858 );
buf ( n194088 , n886 );
xor ( n26812 , n194087 , n194088 );
buf ( n194090 , n26812 );
buf ( n194091 , n194090 );
nand ( n26815 , n194086 , n194091 );
buf ( n194093 , n26815 );
buf ( n194094 , n194093 );
nand ( n26818 , n26808 , n194094 );
buf ( n194096 , n26818 );
buf ( n194097 , n194096 );
not ( n26821 , n194097 );
or ( n26822 , n26799 , n26821 );
buf ( n194100 , n194096 );
buf ( n194101 , n194074 );
or ( n26825 , n194100 , n194101 );
xor ( n26826 , n892 , n853 );
buf ( n194104 , n26826 );
not ( n26828 , n194104 );
buf ( n194106 , n190485 );
not ( n26830 , n194106 );
or ( n26831 , n26828 , n26830 );
buf ( n194109 , n190491 );
buf ( n194110 , n194024 );
nand ( n26834 , n194109 , n194110 );
buf ( n194112 , n26834 );
buf ( n194113 , n194112 );
nand ( n26837 , n26831 , n194113 );
buf ( n194115 , n26837 );
buf ( n194116 , n194115 );
nand ( n26840 , n26825 , n194116 );
buf ( n194118 , n26840 );
buf ( n194119 , n194118 );
nand ( n26843 , n26822 , n194119 );
buf ( n194121 , n26843 );
buf ( n194122 , n194121 );
xor ( n26846 , n194054 , n194122 );
xor ( n26847 , n882 , n863 );
buf ( n194125 , n26847 );
not ( n26849 , n194125 );
buf ( n194127 , n19613 );
not ( n26851 , n194127 );
or ( n26852 , n26849 , n26851 );
buf ( n194130 , n19943 );
buf ( n194131 , n26633 );
nand ( n26855 , n194130 , n194131 );
buf ( n194133 , n26855 );
buf ( n194134 , n194133 );
nand ( n26858 , n26852 , n194134 );
buf ( n194136 , n26858 );
buf ( n194137 , n194136 );
buf ( n194138 , n855 );
buf ( n194139 , n890 );
xor ( n26863 , n194138 , n194139 );
buf ( n194141 , n26863 );
buf ( n194142 , n194141 );
not ( n26866 , n194142 );
buf ( n194144 , n188751 );
not ( n26868 , n194144 );
or ( n26869 , n26866 , n26868 );
buf ( n194147 , n20902 );
xor ( n26871 , n890 , n854 );
buf ( n194149 , n26871 );
nand ( n26873 , n194147 , n194149 );
buf ( n194151 , n26873 );
buf ( n194152 , n194151 );
nand ( n26876 , n26869 , n194152 );
buf ( n194154 , n26876 );
buf ( n194155 , n194154 );
xor ( n26879 , n194137 , n194155 );
xor ( n26880 , n884 , n861 );
buf ( n194158 , n26880 );
not ( n26882 , n194158 );
buf ( n194160 , n192332 );
not ( n26884 , n194160 );
or ( n26885 , n26882 , n26884 );
buf ( n194163 , n192573 );
buf ( n194164 , n26652 );
nand ( n26888 , n194163 , n194164 );
buf ( n194166 , n26888 );
buf ( n194167 , n194166 );
nand ( n26891 , n26885 , n194167 );
buf ( n194169 , n26891 );
buf ( n194170 , n194169 );
and ( n26894 , n26879 , n194170 );
and ( n26895 , n194137 , n194155 );
or ( n26896 , n26894 , n26895 );
buf ( n194174 , n26896 );
buf ( n194175 , n194174 );
and ( n26899 , n26846 , n194175 );
and ( n26900 , n194054 , n194122 );
or ( n26901 , n26899 , n26900 );
buf ( n194179 , n26901 );
buf ( n194180 , n194179 );
and ( n26904 , n26773 , n194180 );
and ( n26905 , n193951 , n194049 );
or ( n26906 , n26904 , n26905 );
buf ( n194184 , n26906 );
buf ( n194185 , n194184 );
xor ( n26909 , n193873 , n194185 );
xor ( n26910 , n193964 , n194000 );
and ( n26911 , n26910 , n194046 );
and ( n26912 , n193964 , n194000 );
or ( n26913 , n26911 , n26912 );
buf ( n194191 , n26913 );
buf ( n194192 , n194191 );
and ( n26916 , n193980 , n193997 );
buf ( n194194 , n26916 );
buf ( n194195 , n194194 );
buf ( n194196 , n855 );
buf ( n194197 , n888 );
xor ( n26921 , n194196 , n194197 );
buf ( n194199 , n26921 );
buf ( n194200 , n194199 );
not ( n26924 , n194200 );
buf ( n194202 , n190454 );
not ( n26926 , n194202 );
or ( n26927 , n26924 , n26926 );
buf ( n194205 , n20396 );
buf ( n194206 , n193733 );
nand ( n26930 , n194205 , n194206 );
buf ( n194208 , n26930 );
buf ( n194209 , n194208 );
nand ( n26933 , n26927 , n194209 );
buf ( n194211 , n26933 );
not ( n26935 , n194034 );
not ( n26936 , n190485 );
or ( n26937 , n26935 , n26936 );
buf ( n194215 , n190128 );
buf ( n194216 , n193754 );
nand ( n26940 , n194215 , n194216 );
buf ( n194218 , n26940 );
nand ( n26942 , n26937 , n194218 );
or ( n26943 , n194211 , n26942 );
buf ( n194221 , n863 );
buf ( n194222 , n880 );
xor ( n26946 , n194221 , n194222 );
buf ( n194224 , n26946 );
buf ( n194225 , n194224 );
not ( n26949 , n194225 );
buf ( n194227 , n186924 );
not ( n26951 , n194227 );
or ( n26952 , n26949 , n26951 );
buf ( n194230 , n18875 );
buf ( n194231 , n193712 );
nand ( n26955 , n194230 , n194231 );
buf ( n194233 , n26955 );
buf ( n194234 , n194233 );
nand ( n26958 , n26952 , n194234 );
buf ( n194236 , n26958 );
nand ( n26960 , n26943 , n194236 );
buf ( n194238 , n26960 );
nand ( n26962 , n26942 , n194211 );
buf ( n194240 , n26962 );
nand ( n26964 , n194238 , n194240 );
buf ( n194242 , n26964 );
buf ( n194243 , n194242 );
xor ( n26967 , n194195 , n194243 );
buf ( n194245 , n857 );
buf ( n194246 , n886 );
xor ( n26970 , n194245 , n194246 );
buf ( n194248 , n26970 );
buf ( n194249 , n194248 );
not ( n26973 , n194249 );
buf ( n194251 , n190337 );
not ( n26975 , n194251 );
or ( n26976 , n26973 , n26975 );
buf ( n194254 , n20558 );
buf ( n194255 , n193699 );
nand ( n26979 , n194254 , n194255 );
buf ( n194257 , n26979 );
buf ( n194258 , n194257 );
nand ( n26982 , n26976 , n194258 );
buf ( n194260 , n26982 );
buf ( n194261 , n194260 );
xor ( n26985 , n890 , n853 );
buf ( n194263 , n26985 );
not ( n26987 , n194263 );
buf ( n194265 , n188751 );
not ( n26989 , n194265 );
or ( n26990 , n26987 , n26989 );
buf ( n194268 , n20902 );
buf ( n194269 , n193800 );
nand ( n26993 , n194268 , n194269 );
buf ( n194271 , n26993 );
buf ( n194272 , n194271 );
nand ( n26996 , n26990 , n194272 );
buf ( n194274 , n26996 );
buf ( n194275 , n194274 );
or ( n26999 , n194261 , n194275 );
buf ( n194277 , n193939 );
not ( n27001 , n194277 );
buf ( n194279 , n192332 );
not ( n27003 , n194279 );
or ( n27004 , n27001 , n27003 );
buf ( n194282 , n192573 );
buf ( n194283 , n193820 );
nand ( n27007 , n194282 , n194283 );
buf ( n194285 , n27007 );
buf ( n194286 , n194285 );
nand ( n27010 , n27004 , n194286 );
buf ( n194288 , n27010 );
buf ( n194289 , n194288 );
nand ( n27013 , n26999 , n194289 );
buf ( n194291 , n27013 );
buf ( n194292 , n194291 );
buf ( n194293 , n194260 );
buf ( n194294 , n194274 );
nand ( n27018 , n194293 , n194294 );
buf ( n194296 , n27018 );
buf ( n194297 , n194296 );
nand ( n27021 , n194292 , n194297 );
buf ( n194299 , n27021 );
buf ( n194300 , n194299 );
xor ( n27024 , n26967 , n194300 );
buf ( n194302 , n27024 );
buf ( n194303 , n194302 );
xor ( n27027 , n194192 , n194303 );
buf ( n194305 , n26871 );
not ( n27029 , n194305 );
buf ( n194307 , n188751 );
not ( n27031 , n194307 );
or ( n27032 , n27029 , n27031 );
buf ( n194310 , n20902 );
buf ( n194311 , n26985 );
nand ( n27035 , n194310 , n194311 );
buf ( n194313 , n27035 );
buf ( n194314 , n194313 );
nand ( n27038 , n27032 , n194314 );
buf ( n194316 , n27038 );
not ( n27040 , n194316 );
buf ( n194318 , n194068 );
not ( n27042 , n194318 );
buf ( n194320 , n190454 );
not ( n27044 , n194320 );
or ( n27045 , n27042 , n27044 );
buf ( n194323 , n20396 );
buf ( n194324 , n194199 );
nand ( n27048 , n194323 , n194324 );
buf ( n194326 , n27048 );
buf ( n194327 , n194326 );
nand ( n27051 , n27045 , n194327 );
buf ( n194329 , n27051 );
not ( n27053 , n194329 );
nand ( n27054 , n27040 , n27053 );
not ( n27055 , n27054 );
buf ( n194333 , n23353 );
buf ( n194334 , n194248 );
nand ( n27058 , n194333 , n194334 );
buf ( n194336 , n27058 );
nand ( n27060 , n20554 , n194090 );
nand ( n27061 , n194336 , n27060 );
not ( n27062 , n27061 );
or ( n27063 , n27055 , n27062 );
buf ( n194341 , n194316 );
buf ( n194342 , n194329 );
nand ( n27066 , n194341 , n194342 );
buf ( n194344 , n27066 );
nand ( n27068 , n27063 , n194344 );
buf ( n194346 , n27068 );
xor ( n27070 , n194211 , n194236 );
xor ( n27071 , n27070 , n26942 );
buf ( n194349 , n27071 );
xor ( n27073 , n194346 , n194349 );
xor ( n27074 , n194274 , n194260 );
xor ( n27075 , n27074 , n194288 );
buf ( n194353 , n27075 );
and ( n27077 , n27073 , n194353 );
and ( n27078 , n194346 , n194349 );
or ( n27079 , n27077 , n27078 );
buf ( n194357 , n27079 );
buf ( n194358 , n194357 );
xor ( n27082 , n27027 , n194358 );
buf ( n194360 , n27082 );
buf ( n194361 , n194360 );
xor ( n27085 , n26909 , n194361 );
buf ( n194363 , n27085 );
buf ( n27087 , n194363 );
xor ( n27088 , n194346 , n194349 );
xor ( n27089 , n27088 , n194353 );
buf ( n194367 , n27089 );
buf ( n194368 , n194367 );
xor ( n27092 , n193909 , n193927 );
xor ( n27093 , n27092 , n193946 );
buf ( n194371 , n27093 );
buf ( n194372 , n194371 );
xor ( n27096 , n27061 , n27040 );
not ( n27097 , n27053 );
xnor ( n27098 , n27096 , n27097 );
buf ( n194376 , n27098 );
xor ( n27100 , n194372 , n194376 );
buf ( n194378 , n193893 );
buf ( n194379 , n26628 );
xor ( n27103 , n194378 , n194379 );
buf ( n194381 , n27103 );
buf ( n194382 , n194381 );
buf ( n194383 , n26571 );
buf ( n194384 , n863 );
and ( n27108 , n194383 , n194384 );
buf ( n194386 , n27108 );
buf ( n194387 , n194386 );
not ( n27111 , n190454 );
xor ( n27112 , n888 , n858 );
not ( n27113 , n27112 );
or ( n27114 , n27111 , n27113 );
buf ( n194392 , n20396 );
buf ( n194393 , n194058 );
nand ( n27117 , n194392 , n194393 );
buf ( n194395 , n27117 );
nand ( n27119 , n27114 , n194395 );
buf ( n194397 , n27119 );
xor ( n27121 , n194387 , n194397 );
buf ( n194399 , n854 );
buf ( n194400 , n892 );
xor ( n27124 , n194399 , n194400 );
buf ( n194402 , n27124 );
buf ( n194403 , n194402 );
not ( n27127 , n194403 );
buf ( n194405 , n190485 );
not ( n27129 , n194405 );
or ( n27130 , n27127 , n27129 );
buf ( n194408 , n190491 );
buf ( n194409 , n26826 );
nand ( n27133 , n194408 , n194409 );
buf ( n194411 , n27133 );
buf ( n194412 , n194411 );
nand ( n27136 , n27130 , n194412 );
buf ( n194414 , n27136 );
buf ( n194415 , n194414 );
and ( n27139 , n27121 , n194415 );
and ( n27140 , n194387 , n194397 );
or ( n27141 , n27139 , n27140 );
buf ( n194419 , n27141 );
buf ( n194420 , n194419 );
xor ( n27144 , n194382 , n194420 );
buf ( n194422 , n852 );
buf ( n194423 , n894 );
xor ( n27147 , n194422 , n194423 );
buf ( n194425 , n27147 );
buf ( n194426 , n194425 );
not ( n27150 , n194426 );
buf ( n194428 , n23321 );
not ( n27152 , n194428 );
or ( n27153 , n27150 , n27152 );
buf ( n194431 , n193877 );
buf ( n194432 , n895 );
nand ( n27156 , n194431 , n194432 );
buf ( n194434 , n27156 );
buf ( n194435 , n194434 );
nand ( n27159 , n27153 , n194435 );
buf ( n194437 , n27159 );
buf ( n194438 , n194437 );
buf ( n194439 , n860 );
buf ( n194440 , n886 );
xor ( n27164 , n194439 , n194440 );
buf ( n194442 , n27164 );
buf ( n194443 , n194442 );
not ( n27167 , n194443 );
buf ( n194445 , n20554 );
not ( n27169 , n194445 );
or ( n27170 , n27167 , n27169 );
buf ( n194448 , n20558 );
buf ( n194449 , n194080 );
nand ( n27173 , n194448 , n194449 );
buf ( n194451 , n27173 );
buf ( n194452 , n194451 );
nand ( n27176 , n27170 , n194452 );
buf ( n194454 , n27176 );
buf ( n194455 , n194454 );
xor ( n27179 , n194438 , n194455 );
xor ( n27180 , n884 , n862 );
buf ( n194458 , n27180 );
not ( n27182 , n194458 );
buf ( n194460 , n192332 );
not ( n27184 , n194460 );
or ( n27185 , n27182 , n27184 );
buf ( n194463 , n192573 );
buf ( n194464 , n26880 );
nand ( n27188 , n194463 , n194464 );
buf ( n194466 , n27188 );
buf ( n194467 , n194466 );
nand ( n27191 , n27185 , n194467 );
buf ( n194469 , n27191 );
buf ( n194470 , n194469 );
and ( n27194 , n27179 , n194470 );
and ( n27195 , n194438 , n194455 );
or ( n27196 , n27194 , n27195 );
buf ( n194474 , n27196 );
buf ( n194475 , n194474 );
and ( n27199 , n27144 , n194475 );
and ( n27200 , n194382 , n194420 );
or ( n27201 , n27199 , n27200 );
buf ( n194479 , n27201 );
buf ( n194480 , n194479 );
and ( n27204 , n27100 , n194480 );
and ( n27205 , n194372 , n194376 );
or ( n27206 , n27204 , n27205 );
buf ( n194484 , n27206 );
buf ( n194485 , n194484 );
xor ( n27209 , n194368 , n194485 );
xor ( n27210 , n193951 , n194049 );
xor ( n27211 , n27210 , n194180 );
buf ( n194489 , n27211 );
buf ( n194490 , n194489 );
xor ( n27214 , n27209 , n194490 );
buf ( n194492 , n27214 );
buf ( n27216 , n194492 );
buf ( n194494 , n190386 );
not ( n27218 , n194494 );
buf ( n194496 , n188751 );
not ( n27220 , n194496 );
or ( n27221 , n27218 , n27220 );
buf ( n194499 , n20902 );
xor ( n27223 , n890 , n856 );
buf ( n194501 , n27223 );
nand ( n27225 , n194499 , n194501 );
buf ( n194503 , n27225 );
buf ( n194504 , n194503 );
nand ( n27228 , n27221 , n194504 );
buf ( n194506 , n27228 );
xor ( n27230 , n884 , n863 );
buf ( n194508 , n27230 );
not ( n27232 , n194508 );
buf ( n194510 , n192332 );
not ( n27234 , n194510 );
or ( n27235 , n27232 , n27234 );
buf ( n194513 , n192573 );
buf ( n194514 , n27180 );
nand ( n27238 , n194513 , n194514 );
buf ( n194516 , n27238 );
buf ( n194517 , n194516 );
nand ( n27241 , n27235 , n194517 );
buf ( n194519 , n27241 );
xor ( n27243 , n194506 , n194519 );
buf ( n194521 , n27243 );
buf ( n194522 , n863 );
buf ( n194523 , n885 );
or ( n27247 , n194522 , n194523 );
buf ( n194525 , n886 );
nand ( n27249 , n27247 , n194525 );
buf ( n194527 , n27249 );
buf ( n194528 , n194527 );
buf ( n194529 , n863 );
buf ( n194530 , n885 );
nand ( n27254 , n194529 , n194530 );
buf ( n194532 , n27254 );
buf ( n194533 , n194532 );
buf ( n194534 , n884 );
nand ( n27258 , n194528 , n194533 , n194534 );
buf ( n194536 , n27258 );
buf ( n194537 , n194536 );
not ( n27261 , n194537 );
buf ( n194539 , n190584 );
not ( n27263 , n194539 );
buf ( n194541 , n190485 );
not ( n27265 , n194541 );
or ( n27266 , n27263 , n27265 );
buf ( n194544 , n190491 );
buf ( n194545 , n194402 );
nand ( n27269 , n194544 , n194545 );
buf ( n194547 , n27269 );
buf ( n194548 , n194547 );
nand ( n27272 , n27266 , n194548 );
buf ( n194550 , n27272 );
buf ( n194551 , n194550 );
not ( n27275 , n194551 );
or ( n27276 , n27261 , n27275 );
buf ( n194554 , n194550 );
buf ( n194555 , n194536 );
or ( n27279 , n194554 , n194555 );
nand ( n27280 , n27276 , n27279 );
buf ( n194558 , n27280 );
buf ( n194559 , n194558 );
xor ( n27283 , n194521 , n194559 );
buf ( n194561 , n27283 );
buf ( n194562 , n194561 );
xor ( n27286 , n190552 , n190573 );
and ( n27287 , n27286 , n190591 );
and ( n27288 , n190552 , n190573 );
or ( n27289 , n27287 , n27288 );
buf ( n194567 , n27289 );
buf ( n194568 , n194567 );
buf ( n194569 , n190392 );
buf ( n194570 , n190371 );
or ( n27294 , n194569 , n194570 );
buf ( n194572 , n190351 );
nand ( n27296 , n27294 , n194572 );
buf ( n194574 , n27296 );
buf ( n194575 , n194574 );
buf ( n194576 , n190392 );
buf ( n194577 , n190371 );
nand ( n27301 , n194576 , n194577 );
buf ( n194579 , n27301 );
buf ( n194580 , n194579 );
nand ( n27304 , n194575 , n194580 );
buf ( n194582 , n27304 );
buf ( n194583 , n194582 );
xor ( n27307 , n194568 , n194583 );
buf ( n194585 , n190364 );
not ( n27309 , n194585 );
buf ( n194587 , n21330 );
not ( n27311 , n194587 );
or ( n27312 , n27309 , n27311 );
buf ( n194590 , n194425 );
buf ( n194591 , n895 );
nand ( n27315 , n194590 , n194591 );
buf ( n194593 , n27315 );
buf ( n194594 , n194593 );
nand ( n27318 , n27312 , n194594 );
buf ( n194596 , n27318 );
buf ( n194597 , n194596 );
buf ( n194598 , n190345 );
not ( n27322 , n194598 );
buf ( n194600 , n20554 );
not ( n27324 , n194600 );
or ( n27325 , n27322 , n27324 );
buf ( n194603 , n20558 );
buf ( n194604 , n194442 );
nand ( n27328 , n194603 , n194604 );
buf ( n194606 , n27328 );
buf ( n194607 , n194606 );
nand ( n27331 , n27325 , n194607 );
buf ( n194609 , n27331 );
buf ( n194610 , n194609 );
xor ( n27334 , n194597 , n194610 );
buf ( n194612 , n190566 );
not ( n27336 , n194612 );
buf ( n194614 , n190454 );
not ( n27338 , n194614 );
or ( n27339 , n27336 , n27338 );
buf ( n194617 , n27112 );
buf ( n194618 , n20396 );
nand ( n27342 , n194617 , n194618 );
buf ( n194620 , n27342 );
buf ( n194621 , n194620 );
nand ( n27345 , n27339 , n194621 );
buf ( n194623 , n27345 );
buf ( n194624 , n194623 );
xor ( n27348 , n27334 , n194624 );
buf ( n194626 , n27348 );
buf ( n194627 , n194626 );
xor ( n27351 , n27307 , n194627 );
buf ( n194629 , n27351 );
buf ( n194630 , n194629 );
xor ( n27354 , n194562 , n194630 );
xor ( n27355 , n190540 , n190594 );
and ( n27356 , n27355 , n190643 );
and ( n27357 , n190540 , n190594 );
or ( n27358 , n27356 , n27357 );
buf ( n194636 , n27358 );
buf ( n194637 , n194636 );
xor ( n27361 , n27354 , n194637 );
buf ( n194639 , n27361 );
buf ( n27363 , n194639 );
buf ( n194641 , n859 );
buf ( n194642 , n892 );
xor ( n27366 , n194641 , n194642 );
buf ( n194644 , n27366 );
not ( n27368 , n194644 );
not ( n27369 , n190485 );
or ( n27370 , n27368 , n27369 );
buf ( n194648 , n190491 );
buf ( n194649 , n858 );
buf ( n194650 , n892 );
xor ( n27374 , n194649 , n194650 );
buf ( n194652 , n27374 );
buf ( n194653 , n194652 );
nand ( n27377 , n194648 , n194653 );
buf ( n194655 , n27377 );
nand ( n27379 , n27370 , n194655 );
buf ( n194657 , n861 );
buf ( n194658 , n890 );
xor ( n27382 , n194657 , n194658 );
buf ( n194660 , n27382 );
not ( n27384 , n194660 );
not ( n27385 , n188751 );
or ( n27386 , n27384 , n27385 );
buf ( n194664 , n20902 );
buf ( n194665 , n860 );
buf ( n194666 , n890 );
xor ( n27390 , n194665 , n194666 );
buf ( n194668 , n27390 );
buf ( n194669 , n194668 );
nand ( n27393 , n194664 , n194669 );
buf ( n194671 , n27393 );
nand ( n27395 , n27386 , n194671 );
xor ( n27396 , n27379 , n27395 );
buf ( n194674 , n863 );
buf ( n194675 , n888 );
xor ( n27399 , n194674 , n194675 );
buf ( n194677 , n27399 );
not ( n27401 , n194677 );
not ( n27402 , n190454 );
or ( n27403 , n27401 , n27402 );
buf ( n27404 , n20396 );
buf ( n194682 , n27404 );
buf ( n194683 , n190449 );
nand ( n27407 , n194682 , n194683 );
buf ( n194685 , n27407 );
nand ( n27409 , n27403 , n194685 );
and ( n27410 , n27396 , n27409 );
and ( n27411 , n27379 , n27395 );
or ( n27412 , n27410 , n27411 );
buf ( n194690 , n190468 );
buf ( n194691 , n190419 );
not ( n27415 , n194691 );
buf ( n194693 , n23157 );
not ( n27417 , n194693 );
or ( n27418 , n27415 , n27417 );
buf ( n194696 , n23157 );
buf ( n194697 , n190419 );
or ( n27421 , n194696 , n194697 );
nand ( n27422 , n27418 , n27421 );
buf ( n194700 , n27422 );
buf ( n194701 , n194700 );
xor ( n27425 , n194690 , n194701 );
buf ( n194703 , n27425 );
not ( n27427 , n194703 );
xor ( n27428 , n27412 , n27427 );
buf ( n194706 , n194668 );
not ( n27430 , n194706 );
buf ( n194708 , n188751 );
not ( n27432 , n194708 );
or ( n27433 , n27430 , n27432 );
buf ( n194711 , n20902 );
buf ( n194712 , n190398 );
nand ( n27436 , n194711 , n194712 );
buf ( n194714 , n27436 );
buf ( n194715 , n194714 );
nand ( n27439 , n27433 , n194715 );
buf ( n194717 , n27439 );
buf ( n194718 , n194652 );
not ( n27442 , n194718 );
buf ( n194720 , n190485 );
not ( n27444 , n194720 );
or ( n27445 , n27442 , n27444 );
buf ( n194723 , n190491 );
buf ( n194724 , n190480 );
nand ( n27448 , n194723 , n194724 );
buf ( n194726 , n27448 );
buf ( n194727 , n194726 );
nand ( n27451 , n27445 , n194727 );
buf ( n194729 , n27451 );
xor ( n27453 , n194717 , n194729 );
buf ( n194731 , n857 );
buf ( n194732 , n894 );
xor ( n27456 , n194731 , n194732 );
buf ( n194734 , n27456 );
buf ( n194735 , n194734 );
not ( n27459 , n194735 );
buf ( n194737 , n23321 );
not ( n27461 , n194737 );
or ( n27462 , n27459 , n27461 );
buf ( n194740 , n190426 );
buf ( n194741 , n895 );
nand ( n27465 , n194740 , n194741 );
buf ( n194743 , n27465 );
buf ( n194744 , n194743 );
nand ( n27468 , n27462 , n194744 );
buf ( n194746 , n27468 );
buf ( n194747 , n194746 );
buf ( n194748 , n863 );
buf ( n194749 , n889 );
or ( n27473 , n194748 , n194749 );
buf ( n194751 , n890 );
nand ( n27475 , n27473 , n194751 );
buf ( n194753 , n27475 );
buf ( n194754 , n194753 );
buf ( n194755 , n863 );
buf ( n194756 , n889 );
nand ( n27480 , n194755 , n194756 );
buf ( n194758 , n27480 );
buf ( n194759 , n194758 );
buf ( n194760 , n888 );
nand ( n27484 , n194754 , n194759 , n194760 );
buf ( n194762 , n27484 );
buf ( n194763 , n194762 );
not ( n27487 , n194763 );
buf ( n194765 , n27487 );
buf ( n194766 , n194765 );
nand ( n27490 , n194747 , n194766 );
buf ( n194768 , n27490 );
buf ( n194769 , n194768 );
not ( n27493 , n194769 );
buf ( n194771 , n27493 );
and ( n27495 , n27453 , n194771 );
not ( n27496 , n27453 );
and ( n27497 , n27496 , n194768 );
or ( n27498 , n27495 , n27497 );
xnor ( n27499 , n27428 , n27498 );
not ( n27500 , n27499 );
buf ( n27501 , n27500 );
buf ( n194779 , n863 );
buf ( n194780 , n893 );
or ( n27504 , n194779 , n194780 );
buf ( n194782 , n894 );
nand ( n27506 , n27504 , n194782 );
buf ( n194784 , n27506 );
buf ( n194785 , n194784 );
buf ( n194786 , n863 );
buf ( n194787 , n893 );
nand ( n27511 , n194786 , n194787 );
buf ( n194789 , n27511 );
buf ( n194790 , n194789 );
buf ( n194791 , n892 );
and ( n27515 , n194785 , n194790 , n194791 );
buf ( n194793 , n27515 );
buf ( n194794 , n194793 );
buf ( n194795 , n861 );
buf ( n194796 , n894 );
xor ( n27520 , n194795 , n194796 );
buf ( n194798 , n27520 );
buf ( n194799 , n194798 );
not ( n27523 , n194799 );
buf ( n194801 , n21330 );
not ( n27525 , n194801 );
or ( n27526 , n27523 , n27525 );
buf ( n194804 , n860 );
buf ( n194805 , n894 );
xor ( n27529 , n194804 , n194805 );
buf ( n194807 , n27529 );
buf ( n194808 , n194807 );
buf ( n194809 , n895 );
nand ( n27533 , n194808 , n194809 );
buf ( n194811 , n27533 );
buf ( n194812 , n194811 );
nand ( n27536 , n27526 , n194812 );
buf ( n194814 , n27536 );
buf ( n194815 , n194814 );
xor ( n27539 , n194794 , n194815 );
buf ( n194817 , n27539 );
buf ( n27541 , n194817 );
xor ( n27542 , n191759 , n192146 );
and ( n27543 , n27542 , n192162 );
and ( n27544 , n191759 , n192146 );
or ( n27545 , n27543 , n27544 );
buf ( n194823 , n27545 );
buf ( n27547 , n194823 );
xor ( n27548 , n194382 , n194420 );
xor ( n27549 , n27548 , n194475 );
buf ( n194827 , n27549 );
buf ( n194828 , n194827 );
xor ( n27552 , n194387 , n194397 );
xor ( n27553 , n27552 , n194415 );
buf ( n194831 , n27553 );
buf ( n194832 , n194831 );
xor ( n27556 , n194438 , n194455 );
xor ( n27557 , n27556 , n194470 );
buf ( n194835 , n27557 );
buf ( n194836 , n194835 );
xor ( n27560 , n194832 , n194836 );
buf ( n194838 , n194519 );
buf ( n194839 , n194506 );
or ( n27563 , n194838 , n194839 );
buf ( n194841 , n27563 );
not ( n27565 , n194841 );
not ( n27566 , n194558 );
or ( n27567 , n27565 , n27566 );
buf ( n194845 , n194506 );
buf ( n194846 , n194519 );
nand ( n27570 , n194845 , n194846 );
buf ( n194848 , n27570 );
nand ( n27572 , n27567 , n194848 );
buf ( n194850 , n27572 );
and ( n27574 , n27560 , n194850 );
and ( n27575 , n194832 , n194836 );
or ( n27576 , n27574 , n27575 );
buf ( n194854 , n27576 );
buf ( n194855 , n194854 );
xor ( n27579 , n194828 , n194855 );
buf ( n27580 , n194115 );
buf ( n194858 , n27580 );
not ( n27582 , n194858 );
xnor ( n27583 , n194096 , n194074 );
buf ( n194861 , n27583 );
not ( n27585 , n194861 );
or ( n27586 , n27582 , n27585 );
buf ( n194864 , n27583 );
buf ( n194865 , n27580 );
or ( n27589 , n194864 , n194865 );
nand ( n27590 , n27586 , n27589 );
buf ( n194868 , n27590 );
buf ( n194869 , n194868 );
xor ( n27593 , n194137 , n194155 );
xor ( n27594 , n27593 , n194170 );
buf ( n194872 , n27594 );
buf ( n194873 , n194872 );
xor ( n27597 , n194869 , n194873 );
buf ( n194875 , n27223 );
not ( n27599 , n194875 );
buf ( n194877 , n188751 );
not ( n27601 , n194877 );
or ( n27602 , n27599 , n27601 );
buf ( n27603 , n20902 );
buf ( n194881 , n27603 );
buf ( n194882 , n194141 );
nand ( n27606 , n194881 , n194882 );
buf ( n194884 , n27606 );
buf ( n194885 , n194884 );
nand ( n27609 , n27602 , n194885 );
buf ( n194887 , n27609 );
buf ( n194888 , n194887 );
buf ( n194889 , n194550 );
not ( n27613 , n194889 );
buf ( n194891 , n194536 );
nor ( n27615 , n27613 , n194891 );
buf ( n194893 , n27615 );
buf ( n194894 , n194893 );
xor ( n27618 , n194888 , n194894 );
xor ( n27619 , n194597 , n194610 );
and ( n27620 , n27619 , n194624 );
and ( n27621 , n194597 , n194610 );
or ( n27622 , n27620 , n27621 );
buf ( n194900 , n27622 );
buf ( n194901 , n194900 );
and ( n27625 , n27618 , n194901 );
and ( n27626 , n194888 , n194894 );
or ( n27627 , n27625 , n27626 );
buf ( n194905 , n27627 );
buf ( n194906 , n194905 );
xor ( n27630 , n27597 , n194906 );
buf ( n194908 , n27630 );
buf ( n194909 , n194908 );
xor ( n27633 , n27579 , n194909 );
buf ( n194911 , n27633 );
buf ( n27635 , n194911 );
buf ( n194913 , n863 );
buf ( n194914 , n877 );
or ( n27638 , n194913 , n194914 );
buf ( n194916 , n878 );
nand ( n27640 , n27638 , n194916 );
buf ( n194918 , n27640 );
buf ( n194919 , n194918 );
buf ( n194920 , n863 );
buf ( n194921 , n877 );
nand ( n27645 , n194920 , n194921 );
buf ( n194923 , n27645 );
buf ( n194924 , n194923 );
buf ( n194925 , n876 );
nand ( n27649 , n194919 , n194924 , n194925 );
buf ( n194927 , n27649 );
buf ( n194928 , n194927 );
not ( n27652 , n194928 );
xor ( n27653 , n894 , n845 );
buf ( n194931 , n27653 );
not ( n27655 , n194931 );
buf ( n194933 , n20165 );
not ( n27657 , n194933 );
or ( n27658 , n27655 , n27657 );
xor ( n27659 , n894 , n844 );
buf ( n194937 , n27659 );
buf ( n194938 , n895 );
nand ( n27662 , n194937 , n194938 );
buf ( n194940 , n27662 );
buf ( n194941 , n194940 );
nand ( n27665 , n27658 , n194941 );
buf ( n194943 , n27665 );
buf ( n194944 , n194943 );
nand ( n27668 , n27652 , n194944 );
buf ( n194946 , n27668 );
buf ( n194947 , n194946 );
not ( n27671 , n194947 );
buf ( n194949 , n856 );
buf ( n194950 , n882 );
xor ( n27674 , n194949 , n194950 );
buf ( n194952 , n27674 );
buf ( n194953 , n194952 );
not ( n27677 , n194953 );
buf ( n194955 , n19613 );
not ( n27679 , n194955 );
or ( n27680 , n27677 , n27679 );
buf ( n194958 , n26571 );
xor ( n27682 , n882 , n855 );
buf ( n194960 , n27682 );
nand ( n27684 , n194958 , n194960 );
buf ( n194962 , n27684 );
buf ( n194963 , n194962 );
nand ( n27687 , n27680 , n194963 );
buf ( n194965 , n27687 );
buf ( n194966 , n194965 );
nor ( n27690 , n27671 , n194966 );
buf ( n194968 , n27690 );
buf ( n194969 , n194968 );
not ( n27693 , n194969 );
buf ( n194971 , n194946 );
not ( n27695 , n194971 );
buf ( n194973 , n194965 );
nand ( n27697 , n27695 , n194973 );
buf ( n194975 , n27697 );
buf ( n194976 , n194975 );
nand ( n27700 , n27693 , n194976 );
buf ( n194978 , n27700 );
buf ( n194979 , n194978 );
buf ( n194980 , n854 );
buf ( n194981 , n884 );
xor ( n27705 , n194980 , n194981 );
buf ( n194983 , n27705 );
buf ( n194984 , n194983 );
not ( n27708 , n194984 );
buf ( n194986 , n192332 );
not ( n27710 , n194986 );
or ( n27711 , n27708 , n27710 );
buf ( n194989 , n192573 );
buf ( n194990 , n853 );
buf ( n194991 , n884 );
xor ( n27715 , n194990 , n194991 );
buf ( n194993 , n27715 );
buf ( n194994 , n194993 );
nand ( n27718 , n194989 , n194994 );
buf ( n194996 , n27718 );
buf ( n194997 , n194996 );
nand ( n27721 , n27711 , n194997 );
buf ( n194999 , n27721 );
buf ( n27723 , n194999 );
not ( n27724 , n27723 );
buf ( n195002 , n27724 );
and ( n27726 , n194979 , n195002 );
not ( n27727 , n194979 );
buf ( n195005 , n27723 );
and ( n27729 , n27727 , n195005 );
nor ( n27730 , n27726 , n27729 );
buf ( n195008 , n27730 );
buf ( n195009 , n195008 );
buf ( n195010 , n194927 );
not ( n27734 , n195010 );
buf ( n195012 , n194943 );
not ( n27736 , n195012 );
or ( n27737 , n27734 , n27736 );
buf ( n195015 , n194943 );
buf ( n195016 , n194927 );
or ( n27740 , n195015 , n195016 );
nand ( n27741 , n27737 , n27740 );
buf ( n195019 , n27741 );
buf ( n195020 , n195019 );
buf ( n195021 , n846 );
buf ( n195022 , n894 );
xor ( n27746 , n195021 , n195022 );
buf ( n195024 , n27746 );
buf ( n195025 , n195024 );
not ( n27749 , n195025 );
buf ( n195027 , n21330 );
not ( n27751 , n195027 );
or ( n27752 , n27749 , n27751 );
buf ( n195030 , n27653 );
buf ( n195031 , n895 );
nand ( n27755 , n195030 , n195031 );
buf ( n195033 , n27755 );
buf ( n195034 , n195033 );
nand ( n27758 , n27752 , n195034 );
buf ( n195036 , n27758 );
buf ( n195037 , n195036 );
buf ( n195038 , n19103 );
buf ( n195039 , n863 );
and ( n27763 , n195038 , n195039 );
buf ( n195041 , n27763 );
buf ( n195042 , n195041 );
xor ( n27766 , n195037 , n195042 );
buf ( n195044 , n190454 );
not ( n27768 , n195044 );
buf ( n195046 , n27768 );
buf ( n195047 , n195046 );
buf ( n195048 , n852 );
buf ( n195049 , n888 );
xnor ( n27773 , n195048 , n195049 );
buf ( n195051 , n27773 );
buf ( n195052 , n195051 );
or ( n27776 , n195047 , n195052 );
buf ( n195054 , n193034 );
buf ( n195055 , n851 );
buf ( n195056 , n888 );
xor ( n27780 , n195055 , n195056 );
buf ( n195058 , n27780 );
buf ( n195059 , n195058 );
not ( n27783 , n195059 );
buf ( n195061 , n27783 );
buf ( n195062 , n195061 );
or ( n27786 , n195054 , n195062 );
nand ( n27787 , n27776 , n27786 );
buf ( n195065 , n27787 );
buf ( n195066 , n195065 );
and ( n27790 , n27766 , n195066 );
and ( n27791 , n195037 , n195042 );
or ( n27792 , n27790 , n27791 );
buf ( n195070 , n27792 );
buf ( n195071 , n195070 );
xor ( n27795 , n195020 , n195071 );
xor ( n27796 , n892 , n848 );
buf ( n195074 , n27796 );
not ( n27798 , n195074 );
buf ( n195076 , n190485 );
not ( n27800 , n195076 );
or ( n27801 , n27798 , n27800 );
buf ( n195079 , n190128 );
xor ( n27803 , n892 , n847 );
buf ( n195081 , n27803 );
nand ( n27805 , n195079 , n195081 );
buf ( n195083 , n27805 );
buf ( n195084 , n195083 );
nand ( n27808 , n27801 , n195084 );
buf ( n195086 , n27808 );
buf ( n195087 , n195086 );
buf ( n195088 , n859 );
buf ( n195089 , n880 );
xor ( n27813 , n195088 , n195089 );
buf ( n195091 , n27813 );
buf ( n195092 , n195091 );
not ( n27816 , n195092 );
buf ( n195094 , n18875 );
not ( n27818 , n195094 );
or ( n27819 , n27816 , n27818 );
buf ( n195097 , n18862 );
buf ( n195098 , n860 );
buf ( n195099 , n880 );
xor ( n27823 , n195098 , n195099 );
buf ( n195101 , n27823 );
buf ( n195102 , n195101 );
nand ( n27826 , n195097 , n195102 );
buf ( n195104 , n27826 );
buf ( n195105 , n195104 );
nand ( n27829 , n27819 , n195105 );
buf ( n195107 , n27829 );
buf ( n195108 , n195107 );
xor ( n27832 , n195087 , n195108 );
buf ( n195110 , n862 );
buf ( n195111 , n878 );
xor ( n27835 , n195110 , n195111 );
buf ( n195113 , n27835 );
buf ( n195114 , n195113 );
not ( n27838 , n195114 );
buf ( n195116 , n186569 );
not ( n27840 , n195116 );
or ( n27841 , n27838 , n27840 );
buf ( n195119 , n186575 );
buf ( n195120 , n861 );
buf ( n195121 , n878 );
xor ( n27845 , n195120 , n195121 );
buf ( n195123 , n27845 );
buf ( n195124 , n195123 );
nand ( n27848 , n195119 , n195124 );
buf ( n195126 , n27848 );
buf ( n195127 , n195126 );
nand ( n27851 , n27841 , n195127 );
buf ( n195129 , n27851 );
buf ( n195130 , n195129 );
and ( n27854 , n27832 , n195130 );
and ( n27855 , n195087 , n195108 );
or ( n27856 , n27854 , n27855 );
buf ( n195134 , n27856 );
buf ( n195135 , n195134 );
and ( n27859 , n27795 , n195135 );
and ( n27860 , n195020 , n195071 );
or ( n27861 , n27859 , n27860 );
buf ( n195139 , n27861 );
buf ( n195140 , n195139 );
xor ( n27864 , n195009 , n195140 );
not ( n27865 , n195058 );
not ( n27866 , n20391 );
or ( n27867 , n27865 , n27866 );
buf ( n195145 , n850 );
buf ( n195146 , n888 );
xor ( n27870 , n195145 , n195146 );
buf ( n195148 , n27870 );
nand ( n27872 , n20396 , n195148 );
nand ( n27873 , n27867 , n27872 );
buf ( n195151 , n195091 );
not ( n27875 , n195151 );
buf ( n195153 , n18862 );
not ( n27877 , n195153 );
or ( n27878 , n27875 , n27877 );
buf ( n195156 , n22304 );
buf ( n195157 , n858 );
buf ( n195158 , n880 );
xor ( n27882 , n195157 , n195158 );
buf ( n195160 , n27882 );
buf ( n195161 , n195160 );
nand ( n27885 , n195156 , n195161 );
buf ( n195163 , n27885 );
buf ( n195164 , n195163 );
nand ( n27888 , n27878 , n195164 );
buf ( n195166 , n27888 );
xor ( n27890 , n27873 , n195166 );
buf ( n195168 , n195123 );
not ( n27892 , n195168 );
buf ( n195170 , n186569 );
not ( n27894 , n195170 );
or ( n27895 , n27892 , n27894 );
buf ( n195173 , n186575 );
buf ( n195174 , n860 );
buf ( n195175 , n878 );
xor ( n27899 , n195174 , n195175 );
buf ( n195177 , n27899 );
buf ( n195178 , n195177 );
nand ( n27902 , n195173 , n195178 );
buf ( n195180 , n27902 );
buf ( n195181 , n195180 );
nand ( n27905 , n27895 , n195181 );
buf ( n195183 , n27905 );
xor ( n27907 , n27890 , n195183 );
buf ( n195185 , n27907 );
buf ( n195186 , n850 );
buf ( n195187 , n890 );
xor ( n27911 , n195186 , n195187 );
buf ( n195189 , n27911 );
buf ( n195190 , n195189 );
not ( n27914 , n195190 );
buf ( n195192 , n188751 );
not ( n27916 , n195192 );
or ( n27917 , n27914 , n27916 );
buf ( n195195 , n20902 );
buf ( n195196 , n849 );
buf ( n195197 , n890 );
xor ( n27921 , n195196 , n195197 );
buf ( n195199 , n27921 );
buf ( n195200 , n195199 );
nand ( n27924 , n195195 , n195200 );
buf ( n195202 , n27924 );
buf ( n195203 , n195202 );
nand ( n27927 , n27917 , n195203 );
buf ( n195205 , n27927 );
not ( n27929 , n195205 );
buf ( n195207 , n854 );
buf ( n195208 , n886 );
xor ( n27932 , n195207 , n195208 );
buf ( n195210 , n27932 );
buf ( n195211 , n195210 );
not ( n27935 , n195211 );
buf ( n195213 , n20554 );
not ( n27937 , n195213 );
or ( n27938 , n27935 , n27937 );
buf ( n195216 , n23353 );
buf ( n195217 , n853 );
buf ( n195218 , n886 );
xor ( n27942 , n195217 , n195218 );
buf ( n195220 , n27942 );
buf ( n195221 , n195220 );
nand ( n27945 , n195216 , n195221 );
buf ( n195223 , n27945 );
buf ( n195224 , n195223 );
nand ( n27948 , n27938 , n195224 );
buf ( n195226 , n27948 );
not ( n27950 , n195226 );
or ( n27951 , n27929 , n27950 );
or ( n27952 , n195205 , n195226 );
buf ( n195230 , n856 );
buf ( n195231 , n884 );
xor ( n27955 , n195230 , n195231 );
buf ( n195233 , n27955 );
buf ( n195234 , n195233 );
not ( n27958 , n195234 );
buf ( n195236 , n192332 );
not ( n27960 , n195236 );
or ( n27961 , n27958 , n27960 );
buf ( n195239 , n190543 );
buf ( n195240 , n855 );
buf ( n195241 , n884 );
xor ( n27965 , n195240 , n195241 );
buf ( n195243 , n27965 );
buf ( n195244 , n195243 );
nand ( n27968 , n195239 , n195244 );
buf ( n195246 , n27968 );
buf ( n195247 , n195246 );
nand ( n27971 , n27961 , n195247 );
buf ( n195249 , n27971 );
nand ( n27973 , n27952 , n195249 );
nand ( n27974 , n27951 , n27973 );
buf ( n195252 , n27974 );
or ( n27976 , n195185 , n195252 );
not ( n27977 , n195199 );
not ( n27978 , n188751 );
or ( n27979 , n27977 , n27978 );
buf ( n195257 , n20902 );
buf ( n195258 , n848 );
buf ( n195259 , n890 );
xor ( n27983 , n195258 , n195259 );
buf ( n195261 , n27983 );
buf ( n195262 , n195261 );
nand ( n27986 , n195257 , n195262 );
buf ( n195264 , n27986 );
nand ( n27988 , n27979 , n195264 );
buf ( n195266 , n27988 );
buf ( n195267 , n857 );
buf ( n195268 , n882 );
xor ( n27992 , n195267 , n195268 );
buf ( n195270 , n27992 );
not ( n27994 , n195270 );
not ( n27995 , n19613 );
or ( n27996 , n27994 , n27995 );
buf ( n195274 , n26571 );
buf ( n195275 , n194952 );
nand ( n27999 , n195274 , n195275 );
buf ( n195277 , n27999 );
nand ( n28001 , n27996 , n195277 );
buf ( n195279 , n28001 );
xor ( n28003 , n195266 , n195279 );
buf ( n195281 , n28003 );
buf ( n195282 , n195281 );
buf ( n195283 , n195243 );
not ( n28007 , n195283 );
buf ( n195285 , n192332 );
not ( n28009 , n195285 );
or ( n28010 , n28007 , n28009 );
buf ( n195288 , n190543 );
buf ( n195289 , n194983 );
nand ( n28013 , n195288 , n195289 );
buf ( n195291 , n28013 );
buf ( n195292 , n195291 );
nand ( n28016 , n28010 , n195292 );
buf ( n195294 , n28016 );
buf ( n195295 , n195294 );
xor ( n28019 , n195282 , n195295 );
buf ( n195297 , n28019 );
buf ( n195298 , n195297 );
nand ( n28022 , n27976 , n195298 );
buf ( n195300 , n28022 );
buf ( n195301 , n195300 );
buf ( n195302 , n27974 );
buf ( n195303 , n27907 );
nand ( n28027 , n195302 , n195303 );
buf ( n195305 , n28027 );
buf ( n195306 , n195305 );
nand ( n28030 , n195301 , n195306 );
buf ( n195308 , n28030 );
buf ( n195309 , n195308 );
and ( n28033 , n27864 , n195309 );
and ( n28034 , n195009 , n195140 );
or ( n28035 , n28033 , n28034 );
buf ( n195313 , n28035 );
buf ( n195314 , n195313 );
buf ( n195315 , n187865 );
buf ( n195316 , n863 );
and ( n28040 , n195315 , n195316 );
buf ( n195318 , n28040 );
buf ( n195319 , n195318 );
buf ( n195320 , n27659 );
not ( n28044 , n195320 );
buf ( n195322 , n23321 );
not ( n28046 , n195322 );
or ( n28047 , n28044 , n28046 );
buf ( n195325 , n843 );
buf ( n195326 , n894 );
xor ( n28050 , n195325 , n195326 );
buf ( n195328 , n28050 );
buf ( n195329 , n195328 );
buf ( n195330 , n895 );
nand ( n28054 , n195329 , n195330 );
buf ( n195332 , n28054 );
buf ( n195333 , n195332 );
nand ( n28057 , n28047 , n195333 );
buf ( n195335 , n28057 );
buf ( n195336 , n195335 );
xor ( n28060 , n195319 , n195336 );
buf ( n195338 , n195148 );
not ( n28062 , n195338 );
buf ( n195340 , n20391 );
not ( n28064 , n195340 );
or ( n28065 , n28062 , n28064 );
buf ( n195343 , n20396 );
buf ( n195344 , n849 );
buf ( n195345 , n888 );
xor ( n28069 , n195344 , n195345 );
buf ( n195347 , n28069 );
buf ( n195348 , n195347 );
nand ( n28072 , n195343 , n195348 );
buf ( n195350 , n28072 );
buf ( n195351 , n195350 );
nand ( n28075 , n28065 , n195351 );
buf ( n195353 , n28075 );
buf ( n195354 , n195353 );
xor ( n28078 , n28060 , n195354 );
buf ( n195356 , n28078 );
buf ( n195357 , n195356 );
buf ( n195358 , n195261 );
not ( n28082 , n195358 );
buf ( n195360 , n188751 );
not ( n28084 , n195360 );
or ( n28085 , n28082 , n28084 );
buf ( n195363 , n20902 );
buf ( n195364 , n847 );
buf ( n195365 , n890 );
xor ( n28089 , n195364 , n195365 );
buf ( n195367 , n28089 );
buf ( n195368 , n195367 );
nand ( n28092 , n195363 , n195368 );
buf ( n195370 , n28092 );
buf ( n195371 , n195370 );
nand ( n28095 , n28085 , n195371 );
buf ( n195373 , n28095 );
buf ( n195374 , n195373 );
buf ( n195375 , n862 );
buf ( n195376 , n876 );
xor ( n28100 , n195375 , n195376 );
buf ( n195378 , n28100 );
buf ( n195379 , n195378 );
not ( n28103 , n195379 );
buf ( n195381 , n19177 );
not ( n28105 , n195381 );
or ( n28106 , n28103 , n28105 );
buf ( n195384 , n19103 );
buf ( n195385 , n861 );
buf ( n195386 , n876 );
xor ( n28110 , n195385 , n195386 );
buf ( n195388 , n28110 );
buf ( n195389 , n195388 );
nand ( n28113 , n195384 , n195389 );
buf ( n195391 , n28113 );
buf ( n195392 , n195391 );
nand ( n28116 , n28106 , n195392 );
buf ( n195394 , n28116 );
buf ( n195395 , n195394 );
xor ( n28119 , n195374 , n195395 );
xor ( n28120 , n886 , n852 );
buf ( n195398 , n28120 );
not ( n28122 , n195398 );
buf ( n195400 , n190337 );
not ( n28124 , n195400 );
or ( n28125 , n28122 , n28124 );
buf ( n195403 , n20558 );
buf ( n195404 , n851 );
buf ( n195405 , n886 );
xor ( n28129 , n195404 , n195405 );
buf ( n195407 , n28129 );
buf ( n195408 , n195407 );
nand ( n28132 , n195403 , n195408 );
buf ( n195410 , n28132 );
buf ( n195411 , n195410 );
nand ( n28135 , n28125 , n195411 );
buf ( n195413 , n28135 );
buf ( n195414 , n195413 );
xor ( n28138 , n28119 , n195414 );
buf ( n195416 , n28138 );
buf ( n195417 , n195416 );
xor ( n28141 , n195357 , n195417 );
buf ( n195419 , n195177 );
not ( n28143 , n195419 );
buf ( n195421 , n186569 );
not ( n28145 , n195421 );
or ( n28146 , n28143 , n28145 );
buf ( n195424 , n186575 );
buf ( n195425 , n859 );
buf ( n195426 , n878 );
xor ( n28150 , n195425 , n195426 );
buf ( n195428 , n28150 );
buf ( n195429 , n195428 );
nand ( n28153 , n195424 , n195429 );
buf ( n195431 , n28153 );
buf ( n195432 , n195431 );
nand ( n28156 , n28146 , n195432 );
buf ( n195434 , n28156 );
buf ( n195435 , n195434 );
not ( n28159 , n195435 );
buf ( n195437 , n195160 );
not ( n28161 , n195437 );
buf ( n195439 , n18862 );
not ( n28163 , n195439 );
or ( n28164 , n28161 , n28163 );
buf ( n195442 , n191227 );
buf ( n195443 , n857 );
buf ( n195444 , n880 );
xor ( n28168 , n195443 , n195444 );
buf ( n195446 , n28168 );
buf ( n195447 , n195446 );
nand ( n28171 , n195442 , n195447 );
buf ( n195449 , n28171 );
buf ( n195450 , n195449 );
nand ( n28174 , n28164 , n195450 );
buf ( n195452 , n28174 );
buf ( n195453 , n195452 );
not ( n28177 , n195453 );
buf ( n195455 , n28177 );
buf ( n195456 , n195455 );
not ( n28180 , n195456 );
or ( n28181 , n28159 , n28180 );
buf ( n195459 , n195434 );
buf ( n195460 , n195455 );
or ( n28184 , n195459 , n195460 );
nand ( n28185 , n28181 , n28184 );
buf ( n195463 , n28185 );
buf ( n195464 , n195463 );
buf ( n195465 , n846 );
buf ( n195466 , n892 );
xor ( n28190 , n195465 , n195466 );
buf ( n195468 , n28190 );
buf ( n195469 , n195468 );
not ( n28193 , n195469 );
buf ( n195471 , n190485 );
not ( n28195 , n195471 );
or ( n28196 , n28193 , n28195 );
buf ( n195474 , n190128 );
buf ( n195475 , n845 );
buf ( n195476 , n892 );
xor ( n28200 , n195475 , n195476 );
buf ( n195478 , n28200 );
buf ( n195479 , n195478 );
nand ( n28203 , n195474 , n195479 );
buf ( n195481 , n28203 );
buf ( n195482 , n195481 );
nand ( n28206 , n28196 , n195482 );
buf ( n195484 , n28206 );
buf ( n195485 , n195484 );
and ( n28209 , n195464 , n195485 );
not ( n28210 , n195464 );
buf ( n195488 , n195484 );
not ( n28212 , n195488 );
buf ( n195490 , n28212 );
buf ( n195491 , n195490 );
and ( n28215 , n28210 , n195491 );
nor ( n28216 , n28209 , n28215 );
buf ( n195494 , n28216 );
buf ( n195495 , n195494 );
xor ( n28219 , n28141 , n195495 );
buf ( n195497 , n28219 );
not ( n28221 , n195497 );
not ( n28222 , n27988 );
not ( n28223 , n28001 );
or ( n28224 , n28222 , n28223 );
or ( n28225 , n27988 , n28001 );
not ( n28226 , n195243 );
not ( n28227 , n192332 );
or ( n28228 , n28226 , n28227 );
nand ( n28229 , n28228 , n195291 );
nand ( n28230 , n28225 , n28229 );
nand ( n28231 , n28224 , n28230 );
buf ( n195509 , n28231 );
xor ( n28233 , n27873 , n195166 );
and ( n28234 , n28233 , n195183 );
and ( n28235 , n27873 , n195166 );
or ( n28236 , n28234 , n28235 );
buf ( n195514 , n28236 );
xor ( n28238 , n195509 , n195514 );
buf ( n195516 , n28238 );
buf ( n195517 , n195516 );
buf ( n195518 , n195220 );
not ( n28242 , n195518 );
buf ( n195520 , n20554 );
not ( n28244 , n195520 );
or ( n28245 , n28242 , n28244 );
buf ( n195523 , n20558 );
buf ( n195524 , n28120 );
nand ( n28248 , n195523 , n195524 );
buf ( n195526 , n28248 );
buf ( n195527 , n195526 );
nand ( n28251 , n28245 , n195527 );
buf ( n195529 , n28251 );
not ( n28253 , n195529 );
buf ( n195531 , n27803 );
not ( n28255 , n195531 );
buf ( n195533 , n190485 );
not ( n28257 , n195533 );
or ( n28258 , n28255 , n28257 );
buf ( n195536 , n190128 );
buf ( n195537 , n195468 );
nand ( n28261 , n195536 , n195537 );
buf ( n195539 , n28261 );
buf ( n195540 , n195539 );
nand ( n28264 , n28258 , n195540 );
buf ( n195542 , n28264 );
not ( n28266 , n195542 );
or ( n28267 , n28253 , n28266 );
buf ( n195545 , n195529 );
buf ( n195546 , n195542 );
or ( n28270 , n195545 , n195546 );
buf ( n195548 , n863 );
buf ( n195549 , n876 );
xor ( n28273 , n195548 , n195549 );
buf ( n195551 , n28273 );
buf ( n195552 , n195551 );
not ( n28276 , n195552 );
buf ( n195554 , n19098 );
not ( n28278 , n195554 );
or ( n28279 , n28276 , n28278 );
buf ( n195557 , n19103 );
buf ( n195558 , n195378 );
nand ( n28282 , n195557 , n195558 );
buf ( n195560 , n28282 );
buf ( n195561 , n195560 );
nand ( n28285 , n28279 , n195561 );
buf ( n195563 , n28285 );
buf ( n195564 , n195563 );
nand ( n28288 , n28270 , n195564 );
buf ( n195566 , n28288 );
nand ( n28290 , n28267 , n195566 );
buf ( n195568 , n28290 );
not ( n28292 , n195568 );
buf ( n195570 , n28292 );
buf ( n195571 , n195570 );
and ( n28295 , n195517 , n195571 );
not ( n28296 , n195517 );
buf ( n195574 , n28290 );
and ( n28298 , n28296 , n195574 );
nor ( n28299 , n28295 , n28298 );
buf ( n195577 , n28299 );
nand ( n28301 , n28221 , n195577 );
not ( n28302 , n28301 );
xor ( n28303 , n195009 , n195140 );
xor ( n28304 , n28303 , n195309 );
buf ( n195582 , n28304 );
not ( n28306 , n195582 );
or ( n28307 , n28302 , n28306 );
buf ( n195585 , n195577 );
not ( n28309 , n195585 );
buf ( n195587 , n195497 );
nand ( n28311 , n28309 , n195587 );
buf ( n195589 , n28311 );
nand ( n28313 , n28307 , n195589 );
buf ( n195591 , n28313 );
xor ( n28315 , n195314 , n195591 );
xor ( n28316 , n195357 , n195417 );
and ( n28317 , n28316 , n195495 );
and ( n28318 , n195357 , n195417 );
or ( n28319 , n28317 , n28318 );
buf ( n195597 , n28319 );
buf ( n195598 , n195597 );
buf ( n195599 , n194968 );
not ( n28323 , n194999 );
buf ( n195601 , n28323 );
or ( n28325 , n195599 , n195601 );
buf ( n195603 , n194975 );
nand ( n28327 , n28325 , n195603 );
buf ( n195605 , n28327 );
buf ( n195606 , n195605 );
buf ( n195607 , n195388 );
not ( n28331 , n195607 );
buf ( n195609 , n19177 );
not ( n28333 , n195609 );
or ( n28334 , n28331 , n28333 );
buf ( n195612 , n20279 );
buf ( n195613 , n860 );
buf ( n195614 , n876 );
xor ( n28338 , n195613 , n195614 );
buf ( n195616 , n28338 );
buf ( n195617 , n195616 );
nand ( n28341 , n195612 , n195617 );
buf ( n195619 , n28341 );
buf ( n195620 , n195619 );
nand ( n28344 , n28334 , n195620 );
buf ( n195622 , n28344 );
buf ( n195623 , n195622 );
not ( n28347 , n195623 );
buf ( n195625 , n28347 );
not ( n28349 , n195407 );
not ( n28350 , n20554 );
or ( n28351 , n28349 , n28350 );
buf ( n195629 , n850 );
buf ( n195630 , n886 );
xor ( n28354 , n195629 , n195630 );
buf ( n195632 , n28354 );
nand ( n28356 , n195632 , n20558 );
nand ( n28357 , n28351 , n28356 );
xor ( n28358 , n195625 , n28357 );
buf ( n195636 , n863 );
buf ( n195637 , n874 );
xor ( n28361 , n195636 , n195637 );
buf ( n195639 , n28361 );
buf ( n195640 , n195639 );
not ( n28364 , n195640 );
buf ( n195642 , n20582 );
not ( n28366 , n195642 );
or ( n28367 , n28364 , n28366 );
buf ( n195645 , n186297 );
xor ( n28369 , n874 , n862 );
buf ( n195647 , n28369 );
nand ( n28371 , n195645 , n195647 );
buf ( n195649 , n28371 );
buf ( n195650 , n195649 );
nand ( n28374 , n28367 , n195650 );
buf ( n195652 , n28374 );
not ( n28376 , n195652 );
xor ( n28377 , n28358 , n28376 );
buf ( n195655 , n28377 );
xor ( n28379 , n195606 , n195655 );
buf ( n195657 , n195446 );
not ( n28381 , n195657 );
buf ( n195659 , n18862 );
not ( n28383 , n195659 );
or ( n28384 , n28381 , n28383 );
buf ( n195662 , n856 );
buf ( n195663 , n880 );
xor ( n28387 , n195662 , n195663 );
buf ( n195665 , n28387 );
buf ( n195666 , n195665 );
buf ( n195667 , n20358 );
nand ( n28391 , n195666 , n195667 );
buf ( n195669 , n28391 );
buf ( n195670 , n195669 );
nand ( n28394 , n28384 , n195670 );
buf ( n195672 , n28394 );
buf ( n195673 , n195672 );
not ( n28397 , n195673 );
buf ( n195675 , n28397 );
buf ( n195676 , n195347 );
not ( n28400 , n195676 );
buf ( n195678 , n20391 );
not ( n28402 , n195678 );
or ( n28403 , n28400 , n28402 );
buf ( n195681 , n20396 );
buf ( n195682 , n848 );
buf ( n195683 , n888 );
xor ( n28407 , n195682 , n195683 );
buf ( n195685 , n28407 );
buf ( n195686 , n195685 );
nand ( n28410 , n195681 , n195686 );
buf ( n195688 , n28410 );
buf ( n195689 , n195688 );
nand ( n28413 , n28403 , n195689 );
buf ( n195691 , n28413 );
xor ( n28415 , n195675 , n195691 );
buf ( n195693 , n195428 );
not ( n28417 , n195693 );
buf ( n195695 , n186569 );
not ( n28419 , n195695 );
or ( n28420 , n28417 , n28419 );
buf ( n195698 , n186575 );
buf ( n195699 , n858 );
buf ( n195700 , n878 );
xor ( n28424 , n195699 , n195700 );
buf ( n195702 , n28424 );
buf ( n195703 , n195702 );
nand ( n28427 , n195698 , n195703 );
buf ( n195705 , n28427 );
buf ( n195706 , n195705 );
nand ( n28430 , n28420 , n195706 );
buf ( n195708 , n28430 );
xnor ( n28432 , n28415 , n195708 );
buf ( n195710 , n28432 );
xor ( n28434 , n28379 , n195710 );
buf ( n195712 , n28434 );
buf ( n195713 , n195712 );
xor ( n28437 , n195598 , n195713 );
buf ( n195715 , n28236 );
not ( n28439 , n195715 );
buf ( n195717 , n28231 );
not ( n28441 , n195717 );
or ( n28442 , n28439 , n28441 );
buf ( n195720 , n28236 );
buf ( n195721 , n28231 );
or ( n28445 , n195720 , n195721 );
buf ( n195723 , n28290 );
nand ( n28447 , n28445 , n195723 );
buf ( n195725 , n28447 );
buf ( n195726 , n195725 );
nand ( n28450 , n28442 , n195726 );
buf ( n195728 , n28450 );
buf ( n195729 , n195728 );
buf ( n195730 , n27682 );
not ( n28454 , n195730 );
buf ( n195732 , n26567 );
not ( n28456 , n195732 );
or ( n28457 , n28454 , n28456 );
buf ( n195735 , n19943 );
buf ( n195736 , n854 );
buf ( n195737 , n882 );
xor ( n28461 , n195736 , n195737 );
buf ( n195739 , n28461 );
buf ( n195740 , n195739 );
nand ( n28464 , n195735 , n195740 );
buf ( n195742 , n28464 );
buf ( n195743 , n195742 );
nand ( n28467 , n28457 , n195743 );
buf ( n195745 , n28467 );
buf ( n195746 , n195745 );
buf ( n195747 , n863 );
buf ( n195748 , n875 );
or ( n28472 , n195747 , n195748 );
buf ( n195750 , n876 );
nand ( n28474 , n28472 , n195750 );
buf ( n195752 , n28474 );
buf ( n195753 , n195752 );
buf ( n195754 , n863 );
buf ( n195755 , n875 );
nand ( n28479 , n195754 , n195755 );
buf ( n195757 , n28479 );
buf ( n195758 , n195757 );
buf ( n195759 , n874 );
and ( n28483 , n195753 , n195758 , n195759 );
buf ( n195761 , n28483 );
buf ( n195762 , n195761 );
buf ( n195763 , n195478 );
not ( n28487 , n195763 );
buf ( n195765 , n190485 );
not ( n28489 , n195765 );
or ( n28490 , n28487 , n28489 );
buf ( n195768 , n190128 );
buf ( n195769 , n844 );
buf ( n195770 , n892 );
xor ( n28494 , n195769 , n195770 );
buf ( n195772 , n28494 );
buf ( n195773 , n195772 );
nand ( n28497 , n195768 , n195773 );
buf ( n195775 , n28497 );
buf ( n195776 , n195775 );
nand ( n28500 , n28490 , n195776 );
buf ( n195778 , n28500 );
buf ( n195779 , n195778 );
xor ( n28503 , n195762 , n195779 );
buf ( n195781 , n28503 );
buf ( n195782 , n195781 );
xor ( n28506 , n195746 , n195782 );
not ( n28507 , n195452 );
not ( n28508 , n195484 );
or ( n28509 , n28507 , n28508 );
not ( n28510 , n195490 );
not ( n28511 , n195455 );
or ( n28512 , n28510 , n28511 );
nand ( n28513 , n28512 , n195434 );
nand ( n28514 , n28509 , n28513 );
buf ( n195792 , n28514 );
xor ( n28516 , n28506 , n195792 );
buf ( n195794 , n28516 );
buf ( n195795 , n195794 );
xor ( n28519 , n195729 , n195795 );
xor ( n28520 , n195319 , n195336 );
and ( n28521 , n28520 , n195354 );
and ( n28522 , n195319 , n195336 );
or ( n28523 , n28521 , n28522 );
buf ( n195801 , n28523 );
buf ( n195802 , n195801 );
xor ( n28526 , n195374 , n195395 );
and ( n28527 , n28526 , n195414 );
and ( n28528 , n195374 , n195395 );
or ( n28529 , n28527 , n28528 );
buf ( n195807 , n28529 );
buf ( n195808 , n195807 );
xor ( n28532 , n195802 , n195808 );
buf ( n195810 , n195328 );
not ( n28534 , n195810 );
buf ( n195812 , n21330 );
not ( n28536 , n195812 );
or ( n28537 , n28534 , n28536 );
buf ( n195815 , n842 );
buf ( n195816 , n894 );
xor ( n28540 , n195815 , n195816 );
buf ( n195818 , n28540 );
buf ( n195819 , n195818 );
buf ( n195820 , n895 );
nand ( n28544 , n195819 , n195820 );
buf ( n195822 , n28544 );
buf ( n195823 , n195822 );
nand ( n28547 , n28537 , n195823 );
buf ( n195825 , n28547 );
buf ( n195826 , n195825 );
buf ( n195827 , n195367 );
not ( n28551 , n195827 );
buf ( n195829 , n188751 );
not ( n28553 , n195829 );
or ( n28554 , n28551 , n28553 );
buf ( n195832 , n20902 );
buf ( n195833 , n846 );
buf ( n195834 , n890 );
xor ( n28558 , n195833 , n195834 );
buf ( n195836 , n28558 );
buf ( n195837 , n195836 );
nand ( n28561 , n195832 , n195837 );
buf ( n195839 , n28561 );
buf ( n195840 , n195839 );
nand ( n28564 , n28554 , n195840 );
buf ( n195842 , n28564 );
buf ( n195843 , n195842 );
xor ( n28567 , n195826 , n195843 );
buf ( n195845 , n194993 );
not ( n28569 , n195845 );
buf ( n195847 , n192332 );
not ( n28571 , n195847 );
or ( n28572 , n28569 , n28571 );
buf ( n195850 , n190543 );
buf ( n195851 , n852 );
buf ( n195852 , n884 );
xor ( n28576 , n195851 , n195852 );
buf ( n195854 , n28576 );
buf ( n195855 , n195854 );
nand ( n28579 , n195850 , n195855 );
buf ( n195857 , n28579 );
buf ( n195858 , n195857 );
nand ( n28582 , n28572 , n195858 );
buf ( n195860 , n28582 );
buf ( n195861 , n195860 );
xor ( n28585 , n28567 , n195861 );
buf ( n195863 , n28585 );
buf ( n195864 , n195863 );
xor ( n28588 , n28532 , n195864 );
buf ( n195866 , n28588 );
buf ( n195867 , n195866 );
xor ( n28591 , n28519 , n195867 );
buf ( n195869 , n28591 );
buf ( n195870 , n195869 );
xor ( n28594 , n28437 , n195870 );
buf ( n195872 , n28594 );
buf ( n195873 , n195872 );
and ( n28597 , n28315 , n195873 );
and ( n28598 , n195314 , n195591 );
or ( n28599 , n28597 , n28598 );
buf ( n195877 , n28599 );
buf ( n28601 , n195877 );
buf ( n195879 , n863 );
buf ( n195880 , n879 );
or ( n28604 , n195879 , n195880 );
buf ( n195882 , n880 );
nand ( n28606 , n28604 , n195882 );
buf ( n195884 , n28606 );
buf ( n195885 , n195884 );
buf ( n195886 , n863 );
buf ( n195887 , n879 );
nand ( n28611 , n195886 , n195887 );
buf ( n195889 , n28611 );
buf ( n195890 , n195889 );
buf ( n195891 , n878 );
and ( n28615 , n195885 , n195890 , n195891 );
buf ( n195893 , n28615 );
buf ( n195894 , n195893 );
buf ( n195895 , n193781 );
not ( n28619 , n195895 );
buf ( n195897 , n22809 );
not ( n28621 , n195897 );
or ( n28622 , n28619 , n28621 );
buf ( n195900 , n195024 );
buf ( n195901 , n895 );
nand ( n28625 , n195900 , n195901 );
buf ( n195903 , n28625 );
buf ( n195904 , n195903 );
nand ( n28628 , n28622 , n195904 );
buf ( n195906 , n28628 );
buf ( n195907 , n195906 );
and ( n28631 , n195894 , n195907 );
buf ( n195909 , n28631 );
buf ( n195910 , n195909 );
not ( n28634 , n195910 );
xor ( n28635 , n882 , n858 );
buf ( n195913 , n28635 );
not ( n28637 , n195913 );
buf ( n195915 , n19613 );
not ( n28639 , n195915 );
or ( n28640 , n28637 , n28639 );
buf ( n195918 , n26571 );
buf ( n195919 , n195270 );
nand ( n28643 , n195918 , n195919 );
buf ( n195921 , n28643 );
buf ( n195922 , n195921 );
nand ( n28646 , n28640 , n195922 );
buf ( n195924 , n28646 );
not ( n28648 , n195924 );
buf ( n195926 , n28648 );
nand ( n28650 , n28634 , n195926 );
buf ( n195928 , n28650 );
buf ( n195929 , n195928 );
not ( n28653 , n195929 );
buf ( n195931 , n193743 );
not ( n28655 , n195931 );
buf ( n195933 , n190454 );
not ( n28657 , n195933 );
or ( n28658 , n28655 , n28657 );
buf ( n195936 , n195051 );
not ( n28660 , n195936 );
buf ( n195938 , n20396 );
nand ( n28662 , n28660 , n195938 );
buf ( n195940 , n28662 );
buf ( n195941 , n195940 );
nand ( n28665 , n28658 , n195941 );
buf ( n195943 , n28665 );
buf ( n195944 , n195943 );
not ( n28668 , n195944 );
buf ( n195946 , n193722 );
not ( n28670 , n195946 );
buf ( n195948 , n186924 );
not ( n28672 , n195948 );
or ( n28673 , n28670 , n28672 );
buf ( n195951 , n22304 );
buf ( n195952 , n195101 );
nand ( n28676 , n195951 , n195952 );
buf ( n195954 , n28676 );
buf ( n195955 , n195954 );
nand ( n28679 , n28673 , n195955 );
buf ( n195957 , n28679 );
buf ( n195958 , n195957 );
not ( n28682 , n195958 );
or ( n28683 , n28668 , n28682 );
buf ( n195961 , n195957 );
buf ( n195962 , n195943 );
or ( n28686 , n195961 , n195962 );
buf ( n195964 , n863 );
buf ( n195965 , n878 );
xor ( n28689 , n195964 , n195965 );
buf ( n195967 , n28689 );
buf ( n195968 , n195967 );
not ( n28692 , n195968 );
buf ( n195970 , n186789 );
not ( n28694 , n195970 );
or ( n28695 , n28692 , n28694 );
buf ( n195973 , n186575 );
buf ( n195974 , n195113 );
nand ( n28698 , n195973 , n195974 );
buf ( n195976 , n28698 );
buf ( n195977 , n195976 );
nand ( n28701 , n28695 , n195977 );
buf ( n195979 , n28701 );
buf ( n195980 , n195979 );
nand ( n28704 , n28686 , n195980 );
buf ( n195982 , n28704 );
buf ( n195983 , n195982 );
nand ( n28707 , n28683 , n195983 );
buf ( n195985 , n28707 );
buf ( n195986 , n195985 );
not ( n28710 , n195986 );
or ( n28711 , n28653 , n28710 );
buf ( n195989 , n195924 );
buf ( n195990 , n195909 );
nand ( n28714 , n195989 , n195990 );
buf ( n195992 , n28714 );
buf ( n195993 , n195992 );
nand ( n28717 , n28711 , n195993 );
buf ( n195995 , n28717 );
buf ( n195996 , n195995 );
xor ( n28720 , n195020 , n195071 );
xor ( n28721 , n28720 , n195135 );
buf ( n195999 , n28721 );
buf ( n196000 , n195999 );
xor ( n28724 , n195996 , n196000 );
buf ( n196002 , n195563 );
buf ( n196003 , n195529 );
xor ( n28727 , n196002 , n196003 );
buf ( n196005 , n28727 );
buf ( n196006 , n196005 );
buf ( n196007 , n195542 );
xor ( n28731 , n196006 , n196007 );
buf ( n196009 , n28731 );
buf ( n196010 , n196009 );
and ( n28734 , n28724 , n196010 );
and ( n28735 , n195996 , n196000 );
or ( n28736 , n28734 , n28735 );
buf ( n196014 , n28736 );
buf ( n196015 , n196014 );
buf ( n196016 , n193853 );
not ( n28740 , n196016 );
buf ( n196018 , n19613 );
not ( n28742 , n196018 );
or ( n28743 , n28740 , n28742 );
buf ( n196021 , n26571 );
buf ( n196022 , n28635 );
nand ( n28746 , n196021 , n196022 );
buf ( n196024 , n28746 );
buf ( n196025 , n196024 );
nand ( n28749 , n28743 , n196025 );
buf ( n196027 , n28749 );
buf ( n196028 , n196027 );
xor ( n28752 , n195894 , n195907 );
buf ( n196030 , n28752 );
buf ( n196031 , n196030 );
or ( n28755 , n196028 , n196031 );
buf ( n196033 , n193830 );
not ( n28757 , n196033 );
buf ( n196035 , n192332 );
not ( n28759 , n196035 );
or ( n28760 , n28757 , n28759 );
buf ( n196038 , n190543 );
buf ( n196039 , n195233 );
nand ( n28763 , n196038 , n196039 );
buf ( n196041 , n28763 );
buf ( n196042 , n196041 );
nand ( n28766 , n28760 , n196042 );
buf ( n196044 , n28766 );
buf ( n196045 , n196044 );
nand ( n28769 , n28755 , n196045 );
buf ( n196047 , n28769 );
buf ( n196048 , n196047 );
buf ( n196049 , n196030 );
buf ( n196050 , n196027 );
nand ( n28774 , n196049 , n196050 );
buf ( n196052 , n28774 );
buf ( n196053 , n196052 );
nand ( n28777 , n196048 , n196053 );
buf ( n196055 , n28777 );
buf ( n196056 , n196055 );
xor ( n28780 , n195087 , n195108 );
xor ( n28781 , n28780 , n195130 );
buf ( n196059 , n28781 );
buf ( n196060 , n196059 );
xor ( n28784 , n196056 , n196060 );
buf ( n196062 , n195909 );
buf ( n196063 , n28648 );
xor ( n28787 , n196062 , n196063 );
buf ( n196065 , n28787 );
buf ( n196066 , n196065 );
not ( n28790 , n196066 );
buf ( n196068 , n195985 );
not ( n28792 , n196068 );
or ( n28793 , n28790 , n28792 );
buf ( n196071 , n195985 );
buf ( n196072 , n196065 );
or ( n28796 , n196071 , n196072 );
nand ( n28797 , n28793 , n28796 );
buf ( n196075 , n28797 );
buf ( n196076 , n196075 );
and ( n28800 , n28784 , n196076 );
and ( n28801 , n196056 , n196060 );
or ( n28802 , n28800 , n28801 );
buf ( n196080 , n28802 );
buf ( n196081 , n196080 );
not ( n28805 , n196081 );
buf ( n196083 , n28805 );
buf ( n196084 , n196083 );
not ( n28808 , n196084 );
buf ( n196086 , n28808 );
buf ( n196087 , n196086 );
not ( n28811 , n196087 );
xor ( n28812 , n195037 , n195042 );
xor ( n28813 , n28812 , n195066 );
buf ( n196091 , n28813 );
buf ( n196092 , n196091 );
buf ( n196093 , n193764 );
not ( n28817 , n196093 );
buf ( n196095 , n190485 );
not ( n28819 , n196095 );
or ( n28820 , n28817 , n28819 );
buf ( n196098 , n190128 );
buf ( n196099 , n27796 );
nand ( n28823 , n196098 , n196099 );
buf ( n196101 , n28823 );
buf ( n196102 , n196101 );
nand ( n28826 , n28820 , n196102 );
buf ( n196104 , n28826 );
not ( n28828 , n196104 );
buf ( n196106 , n28828 );
not ( n28830 , n196106 );
buf ( n196108 , n193810 );
not ( n28832 , n196108 );
buf ( n196110 , n188751 );
not ( n28834 , n196110 );
or ( n28835 , n28832 , n28834 );
buf ( n196113 , n20902 );
buf ( n196114 , n195189 );
nand ( n28838 , n196113 , n196114 );
buf ( n196116 , n28838 );
buf ( n196117 , n196116 );
nand ( n28841 , n28835 , n196117 );
buf ( n196119 , n28841 );
buf ( n196120 , n196119 );
not ( n28844 , n196120 );
buf ( n196122 , n28844 );
buf ( n196123 , n196122 );
not ( n28847 , n196123 );
or ( n28848 , n28830 , n28847 );
buf ( n196126 , n193706 );
not ( n28850 , n196126 );
buf ( n196128 , n190337 );
not ( n28852 , n196128 );
or ( n28853 , n28850 , n28852 );
buf ( n196131 , n20558 );
buf ( n196132 , n195210 );
nand ( n28856 , n196131 , n196132 );
buf ( n196134 , n28856 );
buf ( n196135 , n196134 );
nand ( n28859 , n28853 , n196135 );
buf ( n196137 , n28859 );
buf ( n196138 , n196137 );
nand ( n28862 , n28848 , n196138 );
buf ( n196140 , n28862 );
buf ( n196141 , n196140 );
buf ( n196142 , n196119 );
not ( n28866 , n28828 );
buf ( n196144 , n28866 );
nand ( n28868 , n196142 , n196144 );
buf ( n196146 , n28868 );
buf ( n196147 , n196146 );
nand ( n28871 , n196141 , n196147 );
buf ( n196149 , n28871 );
buf ( n196150 , n196149 );
xor ( n28874 , n196092 , n196150 );
buf ( n196152 , n195249 );
not ( n28876 , n196152 );
buf ( n196154 , n28876 );
buf ( n196155 , n196154 );
not ( n28879 , n196155 );
xor ( n28880 , n195205 , n195226 );
buf ( n196158 , n28880 );
not ( n28882 , n196158 );
or ( n28883 , n28879 , n28882 );
buf ( n196161 , n28880 );
buf ( n196162 , n196154 );
or ( n28886 , n196161 , n196162 );
nand ( n28887 , n28883 , n28886 );
buf ( n196165 , n28887 );
buf ( n196166 , n196165 );
and ( n28890 , n28874 , n196166 );
and ( n28891 , n196092 , n196150 );
or ( n28892 , n28890 , n28891 );
buf ( n196170 , n28892 );
buf ( n196171 , n196170 );
not ( n28895 , n196171 );
or ( n28896 , n28811 , n28895 );
buf ( n196174 , n196170 );
buf ( n196175 , n196086 );
or ( n28899 , n196174 , n196175 );
xor ( n28900 , n27974 , n195297 );
xor ( n28901 , n28900 , n27907 );
buf ( n196179 , n28901 );
nand ( n28903 , n28899 , n196179 );
buf ( n196181 , n28903 );
buf ( n196182 , n196181 );
nand ( n28906 , n28896 , n196182 );
buf ( n196184 , n28906 );
buf ( n196185 , n196184 );
xor ( n28909 , n196015 , n196185 );
buf ( n196187 , n195497 );
not ( n28911 , n196187 );
buf ( n196189 , n195577 );
not ( n28913 , n196189 );
and ( n28914 , n28911 , n28913 );
buf ( n196192 , n195497 );
buf ( n196193 , n195577 );
and ( n28917 , n196192 , n196193 );
nor ( n28918 , n28914 , n28917 );
buf ( n196196 , n28918 );
buf ( n196197 , n196196 );
not ( n28921 , n196197 );
buf ( n196199 , n195582 );
not ( n28923 , n196199 );
or ( n28924 , n28921 , n28923 );
buf ( n196202 , n196196 );
buf ( n196203 , n195582 );
or ( n28927 , n196202 , n196203 );
nand ( n28928 , n28924 , n28927 );
buf ( n196206 , n28928 );
buf ( n196207 , n196206 );
xor ( n28931 , n28909 , n196207 );
buf ( n196209 , n28931 );
buf ( n28933 , n196209 );
xor ( n28934 , n195996 , n196000 );
xor ( n28935 , n28934 , n196010 );
buf ( n196213 , n28935 );
buf ( n196214 , n196213 );
not ( n28938 , n26511 );
nand ( n28939 , n28938 , n26509 );
not ( n28940 , n26510 );
not ( n28941 , n26514 );
or ( n28942 , n28940 , n28941 );
nand ( n28943 , n28942 , n193770 );
nand ( n28944 , n28939 , n28943 );
xor ( n28945 , n193816 , n193836 );
and ( n28946 , n28945 , n193859 );
and ( n28947 , n193816 , n193836 );
or ( n28948 , n28946 , n28947 );
xor ( n28949 , n28944 , n28948 );
buf ( n196227 , n26431 );
not ( n28951 , n196227 );
buf ( n196229 , n193728 );
not ( n28953 , n196229 );
or ( n28954 , n28951 , n28953 );
buf ( n196232 , n26431 );
buf ( n196233 , n193728 );
or ( n28957 , n196232 , n196233 );
buf ( n196235 , n193749 );
nand ( n28959 , n28957 , n196235 );
buf ( n196237 , n28959 );
buf ( n196238 , n196237 );
nand ( n28962 , n28954 , n196238 );
buf ( n196240 , n28962 );
and ( n28964 , n28949 , n196240 );
and ( n28965 , n28944 , n28948 );
or ( n28966 , n28964 , n28965 );
buf ( n196244 , n28966 );
xor ( n28968 , n196092 , n196150 );
xor ( n28969 , n28968 , n196166 );
buf ( n196247 , n28969 );
buf ( n196248 , n196247 );
xor ( n28972 , n196244 , n196248 );
buf ( n28973 , n196044 );
not ( n28974 , n28973 );
xor ( n28975 , n196027 , n196030 );
not ( n28976 , n28975 );
or ( n28977 , n28974 , n28976 );
or ( n28978 , n28975 , n28973 );
nand ( n28979 , n28977 , n28978 );
buf ( n196257 , n28979 );
not ( n28981 , n196257 );
xor ( n28982 , n195957 , n195943 );
xnor ( n28983 , n28982 , n195979 );
buf ( n196261 , n28983 );
not ( n28985 , n196261 );
or ( n28986 , n28981 , n28985 );
xor ( n28987 , n196122 , n196137 );
xnor ( n28988 , n28987 , n28866 );
buf ( n196266 , n28988 );
nand ( n28990 , n28986 , n196266 );
buf ( n196268 , n28990 );
buf ( n196269 , n196268 );
buf ( n196270 , n28983 );
not ( n28994 , n196270 );
not ( n28995 , n28979 );
buf ( n196273 , n28995 );
nand ( n28997 , n28994 , n196273 );
buf ( n196275 , n28997 );
buf ( n196276 , n196275 );
nand ( n29000 , n196269 , n196276 );
buf ( n196278 , n29000 );
buf ( n196279 , n196278 );
and ( n29003 , n28972 , n196279 );
and ( n29004 , n196244 , n196248 );
or ( n29005 , n29003 , n29004 );
buf ( n196283 , n29005 );
buf ( n196284 , n196283 );
xor ( n29008 , n196214 , n196284 );
xor ( n29009 , n196083 , n196170 );
buf ( n196287 , n28901 );
not ( n29011 , n196287 );
buf ( n196289 , n29011 );
and ( n29013 , n29009 , n196289 );
not ( n29014 , n29009 );
and ( n29015 , n29014 , n28901 );
nor ( n29016 , n29013 , n29015 );
buf ( n196294 , n29016 );
and ( n29018 , n29008 , n196294 );
and ( n29019 , n196214 , n196284 );
or ( n29020 , n29018 , n29019 );
buf ( n196298 , n29020 );
buf ( n29022 , n196298 );
buf ( n196300 , n190548 );
not ( n29024 , n196300 );
buf ( n196302 , n22809 );
not ( n29026 , n196302 );
or ( n29027 , n29024 , n29026 );
buf ( n196305 , n862 );
buf ( n196306 , n894 );
xor ( n29030 , n196305 , n196306 );
buf ( n196308 , n29030 );
buf ( n196309 , n196308 );
buf ( n196310 , n895 );
nand ( n29034 , n196309 , n196310 );
buf ( n196312 , n29034 );
buf ( n196313 , n196312 );
nand ( n29037 , n29027 , n196313 );
buf ( n196315 , n29037 );
buf ( n29039 , n196315 );
buf ( n29040 , n177299 );
xor ( n29041 , n866 , n839 );
buf ( n196319 , n29041 );
not ( n29043 , n196319 );
buf ( n196321 , n186241 );
not ( n29045 , n196321 );
or ( n29046 , n29043 , n29045 );
buf ( n196324 , n186254 );
buf ( n196325 , n838 );
buf ( n196326 , n866 );
xor ( n29050 , n196325 , n196326 );
buf ( n196328 , n29050 );
buf ( n196329 , n196328 );
nand ( n29053 , n196324 , n196329 );
buf ( n196331 , n29053 );
buf ( n196332 , n196331 );
nand ( n29056 , n29046 , n196332 );
buf ( n196334 , n29056 );
buf ( n196335 , n196334 );
buf ( n196336 , n835 );
buf ( n196337 , n870 );
xor ( n29061 , n196336 , n196337 );
buf ( n196339 , n29061 );
buf ( n196340 , n196339 );
not ( n29064 , n196340 );
buf ( n196342 , n186435 );
not ( n29066 , n196342 );
or ( n29067 , n29064 , n29066 );
buf ( n196345 , n186444 );
buf ( n196346 , n834 );
buf ( n196347 , n870 );
xor ( n29071 , n196346 , n196347 );
buf ( n196349 , n29071 );
buf ( n196350 , n196349 );
nand ( n29074 , n196345 , n196350 );
buf ( n196352 , n29074 );
buf ( n196353 , n196352 );
nand ( n29077 , n29067 , n196353 );
buf ( n196355 , n29077 );
buf ( n196356 , n196355 );
xor ( n29080 , n196335 , n196356 );
buf ( n196358 , n864 );
buf ( n196359 , n841 );
xor ( n29083 , n196358 , n196359 );
buf ( n196361 , n29083 );
buf ( n196362 , n196361 );
not ( n29086 , n196362 );
buf ( n196364 , n186640 );
not ( n29088 , n196364 );
or ( n29089 , n29086 , n29088 );
buf ( n196367 , n186340 );
buf ( n196368 , n864 );
buf ( n196369 , n840 );
xor ( n29093 , n196368 , n196369 );
buf ( n196371 , n29093 );
buf ( n196372 , n196371 );
nand ( n29096 , n196367 , n196372 );
buf ( n196374 , n29096 );
buf ( n196375 , n196374 );
nand ( n29099 , n29089 , n196375 );
buf ( n196377 , n29099 );
buf ( n196378 , n196377 );
and ( n29102 , n29080 , n196378 );
and ( n29103 , n196335 , n196356 );
or ( n29104 , n29102 , n29103 );
buf ( n196382 , n29104 );
buf ( n196383 , n196382 );
xor ( n29107 , n868 , n837 );
buf ( n196385 , n29107 );
not ( n29109 , n196385 );
buf ( n196387 , n186197 );
not ( n29111 , n196387 );
or ( n29112 , n29109 , n29111 );
buf ( n196390 , n186208 );
buf ( n196391 , n836 );
buf ( n196392 , n868 );
xor ( n29116 , n196391 , n196392 );
buf ( n196394 , n29116 );
buf ( n196395 , n196394 );
nand ( n29119 , n196390 , n196395 );
buf ( n196397 , n29119 );
buf ( n196398 , n196397 );
nand ( n29122 , n29112 , n196398 );
buf ( n196400 , n29122 );
buf ( n196401 , n196400 );
buf ( n196402 , n186294 );
not ( n29126 , n196402 );
buf ( n196404 , n186287 );
not ( n29128 , n196404 );
buf ( n196406 , n29128 );
buf ( n196407 , n196406 );
not ( n29131 , n196407 );
or ( n29132 , n29126 , n29131 );
buf ( n196410 , n874 );
nand ( n29134 , n29132 , n196410 );
buf ( n196412 , n29134 );
buf ( n196413 , n196412 );
xor ( n29137 , n196401 , n196413 );
buf ( n196415 , n833 );
buf ( n196416 , n872 );
xor ( n29140 , n196415 , n196416 );
buf ( n196418 , n29140 );
buf ( n196419 , n196418 );
not ( n29143 , n196419 );
buf ( n196421 , n19260 );
not ( n29145 , n196421 );
or ( n29146 , n29143 , n29145 );
buf ( n196424 , n19265 );
buf ( n196425 , n832 );
buf ( n196426 , n872 );
xor ( n29150 , n196425 , n196426 );
buf ( n196428 , n29150 );
buf ( n196429 , n196428 );
nand ( n29153 , n196424 , n196429 );
buf ( n196431 , n29153 );
buf ( n196432 , n196431 );
nand ( n29156 , n29146 , n196432 );
buf ( n196434 , n29156 );
buf ( n196435 , n196434 );
and ( n29159 , n29137 , n196435 );
and ( n29160 , n196401 , n196413 );
or ( n29161 , n29159 , n29160 );
buf ( n196439 , n29161 );
buf ( n196440 , n196439 );
xor ( n29164 , n196383 , n196440 );
buf ( n196442 , n196328 );
not ( n29166 , n196442 );
buf ( n196444 , n186241 );
not ( n29168 , n196444 );
buf ( n196446 , n29168 );
buf ( n196447 , n196446 );
not ( n29171 , n196447 );
buf ( n196449 , n29171 );
buf ( n196450 , n196449 );
not ( n29174 , n196450 );
or ( n29175 , n29166 , n29174 );
buf ( n196453 , n186254 );
buf ( n196454 , n837 );
buf ( n196455 , n866 );
xor ( n29179 , n196454 , n196455 );
buf ( n196457 , n29179 );
buf ( n196458 , n196457 );
nand ( n29182 , n196453 , n196458 );
buf ( n196460 , n29182 );
buf ( n196461 , n196460 );
nand ( n29185 , n29175 , n196461 );
buf ( n196463 , n29185 );
buf ( n196464 , n196428 );
not ( n29188 , n196464 );
buf ( n196466 , n19260 );
not ( n29190 , n196466 );
or ( n29191 , n29188 , n29190 );
buf ( n196469 , n19264 );
buf ( n196470 , n872 );
nand ( n29194 , n196469 , n196470 );
buf ( n196472 , n29194 );
buf ( n196473 , n196472 );
nand ( n29197 , n29191 , n196473 );
buf ( n196475 , n29197 );
xnor ( n29199 , n196463 , n196475 );
buf ( n196477 , n29199 );
buf ( n196478 , n196371 );
not ( n29202 , n196478 );
buf ( n196480 , n186640 );
not ( n29204 , n196480 );
or ( n29205 , n29202 , n29204 );
buf ( n196483 , n186340 );
buf ( n196484 , n864 );
buf ( n196485 , n839 );
xor ( n29209 , n196484 , n196485 );
buf ( n196487 , n29209 );
buf ( n196488 , n196487 );
nand ( n29212 , n196483 , n196488 );
buf ( n196490 , n29212 );
buf ( n196491 , n196490 );
nand ( n29215 , n29205 , n196491 );
buf ( n196493 , n29215 );
buf ( n196494 , n196493 );
xnor ( n29218 , n196477 , n196494 );
buf ( n196496 , n29218 );
buf ( n196497 , n196496 );
xor ( n29221 , n29164 , n196497 );
buf ( n196499 , n29221 );
buf ( n196500 , n196499 );
and ( n29224 , n196358 , n196359 );
buf ( n196502 , n29224 );
buf ( n196503 , n196502 );
buf ( n196504 , n196394 );
not ( n29228 , n196504 );
buf ( n196506 , n186197 );
not ( n29230 , n196506 );
or ( n29231 , n29228 , n29230 );
buf ( n196509 , n186208 );
buf ( n196510 , n835 );
buf ( n196511 , n868 );
xor ( n29235 , n196510 , n196511 );
buf ( n196513 , n29235 );
buf ( n196514 , n196513 );
nand ( n29238 , n196509 , n196514 );
buf ( n196516 , n29238 );
buf ( n196517 , n196516 );
nand ( n29241 , n29231 , n196517 );
buf ( n196519 , n29241 );
buf ( n196520 , n196519 );
xor ( n29244 , n196503 , n196520 );
buf ( n196522 , n196349 );
not ( n29246 , n196522 );
buf ( n196524 , n186435 );
not ( n29248 , n196524 );
or ( n29249 , n29246 , n29248 );
buf ( n196527 , n186444 );
buf ( n196528 , n870 );
buf ( n196529 , n833 );
xor ( n29253 , n196528 , n196529 );
buf ( n196531 , n29253 );
buf ( n196532 , n196531 );
nand ( n29256 , n196527 , n196532 );
buf ( n196534 , n29256 );
buf ( n196535 , n196534 );
nand ( n29259 , n29249 , n196535 );
buf ( n196537 , n29259 );
buf ( n196538 , n196537 );
not ( n29262 , n196538 );
buf ( n196540 , n29262 );
buf ( n196541 , n196540 );
xor ( n29265 , n29244 , n196541 );
buf ( n196543 , n29265 );
buf ( n196544 , n196543 );
buf ( n196545 , n864 );
buf ( n196546 , n842 );
and ( n29270 , n196545 , n196546 );
buf ( n196548 , n29270 );
buf ( n196549 , n196548 );
buf ( n196550 , n832 );
buf ( n196551 , n874 );
xor ( n29275 , n196550 , n196551 );
buf ( n196553 , n29275 );
buf ( n196554 , n196553 );
not ( n29278 , n196554 );
buf ( n196556 , n186287 );
not ( n29280 , n196556 );
or ( n29281 , n29278 , n29280 );
buf ( n196559 , n186297 );
buf ( n196560 , n874 );
nand ( n29284 , n196559 , n196560 );
buf ( n196562 , n29284 );
buf ( n196563 , n196562 );
nand ( n29287 , n29281 , n196563 );
buf ( n196565 , n29287 );
buf ( n196566 , n196565 );
xor ( n29290 , n196549 , n196566 );
xor ( n29291 , n866 , n840 );
buf ( n196569 , n29291 );
not ( n29293 , n196569 );
buf ( n196571 , n186241 );
not ( n29295 , n196571 );
or ( n29296 , n29293 , n29295 );
buf ( n196574 , n186254 );
buf ( n196575 , n29041 );
nand ( n29299 , n196574 , n196575 );
buf ( n196577 , n29299 );
buf ( n196578 , n196577 );
nand ( n29302 , n29296 , n196578 );
buf ( n196580 , n29302 );
buf ( n196581 , n196580 );
xor ( n29305 , n868 , n838 );
buf ( n196583 , n29305 );
not ( n29307 , n196583 );
buf ( n196585 , n186197 );
not ( n29309 , n196585 );
or ( n29310 , n29307 , n29309 );
buf ( n196588 , n186208 );
buf ( n196589 , n29107 );
nand ( n29313 , n196588 , n196589 );
buf ( n196591 , n29313 );
buf ( n196592 , n196591 );
nand ( n29316 , n29310 , n196592 );
buf ( n196594 , n29316 );
buf ( n196595 , n196594 );
nand ( n29319 , n196581 , n196595 );
buf ( n196597 , n29319 );
buf ( n196598 , n196597 );
buf ( n196599 , n196580 );
buf ( n196600 , n196594 );
or ( n29324 , n196599 , n196600 );
buf ( n196602 , n834 );
buf ( n196603 , n872 );
xor ( n29327 , n196602 , n196603 );
buf ( n196605 , n29327 );
buf ( n196606 , n196605 );
not ( n29330 , n196606 );
buf ( n196608 , n19260 );
not ( n29332 , n196608 );
or ( n29333 , n29330 , n29332 );
buf ( n196611 , n19265 );
buf ( n196612 , n196418 );
nand ( n29336 , n196611 , n196612 );
buf ( n196614 , n29336 );
buf ( n196615 , n196614 );
nand ( n29339 , n29333 , n196615 );
buf ( n196617 , n29339 );
buf ( n196618 , n196617 );
nand ( n29342 , n29324 , n196618 );
buf ( n196620 , n29342 );
buf ( n196621 , n196620 );
nand ( n29345 , n196598 , n196621 );
buf ( n196623 , n29345 );
buf ( n196624 , n196623 );
and ( n29348 , n29290 , n196624 );
and ( n29349 , n196549 , n196566 );
or ( n29350 , n29348 , n29349 );
buf ( n196628 , n29350 );
buf ( n196629 , n196628 );
xor ( n29353 , n196544 , n196629 );
buf ( n196631 , n843 );
buf ( n196632 , n864 );
and ( n29356 , n196631 , n196632 );
buf ( n196634 , n29356 );
buf ( n196635 , n196634 );
xor ( n29359 , n196545 , n196546 );
buf ( n196637 , n29359 );
buf ( n196638 , n196637 );
not ( n29362 , n196638 );
buf ( n196640 , n186640 );
not ( n29364 , n196640 );
or ( n29365 , n29362 , n29364 );
buf ( n196643 , n186340 );
buf ( n196644 , n196361 );
nand ( n29368 , n196643 , n196644 );
buf ( n196646 , n29368 );
buf ( n196647 , n196646 );
nand ( n29371 , n29365 , n196647 );
buf ( n196649 , n29371 );
buf ( n196650 , n196649 );
xor ( n29374 , n196635 , n196650 );
buf ( n196652 , n836 );
buf ( n196653 , n870 );
xor ( n29377 , n196652 , n196653 );
buf ( n196655 , n29377 );
buf ( n196656 , n196655 );
not ( n29380 , n196656 );
buf ( n196658 , n186435 );
not ( n29382 , n196658 );
or ( n29383 , n29380 , n29382 );
buf ( n196661 , n186444 );
buf ( n196662 , n196339 );
nand ( n29386 , n196661 , n196662 );
buf ( n196664 , n29386 );
buf ( n196665 , n196664 );
nand ( n29389 , n29383 , n196665 );
buf ( n196667 , n29389 );
buf ( n196668 , n196667 );
and ( n29392 , n29374 , n196668 );
and ( n29393 , n196635 , n196650 );
or ( n29394 , n29392 , n29393 );
buf ( n196672 , n29394 );
buf ( n196673 , n196672 );
xor ( n29397 , n196401 , n196413 );
xor ( n29398 , n29397 , n196435 );
buf ( n196676 , n29398 );
buf ( n196677 , n196676 );
xor ( n29401 , n196673 , n196677 );
xor ( n29402 , n196335 , n196356 );
xor ( n29403 , n29402 , n196378 );
buf ( n196681 , n29403 );
buf ( n196682 , n196681 );
and ( n29406 , n29401 , n196682 );
and ( n29407 , n196673 , n196677 );
or ( n29408 , n29406 , n29407 );
buf ( n196686 , n29408 );
buf ( n196687 , n196686 );
xor ( n29411 , n29353 , n196687 );
buf ( n196689 , n29411 );
buf ( n196690 , n196689 );
xor ( n29414 , n196500 , n196690 );
xor ( n29415 , n196549 , n196566 );
xor ( n29416 , n29415 , n196624 );
buf ( n196694 , n29416 );
buf ( n196695 , n196694 );
buf ( n196696 , n196565 );
not ( n29420 , n196696 );
buf ( n196698 , n29420 );
buf ( n196699 , n196698 );
buf ( n196700 , n839 );
buf ( n196701 , n868 );
xor ( n29425 , n196700 , n196701 );
buf ( n196703 , n29425 );
buf ( n196704 , n196703 );
not ( n29428 , n196704 );
buf ( n196706 , n186197 );
not ( n29430 , n196706 );
or ( n29431 , n29428 , n29430 );
buf ( n196709 , n186208 );
buf ( n196710 , n29305 );
nand ( n29434 , n196709 , n196710 );
buf ( n196712 , n29434 );
buf ( n196713 , n196712 );
nand ( n29437 , n29431 , n196713 );
buf ( n196715 , n29437 );
buf ( n196716 , n196715 );
and ( n29440 , n193544 , n193545 );
buf ( n196718 , n29440 );
buf ( n196719 , n196718 );
or ( n29443 , n196716 , n196719 );
buf ( n196721 , n835 );
buf ( n196722 , n872 );
xor ( n29446 , n196721 , n196722 );
buf ( n196724 , n29446 );
buf ( n196725 , n196724 );
not ( n29449 , n196725 );
buf ( n196727 , n19260 );
not ( n29451 , n196727 );
or ( n29452 , n29449 , n29451 );
buf ( n196730 , n19265 );
buf ( n196731 , n196605 );
nand ( n29455 , n196730 , n196731 );
buf ( n196733 , n29455 );
buf ( n196734 , n196733 );
nand ( n29458 , n29452 , n196734 );
buf ( n196736 , n29458 );
buf ( n196737 , n196736 );
nand ( n29461 , n29443 , n196737 );
buf ( n196739 , n29461 );
buf ( n196740 , n196739 );
buf ( n196741 , n196715 );
buf ( n196742 , n196718 );
nand ( n29466 , n196741 , n196742 );
buf ( n196744 , n29466 );
buf ( n196745 , n196744 );
nand ( n29469 , n196740 , n196745 );
buf ( n196747 , n29469 );
buf ( n196748 , n196747 );
xor ( n29472 , n196699 , n196748 );
buf ( n196750 , n837 );
buf ( n196751 , n870 );
xor ( n29475 , n196750 , n196751 );
buf ( n196753 , n29475 );
buf ( n196754 , n196753 );
not ( n29478 , n196754 );
buf ( n196756 , n186435 );
not ( n29480 , n196756 );
or ( n29481 , n29478 , n29480 );
buf ( n196759 , n186444 );
buf ( n196760 , n196655 );
nand ( n29484 , n196759 , n196760 );
buf ( n196762 , n29484 );
buf ( n196763 , n196762 );
nand ( n29487 , n29481 , n196763 );
buf ( n196765 , n29487 );
buf ( n196766 , n196765 );
or ( n29490 , n186395 , n19177 );
nand ( n29491 , n29490 , n876 );
buf ( n196769 , n29491 );
xor ( n29493 , n196766 , n196769 );
buf ( n196771 , n833 );
buf ( n196772 , n874 );
xor ( n29496 , n196771 , n196772 );
buf ( n196774 , n29496 );
buf ( n196775 , n196774 );
not ( n29499 , n196775 );
buf ( n196777 , n186287 );
not ( n29501 , n196777 );
or ( n29502 , n29499 , n29501 );
buf ( n196780 , n186297 );
buf ( n196781 , n196553 );
nand ( n29505 , n196780 , n196781 );
buf ( n196783 , n29505 );
buf ( n196784 , n196783 );
nand ( n29508 , n29502 , n196784 );
buf ( n196786 , n29508 );
buf ( n196787 , n196786 );
and ( n29511 , n29493 , n196787 );
and ( n29512 , n196766 , n196769 );
or ( n29513 , n29511 , n29512 );
buf ( n196791 , n29513 );
buf ( n196792 , n196791 );
and ( n29516 , n29472 , n196792 );
and ( n29517 , n196699 , n196748 );
or ( n29518 , n29516 , n29517 );
buf ( n196796 , n29518 );
buf ( n196797 , n196796 );
xor ( n29521 , n196695 , n196797 );
buf ( n196799 , n843 );
buf ( n196800 , n864 );
xor ( n29524 , n196799 , n196800 );
buf ( n196802 , n29524 );
buf ( n196803 , n196802 );
not ( n29527 , n196803 );
buf ( n196805 , n186640 );
not ( n29529 , n196805 );
or ( n29530 , n29527 , n29529 );
buf ( n196808 , n186340 );
buf ( n196809 , n196637 );
nand ( n29533 , n196808 , n196809 );
buf ( n196811 , n29533 );
buf ( n196812 , n196811 );
nand ( n29536 , n29530 , n196812 );
buf ( n196814 , n29536 );
buf ( n196815 , n196814 );
buf ( n196816 , n841 );
buf ( n196817 , n866 );
xor ( n29541 , n196816 , n196817 );
buf ( n196819 , n29541 );
buf ( n196820 , n196819 );
not ( n29544 , n196820 );
buf ( n196822 , n186241 );
not ( n29546 , n196822 );
or ( n29547 , n29544 , n29546 );
buf ( n196825 , n186254 );
buf ( n196826 , n29291 );
nand ( n29550 , n196825 , n196826 );
buf ( n196828 , n29550 );
buf ( n196829 , n196828 );
nand ( n29553 , n29547 , n196829 );
buf ( n196831 , n29553 );
buf ( n196832 , n196831 );
or ( n29556 , n196815 , n196832 );
buf ( n196834 , n26374 );
not ( n29558 , n196834 );
buf ( n196836 , n19177 );
not ( n29560 , n196836 );
or ( n29561 , n29558 , n29560 );
buf ( n196839 , n186395 );
buf ( n196840 , n876 );
nand ( n29564 , n196839 , n196840 );
buf ( n196842 , n29564 );
buf ( n196843 , n196842 );
nand ( n29567 , n29561 , n196843 );
buf ( n196845 , n29567 );
buf ( n196846 , n196845 );
nand ( n29570 , n29556 , n196846 );
buf ( n196848 , n29570 );
buf ( n196849 , n196848 );
buf ( n196850 , n196814 );
buf ( n196851 , n196831 );
nand ( n29575 , n196850 , n196851 );
buf ( n196853 , n29575 );
buf ( n196854 , n196853 );
nand ( n29578 , n196849 , n196854 );
buf ( n196856 , n29578 );
buf ( n196857 , n196856 );
xor ( n29581 , n196635 , n196650 );
xor ( n29582 , n29581 , n196668 );
buf ( n196860 , n29582 );
buf ( n196861 , n196860 );
xor ( n29585 , n196857 , n196861 );
xor ( n29586 , n196580 , n196617 );
buf ( n196864 , n29586 );
buf ( n196865 , n196594 );
xor ( n29589 , n196864 , n196865 );
buf ( n196867 , n29589 );
buf ( n196868 , n196867 );
and ( n29592 , n29585 , n196868 );
and ( n29593 , n196857 , n196861 );
or ( n29594 , n29592 , n29593 );
buf ( n196872 , n29594 );
buf ( n196873 , n196872 );
and ( n29597 , n29521 , n196873 );
and ( n29598 , n196695 , n196797 );
or ( n29599 , n29597 , n29598 );
buf ( n196877 , n29599 );
buf ( n196878 , n196877 );
xor ( n29602 , n29414 , n196878 );
buf ( n196880 , n29602 );
buf ( n29604 , n196880 );
and ( n29605 , n195762 , n195779 );
buf ( n196883 , n29605 );
buf ( n196884 , n196883 );
buf ( n196885 , n195622 );
not ( n29609 , n196885 );
buf ( n196887 , n28357 );
not ( n29611 , n196887 );
or ( n29612 , n29609 , n29611 );
buf ( n196890 , n195625 );
not ( n29614 , n196890 );
buf ( n196892 , n28357 );
not ( n29616 , n196892 );
buf ( n196894 , n29616 );
buf ( n196895 , n196894 );
not ( n29619 , n196895 );
or ( n29620 , n29614 , n29619 );
buf ( n196898 , n195652 );
nand ( n29622 , n29620 , n196898 );
buf ( n196900 , n29622 );
buf ( n196901 , n196900 );
nand ( n29625 , n29612 , n196901 );
buf ( n196903 , n29625 );
buf ( n196904 , n196903 );
xor ( n29628 , n196884 , n196904 );
xor ( n29629 , n195826 , n195843 );
and ( n29630 , n29629 , n195861 );
and ( n29631 , n195826 , n195843 );
or ( n29632 , n29630 , n29631 );
buf ( n196910 , n29632 );
buf ( n196911 , n196910 );
xor ( n29635 , n29628 , n196911 );
buf ( n196913 , n29635 );
buf ( n196914 , n196913 );
xor ( n29638 , n195802 , n195808 );
and ( n29639 , n29638 , n195864 );
and ( n29640 , n195802 , n195808 );
or ( n29641 , n29639 , n29640 );
buf ( n196919 , n29641 );
buf ( n196920 , n196919 );
xor ( n29644 , n196914 , n196920 );
xor ( n29645 , n195606 , n195655 );
and ( n29646 , n29645 , n195710 );
and ( n29647 , n195606 , n195655 );
or ( n29648 , n29646 , n29647 );
buf ( n196926 , n29648 );
buf ( n196927 , n196926 );
xor ( n29651 , n29644 , n196927 );
buf ( n196929 , n29651 );
buf ( n196930 , n196929 );
buf ( n196931 , n195675 );
not ( n29655 , n196931 );
buf ( n196933 , n195691 );
not ( n29657 , n196933 );
buf ( n196935 , n29657 );
buf ( n196936 , n196935 );
not ( n29660 , n196936 );
or ( n29661 , n29655 , n29660 );
buf ( n196939 , n195708 );
nand ( n29663 , n29661 , n196939 );
buf ( n196941 , n29663 );
buf ( n196942 , n196941 );
buf ( n196943 , n195691 );
buf ( n196944 , n195672 );
nand ( n29668 , n196943 , n196944 );
buf ( n196946 , n29668 );
buf ( n196947 , n196946 );
nand ( n29671 , n196942 , n196947 );
buf ( n196949 , n29671 );
buf ( n196950 , n196949 );
buf ( n196951 , n195836 );
not ( n29675 , n196951 );
buf ( n196953 , n188751 );
not ( n29677 , n196953 );
or ( n29678 , n29675 , n29677 );
buf ( n196956 , n20902 );
buf ( n196957 , n845 );
buf ( n196958 , n890 );
xor ( n29682 , n196957 , n196958 );
buf ( n196960 , n29682 );
buf ( n196961 , n196960 );
nand ( n29685 , n196956 , n196961 );
buf ( n196963 , n29685 );
buf ( n196964 , n196963 );
nand ( n29688 , n29678 , n196964 );
buf ( n196966 , n29688 );
buf ( n196967 , n196966 );
buf ( n196968 , n195854 );
not ( n29692 , n196968 );
buf ( n196970 , n20727 );
not ( n29694 , n196970 );
or ( n29695 , n29692 , n29694 );
buf ( n196973 , n188010 );
buf ( n196974 , n851 );
buf ( n196975 , n884 );
xor ( n29699 , n196974 , n196975 );
buf ( n196977 , n29699 );
buf ( n196978 , n196977 );
nand ( n29702 , n196973 , n196978 );
buf ( n196980 , n29702 );
buf ( n196981 , n196980 );
nand ( n29705 , n29695 , n196981 );
buf ( n196983 , n29705 );
buf ( n196984 , n196983 );
xor ( n29708 , n196967 , n196984 );
buf ( n196986 , n195739 );
not ( n29710 , n196986 );
buf ( n196988 , n19613 );
not ( n29712 , n196988 );
or ( n29713 , n29710 , n29712 );
buf ( n196991 , n19943 );
buf ( n196992 , n853 );
buf ( n196993 , n882 );
xor ( n29717 , n196992 , n196993 );
buf ( n196995 , n29717 );
buf ( n196996 , n196995 );
nand ( n29720 , n196991 , n196996 );
buf ( n196998 , n29720 );
buf ( n196999 , n196998 );
nand ( n29723 , n29713 , n196999 );
buf ( n197001 , n29723 );
buf ( n197002 , n197001 );
xor ( n29726 , n29708 , n197002 );
buf ( n197004 , n29726 );
buf ( n197005 , n197004 );
xor ( n29729 , n196950 , n197005 );
buf ( n197007 , n195632 );
not ( n29731 , n197007 );
buf ( n197009 , n21850 );
not ( n29733 , n197009 );
or ( n29734 , n29731 , n29733 );
buf ( n197012 , n20558 );
buf ( n197013 , n849 );
buf ( n197014 , n886 );
xor ( n29738 , n197013 , n197014 );
buf ( n197016 , n29738 );
buf ( n197017 , n197016 );
nand ( n29741 , n197012 , n197017 );
buf ( n197019 , n29741 );
buf ( n197020 , n197019 );
nand ( n29744 , n29734 , n197020 );
buf ( n197022 , n29744 );
not ( n29746 , n195665 );
not ( n29747 , n18862 );
or ( n29748 , n29746 , n29747 );
buf ( n197026 , n20358 );
buf ( n197027 , n855 );
buf ( n197028 , n880 );
xor ( n29752 , n197027 , n197028 );
buf ( n197030 , n29752 );
buf ( n197031 , n197030 );
nand ( n29755 , n197026 , n197031 );
buf ( n197033 , n29755 );
nand ( n29757 , n29748 , n197033 );
xor ( n29758 , n197022 , n29757 );
buf ( n197036 , n195702 );
not ( n29760 , n197036 );
buf ( n197038 , n186569 );
not ( n29762 , n197038 );
or ( n29763 , n29760 , n29762 );
buf ( n197041 , n186575 );
buf ( n197042 , n857 );
buf ( n197043 , n878 );
xor ( n29767 , n197042 , n197043 );
buf ( n197045 , n29767 );
buf ( n197046 , n197045 );
nand ( n29770 , n197041 , n197046 );
buf ( n197048 , n29770 );
buf ( n197049 , n197048 );
nand ( n29773 , n29763 , n197049 );
buf ( n197051 , n29773 );
xor ( n29775 , n29758 , n197051 );
buf ( n197053 , n29775 );
xor ( n29777 , n29729 , n197053 );
buf ( n197055 , n29777 );
buf ( n197056 , n197055 );
and ( n29780 , n19251 , n863 );
buf ( n197058 , n29780 );
buf ( n197059 , n195685 );
not ( n29783 , n197059 );
buf ( n197061 , n20391 );
not ( n29785 , n197061 );
or ( n29786 , n29783 , n29785 );
buf ( n197064 , n847 );
buf ( n197065 , n888 );
xor ( n29789 , n197064 , n197065 );
buf ( n197067 , n29789 );
buf ( n197068 , n197067 );
buf ( n197069 , n20396 );
nand ( n29793 , n197068 , n197069 );
buf ( n197071 , n29793 );
buf ( n197072 , n197071 );
nand ( n29796 , n29786 , n197072 );
buf ( n197074 , n29796 );
buf ( n197075 , n197074 );
xor ( n29799 , n197058 , n197075 );
buf ( n197077 , n195772 );
not ( n29801 , n197077 );
buf ( n197079 , n20632 );
not ( n29803 , n197079 );
or ( n29804 , n29801 , n29803 );
buf ( n197082 , n190128 );
buf ( n197083 , n843 );
buf ( n197084 , n892 );
xor ( n29808 , n197083 , n197084 );
buf ( n197086 , n29808 );
buf ( n197087 , n197086 );
nand ( n29811 , n197082 , n197087 );
buf ( n197089 , n29811 );
buf ( n197090 , n197089 );
nand ( n29814 , n29804 , n197090 );
buf ( n197092 , n29814 );
buf ( n197093 , n197092 );
xor ( n29817 , n29799 , n197093 );
buf ( n197095 , n29817 );
buf ( n197096 , n197095 );
buf ( n197097 , n195818 );
not ( n29821 , n197097 );
buf ( n197099 , n22809 );
not ( n29823 , n197099 );
or ( n29824 , n29821 , n29823 );
buf ( n197102 , n841 );
buf ( n197103 , n894 );
xor ( n29827 , n197102 , n197103 );
buf ( n197105 , n29827 );
buf ( n197106 , n197105 );
buf ( n197107 , n895 );
nand ( n29831 , n197106 , n197107 );
buf ( n197109 , n29831 );
buf ( n197110 , n197109 );
nand ( n29834 , n29824 , n197110 );
buf ( n197112 , n29834 );
buf ( n197113 , n197112 );
buf ( n197114 , n195616 );
not ( n29838 , n197114 );
buf ( n197116 , n19177 );
not ( n29840 , n197116 );
or ( n29841 , n29838 , n29840 );
buf ( n197119 , n20279 );
buf ( n197120 , n859 );
buf ( n197121 , n876 );
xor ( n29845 , n197120 , n197121 );
buf ( n197123 , n29845 );
buf ( n197124 , n197123 );
nand ( n29848 , n197119 , n197124 );
buf ( n197126 , n29848 );
buf ( n197127 , n197126 );
nand ( n29851 , n29841 , n197127 );
buf ( n197129 , n29851 );
buf ( n197130 , n197129 );
xor ( n29854 , n197113 , n197130 );
buf ( n197132 , n28369 );
not ( n29856 , n197132 );
buf ( n197134 , n18992 );
not ( n29858 , n197134 );
or ( n29859 , n29856 , n29858 );
buf ( n197137 , n187865 );
buf ( n197138 , n861 );
buf ( n197139 , n874 );
xor ( n29863 , n197138 , n197139 );
buf ( n197141 , n29863 );
buf ( n197142 , n197141 );
nand ( n29866 , n197137 , n197142 );
buf ( n197144 , n29866 );
buf ( n197145 , n197144 );
nand ( n29869 , n29859 , n197145 );
buf ( n197147 , n29869 );
buf ( n197148 , n197147 );
xor ( n29872 , n29854 , n197148 );
buf ( n197150 , n29872 );
buf ( n197151 , n197150 );
xor ( n29875 , n197096 , n197151 );
xor ( n29876 , n195746 , n195782 );
and ( n29877 , n29876 , n195792 );
and ( n29878 , n195746 , n195782 );
or ( n29879 , n29877 , n29878 );
buf ( n197157 , n29879 );
buf ( n197158 , n197157 );
xor ( n29882 , n29875 , n197158 );
buf ( n197160 , n29882 );
buf ( n197161 , n197160 );
xor ( n29885 , n197056 , n197161 );
xor ( n29886 , n195729 , n195795 );
and ( n29887 , n29886 , n195867 );
and ( n29888 , n195729 , n195795 );
or ( n29889 , n29887 , n29888 );
buf ( n197167 , n29889 );
buf ( n197168 , n197167 );
xor ( n29892 , n29885 , n197168 );
buf ( n197170 , n29892 );
buf ( n197171 , n197170 );
xor ( n29895 , n196930 , n197171 );
xor ( n29896 , n195598 , n195713 );
and ( n29897 , n29896 , n195870 );
and ( n29898 , n195598 , n195713 );
or ( n29899 , n29897 , n29898 );
buf ( n197177 , n29899 );
buf ( n197178 , n197177 );
and ( n29902 , n29895 , n197178 );
and ( n29903 , n196930 , n197171 );
or ( n29904 , n29902 , n29903 );
buf ( n197182 , n29904 );
buf ( n29906 , n197182 );
not ( n29907 , n18559 );
not ( n29908 , n831 );
or ( n29909 , n29907 , n29908 );
buf ( n197187 , n888 );
buf ( n197188 , n9700 );
xor ( n29912 , n197187 , n197188 );
buf ( n197190 , n177131 );
xor ( n29914 , n29912 , n197190 );
buf ( n197192 , n29914 );
buf ( n197193 , n197192 );
buf ( n197194 , n889 );
buf ( n197195 , n177222 );
xor ( n29919 , n197194 , n197195 );
buf ( n197197 , n9820 );
and ( n29921 , n29919 , n197197 );
and ( n29922 , n197194 , n197195 );
or ( n29923 , n29921 , n29922 );
buf ( n197201 , n29923 );
buf ( n197202 , n197201 );
nor ( n29926 , n197193 , n197202 );
buf ( n197204 , n29926 );
buf ( n197205 , n197204 );
not ( n29929 , n197205 );
buf ( n197207 , n29929 );
buf ( n197208 , n197207 );
buf ( n197209 , n891 );
buf ( n197210 , n177360 );
xor ( n29934 , n197209 , n197210 );
buf ( n197212 , n9958 );
xor ( n29936 , n29934 , n197212 );
buf ( n197214 , n29936 );
buf ( n197215 , n197214 );
buf ( n197216 , n892 );
buf ( n197217 , n177398 );
xor ( n29941 , n197216 , n197217 );
buf ( n197219 , n177425 );
and ( n29943 , n29941 , n197219 );
and ( n29944 , n197216 , n197217 );
or ( n29945 , n29943 , n29944 );
buf ( n197223 , n29945 );
buf ( n197224 , n197223 );
nor ( n29948 , n197215 , n197224 );
buf ( n197226 , n29948 );
buf ( n197227 , n197226 );
buf ( n197228 , n890 );
not ( n29952 , n197228 );
not ( n29953 , n9888 );
buf ( n197231 , n29953 );
not ( n29955 , n197231 );
or ( n29956 , n29952 , n29955 );
buf ( n197234 , n890 );
not ( n29958 , n197234 );
buf ( n197236 , n9888 );
nand ( n29960 , n29958 , n197236 );
buf ( n197238 , n29960 );
buf ( n197239 , n197238 );
nand ( n29963 , n29956 , n197239 );
buf ( n197241 , n29963 );
buf ( n197242 , n197241 );
buf ( n197243 , n29040 );
and ( n29967 , n197242 , n197243 );
not ( n29968 , n197242 );
buf ( n197246 , n29040 );
not ( n29970 , n197246 );
buf ( n197248 , n29970 );
buf ( n197249 , n197248 );
and ( n29973 , n29968 , n197249 );
nor ( n29974 , n29967 , n29973 );
buf ( n197252 , n29974 );
buf ( n197253 , n197252 );
xor ( n29977 , n197209 , n197210 );
and ( n29978 , n29977 , n197212 );
and ( n29979 , n197209 , n197210 );
or ( n29980 , n29978 , n29979 );
buf ( n197258 , n29980 );
buf ( n197259 , n197258 );
nor ( n29983 , n197253 , n197259 );
buf ( n197261 , n29983 );
buf ( n197262 , n197261 );
nor ( n29986 , n197227 , n197262 );
buf ( n197264 , n29986 );
buf ( n197265 , n893 );
buf ( n197266 , n177490 );
xor ( n29990 , n197265 , n197266 );
buf ( n197268 , n177484 );
xor ( n29992 , n29990 , n197268 );
buf ( n197270 , n29992 );
buf ( n197271 , n197270 );
and ( n29995 , n168495 , n168500 );
buf ( n197273 , n29995 );
buf ( n197274 , n197273 );
nand ( n29998 , n197271 , n197274 );
buf ( n197276 , n29998 );
buf ( n197277 , n197276 );
not ( n30001 , n197277 );
buf ( n197279 , n30001 );
buf ( n197280 , n197270 );
not ( n30004 , n197280 );
buf ( n197282 , n30004 );
buf ( n197283 , n197282 );
buf ( n197284 , n197273 );
not ( n30008 , n197284 );
buf ( n197286 , n30008 );
buf ( n197287 , n197286 );
and ( n30011 , n197283 , n197287 );
buf ( n197289 , n168486 );
buf ( n197290 , n168503 );
nand ( n30014 , n197289 , n197290 );
buf ( n197292 , n30014 );
buf ( n197293 , n197292 );
buf ( n197294 , n168494 );
and ( n30018 , n197293 , n197294 );
buf ( n197296 , n168485 );
buf ( n197297 , n168502 );
and ( n30021 , n197296 , n197297 );
buf ( n197299 , n30021 );
buf ( n197300 , n197299 );
nor ( n30024 , n30018 , n197300 );
buf ( n197302 , n30024 );
buf ( n197303 , n197302 );
nor ( n30027 , n30011 , n197303 );
buf ( n197305 , n30027 );
or ( n30029 , n197279 , n197305 );
xor ( n30030 , n197216 , n197217 );
xor ( n30031 , n30030 , n197219 );
buf ( n197309 , n30031 );
buf ( n197310 , n197309 );
not ( n30034 , n197310 );
buf ( n197312 , n30034 );
buf ( n197313 , n197312 );
xor ( n30037 , n197265 , n197266 );
and ( n30038 , n30037 , n197268 );
and ( n30039 , n197265 , n197266 );
or ( n30040 , n30038 , n30039 );
buf ( n197318 , n30040 );
buf ( n197319 , n197318 );
not ( n30043 , n197319 );
buf ( n197321 , n30043 );
buf ( n197322 , n197321 );
nand ( n30046 , n197313 , n197322 );
buf ( n197324 , n30046 );
nand ( n30048 , n30029 , n197324 );
buf ( n197326 , n197321 );
not ( n30050 , n197326 );
buf ( n197328 , n197309 );
nand ( n30052 , n30050 , n197328 );
buf ( n197330 , n30052 );
nand ( n30054 , n30048 , n197330 );
nand ( n30055 , n197264 , n30054 );
not ( n30056 , n30055 );
buf ( n197334 , n30056 );
xor ( n30058 , n197194 , n197195 );
xor ( n30059 , n30058 , n197197 );
buf ( n197337 , n30059 );
buf ( n197338 , n197337 );
buf ( n197339 , n9888 );
not ( n30063 , n197339 );
buf ( n197341 , n29040 );
not ( n30065 , n197341 );
or ( n30066 , n30063 , n30065 );
buf ( n197344 , n29040 );
buf ( n197345 , n9888 );
or ( n30069 , n197344 , n197345 );
buf ( n197347 , n890 );
nand ( n30071 , n30069 , n197347 );
buf ( n197349 , n30071 );
buf ( n197350 , n197349 );
nand ( n30074 , n30066 , n197350 );
buf ( n197352 , n30074 );
buf ( n197353 , n197352 );
nor ( n30077 , n197338 , n197353 );
buf ( n197355 , n30077 );
buf ( n197356 , n197355 );
not ( n30080 , n197356 );
buf ( n197358 , n30080 );
buf ( n197359 , n197358 );
nand ( n30083 , n197208 , n197334 , n197359 );
buf ( n197361 , n30083 );
buf ( n197362 , n197361 );
buf ( n197363 , n197207 );
buf ( n197364 , n197252 );
buf ( n197365 , n197258 );
nor ( n30089 , n197364 , n197365 );
buf ( n197367 , n30089 );
buf ( n197368 , n197367 );
buf ( n197369 , n197214 );
buf ( n197370 , n197223 );
nand ( n30094 , n197369 , n197370 );
buf ( n197372 , n30094 );
buf ( n197373 , n197372 );
or ( n30097 , n197368 , n197373 );
buf ( n197375 , n197252 );
buf ( n197376 , n197258 );
nand ( n30100 , n197375 , n197376 );
buf ( n197378 , n30100 );
buf ( n197379 , n197378 );
nand ( n30103 , n30097 , n197379 );
buf ( n197381 , n30103 );
buf ( n197382 , n197381 );
buf ( n197383 , n197358 );
nand ( n30107 , n197363 , n197382 , n197383 );
buf ( n197385 , n30107 );
buf ( n197386 , n197385 );
buf ( n197387 , n197204 );
not ( n30111 , n197387 );
buf ( n197389 , n197337 );
buf ( n197390 , n197352 );
nand ( n30114 , n197389 , n197390 );
buf ( n197392 , n30114 );
buf ( n197393 , n197392 );
not ( n30117 , n197393 );
and ( n30118 , n30111 , n30117 );
buf ( n197396 , n197192 );
buf ( n197397 , n197201 );
and ( n30121 , n197396 , n197397 );
buf ( n197399 , n30121 );
buf ( n197400 , n197399 );
nor ( n30124 , n30118 , n197400 );
buf ( n197402 , n30124 );
buf ( n197403 , n197402 );
nand ( n30127 , n197362 , n197386 , n197403 );
buf ( n197405 , n30127 );
buf ( n197406 , n197405 );
not ( n30130 , n197406 );
buf ( n197408 , n30130 );
buf ( n197409 , n197408 );
not ( n30133 , n197409 );
buf ( n197411 , n30133 );
buf ( n197412 , n197411 );
not ( n30136 , n197412 );
buf ( n197414 , n884 );
buf ( n197415 , n176664 );
xor ( n30139 , n197414 , n197415 );
buf ( n197417 , n176669 );
xor ( n30141 , n30139 , n197417 );
buf ( n197419 , n30141 );
buf ( n197420 , n197419 );
buf ( n197421 , n885 );
buf ( n197422 , n176799 );
xor ( n30146 , n197421 , n197422 );
buf ( n197424 , n176807 );
and ( n30148 , n30146 , n197424 );
and ( n30149 , n197421 , n197422 );
or ( n30150 , n30148 , n30149 );
buf ( n197428 , n30150 );
buf ( n197429 , n197428 );
nor ( n30153 , n197420 , n197429 );
buf ( n197431 , n30153 );
buf ( n197432 , n197431 );
not ( n30156 , n197432 );
buf ( n197434 , n30156 );
buf ( n197435 , n197434 );
xor ( n30159 , n197421 , n197422 );
xor ( n30160 , n30159 , n197424 );
buf ( n197438 , n30160 );
buf ( n197439 , n197438 );
buf ( n197440 , n886 );
buf ( n197441 , n176924 );
xor ( n30165 , n197440 , n197441 );
buf ( n197443 , n176929 );
and ( n30167 , n30165 , n197443 );
and ( n30168 , n197440 , n197441 );
or ( n30169 , n30167 , n30168 );
buf ( n197447 , n30169 );
buf ( n197448 , n197447 );
or ( n30172 , n197439 , n197448 );
buf ( n197450 , n30172 );
buf ( n197451 , n197450 );
buf ( n197452 , n887 );
buf ( n197453 , n177030 );
xor ( n30177 , n197452 , n197453 );
buf ( n197455 , n177035 );
xor ( n30179 , n30177 , n197455 );
buf ( n197457 , n30179 );
not ( n30181 , n197457 );
xor ( n30182 , n197187 , n197188 );
and ( n30183 , n30182 , n197190 );
and ( n30184 , n197187 , n197188 );
or ( n30185 , n30183 , n30184 );
buf ( n197463 , n30185 );
not ( n30187 , n197463 );
and ( n30188 , n30181 , n30187 );
xor ( n30189 , n197440 , n197441 );
xor ( n30190 , n30189 , n197443 );
buf ( n197468 , n30190 );
buf ( n197469 , n197468 );
xor ( n30193 , n197452 , n197453 );
and ( n30194 , n30193 , n197455 );
and ( n30195 , n197452 , n197453 );
or ( n30196 , n30194 , n30195 );
buf ( n197474 , n30196 );
buf ( n197475 , n197474 );
nor ( n30199 , n197469 , n197475 );
buf ( n197477 , n30199 );
nor ( n30201 , n30188 , n197477 );
buf ( n197479 , n30201 );
and ( n30203 , n197435 , n197451 , n197479 );
buf ( n197481 , n30203 );
buf ( n197482 , n197481 );
not ( n30206 , n197482 );
or ( n30207 , n30136 , n30206 );
buf ( n197485 , n197477 );
buf ( n197486 , n197457 );
buf ( n197487 , n197463 );
nand ( n30211 , n197486 , n197487 );
buf ( n197489 , n30211 );
buf ( n197490 , n197489 );
or ( n30214 , n197485 , n197490 );
buf ( n197492 , n197468 );
buf ( n197493 , n197474 );
nand ( n30217 , n197492 , n197493 );
buf ( n197495 , n30217 );
buf ( n197496 , n197495 );
nand ( n30220 , n30214 , n197496 );
buf ( n197498 , n30220 );
buf ( n197499 , n197498 );
not ( n30223 , n197499 );
buf ( n197501 , n197431 );
buf ( n197502 , n197438 );
buf ( n197503 , n197447 );
nor ( n30227 , n197502 , n197503 );
buf ( n197505 , n30227 );
buf ( n197506 , n197505 );
nor ( n30230 , n197501 , n197506 );
buf ( n197508 , n30230 );
buf ( n197509 , n197508 );
not ( n30233 , n197509 );
or ( n30234 , n30223 , n30233 );
buf ( n197512 , n197431 );
not ( n30236 , n197512 );
buf ( n197514 , n197438 );
buf ( n197515 , n197447 );
nand ( n30239 , n197514 , n197515 );
buf ( n197517 , n30239 );
buf ( n197518 , n197517 );
not ( n30242 , n197518 );
and ( n30243 , n30236 , n30242 );
buf ( n197521 , n197419 );
buf ( n197522 , n197428 );
and ( n30246 , n197521 , n197522 );
buf ( n197524 , n30246 );
buf ( n197525 , n197524 );
nor ( n30249 , n30243 , n197525 );
buf ( n197527 , n30249 );
buf ( n197528 , n197527 );
nand ( n30252 , n30234 , n197528 );
buf ( n197530 , n30252 );
buf ( n197531 , n197530 );
not ( n30255 , n197531 );
buf ( n197533 , n30255 );
buf ( n197534 , n197533 );
nand ( n30258 , n30207 , n197534 );
buf ( n197536 , n30258 );
buf ( n197537 , n883 );
buf ( n197538 , n176558 );
xor ( n30262 , n197537 , n197538 );
buf ( n197540 , n176563 );
xor ( n30264 , n30262 , n197540 );
buf ( n197542 , n30264 );
buf ( n197543 , n197542 );
xor ( n30267 , n197414 , n197415 );
and ( n30268 , n30267 , n197417 );
and ( n30269 , n197414 , n197415 );
or ( n30270 , n30268 , n30269 );
buf ( n197548 , n30270 );
buf ( n197549 , n197548 );
nor ( n30273 , n197543 , n197549 );
buf ( n197551 , n30273 );
buf ( n197552 , n197551 );
not ( n30276 , n197552 );
buf ( n197554 , n30276 );
buf ( n197555 , n197554 );
buf ( n197556 , n197542 );
buf ( n197557 , n197548 );
nand ( n30281 , n197556 , n197557 );
buf ( n197559 , n30281 );
buf ( n197560 , n197559 );
buf ( n30284 , n197560 );
buf ( n197562 , n30284 );
buf ( n197563 , n197562 );
nand ( n30287 , n197555 , n197563 );
buf ( n197565 , n30287 );
xnor ( n30289 , n197536 , n197565 );
nand ( n30290 , n30289 , n168462 );
nand ( n30291 , n29909 , n30290 );
buf ( n30292 , n30291 );
or ( n30293 , n197457 , n197463 );
not ( n30294 , n30293 );
nor ( n30295 , n30294 , n197477 , n197505 );
buf ( n197573 , n30295 );
not ( n30297 , n197573 );
buf ( n197575 , n197405 );
buf ( n30299 , n197575 );
buf ( n197577 , n30299 );
buf ( n197578 , n197577 );
not ( n30302 , n197578 );
or ( n30303 , n30297 , n30302 );
buf ( n197581 , n197498 );
not ( n30305 , n197581 );
buf ( n197583 , n197450 );
not ( n30307 , n197583 );
or ( n30308 , n30305 , n30307 );
buf ( n197586 , n197517 );
nand ( n30310 , n30308 , n197586 );
buf ( n197588 , n30310 );
buf ( n197589 , n197588 );
not ( n30313 , n197589 );
buf ( n197591 , n30313 );
buf ( n197592 , n197591 );
nand ( n30316 , n30303 , n197592 );
buf ( n197594 , n30316 );
buf ( n197595 , n197594 );
buf ( n197596 , n197434 );
not ( n30320 , n197596 );
buf ( n197598 , n197524 );
nor ( n30322 , n30320 , n197598 );
buf ( n197600 , n30322 );
buf ( n197601 , n197600 );
and ( n30325 , n197595 , n197601 );
not ( n30326 , n197595 );
buf ( n197604 , n197600 );
not ( n30328 , n197604 );
buf ( n197606 , n30328 );
buf ( n197607 , n197606 );
and ( n30331 , n30326 , n197607 );
nor ( n30332 , n30325 , n30331 );
buf ( n197610 , n30332 );
nand ( n30334 , n197610 , n168462 );
buf ( n197612 , n177589 );
buf ( n197613 , n177150 );
not ( n30337 , n197613 );
buf ( n197615 , n30337 );
buf ( n197616 , n197615 );
or ( n30340 , n177044 , n177040 );
buf ( n197618 , n30340 );
nand ( n30342 , n197616 , n197618 );
buf ( n197620 , n30342 );
buf ( n197621 , n197620 );
nor ( n30345 , n197612 , n197621 );
buf ( n197623 , n30345 );
buf ( n197624 , n197623 );
not ( n30348 , n197624 );
buf ( n197626 , n177559 );
buf ( n30350 , n197626 );
buf ( n197628 , n30350 );
buf ( n197629 , n197628 );
not ( n30353 , n197629 );
or ( n30354 , n30348 , n30353 );
buf ( n197632 , n176940 );
not ( n30356 , n197632 );
buf ( n197634 , n177580 );
not ( n30358 , n197634 );
or ( n30359 , n30356 , n30358 );
buf ( n197637 , n177598 );
nand ( n30361 , n30359 , n197637 );
buf ( n197639 , n30361 );
buf ( n197640 , n197639 );
not ( n30364 , n197640 );
buf ( n197642 , n30364 );
buf ( n197643 , n197642 );
nand ( n30367 , n30354 , n197643 );
buf ( n197645 , n30367 );
buf ( n197646 , n197645 );
not ( n30370 , n176826 );
nor ( n30371 , n30370 , n177607 );
buf ( n197649 , n30371 );
and ( n30373 , n197646 , n197649 );
not ( n30374 , n197646 );
buf ( n197652 , n30371 );
not ( n30376 , n197652 );
buf ( n197654 , n30376 );
buf ( n197655 , n197654 );
and ( n30379 , n30374 , n197655 );
nor ( n30380 , n30373 , n30379 );
buf ( n197658 , n30380 );
nand ( n30382 , n197658 , n831 );
nand ( n30383 , n30334 , n30382 );
buf ( n30384 , n30383 );
not ( n30385 , n831 );
and ( n30386 , n197615 , n177571 );
buf ( n197664 , n30386 );
not ( n30388 , n197664 );
buf ( n197666 , n177562 );
not ( n30390 , n197666 );
or ( n30391 , n30388 , n30390 );
buf ( n197669 , n197628 );
not ( n30393 , n197669 );
buf ( n197671 , n30393 );
buf ( n197672 , n197671 );
buf ( n197673 , n30386 );
or ( n30397 , n197672 , n197673 );
nand ( n30398 , n30391 , n30397 );
buf ( n197676 , n30398 );
not ( n30400 , n197676 );
or ( n30401 , n30385 , n30400 );
buf ( n197679 , n30293 );
buf ( n197680 , n197489 );
and ( n30404 , n197679 , n197680 );
buf ( n197682 , n30404 );
and ( n30406 , n197682 , n197408 );
not ( n30407 , n197682 );
and ( n30408 , n30407 , n197577 );
or ( n30409 , n30406 , n30408 );
nand ( n30410 , n30409 , n168462 );
nand ( n30411 , n30401 , n30410 );
buf ( n30412 , n30411 );
buf ( n197690 , n177307 );
buf ( n30414 , n197690 );
buf ( n197692 , n30414 );
buf ( n197693 , n197692 );
buf ( n197694 , n177453 );
buf ( n197695 , n177445 );
nand ( n30419 , n197694 , n197695 );
buf ( n197697 , n30419 );
buf ( n197698 , n197697 );
buf ( n197699 , n10146 );
not ( n30423 , n197699 );
buf ( n197701 , n30423 );
buf ( n197702 , n197701 );
not ( n30426 , n197702 );
buf ( n197704 , n177453 );
buf ( n197705 , n177470 );
buf ( n30429 , n197705 );
buf ( n197707 , n30429 );
buf ( n197708 , n197707 );
nand ( n30432 , n30426 , n197704 , n197708 );
buf ( n197710 , n30432 );
buf ( n197711 , n197710 );
nand ( n30435 , n197693 , n197698 , n197711 );
buf ( n197713 , n30435 );
buf ( n197714 , n197713 );
not ( n30438 , n197714 );
buf ( n197716 , n177316 );
not ( n30440 , n197716 );
buf ( n197718 , n177234 );
nand ( n30442 , n30440 , n197718 );
buf ( n197720 , n30442 );
buf ( n197721 , n197720 );
not ( n30445 , n197721 );
or ( n30446 , n30438 , n30445 );
buf ( n197724 , n197713 );
buf ( n197725 , n197720 );
or ( n30449 , n197724 , n197725 );
nand ( n30450 , n30446 , n30449 );
buf ( n197728 , n30450 );
and ( n30452 , n831 , n197728 );
not ( n30453 , n831 );
buf ( n197731 , n197399 );
not ( n30455 , n197731 );
buf ( n197733 , n197207 );
nand ( n30457 , n30455 , n197733 );
buf ( n197735 , n30457 );
buf ( n197736 , n197735 );
not ( n30460 , n197736 );
buf ( n197738 , n197392 );
buf ( n197739 , n197337 );
buf ( n197740 , n197352 );
nor ( n30464 , n197739 , n197740 );
buf ( n197742 , n30464 );
buf ( n197743 , n197742 );
not ( n30467 , n197743 );
buf ( n197745 , n197264 );
buf ( n30469 , n197745 );
buf ( n197747 , n30469 );
buf ( n197748 , n197747 );
not ( n30472 , n30054 );
not ( n30473 , n30472 );
buf ( n197751 , n30473 );
nand ( n30475 , n30467 , n197748 , n197751 );
buf ( n197753 , n30475 );
buf ( n197754 , n197753 );
buf ( n197755 , n197381 );
buf ( n197756 , n197742 );
not ( n30480 , n197756 );
buf ( n197758 , n30480 );
buf ( n197759 , n197758 );
nand ( n30483 , n197755 , n197759 );
buf ( n197761 , n30483 );
buf ( n197762 , n197761 );
nand ( n30486 , n197738 , n197754 , n197762 );
buf ( n197764 , n30486 );
buf ( n197765 , n197764 );
not ( n30489 , n197765 );
or ( n30490 , n30460 , n30489 );
buf ( n197768 , n197764 );
buf ( n197769 , n197735 );
or ( n30493 , n197768 , n197769 );
nand ( n30494 , n30490 , n30493 );
buf ( n197772 , n30494 );
and ( n30496 , n30453 , n197772 );
nor ( n30497 , n30452 , n30496 );
not ( n30498 , n30497 );
buf ( n197776 , n30201 );
not ( n30500 , n197776 );
buf ( n197778 , n197405 );
not ( n30502 , n197778 );
or ( n30503 , n30500 , n30502 );
buf ( n197781 , n197498 );
not ( n30505 , n197781 );
buf ( n197783 , n30505 );
buf ( n197784 , n197783 );
nand ( n30508 , n30503 , n197784 );
buf ( n197786 , n30508 );
buf ( n197787 , n197786 );
buf ( n197788 , n197450 );
buf ( n197789 , n197517 );
nand ( n30513 , n197788 , n197789 );
buf ( n197791 , n30513 );
buf ( n197792 , n197791 );
not ( n30516 , n197792 );
buf ( n197794 , n30516 );
buf ( n197795 , n197794 );
and ( n30519 , n197787 , n197795 );
not ( n30520 , n197787 );
buf ( n197798 , n197791 );
and ( n30522 , n30520 , n197798 );
nor ( n30523 , n30519 , n30522 );
buf ( n197801 , n30523 );
and ( n30525 , n168462 , n197801 );
not ( n30526 , n168462 );
buf ( n197804 , n177153 );
not ( n30528 , n197804 );
buf ( n197806 , n177559 );
not ( n30530 , n197806 );
or ( n30531 , n30528 , n30530 );
buf ( n197809 , n177580 );
not ( n30533 , n197809 );
buf ( n197811 , n30533 );
buf ( n197812 , n197811 );
nand ( n30536 , n30531 , n197812 );
buf ( n197814 , n30536 );
buf ( n197815 , n197814 );
buf ( n197816 , n176847 );
not ( n30540 , n197816 );
buf ( n197818 , n176937 );
not ( n30542 , n197818 );
or ( n30543 , n30540 , n30542 );
buf ( n197821 , n177598 );
nand ( n30545 , n30543 , n197821 );
buf ( n197823 , n30545 );
buf ( n197824 , n197823 );
not ( n30548 , n197824 );
buf ( n197826 , n30548 );
buf ( n197827 , n197826 );
and ( n30551 , n197815 , n197827 );
not ( n30552 , n197815 );
buf ( n197830 , n197823 );
and ( n30554 , n30552 , n197830 );
nor ( n30555 , n30551 , n30554 );
buf ( n197833 , n30555 );
and ( n30557 , n30526 , n197833 );
nor ( n30558 , n30525 , n30557 );
not ( n30559 , n168462 );
buf ( n197837 , n30293 );
not ( n30561 , n197837 );
buf ( n197839 , n197405 );
not ( n30563 , n197839 );
or ( n30564 , n30561 , n30563 );
buf ( n197842 , n197489 );
nand ( n30566 , n30564 , n197842 );
buf ( n197844 , n30566 );
buf ( n197845 , n197844 );
buf ( n197846 , n197477 );
not ( n30570 , n197846 );
buf ( n197848 , n197495 );
nand ( n30572 , n30570 , n197848 );
buf ( n197850 , n30572 );
buf ( n197851 , n197850 );
not ( n30575 , n197851 );
buf ( n197853 , n30575 );
buf ( n197854 , n197853 );
and ( n30578 , n197845 , n197854 );
not ( n30579 , n197845 );
buf ( n197857 , n197850 );
and ( n30581 , n30579 , n197857 );
nor ( n30582 , n30578 , n30581 );
buf ( n197860 , n30582 );
not ( n30584 , n197860 );
or ( n30585 , n30559 , n30584 );
buf ( n197863 , n197615 );
not ( n30587 , n197863 );
buf ( n197865 , n177559 );
not ( n30589 , n197865 );
or ( n30590 , n30587 , n30589 );
buf ( n197868 , n177571 );
nand ( n30592 , n30590 , n197868 );
buf ( n197870 , n30592 );
buf ( n197871 , n197870 );
buf ( n197872 , n30340 );
buf ( n197873 , n177577 );
nand ( n30597 , n197872 , n197873 );
buf ( n197875 , n30597 );
buf ( n197876 , n197875 );
not ( n30600 , n197876 );
buf ( n197878 , n30600 );
buf ( n197879 , n197878 );
and ( n30603 , n197871 , n197879 );
not ( n30604 , n197871 );
buf ( n197882 , n197875 );
and ( n30606 , n30604 , n197882 );
nor ( n30607 , n30603 , n30606 );
buf ( n197885 , n30607 );
nand ( n30609 , n197885 , n831 );
nand ( n30610 , n30585 , n30609 );
not ( n30611 , n831 );
buf ( n197889 , n177539 );
buf ( n197890 , n177548 );
nand ( n30614 , n197889 , n197890 );
buf ( n197892 , n30614 );
buf ( n197893 , n197892 );
buf ( n197894 , n177523 );
not ( n30618 , n197894 );
buf ( n197896 , n30618 );
buf ( n197897 , n197896 );
and ( n30621 , n197893 , n197897 );
not ( n30622 , n197893 );
buf ( n197900 , n177523 );
and ( n30624 , n30622 , n197900 );
nor ( n30625 , n30621 , n30624 );
buf ( n197903 , n30625 );
not ( n30627 , n197903 );
or ( n30628 , n30611 , n30627 );
buf ( n197906 , n197324 );
buf ( n197907 , n197330 );
nand ( n30631 , n197906 , n197907 );
buf ( n197909 , n30631 );
buf ( n197910 , n197909 );
buf ( n197911 , n197305 );
not ( n30635 , n197911 );
buf ( n197913 , n197276 );
nand ( n30637 , n30635 , n197913 );
buf ( n197915 , n30637 );
buf ( n197916 , n197915 );
xnor ( n30640 , n197910 , n197916 );
buf ( n197918 , n30640 );
nand ( n30642 , n197918 , n168462 );
nand ( n30643 , n30628 , n30642 );
not ( n30644 , n831 );
buf ( n197922 , n177499 );
not ( n30646 , n197922 );
buf ( n197924 , n177520 );
nand ( n30648 , n30646 , n197924 );
buf ( n197926 , n30648 );
xor ( n30650 , n197926 , n10108 );
not ( n30651 , n30650 );
or ( n30652 , n30644 , n30651 );
buf ( n197930 , n197302 );
buf ( n197931 , n197286 );
not ( n30655 , n197931 );
buf ( n197933 , n197282 );
not ( n30657 , n197933 );
or ( n30658 , n30655 , n30657 );
buf ( n197936 , n197276 );
nand ( n30660 , n30658 , n197936 );
buf ( n197938 , n30660 );
buf ( n197939 , n197938 );
xor ( n30663 , n197930 , n197939 );
buf ( n197941 , n30663 );
nand ( n30665 , n197941 , n168462 );
nand ( n30666 , n30652 , n30665 );
not ( n30667 , n831 );
buf ( n197945 , n8773 );
not ( n30669 , n197945 );
buf ( n197947 , n175724 );
nor ( n30671 , n30669 , n197947 );
buf ( n197949 , n30671 );
buf ( n197950 , n197949 );
not ( n30674 , n197950 );
buf ( n197952 , n18819 );
not ( n30676 , n197952 );
or ( n30677 , n30674 , n30676 );
buf ( n197955 , n186122 );
buf ( n197956 , n186130 );
and ( n30680 , n197955 , n197956 );
buf ( n197958 , n176098 );
nor ( n30682 , n30680 , n197958 );
buf ( n197960 , n30682 );
buf ( n197961 , n197960 );
nand ( n30685 , n30677 , n197961 );
buf ( n197963 , n30685 );
buf ( n197964 , n197963 );
buf ( n197965 , n176087 );
not ( n30689 , n197965 );
buf ( n197967 , n176104 );
nor ( n30691 , n30689 , n197967 );
buf ( n197969 , n30691 );
buf ( n197970 , n197969 );
and ( n30694 , n197964 , n197970 );
not ( n30695 , n197964 );
buf ( n197973 , n197969 );
not ( n30697 , n197973 );
buf ( n197975 , n30697 );
buf ( n197976 , n197975 );
and ( n30700 , n30695 , n197976 );
nor ( n30701 , n30694 , n30700 );
buf ( n197979 , n30701 );
not ( n30703 , n197979 );
or ( n30704 , n30667 , n30703 );
buf ( n197982 , n878 );
buf ( n197983 , n175711 );
xor ( n30707 , n197982 , n197983 );
buf ( n197985 , n175716 );
xor ( n30709 , n30707 , n197985 );
buf ( n197987 , n30709 );
not ( n30711 , n197987 );
buf ( n197989 , n879 );
buf ( n197990 , n176047 );
xor ( n30714 , n197989 , n197990 );
buf ( n197992 , n176052 );
and ( n30716 , n30714 , n197992 );
and ( n30717 , n197989 , n197990 );
or ( n30718 , n30716 , n30717 );
buf ( n197996 , n30718 );
not ( n30720 , n197996 );
and ( n30721 , n30711 , n30720 );
buf ( n197999 , n880 );
buf ( n198000 , n176016 );
xor ( n30724 , n197999 , n198000 );
buf ( n198002 , n176035 );
and ( n30726 , n30724 , n198002 );
and ( n30727 , n197999 , n198000 );
or ( n30728 , n30726 , n30727 );
buf ( n198006 , n30728 );
xor ( n30730 , n197989 , n197990 );
xor ( n30731 , n30730 , n197992 );
buf ( n198009 , n30731 );
nor ( n30733 , n198006 , n198009 );
nor ( n30734 , n30721 , n30733 );
buf ( n198012 , n877 );
buf ( n198013 , n175469 );
xor ( n30737 , n198012 , n198013 );
buf ( n198015 , n8040 );
xor ( n30739 , n30737 , n198015 );
buf ( n198017 , n30739 );
buf ( n198018 , n198017 );
xor ( n30742 , n197982 , n197983 );
and ( n30743 , n30742 , n197985 );
and ( n30744 , n197982 , n197983 );
or ( n30745 , n30743 , n30744 );
buf ( n198023 , n30745 );
buf ( n198024 , n198023 );
nor ( n30748 , n198018 , n198024 );
buf ( n198026 , n30748 );
buf ( n198027 , n198026 );
not ( n30751 , n198027 );
buf ( n198029 , n30751 );
and ( n30753 , n30734 , n198029 );
buf ( n198031 , n30753 );
not ( n30755 , n198031 );
buf ( n198033 , n881 );
buf ( n198034 , n176288 );
xor ( n30758 , n198033 , n198034 );
buf ( n198036 , n176293 );
and ( n30760 , n30758 , n198036 );
and ( n30761 , n198033 , n198034 );
or ( n30762 , n30760 , n30761 );
buf ( n198040 , n30762 );
buf ( n198041 , n198040 );
not ( n30765 , n198041 );
xor ( n30766 , n197999 , n198000 );
xor ( n30767 , n30766 , n198002 );
buf ( n198045 , n30767 );
buf ( n198046 , n198045 );
not ( n30770 , n198046 );
buf ( n198048 , n30770 );
buf ( n198049 , n198048 );
nand ( n30773 , n30765 , n198049 );
buf ( n198051 , n30773 );
buf ( n198052 , n198051 );
buf ( n198053 , n197551 );
xor ( n30777 , n197537 , n197538 );
and ( n30778 , n30777 , n197540 );
and ( n30779 , n197537 , n197538 );
or ( n30780 , n30778 , n30779 );
buf ( n198058 , n30780 );
buf ( n198059 , n198058 );
buf ( n198060 , n882 );
buf ( n198061 , n176433 );
xor ( n30785 , n198060 , n198061 );
buf ( n198063 , n176438 );
xor ( n30787 , n30785 , n198063 );
buf ( n198065 , n30787 );
buf ( n198066 , n198065 );
nor ( n30790 , n198059 , n198066 );
buf ( n198068 , n30790 );
buf ( n198069 , n198068 );
nor ( n30793 , n198053 , n198069 );
buf ( n198071 , n30793 );
buf ( n198072 , n198071 );
xor ( n30796 , n198033 , n198034 );
xor ( n30797 , n30796 , n198036 );
buf ( n198075 , n30797 );
buf ( n198076 , n198075 );
xor ( n30800 , n198060 , n198061 );
and ( n30801 , n30800 , n198063 );
and ( n30802 , n198060 , n198061 );
or ( n30803 , n30801 , n30802 );
buf ( n198081 , n30803 );
buf ( n198082 , n198081 );
nor ( n30806 , n198076 , n198082 );
buf ( n198084 , n30806 );
buf ( n198085 , n198084 );
not ( n30809 , n198085 );
buf ( n198087 , n30809 );
buf ( n198088 , n198087 );
and ( n30812 , n198052 , n198072 , n198088 );
buf ( n198090 , n30812 );
buf ( n198091 , n198090 );
not ( n30815 , n198091 );
buf ( n198093 , n197536 );
not ( n30817 , n198093 );
or ( n30818 , n30815 , n30817 );
buf ( n198096 , n198065 );
buf ( n198097 , n198058 );
nor ( n30821 , n198096 , n198097 );
buf ( n198099 , n30821 );
buf ( n198100 , n198099 );
buf ( n198101 , n197559 );
or ( n30825 , n198100 , n198101 );
buf ( n198103 , n198065 );
buf ( n198104 , n198058 );
nand ( n30828 , n198103 , n198104 );
buf ( n198106 , n30828 );
buf ( n198107 , n198106 );
nand ( n30831 , n30825 , n198107 );
buf ( n198109 , n30831 );
buf ( n198110 , n198109 );
not ( n30834 , n198110 );
buf ( n198112 , n198040 );
buf ( n198113 , n198045 );
nor ( n30837 , n198112 , n198113 );
buf ( n198115 , n30837 );
buf ( n198116 , n198115 );
buf ( n198117 , n198084 );
nor ( n30841 , n198116 , n198117 );
buf ( n198119 , n30841 );
buf ( n198120 , n198119 );
not ( n30844 , n198120 );
or ( n30845 , n30834 , n30844 );
buf ( n198123 , n198051 );
buf ( n198124 , n198075 );
buf ( n198125 , n198081 );
and ( n30849 , n198124 , n198125 );
buf ( n198127 , n30849 );
buf ( n198128 , n198127 );
and ( n30852 , n198123 , n198128 );
buf ( n198130 , n198040 );
not ( n30854 , n198130 );
buf ( n198132 , n198048 );
nor ( n30856 , n30854 , n198132 );
buf ( n198134 , n30856 );
buf ( n198135 , n198134 );
nor ( n30859 , n30852 , n198135 );
buf ( n198137 , n30859 );
buf ( n198138 , n198137 );
nand ( n30862 , n30845 , n198138 );
buf ( n198140 , n30862 );
buf ( n198141 , n198140 );
not ( n30865 , n198141 );
buf ( n198143 , n30865 );
buf ( n198144 , n198143 );
nand ( n30868 , n30818 , n198144 );
buf ( n198146 , n30868 );
buf ( n198147 , n198146 );
not ( n30871 , n198147 );
or ( n30872 , n30755 , n30871 );
buf ( n198150 , n198006 );
buf ( n198151 , n198009 );
nand ( n30875 , n198150 , n198151 );
buf ( n198153 , n30875 );
buf ( n198154 , n197987 );
buf ( n198155 , n197996 );
nand ( n30879 , n198154 , n198155 );
buf ( n198157 , n30879 );
and ( n30881 , n198153 , n198157 );
buf ( n198159 , n197987 );
not ( n30883 , n198159 );
buf ( n198161 , n30883 );
buf ( n198162 , n198161 );
buf ( n198163 , n197996 );
not ( n30887 , n198163 );
buf ( n198165 , n30887 );
buf ( n198166 , n198165 );
nand ( n30890 , n198162 , n198166 );
buf ( n198168 , n30890 );
not ( n30892 , n198168 );
nor ( n30893 , n30881 , n30892 );
buf ( n30894 , n30893 );
and ( n30895 , n198029 , n30894 );
buf ( n198173 , n198017 );
not ( n30897 , n198173 );
buf ( n198175 , n30897 );
buf ( n198176 , n198175 );
buf ( n198177 , n198023 );
not ( n30901 , n198177 );
buf ( n198179 , n30901 );
buf ( n198180 , n198179 );
nor ( n30904 , n198176 , n198180 );
buf ( n198182 , n30904 );
buf ( n198183 , n198182 );
buf ( n30907 , n198183 );
buf ( n198185 , n30907 );
nor ( n30909 , n30895 , n198185 );
buf ( n198187 , n30909 );
nand ( n30911 , n30872 , n198187 );
buf ( n198189 , n30911 );
buf ( n198190 , n198189 );
xor ( n30914 , n198012 , n198013 );
and ( n30915 , n30914 , n198015 );
and ( n30916 , n198012 , n198013 );
or ( n30917 , n30915 , n30916 );
buf ( n198195 , n30917 );
buf ( n198196 , n198195 );
not ( n30920 , n198196 );
buf ( n198198 , n876 );
buf ( n198199 , n7818 );
xor ( n30923 , n198198 , n198199 );
buf ( n198201 , n7822 );
xor ( n30925 , n30923 , n198201 );
buf ( n198203 , n30925 );
buf ( n198204 , n198203 );
not ( n30928 , n198204 );
buf ( n198206 , n30928 );
buf ( n198207 , n198206 );
nand ( n30931 , n30920 , n198207 );
buf ( n198209 , n30931 );
buf ( n198210 , n198209 );
not ( n30934 , n198210 );
buf ( n198212 , n30934 );
buf ( n198213 , n198212 );
not ( n30937 , n198213 );
buf ( n198215 , n30937 );
buf ( n198216 , n198215 );
buf ( n198217 , n198203 );
buf ( n198218 , n198195 );
buf ( n30942 , n198218 );
buf ( n198220 , n30942 );
buf ( n198221 , n198220 );
nand ( n30945 , n198217 , n198221 );
buf ( n198223 , n30945 );
buf ( n198224 , n198223 );
and ( n30948 , n198216 , n198224 );
buf ( n198226 , n30948 );
buf ( n198227 , n198226 );
and ( n30951 , n198190 , n198227 );
not ( n30952 , n198190 );
buf ( n198230 , n198226 );
not ( n30954 , n198230 );
buf ( n198232 , n30954 );
buf ( n198233 , n198232 );
and ( n30957 , n30952 , n198233 );
nor ( n30958 , n30951 , n30957 );
buf ( n198236 , n30958 );
nand ( n30960 , n198236 , n168462 );
nand ( n30961 , n30704 , n30960 );
buf ( n30962 , n30961 );
not ( n30963 , n831 );
buf ( n198241 , n176193 );
not ( n30965 , n198241 );
buf ( n198243 , n30965 );
buf ( n198244 , n198243 );
buf ( n198245 , n176058 );
nand ( n30969 , n198244 , n198245 );
buf ( n198247 , n30969 );
buf ( n198248 , n198247 );
not ( n30972 , n198248 );
buf ( n198250 , n18819 );
not ( n30974 , n198250 );
buf ( n198252 , n30974 );
buf ( n198253 , n198252 );
not ( n30977 , n198253 );
buf ( n198255 , n30977 );
buf ( n198256 , n198255 );
not ( n30980 , n198256 );
or ( n30981 , n30972 , n30980 );
buf ( n198259 , n198252 );
not ( n30983 , n198259 );
buf ( n198261 , n30983 );
buf ( n198262 , n198261 );
buf ( n198263 , n198247 );
or ( n30987 , n198262 , n198263 );
nand ( n30988 , n30981 , n30987 );
buf ( n198266 , n30988 );
not ( n30990 , n198266 );
or ( n30991 , n30963 , n30990 );
not ( n30992 , n30733 );
and ( n30993 , n198153 , n30992 );
xor ( n30994 , n30993 , n198146 );
nand ( n30995 , n30994 , n168462 );
nand ( n30996 , n30991 , n30995 );
buf ( n30997 , n30996 );
nand ( n30998 , n182581 , n182251 );
buf ( n198276 , n30998 );
buf ( n198277 , n182944 );
buf ( n198278 , n182642 );
xor ( n31002 , n198277 , n198278 );
buf ( n198280 , n31002 );
buf ( n198281 , n198280 );
not ( n31005 , n198281 );
buf ( n198283 , n31005 );
buf ( n198284 , n198283 );
nand ( n31008 , n198276 , n198284 );
buf ( n198286 , n31008 );
buf ( n198287 , n198286 );
not ( n31011 , n198287 );
buf ( n198289 , n181436 );
buf ( n198290 , n181431 );
nand ( n31014 , n198289 , n198290 );
buf ( n198292 , n31014 );
buf ( n198293 , n198292 );
not ( n31017 , n198293 );
buf ( n198295 , n31017 );
not ( n31019 , n198295 );
buf ( n198297 , n181820 );
buf ( n198298 , n181810 );
xor ( n31022 , n198297 , n198298 );
buf ( n198300 , n31022 );
not ( n31024 , n198300 );
and ( n31025 , n31019 , n31024 );
buf ( n198303 , n181436 );
not ( n31027 , n198303 );
buf ( n198305 , n14477 );
not ( n31029 , n198305 );
or ( n31030 , n31027 , n31029 );
buf ( n198308 , n181844 );
buf ( n198309 , n181431 );
nand ( n31033 , n198308 , n198309 );
buf ( n198311 , n31033 );
buf ( n198312 , n198311 );
nand ( n31036 , n31030 , n198312 );
buf ( n198314 , n31036 );
buf ( n198315 , n198314 );
and ( n31039 , n180586 , n180968 );
buf ( n198317 , n31039 );
nor ( n31041 , n198315 , n198317 );
buf ( n198319 , n31041 );
nor ( n31043 , n31025 , n198319 );
and ( n31044 , n198297 , n198298 );
buf ( n198322 , n31044 );
buf ( n198323 , n198322 );
not ( n31047 , n198323 );
buf ( n198325 , n31047 );
buf ( n198326 , n198325 );
xnor ( n31050 , n182600 , n182594 );
buf ( n198328 , n31050 );
nand ( n31052 , n198326 , n198328 );
buf ( n198330 , n31052 );
buf ( n198331 , n182594 );
buf ( n198332 , n182600 );
nand ( n31056 , n198331 , n198332 );
buf ( n198334 , n31056 );
buf ( n198335 , n198334 );
xnor ( n31059 , n182251 , n182581 );
buf ( n198337 , n31059 );
nand ( n31061 , n198335 , n198337 );
buf ( n198339 , n31061 );
nand ( n31063 , n198330 , n198339 );
not ( n31064 , n31063 );
nand ( n31065 , n31043 , n31064 );
not ( n31066 , n31065 );
buf ( n198344 , n31066 );
not ( n31068 , n198344 );
buf ( n198346 , n31068 );
buf ( n198347 , n198346 );
nor ( n31071 , n31011 , n198347 );
buf ( n198349 , n31071 );
buf ( n198350 , n864 );
buf ( n198351 , n170630 );
xor ( n31075 , n198350 , n198351 );
buf ( n198353 , n171093 );
and ( n31077 , n31075 , n198353 );
and ( n31078 , n198350 , n198351 );
or ( n31079 , n31077 , n31078 );
buf ( n198357 , n31079 );
buf ( n198358 , n198357 );
buf ( n198359 , n171104 );
not ( n31083 , n198359 );
buf ( n198361 , n171638 );
not ( n31085 , n198361 );
or ( n31086 , n31083 , n31085 );
buf ( n198364 , n171635 );
buf ( n198365 , n171645 );
nand ( n31089 , n198364 , n198365 );
buf ( n198367 , n31089 );
buf ( n198368 , n198367 );
nand ( n31092 , n31086 , n198368 );
buf ( n198370 , n31092 );
buf ( n198371 , n198370 );
nor ( n31095 , n198358 , n198371 );
buf ( n198373 , n31095 );
not ( n31097 , n181029 );
not ( n31098 , n13682 );
or ( n31099 , n31097 , n31098 );
buf ( n198377 , n13656 );
buf ( n198378 , n181056 );
nand ( n31102 , n198377 , n198378 );
buf ( n198380 , n31102 );
nand ( n31104 , n31099 , n198380 );
buf ( n198382 , n31104 );
buf ( n198383 , n171635 );
buf ( n198384 , n171104 );
and ( n31108 , n198383 , n198384 );
buf ( n198386 , n31108 );
buf ( n198387 , n198386 );
nor ( n31111 , n198382 , n198387 );
buf ( n198389 , n31111 );
nor ( n31113 , n198373 , n198389 );
buf ( n198391 , n13649 );
not ( n31115 , n198391 );
buf ( n198393 , n13627 );
not ( n31117 , n198393 );
or ( n31118 , n31115 , n31117 );
buf ( n198396 , n13628 );
buf ( n198397 , n13652 );
nand ( n31121 , n198396 , n198397 );
buf ( n198399 , n31121 );
buf ( n198400 , n198399 );
nand ( n31124 , n31118 , n198400 );
buf ( n198402 , n31124 );
not ( n31126 , n198402 );
and ( n31127 , n13656 , n181029 );
not ( n31128 , n31127 );
and ( n31129 , n31126 , n31128 );
not ( n31130 , n12649 );
buf ( n198408 , n31130 );
not ( n31132 , n198408 );
buf ( n198410 , n180112 );
not ( n31134 , n198410 );
or ( n31135 , n31132 , n31134 );
not ( n31136 , n180112 );
nand ( n31137 , n31136 , n12649 );
buf ( n198415 , n31137 );
nand ( n31139 , n31135 , n198415 );
buf ( n198417 , n31139 );
buf ( n198418 , n198417 );
and ( n31142 , n13628 , n13649 );
buf ( n198420 , n31142 );
nor ( n31144 , n198418 , n198420 );
buf ( n198422 , n31144 );
nor ( n31146 , n31129 , n198422 );
nand ( n31147 , n31113 , n31146 );
not ( n31148 , n31147 );
and ( n31149 , n179706 , n179884 );
buf ( n198427 , n31149 );
not ( n31151 , n198427 );
buf ( n198429 , n180125 );
not ( n31153 , n198429 );
buf ( n198431 , n13167 );
not ( n31155 , n198431 );
or ( n31156 , n31153 , n31155 );
buf ( n198434 , n180546 );
buf ( n198435 , n13166 );
nand ( n31159 , n198434 , n198435 );
buf ( n198437 , n31159 );
buf ( n198438 , n198437 );
nand ( n31162 , n31156 , n198438 );
buf ( n198440 , n31162 );
buf ( n198441 , n198440 );
not ( n31165 , n198441 );
buf ( n198443 , n31165 );
buf ( n198444 , n198443 );
nand ( n31168 , n31151 , n198444 );
buf ( n198446 , n31168 );
buf ( n198447 , n198446 );
buf ( n198448 , n180509 );
not ( n31172 , n198448 );
buf ( n198450 , n180525 );
not ( n31174 , n198450 );
or ( n31175 , n31172 , n31174 );
buf ( n198453 , n180583 );
nand ( n31177 , n31175 , n198453 );
buf ( n198455 , n31177 );
not ( n31179 , n198455 );
not ( n31180 , n180971 );
or ( n31181 , n31179 , n31180 );
buf ( n198459 , n180968 );
buf ( n198460 , n13214 );
nand ( n31184 , n198459 , n198460 );
buf ( n198462 , n31184 );
nand ( n31186 , n31181 , n198462 );
buf ( n198464 , n13166 );
buf ( n198465 , n180125 );
and ( n31189 , n198464 , n198465 );
buf ( n198467 , n31189 );
nor ( n31191 , n31186 , n198467 );
buf ( n198469 , n12631 );
buf ( n198470 , n180014 );
xor ( n31194 , n198469 , n198470 );
buf ( n198472 , n31194 );
buf ( n198473 , n12649 );
buf ( n198474 , n180112 );
and ( n31198 , n198473 , n198474 );
buf ( n198476 , n31198 );
nor ( n31200 , n198472 , n198476 );
nor ( n31201 , n31191 , n31200 );
buf ( n198479 , n31201 );
and ( n31203 , n198469 , n198470 );
buf ( n198481 , n31203 );
not ( n31205 , n198481 );
xnor ( n31206 , n179706 , n179884 );
nand ( n31207 , n31205 , n31206 );
buf ( n198485 , n31207 );
nand ( n31209 , n198447 , n198479 , n198485 );
buf ( n198487 , n31209 );
buf ( n198488 , n198487 );
not ( n31212 , n198488 );
buf ( n198490 , n31212 );
nand ( n31214 , n31148 , n198490 );
not ( n31215 , n31214 );
and ( n31216 , n198349 , n31215 );
buf ( n198494 , n31216 );
not ( n31218 , n198494 );
buf ( n198496 , n870 );
buf ( n198497 , n173623 );
xor ( n31221 , n198496 , n198497 );
buf ( n198499 , n173628 );
xor ( n31223 , n31221 , n198499 );
buf ( n198501 , n31223 );
buf ( n198502 , n198501 );
buf ( n198503 , n871 );
buf ( n198504 , n174067 );
xor ( n31228 , n198503 , n198504 );
buf ( n198506 , n174072 );
and ( n31230 , n31228 , n198506 );
and ( n31231 , n198503 , n198504 );
or ( n31232 , n31230 , n31231 );
buf ( n198510 , n31232 );
buf ( n198511 , n198510 );
nor ( n31235 , n198502 , n198511 );
buf ( n198513 , n31235 );
buf ( n198514 , n198513 );
xor ( n31238 , n198503 , n198504 );
xor ( n31239 , n31238 , n198506 );
buf ( n198517 , n31239 );
buf ( n198518 , n198517 );
buf ( n198519 , n872 );
buf ( n198520 , n174151 );
xor ( n31244 , n198519 , n198520 );
buf ( n198522 , n174156 );
and ( n31246 , n31244 , n198522 );
and ( n31247 , n198519 , n198520 );
or ( n31248 , n31246 , n31247 );
buf ( n198526 , n31248 );
buf ( n198527 , n198526 );
nor ( n31251 , n198518 , n198527 );
buf ( n198529 , n31251 );
buf ( n198530 , n198529 );
nor ( n31254 , n198514 , n198530 );
buf ( n198532 , n31254 );
buf ( n198533 , n198532 );
not ( n31257 , n198533 );
buf ( n198535 , n31257 );
buf ( n198536 , n198535 );
not ( n31260 , n198536 );
buf ( n198538 , n31260 );
buf ( n198539 , n867 );
buf ( n198540 , n172802 );
xor ( n31264 , n198539 , n198540 );
buf ( n198542 , n172797 );
and ( n31266 , n31264 , n198542 );
and ( n31267 , n198539 , n198540 );
or ( n31268 , n31266 , n31267 );
buf ( n198546 , n31268 );
buf ( n198547 , n198546 );
not ( n31271 , n198547 );
buf ( n198549 , n866 );
buf ( n198550 , n172449 );
xor ( n31274 , n198549 , n198550 );
buf ( n198552 , n172478 );
xor ( n31276 , n31274 , n198552 );
buf ( n198554 , n31276 );
buf ( n198555 , n198554 );
not ( n31279 , n198555 );
buf ( n198557 , n31279 );
buf ( n198558 , n198557 );
nand ( n31282 , n31271 , n198558 );
buf ( n198560 , n31282 );
buf ( n198561 , n198560 );
buf ( n198562 , n868 );
buf ( n198563 , n173170 );
xor ( n31287 , n198562 , n198563 );
buf ( n198565 , n173175 );
and ( n31289 , n31287 , n198565 );
and ( n31290 , n198562 , n198563 );
or ( n31291 , n31289 , n31290 );
buf ( n198569 , n31291 );
buf ( n198570 , n198569 );
not ( n31294 , n198570 );
xor ( n31295 , n198539 , n198540 );
xor ( n31296 , n31295 , n198542 );
buf ( n198574 , n31296 );
buf ( n198575 , n198574 );
not ( n31299 , n198575 );
buf ( n198577 , n31299 );
buf ( n198578 , n198577 );
nand ( n31302 , n31294 , n198578 );
buf ( n198580 , n31302 );
buf ( n198581 , n198580 );
and ( n31305 , n198561 , n198581 );
buf ( n198583 , n31305 );
buf ( n198584 , n198212 );
not ( n31308 , n198584 );
buf ( n198586 , n198029 );
buf ( n198587 , n30734 );
nand ( n31311 , n31308 , n198586 , n198587 );
buf ( n198589 , n31311 );
buf ( n198590 , n198589 );
not ( n31314 , n198590 );
buf ( n198592 , n31314 );
and ( n31316 , n198538 , n198583 , n198592 );
xor ( n31317 , n198562 , n198563 );
xor ( n31318 , n31317 , n198565 );
buf ( n198596 , n31318 );
buf ( n198597 , n198596 );
buf ( n198598 , n869 );
buf ( n198599 , n173498 );
xor ( n31323 , n198598 , n198599 );
buf ( n198601 , n173503 );
and ( n31325 , n31323 , n198601 );
and ( n31326 , n198598 , n198599 );
or ( n31327 , n31325 , n31326 );
buf ( n198605 , n31327 );
buf ( n198606 , n198605 );
nor ( n31330 , n198597 , n198606 );
buf ( n198608 , n31330 );
buf ( n198609 , n198608 );
xor ( n31333 , n198598 , n198599 );
xor ( n31334 , n31333 , n198601 );
buf ( n198612 , n31334 );
buf ( n198613 , n198612 );
xor ( n31337 , n198496 , n198497 );
and ( n31338 , n31337 , n198499 );
and ( n31339 , n198496 , n198497 );
or ( n31340 , n31338 , n31339 );
buf ( n198618 , n31340 );
buf ( n198619 , n198618 );
nor ( n31343 , n198613 , n198619 );
buf ( n198621 , n31343 );
buf ( n198622 , n198621 );
nor ( n31346 , n198609 , n198622 );
buf ( n198624 , n31346 );
buf ( n198625 , n198624 );
buf ( n31349 , n198625 );
buf ( n198627 , n31349 );
buf ( n198628 , n198146 );
buf ( n31352 , n198628 );
buf ( n198630 , n31352 );
buf ( n198631 , n873 );
buf ( n198632 , n174438 );
xor ( n31356 , n198631 , n198632 );
buf ( n198634 , n174443 );
and ( n31358 , n31356 , n198634 );
and ( n31359 , n198631 , n198632 );
or ( n31360 , n31358 , n31359 );
buf ( n198638 , n31360 );
buf ( n198639 , n198638 );
xor ( n31363 , n198519 , n198520 );
xor ( n31364 , n31363 , n198522 );
buf ( n198642 , n31364 );
buf ( n198643 , n198642 );
nor ( n31367 , n198639 , n198643 );
buf ( n198645 , n31367 );
buf ( n198646 , n198645 );
buf ( n198647 , n874 );
buf ( n198648 , n7305 );
xor ( n31372 , n198647 , n198648 );
buf ( n198650 , n174761 );
and ( n31374 , n31372 , n198650 );
and ( n31375 , n198647 , n198648 );
or ( n31376 , n31374 , n31375 );
buf ( n198654 , n31376 );
buf ( n198655 , n198654 );
xor ( n31379 , n198631 , n198632 );
xor ( n31380 , n31379 , n198634 );
buf ( n198658 , n31380 );
buf ( n198659 , n198658 );
nor ( n31383 , n198655 , n198659 );
buf ( n198661 , n31383 );
buf ( n198662 , n198661 );
nor ( n31386 , n198646 , n198662 );
buf ( n198664 , n31386 );
buf ( n198665 , n198664 );
buf ( n198666 , n875 );
buf ( n198667 , n7577 );
xor ( n31391 , n198666 , n198667 );
buf ( n198669 , n7584 );
and ( n31393 , n31391 , n198669 );
and ( n31394 , n198666 , n198667 );
or ( n31395 , n31393 , n31394 );
buf ( n198673 , n31395 );
not ( n31397 , n198673 );
not ( n31398 , n31397 );
xor ( n31399 , n198647 , n198648 );
xor ( n31400 , n31399 , n198650 );
buf ( n198678 , n31400 );
buf ( n198679 , n198678 );
not ( n31403 , n198679 );
buf ( n198681 , n31403 );
not ( n31405 , n198681 );
or ( n31406 , n31398 , n31405 );
xor ( n31407 , n198666 , n198667 );
xor ( n31408 , n31407 , n198669 );
buf ( n198686 , n31408 );
buf ( n198687 , n198686 );
not ( n31411 , n198687 );
buf ( n198689 , n31411 );
xor ( n31413 , n198198 , n198199 );
and ( n31414 , n31413 , n198201 );
and ( n31415 , n198198 , n198199 );
or ( n31416 , n31414 , n31415 );
buf ( n198694 , n31416 );
buf ( n198695 , n198694 );
not ( n31419 , n198695 );
buf ( n198697 , n31419 );
nand ( n31421 , n198689 , n198697 );
nand ( n31422 , n31406 , n31421 );
not ( n31423 , n31422 );
buf ( n198701 , n31423 );
nand ( n31425 , n198665 , n198701 );
buf ( n198703 , n31425 );
buf ( n198704 , n198703 );
not ( n31428 , n198704 );
buf ( n198706 , n31428 );
and ( n31430 , n198627 , n198630 , n198706 );
buf ( n198708 , n865 );
buf ( n198709 , n172152 );
xor ( n31433 , n198708 , n198709 );
buf ( n198711 , n171675 );
and ( n31435 , n31433 , n198711 );
and ( n31436 , n198708 , n198709 );
or ( n31437 , n31435 , n31436 );
buf ( n198715 , n31437 );
buf ( n198716 , n198715 );
xor ( n31440 , n198350 , n198351 );
xor ( n31441 , n31440 , n198353 );
buf ( n198719 , n31441 );
buf ( n198720 , n198719 );
nor ( n31444 , n198716 , n198720 );
buf ( n198722 , n31444 );
xor ( n31446 , n198708 , n198709 );
xor ( n31447 , n31446 , n198711 );
buf ( n198725 , n31447 );
xor ( n31449 , n198549 , n198550 );
and ( n31450 , n31449 , n198552 );
and ( n31451 , n198549 , n198550 );
or ( n31452 , n31450 , n31451 );
buf ( n198730 , n31452 );
nor ( n31454 , n198725 , n198730 );
nor ( n31455 , n198722 , n31454 );
buf ( n198733 , n31455 );
buf ( n31457 , n198733 );
buf ( n198735 , n31457 );
nand ( n31459 , n31316 , n31430 , n198735 );
buf ( n198737 , n198722 );
not ( n31461 , n198737 );
buf ( n198739 , n31461 );
buf ( n198740 , n198608 );
buf ( n31464 , n198740 );
buf ( n198742 , n31464 );
buf ( n198743 , n198742 );
not ( n31467 , n198743 );
buf ( n198745 , n31467 );
or ( n31469 , n198725 , n198730 );
and ( n31470 , n198739 , n198745 , n31469 );
buf ( n198748 , n198608 );
not ( n31472 , n198748 );
buf ( n198750 , n198612 );
buf ( n198751 , n198618 );
nand ( n31475 , n198750 , n198751 );
buf ( n198753 , n31475 );
buf ( n198754 , n198753 );
not ( n31478 , n198754 );
and ( n31479 , n31472 , n31478 );
buf ( n198757 , n198596 );
buf ( n198758 , n198605 );
and ( n31482 , n198757 , n198758 );
buf ( n198760 , n31482 );
buf ( n198761 , n198760 );
nor ( n31485 , n31479 , n198761 );
buf ( n198763 , n31485 );
buf ( n198764 , n198763 );
not ( n31488 , n198764 );
buf ( n198766 , n31488 );
buf ( n198767 , n198766 );
not ( n31491 , n198767 );
buf ( n198769 , n198664 );
not ( n31493 , n198769 );
buf ( n198771 , n198686 );
buf ( n198772 , n198694 );
nand ( n31496 , n198771 , n198772 );
buf ( n198774 , n31496 );
buf ( n198775 , n198774 );
not ( n31499 , n198775 );
buf ( n198777 , n31499 );
buf ( n198778 , n198777 );
not ( n31502 , n198778 );
nand ( n31503 , n198681 , n31397 );
buf ( n198781 , n31503 );
not ( n31505 , n198781 );
or ( n31506 , n31502 , n31505 );
buf ( n198784 , n198681 );
not ( n31508 , n198784 );
buf ( n198786 , n198673 );
nand ( n31510 , n31508 , n198786 );
buf ( n198788 , n31510 );
buf ( n198789 , n198788 );
nand ( n31513 , n31506 , n198789 );
buf ( n198791 , n31513 );
buf ( n198792 , n198791 );
not ( n31516 , n198792 );
or ( n31517 , n31493 , n31516 );
buf ( n198795 , n198645 );
not ( n31519 , n198795 );
buf ( n198797 , n31519 );
buf ( n198798 , n198797 );
buf ( n198799 , n198658 );
buf ( n198800 , n198654 );
and ( n31524 , n198799 , n198800 );
buf ( n198802 , n31524 );
buf ( n198803 , n198802 );
and ( n31527 , n198798 , n198803 );
buf ( n198805 , n198642 );
buf ( n198806 , n198638 );
nand ( n31530 , n198805 , n198806 );
buf ( n198808 , n31530 );
buf ( n198809 , n198808 );
not ( n31533 , n198809 );
buf ( n198811 , n31533 );
buf ( n198812 , n198811 );
nor ( n31536 , n31527 , n198812 );
buf ( n198814 , n31536 );
buf ( n198815 , n198814 );
nand ( n31539 , n31517 , n198815 );
buf ( n198817 , n31539 );
buf ( n198818 , n198817 );
buf ( n198819 , n198517 );
buf ( n198820 , n198526 );
nand ( n31544 , n198819 , n198820 );
buf ( n198822 , n31544 );
buf ( n198823 , n198822 );
not ( n31547 , n198823 );
buf ( n198825 , n31547 );
buf ( n198826 , n198825 );
not ( n31550 , n198826 );
buf ( n198828 , n198513 );
not ( n31552 , n198828 );
buf ( n198830 , n31552 );
buf ( n198831 , n198830 );
not ( n31555 , n198831 );
or ( n31556 , n31550 , n31555 );
buf ( n198834 , n198501 );
buf ( n31558 , n198834 );
buf ( n198836 , n31558 );
buf ( n198837 , n198836 );
buf ( n198838 , n198510 );
nand ( n31562 , n198837 , n198838 );
buf ( n198840 , n31562 );
buf ( n198841 , n198840 );
nand ( n31565 , n31556 , n198841 );
buf ( n198843 , n31565 );
buf ( n198844 , n198843 );
nor ( n31568 , n198818 , n198844 );
buf ( n198846 , n31568 );
buf ( n198847 , n198846 );
buf ( n198848 , n198706 );
nor ( n31572 , n198212 , n198026 );
not ( n31573 , n31572 );
not ( n31574 , n30893 );
or ( n31575 , n31573 , n31574 );
not ( n31576 , n198182 );
not ( n31577 , n198209 );
or ( n31578 , n31576 , n31577 );
nand ( n31579 , n31578 , n198223 );
not ( n31580 , n31579 );
nand ( n31581 , n31575 , n31580 );
buf ( n198859 , n31581 );
nand ( n31583 , n198848 , n198859 );
buf ( n198861 , n31583 );
buf ( n198862 , n198861 );
nand ( n31586 , n31491 , n198847 , n198862 );
buf ( n198864 , n31586 );
buf ( n198865 , n198766 );
not ( n31589 , n198865 );
buf ( n198867 , n198843 );
buf ( n198868 , n198538 );
nor ( n31592 , n198867 , n198868 );
buf ( n198870 , n31592 );
buf ( n198871 , n198870 );
nand ( n31595 , n31589 , n198871 );
buf ( n198873 , n31595 );
buf ( n198874 , n198760 );
not ( n31598 , n198874 );
buf ( n198876 , n31598 );
buf ( n198877 , n198876 );
buf ( n198878 , n198621 );
nand ( n31602 , n198877 , n198878 );
buf ( n198880 , n31602 );
buf ( n198881 , n198880 );
buf ( n198882 , n198560 );
not ( n31606 , n198882 );
buf ( n198884 , n31606 );
buf ( n198885 , n198884 );
buf ( n198886 , n198580 );
not ( n31610 , n198886 );
buf ( n198888 , n31610 );
buf ( n198889 , n198888 );
nor ( n31613 , n198885 , n198889 );
buf ( n198891 , n31613 );
buf ( n198892 , n198891 );
and ( n31616 , n198881 , n198892 );
buf ( n198894 , n31616 );
nand ( n31618 , n31470 , n198864 , n198873 , n198894 );
not ( n31619 , n31455 );
buf ( n198897 , n198546 );
not ( n31621 , n198897 );
buf ( n198899 , n198557 );
nand ( n31623 , n31621 , n198899 );
buf ( n198901 , n31623 );
buf ( n198902 , n198901 );
not ( n31626 , n198902 );
buf ( n198904 , n198574 );
buf ( n198905 , n198569 );
nand ( n31629 , n198904 , n198905 );
buf ( n198907 , n31629 );
buf ( n198908 , n198907 );
not ( n31632 , n198908 );
buf ( n198910 , n31632 );
buf ( n198911 , n198910 );
not ( n31635 , n198911 );
or ( n31636 , n31626 , n31635 );
buf ( n198914 , n198546 );
buf ( n198915 , n198554 );
buf ( n31639 , n198915 );
buf ( n198917 , n31639 );
buf ( n198918 , n198917 );
nand ( n31642 , n198914 , n198918 );
buf ( n198920 , n31642 );
buf ( n198921 , n198920 );
nand ( n31645 , n31636 , n198921 );
buf ( n198923 , n31645 );
not ( n31647 , n198923 );
or ( n31648 , n31619 , n31647 );
buf ( n198926 , n198725 );
buf ( n198927 , n198730 );
nand ( n31651 , n198926 , n198927 );
buf ( n198929 , n31651 );
not ( n31653 , n198929 );
not ( n31654 , n198722 );
and ( n31655 , n31653 , n31654 );
buf ( n198933 , n198719 );
buf ( n31657 , n198933 );
buf ( n198935 , n31657 );
and ( n31659 , n198935 , n198715 );
nor ( n31660 , n31655 , n31659 );
nand ( n31661 , n31648 , n31660 );
not ( n31662 , n31661 );
nand ( n31663 , n31459 , n31618 , n31662 );
not ( n31664 , n31663 );
not ( n31665 , n31664 );
buf ( n198943 , n31665 );
not ( n31667 , n198943 );
or ( n31668 , n31218 , n31667 );
buf ( n198946 , n198349 );
not ( n31670 , n198946 );
buf ( n198948 , n198417 );
buf ( n198949 , n31142 );
nand ( n31673 , n198948 , n198949 );
buf ( n198951 , n31673 );
buf ( n198952 , n198951 );
buf ( n198953 , n198402 );
buf ( n198954 , n31127 );
nand ( n31678 , n198953 , n198954 );
buf ( n198956 , n31678 );
buf ( n198957 , n198956 );
and ( n31681 , n198952 , n198957 );
buf ( n198959 , n31681 );
buf ( n198960 , n198959 );
not ( n31684 , n198960 );
nand ( n31685 , n31104 , n198386 );
nand ( n31686 , n198370 , n31104 , n198357 );
nand ( n31687 , n31685 , n31686 );
nand ( n31688 , n31128 , n31126 );
nand ( n31689 , n31687 , n31688 );
buf ( n198967 , n31689 );
not ( n31691 , n198967 );
or ( n31692 , n31684 , n31691 );
buf ( n198970 , n198487 );
buf ( n198971 , n198417 );
buf ( n198972 , n31142 );
nor ( n31696 , n198971 , n198972 );
buf ( n198974 , n31696 );
buf ( n198975 , n198974 );
nor ( n31699 , n198970 , n198975 );
buf ( n198977 , n31699 );
buf ( n198978 , n198977 );
nand ( n31702 , n31692 , n198978 );
buf ( n198980 , n31702 );
buf ( n198981 , n31191 );
buf ( n31705 , n198981 );
buf ( n198983 , n31705 );
buf ( n198984 , n198983 );
buf ( n198985 , n198440 );
buf ( n198986 , n31149 );
nand ( n31710 , n198985 , n198986 );
buf ( n198988 , n31710 );
buf ( n198989 , n198988 );
or ( n31713 , n198984 , n198989 );
buf ( n198991 , n31186 );
buf ( n31715 , n198991 );
buf ( n198993 , n31715 );
buf ( n198994 , n198993 );
buf ( n198995 , n198467 );
buf ( n31719 , n198995 );
buf ( n198997 , n31719 );
buf ( n198998 , n198997 );
nand ( n31722 , n198994 , n198998 );
buf ( n199000 , n31722 );
buf ( n199001 , n199000 );
nand ( n31725 , n31713 , n199001 );
buf ( n199003 , n31725 );
not ( n31727 , n199003 );
buf ( n199005 , n198472 );
buf ( n199006 , n198476 );
and ( n31730 , n199005 , n199006 );
buf ( n199008 , n31730 );
buf ( n199009 , n199008 );
not ( n31733 , n199009 );
buf ( n199011 , n31207 );
not ( n31735 , n199011 );
or ( n31736 , n31733 , n31735 );
buf ( n199014 , n31206 );
not ( n31738 , n199014 );
buf ( n199016 , n198481 );
nand ( n31740 , n31738 , n199016 );
buf ( n199018 , n31740 );
buf ( n199019 , n199018 );
nand ( n31743 , n31736 , n199019 );
buf ( n199021 , n31743 );
not ( n31745 , n31149 );
not ( n31746 , n198440 );
and ( n31747 , n31745 , n31746 );
nor ( n31748 , n31747 , n198983 );
nand ( n31749 , n199021 , n31748 );
nand ( n31750 , n31727 , n31749 );
buf ( n199028 , n31750 );
not ( n31752 , n199028 );
buf ( n199030 , n31752 );
nand ( n31754 , n198980 , n199030 );
buf ( n199032 , n31754 );
not ( n31756 , n199032 );
or ( n31757 , n31670 , n31756 );
buf ( n199035 , n198286 );
not ( n31759 , n199035 );
not ( n31760 , n198300 );
nand ( n31761 , n31760 , n198292 );
buf ( n199039 , n31761 );
not ( n31763 , n199039 );
buf ( n199041 , n198314 );
buf ( n199042 , n31039 );
and ( n31766 , n199041 , n199042 );
buf ( n199044 , n31766 );
buf ( n199045 , n199044 );
not ( n31769 , n199045 );
or ( n31770 , n31763 , n31769 );
buf ( n199048 , n198295 );
buf ( n199049 , n198300 );
nand ( n31773 , n199048 , n199049 );
buf ( n199051 , n31773 );
buf ( n199052 , n199051 );
nand ( n31776 , n31770 , n199052 );
buf ( n199054 , n31776 );
buf ( n199055 , n199054 );
buf ( n199056 , n31064 );
nand ( n31780 , n199055 , n199056 );
buf ( n199058 , n31780 );
buf ( n199059 , n199058 );
not ( n31783 , n198339 );
buf ( n199061 , n198325 );
buf ( n199062 , n31050 );
nor ( n31786 , n199061 , n199062 );
buf ( n199064 , n31786 );
not ( n31788 , n199064 );
or ( n31789 , n31783 , n31788 );
or ( n31790 , n31059 , n198334 );
nand ( n31791 , n31789 , n31790 );
not ( n31792 , n31791 );
buf ( n199070 , n31792 );
nand ( n31794 , n199059 , n199070 );
buf ( n199072 , n31794 );
buf ( n199073 , n199072 );
not ( n31797 , n199073 );
or ( n31798 , n31759 , n31797 );
nor ( n31799 , n30998 , n198283 );
buf ( n199077 , n31799 );
not ( n31801 , n199077 );
buf ( n199079 , n31801 );
buf ( n199080 , n199079 );
nand ( n31804 , n31798 , n199080 );
buf ( n199082 , n31804 );
buf ( n199083 , n199082 );
not ( n31807 , n199083 );
buf ( n199085 , n31807 );
buf ( n199086 , n199085 );
nand ( n31810 , n31757 , n199086 );
buf ( n199088 , n31810 );
buf ( n199089 , n199088 );
not ( n31813 , n199089 );
buf ( n199091 , n31813 );
buf ( n199092 , n199091 );
nand ( n31816 , n31668 , n199092 );
buf ( n199094 , n31816 );
buf ( n199095 , n199094 );
not ( n31819 , n183233 );
not ( n31820 , n182960 );
or ( n31821 , n31819 , n31820 );
buf ( n199099 , n183240 );
buf ( n199100 , n183230 );
nand ( n31824 , n199099 , n199100 );
buf ( n199102 , n31824 );
nand ( n31826 , n31821 , n199102 );
and ( n31827 , n198277 , n198278 );
buf ( n199105 , n31827 );
or ( n31829 , n31826 , n199105 );
buf ( n199107 , n31829 );
nand ( n31831 , n199105 , n31826 );
buf ( n199109 , n31831 );
nand ( n31833 , n199107 , n199109 );
buf ( n199111 , n31833 );
buf ( n199112 , n199111 );
not ( n31836 , n199112 );
buf ( n199114 , n31836 );
buf ( n199115 , n199114 );
and ( n31839 , n199095 , n199115 );
not ( n31840 , n199095 );
buf ( n199118 , n199111 );
and ( n31842 , n31840 , n199118 );
nor ( n31843 , n31839 , n31842 );
buf ( n199121 , n31843 );
and ( n31845 , n168462 , n199121 );
not ( n31846 , n168462 );
and ( n31847 , n31846 , n184086 );
nor ( n31848 , n31845 , n31847 );
nand ( n31849 , n185731 , n831 );
buf ( n31850 , n31663 );
nor ( n31851 , n31214 , n198346 );
and ( n31852 , n31850 , n31851 );
buf ( n199130 , n31066 );
not ( n31854 , n199130 );
buf ( n199132 , n31754 );
not ( n31856 , n199132 );
or ( n31857 , n31854 , n31856 );
buf ( n199135 , n199072 );
not ( n31859 , n199135 );
buf ( n199137 , n31859 );
buf ( n199138 , n199137 );
nand ( n31862 , n31857 , n199138 );
buf ( n199140 , n31862 );
nor ( n31864 , n31852 , n199140 );
buf ( n199142 , n31864 );
buf ( n199143 , n198286 );
buf ( n199144 , n199079 );
nand ( n31868 , n199143 , n199144 );
buf ( n199146 , n31868 );
not ( n31870 , n199146 );
nand ( n31871 , n31870 , n168462 );
buf ( n199149 , n31871 );
and ( n31873 , n199142 , n199149 );
not ( n31874 , n199142 );
nand ( n31875 , n199146 , n168462 );
buf ( n199153 , n31875 );
and ( n31877 , n31874 , n199153 );
or ( n31878 , n31873 , n31877 );
buf ( n199156 , n31878 );
nand ( n31880 , n31849 , n199156 );
buf ( n199158 , n176204 );
not ( n31882 , n199158 );
buf ( n199160 , n177669 );
not ( n31884 , n199160 );
or ( n31885 , n31882 , n31884 );
not ( n31886 , n8307 );
not ( n31887 , n176082 );
or ( n31888 , n31886 , n31887 );
nand ( n31889 , n31888 , n176107 );
buf ( n199167 , n31889 );
not ( n31891 , n199167 );
buf ( n199169 , n31891 );
buf ( n199170 , n199169 );
nand ( n31894 , n31885 , n199170 );
buf ( n199172 , n31894 );
nand ( n31896 , n18433 , n18437 );
not ( n31897 , n31896 );
and ( n31898 , n199172 , n31897 );
not ( n31899 , n199172 );
and ( n31900 , n31899 , n31896 );
nor ( n31901 , n31898 , n31900 );
nand ( n31902 , n31901 , n831 );
buf ( n199180 , n198592 );
not ( n31904 , n199180 );
buf ( n199182 , n198090 );
not ( n31906 , n199182 );
buf ( n199184 , n197536 );
not ( n31908 , n199184 );
or ( n31909 , n31906 , n31908 );
buf ( n199187 , n198143 );
nand ( n31911 , n31909 , n199187 );
buf ( n199189 , n31911 );
buf ( n199190 , n199189 );
not ( n31914 , n199190 );
or ( n31915 , n31904 , n31914 );
buf ( n199193 , n31581 );
not ( n31917 , n199193 );
buf ( n199195 , n31917 );
buf ( n199196 , n199195 );
nand ( n31920 , n31915 , n199196 );
buf ( n199198 , n31920 );
buf ( n199199 , n199198 );
buf ( n199200 , n31421 );
buf ( n31924 , n199200 );
buf ( n199202 , n31924 );
buf ( n199203 , n199202 );
buf ( n199204 , n198774 );
buf ( n31928 , n199204 );
buf ( n199206 , n31928 );
buf ( n199207 , n199206 );
nand ( n31931 , n199203 , n199207 );
buf ( n199209 , n31931 );
buf ( n199210 , n199209 );
not ( n31934 , n199210 );
buf ( n199212 , n31934 );
buf ( n199213 , n199212 );
and ( n31937 , n199199 , n199213 );
not ( n31938 , n199199 );
buf ( n199216 , n199209 );
and ( n31940 , n31938 , n199216 );
nor ( n31941 , n31937 , n31940 );
buf ( n199219 , n31941 );
nand ( n31943 , n199219 , n168462 );
nand ( n31944 , n31902 , n31943 );
not ( n31945 , n168462 );
not ( n31946 , n30992 );
not ( n31947 , n199189 );
or ( n31948 , n31946 , n31947 );
nand ( n31949 , n31948 , n198153 );
buf ( n199227 , n31949 );
buf ( n199228 , n198168 );
buf ( n199229 , n198157 );
nand ( n31953 , n199228 , n199229 );
buf ( n199231 , n31953 );
buf ( n199232 , n199231 );
not ( n31956 , n199232 );
buf ( n199234 , n31956 );
buf ( n199235 , n199234 );
and ( n31959 , n199227 , n199235 );
not ( n31960 , n199227 );
buf ( n199238 , n199231 );
and ( n31962 , n31960 , n199238 );
nor ( n31963 , n31959 , n31962 );
buf ( n199241 , n31963 );
not ( n31965 , n199241 );
or ( n31966 , n31945 , n31965 );
buf ( n199244 , n198243 );
not ( n31968 , n199244 );
buf ( n199246 , n18819 );
not ( n31970 , n199246 );
or ( n31971 , n31968 , n31970 );
buf ( n199249 , n176058 );
nand ( n31973 , n31971 , n199249 );
buf ( n199251 , n31973 );
buf ( n199252 , n199251 );
buf ( n199253 , n8652 );
buf ( n199254 , n176072 );
nand ( n31978 , n199253 , n199254 );
buf ( n199256 , n31978 );
buf ( n199257 , n199256 );
not ( n31981 , n199257 );
buf ( n199259 , n31981 );
buf ( n199260 , n199259 );
and ( n31984 , n199252 , n199260 );
not ( n31985 , n199252 );
buf ( n199263 , n199256 );
and ( n31987 , n31985 , n199263 );
nor ( n31988 , n31984 , n31987 );
buf ( n199266 , n31988 );
nand ( n31990 , n199266 , n831 );
nand ( n31991 , n31966 , n31990 );
buf ( n199269 , n31148 );
not ( n31993 , n199269 );
buf ( n199271 , n31459 );
buf ( n199272 , n31618 );
buf ( n199273 , n31662 );
nand ( n31997 , n199271 , n199272 , n199273 );
buf ( n199275 , n31997 );
buf ( n199276 , n199275 );
buf ( n32000 , n199276 );
buf ( n199278 , n32000 );
buf ( n199279 , n199278 );
not ( n32003 , n199279 );
or ( n32004 , n31993 , n32003 );
and ( n32005 , n31126 , n31128 );
nor ( n32006 , n32005 , n198422 );
not ( n32007 , n32006 );
not ( n32008 , n31687 );
or ( n32009 , n32007 , n32008 );
not ( n32010 , n198956 );
not ( n32011 , n198974 );
and ( n32012 , n32010 , n32011 );
not ( n32013 , n198951 );
nor ( n32014 , n32012 , n32013 );
nand ( n32015 , n32009 , n32014 );
buf ( n199293 , n32015 );
not ( n32017 , n199293 );
buf ( n199295 , n32017 );
buf ( n199296 , n199295 );
nand ( n32020 , n32004 , n199296 );
buf ( n199298 , n32020 );
buf ( n199299 , n199298 );
buf ( n32023 , n31200 );
not ( n32024 , n32023 );
buf ( n32025 , n199008 );
buf ( n199303 , n32025 );
not ( n32027 , n199303 );
buf ( n199305 , n32027 );
nand ( n32029 , n32024 , n199305 );
buf ( n199307 , n32029 );
not ( n32031 , n199307 );
buf ( n199309 , n32031 );
buf ( n199310 , n199309 );
and ( n32034 , n199299 , n199310 );
not ( n32035 , n199299 );
buf ( n199313 , n32029 );
and ( n32037 , n32035 , n199313 );
nor ( n32038 , n32034 , n32037 );
buf ( n199316 , n32038 );
nand ( n32040 , n199316 , n168462 );
or ( n32041 , n177380 , n177430 );
buf ( n199319 , n32041 );
not ( n32043 , n199319 );
buf ( n199321 , n10146 );
not ( n32045 , n199321 );
or ( n32046 , n32043 , n32045 );
buf ( n199324 , n177433 );
nand ( n32048 , n32046 , n199324 );
buf ( n199326 , n32048 );
buf ( n199327 , n199326 );
buf ( n199328 , n177442 );
buf ( n199329 , n177376 );
not ( n32053 , n199329 );
buf ( n199331 , n32053 );
buf ( n199332 , n199331 );
nand ( n32056 , n199328 , n199332 );
buf ( n199334 , n32056 );
buf ( n199335 , n199334 );
not ( n32059 , n199335 );
buf ( n199337 , n32059 );
buf ( n199338 , n199337 );
and ( n32062 , n199327 , n199338 );
not ( n32063 , n199327 );
buf ( n199341 , n199334 );
and ( n32065 , n32063 , n199341 );
nor ( n32066 , n32062 , n32065 );
buf ( n199344 , n32066 );
nand ( n32068 , n199344 , n831 );
nand ( n32069 , n18813 , n831 );
buf ( n199347 , n30472 );
buf ( n199348 , n197226 );
not ( n32072 , n199348 );
buf ( n199350 , n32072 );
buf ( n199351 , n199350 );
buf ( n199352 , n197372 );
nand ( n32076 , n199351 , n199352 );
buf ( n199354 , n32076 );
buf ( n199355 , n199354 );
and ( n32079 , n199347 , n199355 );
not ( n32080 , n199347 );
buf ( n199358 , n199354 );
not ( n32082 , n199358 );
buf ( n199360 , n32082 );
buf ( n199361 , n199360 );
and ( n32085 , n32080 , n199361 );
nor ( n32086 , n32079 , n32085 );
buf ( n199364 , n32086 );
nand ( n32088 , n199364 , n168462 );
nand ( n32089 , n184019 , n831 );
nand ( n32090 , n185951 , n831 );
not ( n32091 , n30734 );
not ( n32092 , n199189 );
or ( n32093 , n32091 , n32092 );
not ( n32094 , n30894 );
nand ( n32095 , n32093 , n32094 );
buf ( n199373 , n32095 );
buf ( n199374 , n198185 );
not ( n32098 , n199374 );
buf ( n199376 , n198029 );
nand ( n32100 , n32098 , n199376 );
buf ( n199378 , n32100 );
buf ( n199379 , n199378 );
not ( n32103 , n199379 );
buf ( n199381 , n32103 );
buf ( n199382 , n199381 );
and ( n32106 , n199373 , n199382 );
not ( n32107 , n199373 );
buf ( n199385 , n199378 );
and ( n32109 , n32107 , n199385 );
nor ( n32110 , n32106 , n32109 );
buf ( n199388 , n32110 );
nand ( n32112 , n199388 , n168462 );
not ( n32113 , n31754 );
buf ( n199391 , n198624 );
not ( n32115 , n199391 );
buf ( n199393 , n198843 );
not ( n32117 , n199393 );
or ( n32118 , n32115 , n32117 );
buf ( n199396 , n198763 );
nand ( n32120 , n32118 , n199396 );
buf ( n199398 , n32120 );
buf ( n199399 , n199398 );
buf ( n32123 , n199399 );
buf ( n199401 , n32123 );
nor ( n32125 , n31661 , n199401 );
not ( n32126 , n32125 );
or ( n32127 , n198817 , n198706 );
buf ( n199405 , n198624 );
buf ( n199406 , n198532 );
and ( n32130 , n199405 , n199406 );
buf ( n199408 , n32130 );
buf ( n199409 , n199408 );
buf ( n32133 , n199409 );
buf ( n199411 , n32133 );
buf ( n199412 , n198630 );
buf ( n199413 , n198592 );
nand ( n32137 , n199412 , n199413 );
buf ( n199415 , n32137 );
buf ( n199416 , n199415 );
buf ( n199417 , n198817 );
not ( n32141 , n199417 );
buf ( n199419 , n32141 );
buf ( n199420 , n199419 );
buf ( n199421 , n199195 );
nand ( n32145 , n199416 , n199420 , n199421 );
buf ( n199423 , n32145 );
nand ( n32147 , n32127 , n199411 , n199423 );
not ( n32148 , n32147 );
or ( n32149 , n32126 , n32148 );
nand ( n32150 , n31469 , n198739 );
not ( n32151 , n32150 );
buf ( n32152 , n198891 );
nand ( n32153 , n32151 , n32152 );
and ( n32154 , n32153 , n31662 );
nor ( n32155 , n32154 , n31214 );
nand ( n32156 , n32149 , n32155 );
nand ( n32157 , n32113 , n32156 );
buf ( n199435 , n32157 );
buf ( n199436 , n198319 );
not ( n32160 , n199436 );
buf ( n199438 , n32160 );
buf ( n199439 , n199438 );
buf ( n199440 , n199044 );
not ( n32164 , n199440 );
buf ( n199442 , n32164 );
buf ( n199443 , n199442 );
nand ( n32167 , n199439 , n199443 );
buf ( n199445 , n32167 );
buf ( n199446 , n199445 );
xnor ( n32170 , n199435 , n199446 );
buf ( n199448 , n32170 );
nand ( n32172 , n199448 , n168462 );
buf ( n32173 , n31207 );
not ( n32174 , n32173 );
nor ( n32175 , n32174 , n32023 );
buf ( n199453 , n32175 );
buf ( n199454 , n198446 );
buf ( n32178 , n199454 );
buf ( n199456 , n32178 );
buf ( n199457 , n199456 );
nand ( n32181 , n199453 , n199457 );
buf ( n199459 , n32181 );
buf ( n199460 , n199459 );
buf ( n199461 , n31147 );
nor ( n32185 , n199460 , n199461 );
buf ( n199463 , n32185 );
buf ( n199464 , n199463 );
not ( n32188 , n199464 );
buf ( n199466 , n31665 );
not ( n32190 , n199466 );
or ( n32191 , n32188 , n32190 );
buf ( n199469 , n32015 );
not ( n32193 , n199469 );
not ( n32194 , n199459 );
buf ( n199472 , n32194 );
not ( n32196 , n199472 );
or ( n32197 , n32193 , n32196 );
buf ( n199475 , n199456 );
not ( n32199 , n199475 );
buf ( n199477 , n199021 );
buf ( n32201 , n199477 );
buf ( n199479 , n32201 );
buf ( n199480 , n199479 );
not ( n32204 , n199480 );
or ( n32205 , n32199 , n32204 );
buf ( n199483 , n198988 );
nand ( n32207 , n32205 , n199483 );
buf ( n199485 , n32207 );
buf ( n199486 , n199485 );
not ( n32210 , n199486 );
buf ( n199488 , n32210 );
buf ( n199489 , n199488 );
nand ( n32213 , n32197 , n199489 );
buf ( n199491 , n32213 );
buf ( n199492 , n199491 );
not ( n32216 , n199492 );
buf ( n199494 , n32216 );
buf ( n199495 , n199494 );
nand ( n32219 , n32191 , n199495 );
buf ( n199497 , n32219 );
buf ( n199498 , n199497 );
buf ( n199499 , n198983 );
not ( n32223 , n199499 );
buf ( n199501 , n199000 );
nand ( n32225 , n32223 , n199501 );
buf ( n199503 , n32225 );
buf ( n199504 , n199503 );
not ( n32228 , n199504 );
buf ( n199506 , n32228 );
buf ( n199507 , n199506 );
and ( n32231 , n199498 , n199507 );
not ( n32232 , n199498 );
buf ( n199510 , n199503 );
and ( n32234 , n32232 , n199510 );
nor ( n32235 , n32231 , n32234 );
buf ( n199513 , n32235 );
nand ( n32237 , n199513 , n168462 );
xor ( n32238 , n187025 , n187070 );
xor ( n32239 , n32238 , n187082 );
buf ( n199517 , n32239 );
buf ( n199518 , n187107 );
buf ( n199519 , n844 );
buf ( n199520 , n870 );
xor ( n32244 , n199519 , n199520 );
buf ( n199522 , n32244 );
buf ( n199523 , n199522 );
not ( n32247 , n199523 );
buf ( n199525 , n186435 );
not ( n32249 , n199525 );
or ( n32250 , n32247 , n32249 );
buf ( n199528 , n186444 );
buf ( n199529 , n19835 );
nand ( n32253 , n199528 , n199529 );
buf ( n199531 , n32253 );
buf ( n199532 , n199531 );
nand ( n32256 , n32250 , n199532 );
buf ( n199534 , n32256 );
buf ( n199535 , n199534 );
xor ( n32259 , n199518 , n199535 );
buf ( n199537 , n851 );
buf ( n199538 , n864 );
xor ( n32262 , n199537 , n199538 );
buf ( n199540 , n32262 );
buf ( n199541 , n199540 );
not ( n32265 , n199541 );
buf ( n199543 , n19031 );
not ( n32267 , n199543 );
or ( n32268 , n32265 , n32267 );
buf ( n199546 , n186340 );
buf ( n199547 , n187278 );
nand ( n32271 , n199546 , n199547 );
buf ( n199549 , n32271 );
buf ( n199550 , n199549 );
nand ( n32274 , n32268 , n199550 );
buf ( n199552 , n32274 );
buf ( n199553 , n199552 );
not ( n32277 , n199553 );
buf ( n199555 , n835 );
buf ( n199556 , n880 );
xor ( n32280 , n199555 , n199556 );
buf ( n199558 , n32280 );
buf ( n199559 , n199558 );
not ( n32283 , n199559 );
buf ( n199561 , n18862 );
not ( n32285 , n199561 );
or ( n32286 , n32283 , n32285 );
buf ( n199564 , n18875 );
buf ( n199565 , n187100 );
nand ( n32289 , n199564 , n199565 );
buf ( n199567 , n32289 );
buf ( n199568 , n199567 );
nand ( n32292 , n32286 , n199568 );
buf ( n199570 , n32292 );
buf ( n199571 , n199570 );
not ( n32295 , n199571 );
or ( n32296 , n32277 , n32295 );
buf ( n199574 , n199570 );
buf ( n199575 , n199552 );
or ( n32299 , n199574 , n199575 );
buf ( n199577 , n849 );
buf ( n199578 , n866 );
xor ( n32302 , n199577 , n199578 );
buf ( n199580 , n32302 );
buf ( n199581 , n199580 );
not ( n32305 , n199581 );
buf ( n199583 , n186241 );
not ( n32307 , n199583 );
or ( n32308 , n32305 , n32307 );
buf ( n199586 , n186254 );
buf ( n199587 , n187156 );
nand ( n32311 , n199586 , n199587 );
buf ( n199589 , n32311 );
buf ( n199590 , n199589 );
nand ( n32314 , n32308 , n199590 );
buf ( n199592 , n32314 );
buf ( n199593 , n199592 );
nand ( n32317 , n32299 , n199593 );
buf ( n199595 , n32317 );
buf ( n199596 , n199595 );
nand ( n32320 , n32296 , n199596 );
buf ( n199598 , n32320 );
buf ( n199599 , n199598 );
and ( n32323 , n32259 , n199599 );
and ( n32324 , n199518 , n199535 );
or ( n32325 , n32323 , n32324 );
buf ( n199603 , n32325 );
buf ( n199604 , n199603 );
xor ( n32328 , n187111 , n187125 );
xor ( n32329 , n32328 , n187143 );
buf ( n199607 , n32329 );
buf ( n199608 , n199607 );
xor ( n32332 , n199604 , n199608 );
buf ( n199610 , n852 );
buf ( n199611 , n864 );
and ( n32335 , n199610 , n199611 );
buf ( n199613 , n32335 );
buf ( n199614 , n199613 );
buf ( n199615 , n843 );
buf ( n199616 , n872 );
xor ( n32340 , n199615 , n199616 );
buf ( n199618 , n32340 );
buf ( n199619 , n199618 );
not ( n32343 , n199619 );
buf ( n199621 , n19260 );
not ( n32345 , n199621 );
or ( n32346 , n32343 , n32345 );
buf ( n199624 , n19265 );
buf ( n199625 , n187232 );
nand ( n32349 , n199624 , n199625 );
buf ( n199627 , n32349 );
buf ( n199628 , n199627 );
nand ( n32352 , n32346 , n199628 );
buf ( n199630 , n32352 );
buf ( n199631 , n199630 );
xor ( n32355 , n199614 , n199631 );
buf ( n199633 , n841 );
buf ( n199634 , n874 );
xor ( n32358 , n199633 , n199634 );
buf ( n199636 , n32358 );
buf ( n199637 , n199636 );
not ( n32361 , n199637 );
buf ( n199639 , n186287 );
not ( n32363 , n199639 );
or ( n32364 , n32361 , n32363 );
buf ( n199642 , n186297 );
buf ( n199643 , n187296 );
nand ( n32367 , n199642 , n199643 );
buf ( n199645 , n32367 );
buf ( n199646 , n199645 );
nand ( n32370 , n32364 , n199646 );
buf ( n199648 , n32370 );
buf ( n199649 , n199648 );
and ( n32373 , n32355 , n199649 );
and ( n32374 , n199614 , n199631 );
or ( n32375 , n32373 , n32374 );
buf ( n199653 , n32375 );
buf ( n199654 , n199653 );
buf ( n199655 , n847 );
buf ( n199656 , n868 );
xor ( n32380 , n199655 , n199656 );
buf ( n199658 , n32380 );
buf ( n199659 , n199658 );
not ( n32383 , n199659 );
buf ( n199661 , n186197 );
not ( n32385 , n199661 );
or ( n32386 , n32383 , n32385 );
buf ( n199664 , n18907 );
buf ( n199665 , n19893 );
nand ( n32389 , n199664 , n199665 );
buf ( n199667 , n32389 );
buf ( n199668 , n199667 );
nand ( n32392 , n32386 , n199668 );
buf ( n199670 , n32392 );
buf ( n199671 , n199670 );
buf ( n199672 , n839 );
buf ( n199673 , n876 );
xor ( n32397 , n199672 , n199673 );
buf ( n199675 , n32397 );
buf ( n199676 , n199675 );
not ( n32400 , n199676 );
buf ( n199678 , n19098 );
not ( n32402 , n199678 );
or ( n32403 , n32400 , n32402 );
buf ( n199681 , n186395 );
buf ( n199682 , n19908 );
nand ( n32406 , n199681 , n199682 );
buf ( n199684 , n32406 );
buf ( n199685 , n199684 );
nand ( n32409 , n32403 , n199685 );
buf ( n199687 , n32409 );
buf ( n199688 , n199687 );
xor ( n32412 , n199671 , n199688 );
buf ( n199690 , n845 );
buf ( n199691 , n870 );
xor ( n32415 , n199690 , n199691 );
buf ( n199693 , n32415 );
buf ( n199694 , n199693 );
not ( n32418 , n199694 );
buf ( n199696 , n186435 );
not ( n32420 , n199696 );
or ( n32421 , n32418 , n32420 );
buf ( n199699 , n186444 );
buf ( n199700 , n199522 );
nand ( n32424 , n199699 , n199700 );
buf ( n199702 , n32424 );
buf ( n199703 , n199702 );
nand ( n32427 , n32421 , n199703 );
buf ( n199705 , n32427 );
buf ( n199706 , n199705 );
and ( n32430 , n32412 , n199706 );
and ( n32431 , n199671 , n199688 );
or ( n32432 , n32430 , n32431 );
buf ( n199710 , n32432 );
buf ( n199711 , n199710 );
xor ( n32435 , n199654 , n199711 );
buf ( n199713 , n192332 );
buf ( n199714 , n192573 );
or ( n32438 , n199713 , n199714 );
buf ( n199716 , n884 );
nand ( n32440 , n32438 , n199716 );
buf ( n199718 , n32440 );
buf ( n199719 , n199718 );
xor ( n32443 , n882 , n833 );
buf ( n199721 , n32443 );
not ( n32445 , n199721 );
buf ( n199723 , n26567 );
not ( n32447 , n199723 );
or ( n32448 , n32445 , n32447 );
buf ( n199726 , n19943 );
buf ( n199727 , n187207 );
nand ( n32451 , n199726 , n199727 );
buf ( n199729 , n32451 );
buf ( n199730 , n199729 );
nand ( n32454 , n32448 , n199730 );
buf ( n199732 , n32454 );
buf ( n199733 , n199732 );
xor ( n32457 , n199719 , n199733 );
buf ( n199735 , n837 );
buf ( n199736 , n878 );
xor ( n32460 , n199735 , n199736 );
buf ( n199738 , n32460 );
buf ( n199739 , n199738 );
not ( n32463 , n199739 );
buf ( n199741 , n186789 );
not ( n32465 , n199741 );
or ( n32466 , n32463 , n32465 );
buf ( n199744 , n186575 );
buf ( n199745 , n187250 );
nand ( n32469 , n199744 , n199745 );
buf ( n199747 , n32469 );
buf ( n199748 , n199747 );
nand ( n32472 , n32466 , n199748 );
buf ( n199750 , n32472 );
buf ( n199751 , n199750 );
and ( n32475 , n32457 , n199751 );
and ( n32476 , n199719 , n199733 );
or ( n32477 , n32475 , n32476 );
buf ( n199755 , n32477 );
buf ( n199756 , n199755 );
and ( n32480 , n32435 , n199756 );
and ( n32481 , n199654 , n199711 );
or ( n32482 , n32480 , n32481 );
buf ( n199760 , n32482 );
buf ( n199761 , n199760 );
and ( n32485 , n32332 , n199761 );
and ( n32486 , n199604 , n199608 );
or ( n32487 , n32485 , n32486 );
buf ( n199765 , n32487 );
xor ( n32489 , n187148 , n187151 );
xor ( n32490 , n32489 , n187319 );
buf ( n199768 , n32490 );
xor ( n32492 , n199765 , n199768 );
xor ( n32493 , n187228 , n187245 );
xor ( n32494 , n32493 , n187263 );
buf ( n199772 , n32494 );
buf ( n199773 , n199772 );
xor ( n32497 , n187169 , n187183 );
xor ( n32498 , n32497 , n187198 );
buf ( n199776 , n32498 );
buf ( n199777 , n199776 );
or ( n32501 , n199773 , n199777 );
xor ( n32502 , n187274 , n187291 );
xor ( n32503 , n32502 , n187309 );
buf ( n199781 , n32503 );
buf ( n199782 , n199781 );
nand ( n32506 , n32501 , n199782 );
buf ( n199784 , n32506 );
buf ( n199785 , n199784 );
buf ( n199786 , n199772 );
buf ( n199787 , n199776 );
nand ( n32511 , n199786 , n199787 );
buf ( n199789 , n32511 );
buf ( n199790 , n199789 );
nand ( n32514 , n199785 , n199790 );
buf ( n199792 , n32514 );
buf ( n199793 , n199792 );
xor ( n32517 , n187203 , n187268 );
xor ( n32518 , n32517 , n187314 );
buf ( n199796 , n32518 );
buf ( n199797 , n199796 );
xor ( n32521 , n199793 , n199797 );
xor ( n32522 , n20050 , n187330 );
xor ( n32523 , n32522 , n187351 );
buf ( n199801 , n32523 );
and ( n32525 , n32521 , n199801 );
and ( n32526 , n199793 , n199797 );
or ( n32527 , n32525 , n32526 );
buf ( n199805 , n32527 );
and ( n32529 , n32492 , n199805 );
and ( n32530 , n199765 , n199768 );
or ( n32531 , n32529 , n32530 );
xor ( n32532 , n199517 , n32531 );
xor ( n32533 , n187095 , n187324 );
xor ( n32534 , n32533 , n187398 );
buf ( n199812 , n32534 );
and ( n32536 , n32532 , n199812 );
and ( n32537 , n199517 , n32531 );
or ( n32538 , n32536 , n32537 );
not ( n32539 , n32538 );
not ( n32540 , n187405 );
nand ( n32541 , n32539 , n32540 );
xor ( n32542 , n186711 , n187090 );
and ( n32543 , n32542 , n187403 );
and ( n32544 , n186711 , n187090 );
or ( n32545 , n32543 , n32544 );
buf ( n199823 , n32545 );
not ( n32547 , n199823 );
not ( n32548 , n193688 );
nand ( n32549 , n32547 , n32548 );
nand ( n32550 , n32541 , n32549 );
xor ( n32551 , n193526 , n193679 );
and ( n32552 , n32551 , n193686 );
and ( n32553 , n193526 , n193679 );
or ( n32554 , n32552 , n32553 );
buf ( n199832 , n32554 );
not ( n32556 , n199832 );
xor ( n32557 , n193499 , n193505 );
and ( n32558 , n32557 , n193523 );
and ( n32559 , n193499 , n193505 );
or ( n32560 , n32558 , n32559 );
buf ( n199838 , n32560 );
buf ( n199839 , n199838 );
xor ( n32563 , n193537 , n193554 );
and ( n32564 , n32563 , n193572 );
and ( n32565 , n193537 , n193554 );
or ( n32566 , n32564 , n32565 );
buf ( n199844 , n32566 );
buf ( n199845 , n199844 );
xor ( n32569 , n193592 , n193609 );
and ( n32570 , n32569 , n193627 );
and ( n32571 , n193592 , n193609 );
or ( n32572 , n32570 , n32571 );
buf ( n199850 , n32572 );
buf ( n199851 , n199850 );
xor ( n32575 , n199845 , n199851 );
buf ( n199853 , n193585 );
not ( n32577 , n199853 );
buf ( n199855 , n186241 );
not ( n32579 , n199855 );
or ( n32580 , n32577 , n32579 );
buf ( n199858 , n186254 );
buf ( n199859 , n196819 );
nand ( n32583 , n199858 , n199859 );
buf ( n199861 , n32583 );
buf ( n199862 , n199861 );
nand ( n32586 , n32580 , n199862 );
buf ( n199864 , n32586 );
buf ( n199865 , n199864 );
buf ( n199866 , n26361 );
not ( n32590 , n199866 );
buf ( n199868 , n19260 );
not ( n32592 , n199868 );
or ( n32593 , n32590 , n32592 );
buf ( n199871 , n19265 );
buf ( n199872 , n196724 );
nand ( n32596 , n199871 , n199872 );
buf ( n199874 , n32596 );
buf ( n199875 , n199874 );
nand ( n32599 , n32593 , n199875 );
buf ( n199877 , n32599 );
buf ( n199878 , n199877 );
xor ( n32602 , n199865 , n199878 );
buf ( n199880 , n193620 );
not ( n32604 , n199880 );
buf ( n199882 , n186197 );
not ( n32606 , n199882 );
or ( n32607 , n32604 , n32606 );
buf ( n199885 , n186208 );
buf ( n199886 , n196703 );
nand ( n32610 , n199885 , n199886 );
buf ( n199888 , n32610 );
buf ( n199889 , n199888 );
nand ( n32613 , n32607 , n199889 );
buf ( n199891 , n32613 );
buf ( n199892 , n199891 );
xor ( n32616 , n32602 , n199892 );
buf ( n199894 , n32616 );
buf ( n199895 , n199894 );
xor ( n32619 , n32575 , n199895 );
buf ( n199897 , n32619 );
buf ( n199898 , n199897 );
xor ( n32622 , n193575 , n193630 );
and ( n32623 , n32622 , n193666 );
and ( n32624 , n193575 , n193630 );
or ( n32625 , n32623 , n32624 );
buf ( n199903 , n32625 );
buf ( n199904 , n199903 );
xor ( n32628 , n199898 , n199904 );
buf ( n199906 , n845 );
buf ( n199907 , n864 );
and ( n32631 , n199906 , n199907 );
buf ( n199909 , n32631 );
buf ( n199910 , n199909 );
buf ( n199911 , n193565 );
not ( n32635 , n199911 );
buf ( n199913 , n186435 );
not ( n32637 , n199913 );
or ( n32638 , n32635 , n32637 );
buf ( n199916 , n186444 );
buf ( n199917 , n196753 );
nand ( n32641 , n199916 , n199917 );
buf ( n199919 , n32641 );
buf ( n199920 , n199919 );
nand ( n32644 , n32638 , n199920 );
buf ( n199922 , n32644 );
buf ( n199923 , n199922 );
xor ( n32647 , n199910 , n199923 );
buf ( n199925 , n193602 );
not ( n32649 , n199925 );
buf ( n199927 , n186287 );
not ( n32651 , n199927 );
or ( n32652 , n32649 , n32651 );
buf ( n199930 , n186297 );
buf ( n199931 , n196774 );
nand ( n32655 , n199930 , n199931 );
buf ( n199933 , n32655 );
buf ( n199934 , n199933 );
nand ( n32658 , n32652 , n199934 );
buf ( n199936 , n32658 );
buf ( n199937 , n199936 );
xor ( n32661 , n32647 , n199937 );
buf ( n199939 , n32661 );
buf ( n199940 , n199939 );
buf ( n199941 , n196845 );
not ( n32665 , n199941 );
buf ( n199943 , n32665 );
buf ( n199944 , n199943 );
buf ( n199945 , n193547 );
not ( n32669 , n199945 );
buf ( n199947 , n186640 );
not ( n32671 , n199947 );
or ( n32672 , n32669 , n32671 );
buf ( n199950 , n186340 );
buf ( n199951 , n196802 );
nand ( n32675 , n199950 , n199951 );
buf ( n199953 , n32675 );
buf ( n199954 , n199953 );
nand ( n32678 , n32672 , n199954 );
buf ( n199956 , n32678 );
buf ( n199957 , n199956 );
xor ( n32681 , n199944 , n199957 );
buf ( n199959 , n193657 );
buf ( n199960 , n193644 );
or ( n32684 , n199959 , n199960 );
buf ( n199962 , n193664 );
nand ( n32686 , n32684 , n199962 );
buf ( n199964 , n32686 );
buf ( n199965 , n199964 );
buf ( n199966 , n193657 );
buf ( n199967 , n193644 );
nand ( n32691 , n199966 , n199967 );
buf ( n199969 , n32691 );
buf ( n199970 , n199969 );
nand ( n32694 , n199965 , n199970 );
buf ( n199972 , n32694 );
buf ( n199973 , n199972 );
xor ( n32697 , n32681 , n199973 );
buf ( n199975 , n32697 );
buf ( n199976 , n199975 );
xor ( n32700 , n199940 , n199976 );
xor ( n32701 , n193507 , n193513 );
and ( n32702 , n32701 , n193520 );
and ( n32703 , n193507 , n193513 );
or ( n32704 , n32702 , n32703 );
buf ( n199982 , n32704 );
buf ( n199983 , n199982 );
xor ( n32707 , n32700 , n199983 );
buf ( n199985 , n32707 );
buf ( n199986 , n199985 );
xor ( n32710 , n32628 , n199986 );
buf ( n199988 , n32710 );
buf ( n199989 , n199988 );
xor ( n32713 , n199839 , n199989 );
xor ( n32714 , n193532 , n193669 );
and ( n32715 , n32714 , n193676 );
and ( n32716 , n193532 , n193669 );
or ( n32717 , n32715 , n32716 );
buf ( n199995 , n32717 );
buf ( n199996 , n199995 );
xor ( n32720 , n32713 , n199996 );
buf ( n199998 , n32720 );
not ( n32722 , n199998 );
nand ( n32723 , n32556 , n32722 );
buf ( n200001 , n196715 );
buf ( n200002 , n196718 );
xor ( n32726 , n200001 , n200002 );
buf ( n200004 , n32726 );
buf ( n200005 , n200004 );
buf ( n200006 , n196736 );
xor ( n32730 , n200005 , n200006 );
buf ( n200008 , n32730 );
buf ( n200009 , n200008 );
xor ( n32733 , n196814 , n196831 );
buf ( n200011 , n32733 );
buf ( n200012 , n196845 );
and ( n32736 , n200011 , n200012 );
not ( n32737 , n200011 );
buf ( n200015 , n199943 );
and ( n32739 , n32737 , n200015 );
nor ( n32740 , n32736 , n32739 );
buf ( n200018 , n32740 );
buf ( n200019 , n200018 );
xor ( n32743 , n200009 , n200019 );
xor ( n32744 , n199944 , n199957 );
and ( n32745 , n32744 , n199973 );
and ( n32746 , n199944 , n199957 );
or ( n32747 , n32745 , n32746 );
buf ( n200025 , n32747 );
buf ( n200026 , n200025 );
xor ( n32750 , n32743 , n200026 );
buf ( n200028 , n32750 );
buf ( n200029 , n200028 );
xor ( n32753 , n199845 , n199851 );
and ( n32754 , n32753 , n199895 );
and ( n32755 , n199845 , n199851 );
or ( n32756 , n32754 , n32755 );
buf ( n200034 , n32756 );
buf ( n200035 , n200034 );
xor ( n32759 , n199910 , n199923 );
and ( n32760 , n32759 , n199937 );
and ( n32761 , n199910 , n199923 );
or ( n32762 , n32760 , n32761 );
buf ( n200040 , n32762 );
buf ( n200041 , n200040 );
xor ( n32765 , n199865 , n199878 );
and ( n32766 , n32765 , n199892 );
and ( n32767 , n199865 , n199878 );
or ( n32768 , n32766 , n32767 );
buf ( n200046 , n32768 );
buf ( n200047 , n200046 );
xor ( n32771 , n200041 , n200047 );
xor ( n32772 , n196766 , n196769 );
xor ( n32773 , n32772 , n196787 );
buf ( n200051 , n32773 );
buf ( n200052 , n200051 );
xor ( n32776 , n32771 , n200052 );
buf ( n200054 , n32776 );
buf ( n200055 , n200054 );
xor ( n32779 , n200035 , n200055 );
xor ( n32780 , n199940 , n199976 );
and ( n32781 , n32780 , n199983 );
and ( n32782 , n199940 , n199976 );
or ( n32783 , n32781 , n32782 );
buf ( n200061 , n32783 );
buf ( n200062 , n200061 );
xor ( n32786 , n32779 , n200062 );
buf ( n200064 , n32786 );
buf ( n200065 , n200064 );
xor ( n32789 , n200029 , n200065 );
xor ( n32790 , n199898 , n199904 );
and ( n32791 , n32790 , n199986 );
and ( n32792 , n199898 , n199904 );
or ( n32793 , n32791 , n32792 );
buf ( n200071 , n32793 );
buf ( n200072 , n200071 );
xor ( n32796 , n32789 , n200072 );
buf ( n200074 , n32796 );
not ( n32798 , n200074 );
xor ( n32799 , n199839 , n199989 );
and ( n32800 , n32799 , n199996 );
and ( n32801 , n199839 , n199989 );
or ( n32802 , n32800 , n32801 );
buf ( n200080 , n32802 );
not ( n32804 , n200080 );
nand ( n32805 , n32798 , n32804 );
nand ( n32806 , n32723 , n32805 );
nor ( n32807 , n32550 , n32806 );
not ( n32808 , n32807 );
xor ( n32809 , n200009 , n200019 );
and ( n32810 , n32809 , n200026 );
and ( n32811 , n200009 , n200019 );
or ( n32812 , n32810 , n32811 );
buf ( n200090 , n32812 );
buf ( n200091 , n200090 );
xor ( n32815 , n196699 , n196748 );
xor ( n32816 , n32815 , n196792 );
buf ( n200094 , n32816 );
buf ( n200095 , n200094 );
xor ( n32819 , n200041 , n200047 );
and ( n32820 , n32819 , n200052 );
and ( n32821 , n200041 , n200047 );
or ( n32822 , n32820 , n32821 );
buf ( n200100 , n32822 );
buf ( n200101 , n200100 );
xor ( n32825 , n200095 , n200101 );
xor ( n32826 , n196857 , n196861 );
xor ( n32827 , n32826 , n196868 );
buf ( n200105 , n32827 );
buf ( n200106 , n200105 );
xor ( n32830 , n32825 , n200106 );
buf ( n200108 , n32830 );
buf ( n200109 , n200108 );
xor ( n32833 , n200091 , n200109 );
xor ( n32834 , n200035 , n200055 );
and ( n32835 , n32834 , n200062 );
and ( n32836 , n200035 , n200055 );
or ( n32837 , n32835 , n32836 );
buf ( n200115 , n32837 );
buf ( n200116 , n200115 );
and ( n32840 , n32833 , n200116 );
and ( n32841 , n200091 , n200109 );
or ( n32842 , n32840 , n32841 );
buf ( n200120 , n32842 );
xor ( n32844 , n196673 , n196677 );
xor ( n32845 , n32844 , n196682 );
buf ( n200123 , n32845 );
buf ( n200124 , n200123 );
xor ( n32848 , n196695 , n196797 );
xor ( n32849 , n32848 , n196873 );
buf ( n200127 , n32849 );
buf ( n200128 , n200127 );
xor ( n32852 , n200124 , n200128 );
xor ( n32853 , n200095 , n200101 );
and ( n32854 , n32853 , n200106 );
and ( n32855 , n200095 , n200101 );
or ( n32856 , n32854 , n32855 );
buf ( n200134 , n32856 );
buf ( n200135 , n200134 );
xor ( n32859 , n32852 , n200135 );
buf ( n200137 , n32859 );
or ( n32861 , n200120 , n200137 );
xor ( n32862 , n200091 , n200109 );
xor ( n32863 , n32862 , n200116 );
buf ( n200141 , n32863 );
xor ( n32865 , n200029 , n200065 );
and ( n32866 , n32865 , n200072 );
and ( n32867 , n200029 , n200065 );
or ( n32868 , n32866 , n32867 );
buf ( n200146 , n32868 );
or ( n32870 , n200141 , n200146 );
nand ( n32871 , n32861 , n32870 );
nor ( n32872 , n32808 , n32871 );
not ( n32873 , n32872 );
xor ( n32874 , n199614 , n199631 );
xor ( n32875 , n32874 , n199649 );
buf ( n200153 , n32875 );
buf ( n200154 , n200153 );
not ( n32878 , n200154 );
buf ( n200156 , n32878 );
buf ( n200157 , n200156 );
not ( n32881 , n200157 );
xor ( n32882 , n199552 , n199592 );
xnor ( n32883 , n32882 , n199570 );
buf ( n200161 , n32883 );
not ( n32885 , n200161 );
or ( n32886 , n32881 , n32885 );
buf ( n200164 , n192179 );
not ( n32888 , n200164 );
buf ( n200166 , n186241 );
not ( n32890 , n200166 );
or ( n32891 , n32888 , n32890 );
buf ( n200169 , n186254 );
buf ( n200170 , n199580 );
nand ( n32894 , n200169 , n200170 );
buf ( n200172 , n32894 );
buf ( n200173 , n200172 );
nand ( n32897 , n32891 , n200173 );
buf ( n200175 , n32897 );
buf ( n200176 , n200175 );
buf ( n200177 , n192364 );
not ( n32901 , n200177 );
buf ( n200179 , n19031 );
not ( n32903 , n200179 );
or ( n32904 , n32901 , n32903 );
buf ( n200182 , n186340 );
buf ( n200183 , n199540 );
nand ( n32907 , n200182 , n200183 );
buf ( n200185 , n32907 );
buf ( n200186 , n200185 );
nand ( n32910 , n32904 , n200186 );
buf ( n200188 , n32910 );
buf ( n200189 , n200188 );
xor ( n32913 , n200176 , n200189 );
buf ( n200191 , n192386 );
not ( n32915 , n200191 );
buf ( n200193 , n19177 );
not ( n32917 , n200193 );
or ( n32918 , n32915 , n32917 );
buf ( n32919 , n20279 );
buf ( n200197 , n32919 );
buf ( n200198 , n199675 );
nand ( n32922 , n200197 , n200198 );
buf ( n200200 , n32922 );
buf ( n200201 , n200200 );
nand ( n32925 , n32918 , n200201 );
buf ( n200203 , n32925 );
buf ( n200204 , n200203 );
and ( n32928 , n32913 , n200204 );
and ( n32929 , n200176 , n200189 );
or ( n32930 , n32928 , n32929 );
buf ( n200208 , n32930 );
buf ( n200209 , n200208 );
nand ( n32933 , n32886 , n200209 );
buf ( n200211 , n32933 );
buf ( n200212 , n200211 );
not ( n32936 , n32883 );
nand ( n32937 , n32936 , n200153 );
buf ( n200215 , n32937 );
nand ( n32939 , n200212 , n200215 );
buf ( n200217 , n32939 );
buf ( n200218 , n200217 );
buf ( n200219 , n192266 );
not ( n32943 , n200219 );
buf ( n200221 , n25318 );
not ( n32945 , n200221 );
or ( n32946 , n32943 , n32945 );
buf ( n200224 , n19264 );
buf ( n200225 , n199618 );
nand ( n32949 , n200224 , n200225 );
buf ( n200227 , n32949 );
buf ( n200228 , n200227 );
nand ( n32952 , n32946 , n200228 );
buf ( n200230 , n32952 );
buf ( n200231 , n200230 );
buf ( n200232 , n192407 );
not ( n32956 , n200232 );
buf ( n200234 , n186287 );
not ( n32958 , n200234 );
or ( n32959 , n32956 , n32958 );
buf ( n200237 , n186297 );
buf ( n200238 , n199636 );
nand ( n32962 , n200237 , n200238 );
buf ( n200240 , n32962 );
buf ( n200241 , n200240 );
nand ( n32965 , n32959 , n200241 );
buf ( n200243 , n32965 );
buf ( n200244 , n200243 );
xor ( n32968 , n200231 , n200244 );
buf ( n200246 , n192220 );
not ( n32970 , n200246 );
buf ( n200248 , n19613 );
not ( n32972 , n200248 );
or ( n32973 , n32970 , n32972 );
buf ( n200251 , n26571 );
buf ( n200252 , n32443 );
nand ( n32976 , n200251 , n200252 );
buf ( n200254 , n32976 );
buf ( n200255 , n200254 );
nand ( n32979 , n32973 , n200255 );
buf ( n200257 , n32979 );
buf ( n200258 , n200257 );
not ( n32982 , n200258 );
buf ( n200260 , n32982 );
buf ( n200261 , n200260 );
and ( n32985 , n32968 , n200261 );
and ( n32986 , n200231 , n200244 );
or ( n32987 , n32985 , n32986 );
buf ( n200265 , n32987 );
buf ( n200266 , n200265 );
xor ( n32990 , n199671 , n199688 );
xor ( n32991 , n32990 , n199706 );
buf ( n200269 , n32991 );
buf ( n200270 , n200269 );
xor ( n32994 , n200266 , n200270 );
xor ( n32995 , n199719 , n199733 );
xor ( n32996 , n32995 , n199751 );
buf ( n200274 , n32996 );
buf ( n200275 , n200274 );
and ( n32999 , n32994 , n200275 );
and ( n33000 , n200266 , n200270 );
or ( n33001 , n32999 , n33000 );
buf ( n200279 , n33001 );
buf ( n200280 , n200279 );
xor ( n33004 , n200218 , n200280 );
xor ( n33005 , n199776 , n199772 );
buf ( n200283 , n33005 );
buf ( n200284 , n199781 );
xor ( n33008 , n200283 , n200284 );
buf ( n200286 , n33008 );
buf ( n200287 , n200286 );
xor ( n33011 , n33004 , n200287 );
buf ( n200289 , n33011 );
buf ( n200290 , n200289 );
xor ( n33014 , n192414 , n192431 );
and ( n33015 , n33014 , n192493 );
and ( n33016 , n192414 , n192431 );
or ( n33017 , n33015 , n33016 );
buf ( n200295 , n33017 );
buf ( n200296 , n200295 );
not ( n33020 , n192185 );
not ( n33021 , n192226 );
or ( n33022 , n33020 , n33021 );
buf ( n200300 , n192226 );
buf ( n200301 , n192185 );
nor ( n33025 , n200300 , n200301 );
buf ( n200303 , n33025 );
buf ( n200304 , n192205 );
not ( n33028 , n200304 );
buf ( n200306 , n33028 );
or ( n33030 , n200303 , n200306 );
nand ( n33031 , n33022 , n33030 );
buf ( n200309 , n33031 );
buf ( n200310 , n25046 );
not ( n33034 , n200310 );
buf ( n200312 , n25030 );
not ( n33036 , n200312 );
or ( n33037 , n33034 , n33036 );
not ( n33038 , n25030 );
not ( n33039 , n33038 );
not ( n33040 , n25046 );
not ( n33041 , n33040 );
or ( n33042 , n33039 , n33041 );
nand ( n33043 , n33042 , n25066 );
buf ( n200321 , n33043 );
nand ( n33045 , n33037 , n200321 );
buf ( n200323 , n33045 );
buf ( n200324 , n200323 );
xor ( n33048 , n200309 , n200324 );
xor ( n33049 , n192350 , n192371 );
and ( n33050 , n33049 , n192393 );
and ( n33051 , n192350 , n192371 );
or ( n33052 , n33050 , n33051 );
buf ( n200330 , n33052 );
buf ( n200331 , n200330 );
xor ( n33055 , n33048 , n200331 );
buf ( n200333 , n33055 );
buf ( n200334 , n200333 );
xor ( n33058 , n200296 , n200334 );
not ( n33059 , n24954 );
nand ( n33060 , n33059 , n25067 );
nand ( n33061 , n33059 , n192297 );
nand ( n33062 , n25067 , n192297 );
nand ( n33063 , n33060 , n33061 , n33062 );
buf ( n200341 , n33063 );
and ( n33065 , n33058 , n200341 );
and ( n33066 , n200296 , n200334 );
or ( n33067 , n33065 , n33066 );
buf ( n200345 , n33067 );
buf ( n200346 , n200345 );
xor ( n33070 , n200309 , n200324 );
and ( n33071 , n33070 , n200331 );
and ( n33072 , n200309 , n200324 );
or ( n33073 , n33071 , n33072 );
buf ( n200351 , n33073 );
buf ( n200352 , n200351 );
buf ( n200353 , n200257 );
buf ( n200354 , n853 );
buf ( n200355 , n864 );
and ( n33079 , n200354 , n200355 );
buf ( n200357 , n33079 );
buf ( n200358 , n200357 );
buf ( n200359 , n192319 );
not ( n33083 , n200359 );
buf ( n200361 , n186924 );
not ( n33085 , n200361 );
or ( n33086 , n33083 , n33085 );
buf ( n200364 , n18875 );
buf ( n200365 , n199558 );
nand ( n33089 , n200364 , n200365 );
buf ( n200367 , n33089 );
buf ( n200368 , n200367 );
nand ( n33092 , n33086 , n200368 );
buf ( n200370 , n33092 );
buf ( n200371 , n200370 );
xor ( n33095 , n200358 , n200371 );
buf ( n200373 , n192339 );
not ( n33097 , n200373 );
buf ( n200375 , n192332 );
not ( n33099 , n200375 );
or ( n33100 , n33097 , n33099 );
buf ( n200378 , n192573 );
buf ( n200379 , n884 );
nand ( n33103 , n200378 , n200379 );
buf ( n200381 , n33103 );
buf ( n200382 , n200381 );
nand ( n33106 , n33100 , n200382 );
buf ( n200384 , n33106 );
buf ( n200385 , n200384 );
and ( n33109 , n33095 , n200385 );
and ( n33110 , n200358 , n200371 );
or ( n33111 , n33109 , n33110 );
buf ( n200389 , n33111 );
buf ( n200390 , n200389 );
xor ( n33114 , n200353 , n200390 );
buf ( n200392 , n192245 );
not ( n33116 , n200392 );
buf ( n200394 , n186432 );
not ( n33118 , n200394 );
or ( n33119 , n33116 , n33118 );
buf ( n200397 , n186441 );
buf ( n200398 , n199693 );
nand ( n33122 , n200397 , n200398 );
buf ( n200400 , n33122 );
buf ( n200401 , n200400 );
nand ( n33125 , n33119 , n200401 );
buf ( n200403 , n33125 );
buf ( n200404 , n200403 );
buf ( n200405 , n192288 );
not ( n33129 , n200405 );
buf ( n200407 , n186789 );
not ( n33131 , n200407 );
or ( n33132 , n33129 , n33131 );
buf ( n200410 , n186575 );
buf ( n200411 , n199738 );
nand ( n33135 , n200410 , n200411 );
buf ( n200413 , n33135 );
buf ( n200414 , n200413 );
nand ( n33138 , n33132 , n200414 );
buf ( n200416 , n33138 );
buf ( n200417 , n200416 );
xor ( n33141 , n200404 , n200417 );
buf ( n200419 , n192199 );
not ( n33143 , n200419 );
buf ( n200421 , n186197 );
not ( n33145 , n200421 );
or ( n33146 , n33143 , n33145 );
buf ( n200424 , n19494 );
buf ( n200425 , n199658 );
nand ( n33149 , n200424 , n200425 );
buf ( n200427 , n33149 );
buf ( n200428 , n200427 );
nand ( n33152 , n33146 , n200428 );
buf ( n200430 , n33152 );
buf ( n200431 , n200430 );
and ( n33155 , n33141 , n200431 );
and ( n33156 , n200404 , n200417 );
or ( n33157 , n33155 , n33156 );
buf ( n200435 , n33157 );
buf ( n200436 , n200435 );
xor ( n33160 , n33114 , n200436 );
buf ( n200438 , n33160 );
buf ( n200439 , n200438 );
xor ( n33163 , n200352 , n200439 );
xor ( n33164 , n200358 , n200371 );
xor ( n33165 , n33164 , n200385 );
buf ( n200443 , n33165 );
buf ( n200444 , n200443 );
xor ( n33168 , n192252 , n192273 );
and ( n33169 , n33168 , n192295 );
and ( n33170 , n192252 , n192273 );
or ( n33171 , n33169 , n33170 );
buf ( n200449 , n33171 );
buf ( n200450 , n200449 );
xor ( n33174 , n200444 , n200450 );
xor ( n33175 , n200404 , n200417 );
xor ( n33176 , n33175 , n200431 );
buf ( n200454 , n33176 );
buf ( n200455 , n200454 );
and ( n33179 , n33174 , n200455 );
and ( n33180 , n200444 , n200450 );
or ( n33181 , n33179 , n33180 );
buf ( n200459 , n33181 );
buf ( n200460 , n200459 );
xor ( n33184 , n33163 , n200460 );
buf ( n200462 , n33184 );
buf ( n200463 , n200462 );
xor ( n33187 , n200346 , n200463 );
xor ( n33188 , n200444 , n200450 );
xor ( n33189 , n33188 , n200455 );
buf ( n200467 , n33189 );
buf ( n200468 , n200467 );
xor ( n33192 , n200176 , n200189 );
xor ( n33193 , n33192 , n200204 );
buf ( n200471 , n33193 );
buf ( n200472 , n200471 );
xor ( n33196 , n200231 , n200244 );
xor ( n33197 , n33196 , n200261 );
buf ( n200475 , n33197 );
buf ( n200476 , n200475 );
xor ( n33200 , n200472 , n200476 );
xor ( n33201 , n193394 , n193400 );
and ( n33202 , n33201 , n193442 );
and ( n33203 , n193394 , n193400 );
or ( n33204 , n33202 , n33203 );
buf ( n200482 , n33204 );
buf ( n200483 , n200482 );
xor ( n33207 , n33200 , n200483 );
buf ( n200485 , n33207 );
buf ( n200486 , n200485 );
xor ( n33210 , n200468 , n200486 );
xor ( n33211 , n192396 , n192496 );
and ( n33212 , n33211 , n192660 );
and ( n33213 , n192396 , n192496 );
or ( n33214 , n33212 , n33213 );
buf ( n200492 , n33214 );
buf ( n200493 , n200492 );
and ( n33217 , n33210 , n200493 );
and ( n33218 , n200468 , n200486 );
or ( n33219 , n33217 , n33218 );
buf ( n200497 , n33219 );
buf ( n200498 , n200497 );
and ( n33222 , n33187 , n200498 );
and ( n33223 , n200346 , n200463 );
or ( n33224 , n33222 , n33223 );
buf ( n200502 , n33224 );
buf ( n200503 , n200502 );
xor ( n33227 , n200290 , n200503 );
xor ( n33228 , n200352 , n200439 );
and ( n33229 , n33228 , n200460 );
and ( n33230 , n200352 , n200439 );
or ( n33231 , n33229 , n33230 );
buf ( n200509 , n33231 );
buf ( n200510 , n200509 );
xor ( n33234 , n199518 , n199535 );
xor ( n33235 , n33234 , n199599 );
buf ( n200513 , n33235 );
buf ( n200514 , n200513 );
xor ( n33238 , n200353 , n200390 );
and ( n33239 , n33238 , n200436 );
and ( n33240 , n200353 , n200390 );
or ( n33241 , n33239 , n33240 );
buf ( n200519 , n33241 );
buf ( n200520 , n200519 );
xor ( n33244 , n200514 , n200520 );
xor ( n33245 , n199654 , n199711 );
xor ( n33246 , n33245 , n199756 );
buf ( n200524 , n33246 );
buf ( n200525 , n200524 );
xor ( n33249 , n33244 , n200525 );
buf ( n200527 , n33249 );
buf ( n200528 , n200527 );
xor ( n33252 , n200510 , n200528 );
xor ( n33253 , n200266 , n200270 );
xor ( n33254 , n33253 , n200275 );
buf ( n200532 , n33254 );
buf ( n200533 , n200532 );
not ( n33257 , n200533 );
buf ( n200535 , n33257 );
buf ( n200536 , n200535 );
not ( n33260 , n200536 );
xor ( n33261 , n200153 , n200208 );
xor ( n33262 , n33261 , n32883 );
buf ( n200540 , n33262 );
not ( n33264 , n200540 );
or ( n33265 , n33260 , n33264 );
xor ( n33266 , n200472 , n200476 );
and ( n33267 , n33266 , n200483 );
and ( n33268 , n200472 , n200476 );
or ( n33269 , n33267 , n33268 );
buf ( n200547 , n33269 );
buf ( n200548 , n200547 );
nand ( n33272 , n33265 , n200548 );
buf ( n200550 , n33272 );
buf ( n200551 , n200550 );
buf ( n200552 , n200532 );
buf ( n200553 , n33262 );
not ( n33277 , n200553 );
buf ( n200555 , n33277 );
buf ( n200556 , n200555 );
nand ( n33280 , n200552 , n200556 );
buf ( n200558 , n33280 );
buf ( n200559 , n200558 );
nand ( n33283 , n200551 , n200559 );
buf ( n200561 , n33283 );
buf ( n200562 , n200561 );
xor ( n33286 , n33252 , n200562 );
buf ( n200564 , n33286 );
buf ( n200565 , n200564 );
xor ( n33289 , n33227 , n200565 );
buf ( n200567 , n33289 );
not ( n33291 , n200567 );
buf ( n200569 , n200555 );
not ( n33293 , n200569 );
buf ( n200571 , n200535 );
not ( n33295 , n200571 );
or ( n33296 , n33293 , n33295 );
buf ( n200574 , n200532 );
buf ( n200575 , n33262 );
nand ( n33299 , n200574 , n200575 );
buf ( n200577 , n33299 );
buf ( n200578 , n200577 );
nand ( n33302 , n33296 , n200578 );
buf ( n200580 , n33302 );
buf ( n200581 , n200580 );
buf ( n200582 , n200547 );
and ( n33306 , n200581 , n200582 );
not ( n33307 , n200581 );
buf ( n200585 , n200547 );
not ( n33309 , n200585 );
buf ( n200587 , n33309 );
buf ( n200588 , n200587 );
and ( n33312 , n33307 , n200588 );
nor ( n33313 , n33306 , n33312 );
buf ( n200591 , n33313 );
buf ( n200592 , n200591 );
xor ( n33316 , n200296 , n200334 );
xor ( n33317 , n33316 , n200341 );
buf ( n200595 , n33317 );
buf ( n200596 , n200595 );
xor ( n33320 , n193342 , n193445 );
and ( n33321 , n33320 , n193467 );
and ( n33322 , n193342 , n193445 );
or ( n33323 , n33321 , n33322 );
buf ( n200601 , n33323 );
buf ( n200602 , n200601 );
xor ( n33326 , n200596 , n200602 );
nand ( n33327 , n25068 , n192662 );
nand ( n33328 , n25068 , n192895 );
nand ( n33329 , n192662 , n192895 );
nand ( n33330 , n33327 , n33328 , n33329 );
buf ( n200608 , n33330 );
and ( n33332 , n33326 , n200608 );
and ( n33333 , n200596 , n200602 );
or ( n33334 , n33332 , n33333 );
buf ( n200612 , n33334 );
buf ( n200613 , n200612 );
xor ( n33337 , n200592 , n200613 );
xor ( n33338 , n200346 , n200463 );
xor ( n33339 , n33338 , n200498 );
buf ( n200617 , n33339 );
buf ( n200618 , n200617 );
and ( n33342 , n33337 , n200618 );
and ( n33343 , n200592 , n200613 );
or ( n33344 , n33342 , n33343 );
buf ( n200622 , n33344 );
not ( n33346 , n200622 );
nand ( n33347 , n33291 , n33346 );
xor ( n33348 , n200218 , n200280 );
and ( n33349 , n33348 , n200287 );
and ( n33350 , n200218 , n200280 );
or ( n33351 , n33349 , n33350 );
buf ( n200629 , n33351 );
buf ( n200630 , n200629 );
xor ( n33354 , n200510 , n200528 );
and ( n33355 , n33354 , n200562 );
and ( n33356 , n200510 , n200528 );
or ( n33357 , n33355 , n33356 );
buf ( n200635 , n33357 );
buf ( n200636 , n200635 );
xor ( n33360 , n200630 , n200636 );
xor ( n33361 , n199604 , n199608 );
xor ( n33362 , n33361 , n199761 );
buf ( n200640 , n33362 );
buf ( n200641 , n200640 );
xor ( n33365 , n200514 , n200520 );
and ( n33366 , n33365 , n200525 );
and ( n33367 , n200514 , n200520 );
or ( n33368 , n33366 , n33367 );
buf ( n200646 , n33368 );
buf ( n200647 , n200646 );
xor ( n33371 , n200641 , n200647 );
xor ( n33372 , n199793 , n199797 );
xor ( n33373 , n33372 , n199801 );
buf ( n200651 , n33373 );
buf ( n200652 , n200651 );
xor ( n33376 , n33371 , n200652 );
buf ( n200654 , n33376 );
buf ( n200655 , n200654 );
xor ( n33379 , n33360 , n200655 );
buf ( n200657 , n33379 );
not ( n33381 , n200657 );
xor ( n33382 , n200290 , n200503 );
and ( n33383 , n33382 , n200565 );
and ( n33384 , n200290 , n200503 );
or ( n33385 , n33383 , n33384 );
buf ( n200663 , n33385 );
not ( n33387 , n200663 );
nand ( n33388 , n33381 , n33387 );
nand ( n33389 , n33347 , n33388 );
xor ( n33390 , n200630 , n200636 );
and ( n33391 , n33390 , n200655 );
and ( n33392 , n200630 , n200636 );
or ( n33393 , n33391 , n33392 );
buf ( n200671 , n33393 );
not ( n33395 , n200671 );
buf ( n200673 , n187383 );
not ( n33397 , n200673 );
buf ( n200675 , n20077 );
not ( n33399 , n200675 );
or ( n33400 , n33397 , n33399 );
buf ( n200678 , n20077 );
buf ( n200679 , n187383 );
or ( n33403 , n200678 , n200679 );
nand ( n33404 , n33400 , n33403 );
buf ( n200682 , n33404 );
xor ( n33406 , n20086 , n200682 );
xor ( n33407 , n199765 , n199768 );
xor ( n33408 , n33407 , n199805 );
xor ( n33409 , n33406 , n33408 );
xor ( n33410 , n200641 , n200647 );
and ( n33411 , n33410 , n200652 );
and ( n33412 , n200641 , n200647 );
or ( n33413 , n33411 , n33412 );
buf ( n200691 , n33413 );
xor ( n33415 , n33409 , n200691 );
not ( n33416 , n33415 );
nand ( n33417 , n33395 , n33416 );
xor ( n33418 , n199517 , n32531 );
xor ( n33419 , n33418 , n199812 );
not ( n33420 , n33419 );
xor ( n33421 , n33406 , n33408 );
and ( n33422 , n33421 , n200691 );
and ( n33423 , n33406 , n33408 );
or ( n33424 , n33422 , n33423 );
not ( n33425 , n33424 );
nand ( n33426 , n33420 , n33425 );
nand ( n33427 , n33417 , n33426 );
nor ( n33428 , n33389 , n33427 );
not ( n33429 , n33428 );
xor ( n33430 , n200592 , n200613 );
xor ( n33431 , n33430 , n200618 );
buf ( n200709 , n33431 );
not ( n33433 , n200709 );
xor ( n33434 , n200468 , n200486 );
xor ( n33435 , n33434 , n200493 );
buf ( n200713 , n33435 );
buf ( n200714 , n200713 );
xor ( n33438 , n193336 , n193470 );
and ( n33439 , n33438 , n193487 );
and ( n33440 , n193336 , n193470 );
or ( n33441 , n33439 , n33440 );
buf ( n200719 , n33441 );
buf ( n200720 , n200719 );
xor ( n33444 , n200714 , n200720 );
xor ( n33445 , n200596 , n200602 );
xor ( n33446 , n33445 , n200608 );
buf ( n200724 , n33446 );
buf ( n200725 , n200724 );
and ( n33449 , n33444 , n200725 );
and ( n33450 , n200714 , n200720 );
or ( n33451 , n33449 , n33450 );
buf ( n200729 , n33451 );
not ( n33453 , n200729 );
nand ( n33454 , n33433 , n33453 );
not ( n33455 , n193694 );
xor ( n33456 , n200714 , n200720 );
xor ( n33457 , n33456 , n200725 );
buf ( n200735 , n33457 );
not ( n33459 , n200735 );
nand ( n33460 , n33455 , n33459 );
nand ( n33461 , n33454 , n33460 );
not ( n33462 , n33461 );
not ( n33463 , n33462 );
xor ( n33464 , n193474 , n193477 );
xor ( n33465 , n33464 , n193483 );
buf ( n200743 , n33465 );
xor ( n33467 , n193147 , n193186 );
xor ( n33468 , n33467 , n193324 );
buf ( n200746 , n33468 );
buf ( n200747 , n200746 );
xor ( n33471 , n200743 , n200747 );
xor ( n33472 , n191146 , n23903 );
and ( n33473 , n33472 , n191241 );
and ( n33474 , n191146 , n23903 );
or ( n33475 , n33473 , n33474 );
buf ( n200753 , n33475 );
xor ( n33477 , n193157 , n193161 );
xor ( n33478 , n33477 , n193171 );
buf ( n200756 , n33478 );
buf ( n200757 , n200756 );
xor ( n33481 , n200753 , n200757 );
xor ( n33482 , n191250 , n191301 );
and ( n33483 , n33482 , n191308 );
and ( n33484 , n191250 , n191301 );
or ( n33485 , n33483 , n33484 );
buf ( n200763 , n33485 );
buf ( n200764 , n200763 );
and ( n33488 , n33481 , n200764 );
and ( n33489 , n200753 , n200757 );
or ( n33490 , n33488 , n33489 );
buf ( n200768 , n33490 );
buf ( n200769 , n200768 );
xor ( n33493 , n193151 , n193176 );
xor ( n33494 , n33493 , n193181 );
buf ( n200772 , n33494 );
buf ( n200773 , n200772 );
xor ( n33497 , n200769 , n200773 );
xor ( n33498 , n193248 , n193298 );
xor ( n33499 , n33498 , n193319 );
buf ( n200777 , n33499 );
buf ( n200778 , n200777 );
and ( n33502 , n33497 , n200778 );
and ( n33503 , n200769 , n200773 );
or ( n33504 , n33502 , n33503 );
buf ( n200782 , n33504 );
buf ( n200783 , n200782 );
xor ( n33507 , n33471 , n200783 );
buf ( n200785 , n33507 );
not ( n33509 , n200785 );
xor ( n33510 , n193203 , n193206 );
xor ( n33511 , n33510 , n193243 );
buf ( n200789 , n33511 );
buf ( n200790 , n200789 );
xor ( n33514 , n23515 , n190854 );
and ( n33515 , n33514 , n23715 );
and ( n33516 , n23515 , n190854 );
or ( n33517 , n33515 , n33516 );
buf ( n200795 , n33517 );
xor ( n33519 , n200790 , n200795 );
xor ( n33520 , n193254 , n193263 );
xor ( n33521 , n33520 , n193293 );
buf ( n200799 , n33521 );
buf ( n200800 , n200799 );
and ( n33524 , n33519 , n200800 );
and ( n33525 , n200790 , n200795 );
or ( n33526 , n33524 , n33525 );
buf ( n200804 , n33526 );
buf ( n200805 , n200804 );
xor ( n33529 , n191104 , n191243 );
and ( n33530 , n33529 , n191311 );
and ( n33531 , n191104 , n191243 );
or ( n33532 , n33530 , n33531 );
buf ( n200810 , n33532 );
buf ( n200811 , n200810 );
xor ( n33535 , n200753 , n200757 );
xor ( n33536 , n33535 , n200764 );
buf ( n200814 , n33536 );
buf ( n200815 , n200814 );
xor ( n33539 , n200811 , n200815 );
xor ( n33540 , n200790 , n200795 );
xor ( n33541 , n33540 , n200800 );
buf ( n200819 , n33541 );
buf ( n200820 , n200819 );
and ( n33544 , n33539 , n200820 );
and ( n33545 , n200811 , n200815 );
or ( n33546 , n33544 , n33545 );
buf ( n200824 , n33546 );
buf ( n200825 , n200824 );
xor ( n33549 , n200805 , n200825 );
xor ( n33550 , n200769 , n200773 );
xor ( n33551 , n33550 , n200778 );
buf ( n200829 , n33551 );
buf ( n200830 , n200829 );
and ( n33554 , n33549 , n200830 );
and ( n33555 , n200805 , n200825 );
or ( n33556 , n33554 , n33555 );
buf ( n200834 , n33556 );
not ( n33558 , n200834 );
nor ( n33559 , n33509 , n33558 );
not ( n33560 , n33559 );
not ( n33561 , n193492 );
xor ( n33562 , n200743 , n200747 );
and ( n33563 , n33562 , n200783 );
and ( n33564 , n200743 , n200747 );
or ( n33565 , n33563 , n33564 );
buf ( n200843 , n33565 );
not ( n33567 , n200843 );
nand ( n33568 , n33561 , n33567 );
not ( n33569 , n33568 );
or ( n33570 , n33560 , n33569 );
not ( n33571 , n33567 );
not ( n33572 , n33561 );
nand ( n33573 , n33571 , n33572 );
nand ( n33574 , n33570 , n33573 );
not ( n33575 , n33574 );
or ( n33576 , n33463 , n33575 );
nor ( n33577 , n200709 , n200729 );
not ( n33578 , n33577 );
nand ( n33579 , n193694 , n200735 );
not ( n33580 , n33579 );
and ( n33581 , n33578 , n33580 );
nand ( n33582 , n200709 , n200729 );
not ( n33583 , n33582 );
nor ( n33584 , n33581 , n33583 );
nand ( n33585 , n33576 , n33584 );
not ( n33586 , n33585 );
or ( n33587 , n33429 , n33586 );
not ( n33588 , n33427 );
not ( n33589 , n33388 );
not ( n33590 , n33346 );
buf ( n33591 , n200567 );
nand ( n33592 , n33590 , n33591 );
or ( n33593 , n33589 , n33592 );
not ( n33594 , n33387 );
nand ( n33595 , n33594 , n200657 );
nand ( n33596 , n33593 , n33595 );
and ( n33597 , n33588 , n33596 );
not ( n33598 , n33426 );
nand ( n33599 , n200671 , n33415 );
or ( n33600 , n33598 , n33599 );
or ( n33601 , n33420 , n33425 );
nand ( n33602 , n33600 , n33601 );
nor ( n33603 , n33597 , n33602 );
nand ( n33604 , n33587 , n33603 );
not ( n33605 , n33604 );
xor ( n33606 , n191318 , n191327 );
xor ( n33607 , n33606 , n191332 );
buf ( n200885 , n33607 );
buf ( n200886 , n200885 );
xor ( n33610 , n189439 , n189778 );
and ( n33611 , n33610 , n189821 );
and ( n33612 , n189439 , n189778 );
or ( n33613 , n33611 , n33612 );
buf ( n200891 , n33613 );
buf ( n200892 , n200891 );
xor ( n33616 , n200886 , n200892 );
not ( n33617 , n191349 );
not ( n33618 , n24077 );
or ( n33619 , n33617 , n33618 );
nand ( n33620 , n24075 , n191343 );
nand ( n33621 , n33619 , n33620 );
and ( n33622 , n33621 , n191378 );
not ( n33623 , n33621 );
not ( n33624 , n191378 );
and ( n33625 , n33623 , n33624 );
nor ( n33626 , n33622 , n33625 );
buf ( n200904 , n33626 );
and ( n33628 , n33616 , n200904 );
and ( n33629 , n200886 , n200892 );
or ( n33630 , n33628 , n33629 );
buf ( n200908 , n33630 );
not ( n33632 , n200908 );
not ( n33633 , n33632 );
not ( n33634 , n33633 );
xor ( n33635 , n23775 , n24103 );
xor ( n33636 , n33635 , n24060 );
buf ( n33637 , n33636 );
not ( n33638 , n33637 );
or ( n33639 , n33634 , n33638 );
not ( n33640 , n33636 );
not ( n33641 , n33640 );
not ( n33642 , n33632 );
or ( n33643 , n33641 , n33642 );
xor ( n33644 , n200886 , n200892 );
xor ( n33645 , n33644 , n200904 );
buf ( n200923 , n33645 );
and ( n33647 , n200923 , n189835 );
nand ( n33648 , n33643 , n33647 );
nand ( n33649 , n33639 , n33648 );
buf ( n33650 , n189411 );
buf ( n200928 , n33650 );
not ( n33652 , n200928 );
not ( n33653 , n22129 );
not ( n33654 , n21948 );
or ( n33655 , n33653 , n33654 );
or ( n33656 , n22129 , n21948 );
nand ( n33657 , n33655 , n33656 );
buf ( n200935 , n33657 );
not ( n33659 , n200935 );
or ( n33660 , n33652 , n33659 );
buf ( n200938 , n33650 );
buf ( n200939 , n33657 );
or ( n33663 , n200938 , n200939 );
nand ( n33664 , n33660 , n33663 );
buf ( n200942 , n33664 );
buf ( n200943 , n200942 );
xor ( n33667 , n192150 , n192154 );
and ( n33668 , n33667 , n192159 );
and ( n33669 , n192150 , n192154 );
or ( n33670 , n33668 , n33669 );
buf ( n200948 , n33670 );
buf ( n200949 , n200948 );
xor ( n33673 , n200943 , n200949 );
xor ( n33674 , n190055 , n190058 );
xor ( n33675 , n33674 , n190317 );
buf ( n200953 , n33675 );
buf ( n200954 , n200953 );
xor ( n33678 , n33673 , n200954 );
buf ( n200956 , n33678 );
not ( n33680 , n200956 );
not ( n33681 , n194823 );
nand ( n33682 , n33680 , n33681 );
xor ( n33683 , n191401 , n191618 );
xor ( n33684 , n33683 , n191754 );
buf ( n200962 , n33684 );
buf ( n200963 , n200962 );
xor ( n33687 , n191632 , n191745 );
xor ( n33688 , n33687 , n191749 );
buf ( n200966 , n33688 );
buf ( n200967 , n200966 );
xor ( n33691 , n191405 , n191577 );
xor ( n33692 , n33691 , n191613 );
buf ( n200970 , n33692 );
buf ( n200971 , n200970 );
xor ( n33695 , n200967 , n200971 );
xor ( n33696 , n24313 , n191600 );
xor ( n33697 , n33696 , n191609 );
buf ( n200975 , n33697 );
not ( n33699 , n24455 );
not ( n33700 , n33699 );
not ( n33701 , n191704 );
not ( n33702 , n20727 );
or ( n33703 , n33701 , n33702 );
nand ( n33704 , n33703 , n191713 );
xor ( n33705 , n33704 , n191698 );
not ( n33706 , n33705 );
or ( n33707 , n33700 , n33706 );
or ( n33708 , n33699 , n33705 );
nand ( n33709 , n33707 , n33708 );
buf ( n200987 , n849 );
buf ( n200988 , n882 );
xor ( n33712 , n200987 , n200988 );
buf ( n200990 , n33712 );
buf ( n200991 , n200990 );
not ( n33715 , n200991 );
buf ( n200993 , n19613 );
not ( n33717 , n200993 );
or ( n33718 , n33715 , n33717 );
buf ( n200996 , n26571 );
buf ( n200997 , n191636 );
nand ( n33721 , n200996 , n200997 );
buf ( n200999 , n33721 );
buf ( n201000 , n200999 );
nand ( n33724 , n33718 , n201000 );
buf ( n201002 , n33724 );
not ( n33726 , n201002 );
not ( n33727 , n24521 );
not ( n33728 , n24509 );
or ( n33729 , n33727 , n33728 );
or ( n33730 , n24509 , n24521 );
nand ( n33731 , n33729 , n33730 );
not ( n33732 , n33731 );
not ( n33733 , n33732 );
or ( n33734 , n33726 , n33733 );
buf ( n201012 , n201002 );
not ( n33736 , n201012 );
buf ( n201014 , n33736 );
buf ( n201015 , n201014 );
not ( n33739 , n201015 );
buf ( n201017 , n33731 );
not ( n33741 , n201017 );
or ( n33742 , n33739 , n33741 );
buf ( n201020 , n18907 );
buf ( n201021 , n863 );
and ( n33745 , n201020 , n201021 );
buf ( n201023 , n33745 );
buf ( n201024 , n201023 );
xor ( n33748 , n888 , n844 );
buf ( n201026 , n33748 );
not ( n33750 , n201026 );
buf ( n201028 , n190454 );
not ( n33752 , n201028 );
or ( n33753 , n33750 , n33752 );
buf ( n201031 , n20396 );
buf ( n201032 , n191819 );
nand ( n33756 , n201031 , n201032 );
buf ( n201034 , n33756 );
buf ( n201035 , n201034 );
nand ( n33759 , n33753 , n201035 );
buf ( n201037 , n33759 );
buf ( n201038 , n201037 );
xor ( n33762 , n201024 , n201038 );
xor ( n33763 , n892 , n840 );
buf ( n201041 , n33763 );
not ( n33765 , n201041 );
buf ( n201043 , n190485 );
not ( n33767 , n201043 );
or ( n33768 , n33765 , n33767 );
buf ( n201046 , n190128 );
buf ( n201047 , n191778 );
nand ( n33771 , n201046 , n201047 );
buf ( n201049 , n33771 );
buf ( n201050 , n201049 );
nand ( n33774 , n33768 , n201050 );
buf ( n201052 , n33774 );
buf ( n201053 , n201052 );
and ( n33777 , n33762 , n201053 );
and ( n33778 , n201024 , n201038 );
or ( n33779 , n33777 , n33778 );
buf ( n201057 , n33779 );
buf ( n201058 , n201057 );
nand ( n33782 , n33742 , n201058 );
buf ( n201060 , n33782 );
nand ( n33784 , n33734 , n201060 );
xor ( n33785 , n33709 , n33784 );
buf ( n201063 , n852 );
buf ( n201064 , n880 );
xor ( n33788 , n201063 , n201064 );
buf ( n201066 , n33788 );
buf ( n201067 , n201066 );
not ( n33791 , n201067 );
buf ( n201069 , n18862 );
not ( n33793 , n201069 );
or ( n33794 , n33791 , n33793 );
buf ( n201072 , n18875 );
buf ( n201073 , n191809 );
nand ( n33797 , n201072 , n201073 );
buf ( n201075 , n33797 );
buf ( n201076 , n201075 );
nand ( n33800 , n33794 , n201076 );
buf ( n201078 , n33800 );
buf ( n201079 , n846 );
buf ( n201080 , n886 );
xor ( n33804 , n201079 , n201080 );
buf ( n201082 , n33804 );
buf ( n201083 , n201082 );
not ( n33807 , n201083 );
buf ( n201085 , n20554 );
not ( n33809 , n201085 );
or ( n33810 , n33807 , n33809 );
buf ( n201088 , n20558 );
buf ( n201089 , n191863 );
nand ( n33813 , n201088 , n201089 );
buf ( n201091 , n33813 );
buf ( n201092 , n201091 );
nand ( n33816 , n33810 , n201092 );
buf ( n201094 , n33816 );
or ( n33818 , n201078 , n201094 );
buf ( n201096 , n854 );
buf ( n201097 , n878 );
xor ( n33821 , n201096 , n201097 );
buf ( n201099 , n33821 );
buf ( n201100 , n201099 );
not ( n33824 , n201100 );
buf ( n201102 , n186569 );
not ( n33826 , n201102 );
or ( n33827 , n33824 , n33826 );
buf ( n201105 , n186575 );
buf ( n201106 , n191840 );
nand ( n33830 , n201105 , n201106 );
buf ( n201108 , n33830 );
buf ( n201109 , n201108 );
nand ( n33833 , n33827 , n201109 );
buf ( n201111 , n33833 );
nand ( n33835 , n33818 , n201111 );
buf ( n201113 , n201094 );
buf ( n201114 , n201078 );
nand ( n33838 , n201113 , n201114 );
buf ( n201116 , n33838 );
nand ( n33840 , n33835 , n201116 );
not ( n33841 , n33840 );
xor ( n33842 , n872 , n860 );
buf ( n201120 , n33842 );
not ( n33844 , n201120 );
buf ( n201122 , n20244 );
not ( n33846 , n201122 );
or ( n33847 , n33844 , n33846 );
buf ( n201125 , n19264 );
buf ( n201126 , n24753 );
nand ( n33850 , n201125 , n201126 );
buf ( n201128 , n33850 );
buf ( n201129 , n201128 );
nand ( n33853 , n33847 , n201129 );
buf ( n201131 , n33853 );
buf ( n201132 , n201131 );
buf ( n201133 , n848 );
buf ( n201134 , n884 );
xor ( n33858 , n201133 , n201134 );
buf ( n201136 , n33858 );
buf ( n201137 , n201136 );
not ( n33861 , n201137 );
buf ( n201139 , n20727 );
not ( n33863 , n201139 );
or ( n33864 , n33861 , n33863 );
buf ( n201142 , n190543 );
buf ( n201143 , n192015 );
nand ( n33867 , n201142 , n201143 );
buf ( n201145 , n33867 );
buf ( n201146 , n201145 );
nand ( n33870 , n33864 , n201146 );
buf ( n201148 , n33870 );
buf ( n201149 , n201148 );
xor ( n33873 , n201132 , n201149 );
buf ( n201151 , n862 );
buf ( n201152 , n870 );
xor ( n33876 , n201151 , n201152 );
buf ( n201154 , n33876 );
buf ( n201155 , n201154 );
not ( n33879 , n201155 );
buf ( n201157 , n186432 );
not ( n33881 , n201157 );
or ( n33882 , n33879 , n33881 );
buf ( n201160 , n186444 );
buf ( n201161 , n192092 );
nand ( n33885 , n201160 , n201161 );
buf ( n201163 , n33885 );
buf ( n201164 , n201163 );
nand ( n33888 , n33882 , n201164 );
buf ( n201166 , n33888 );
buf ( n201167 , n201166 );
and ( n33891 , n33873 , n201167 );
and ( n33892 , n201132 , n201149 );
or ( n33893 , n33891 , n33892 );
buf ( n201171 , n33893 );
not ( n33895 , n201171 );
or ( n33896 , n33841 , n33895 );
nor ( n33897 , n33840 , n201171 );
buf ( n201175 , n838 );
buf ( n201176 , n894 );
xor ( n33900 , n201175 , n201176 );
buf ( n201178 , n33900 );
buf ( n201179 , n201178 );
not ( n33903 , n201179 );
buf ( n201181 , n21330 );
not ( n33905 , n201181 );
or ( n33906 , n33903 , n33905 );
buf ( n201184 , n191998 );
buf ( n201185 , n895 );
nand ( n33909 , n201184 , n201185 );
buf ( n201187 , n33909 );
buf ( n201188 , n201187 );
nand ( n33912 , n33906 , n201188 );
buf ( n201190 , n33912 );
buf ( n201191 , n201190 );
xor ( n33915 , n858 , n874 );
not ( n33916 , n33915 );
not ( n33917 , n18992 );
or ( n33918 , n33916 , n33917 );
nand ( n33919 , n191903 , n188823 );
nand ( n33920 , n33918 , n33919 );
buf ( n201198 , n33920 );
xor ( n33922 , n201191 , n201198 );
buf ( n201200 , n856 );
buf ( n201201 , n876 );
xor ( n33925 , n201200 , n201201 );
buf ( n201203 , n33925 );
not ( n33927 , n201203 );
not ( n33928 , n19177 );
or ( n33929 , n33927 , n33928 );
nand ( n33930 , n191880 , n19103 );
nand ( n33931 , n33929 , n33930 );
buf ( n201209 , n33931 );
and ( n33933 , n33922 , n201209 );
and ( n33934 , n201191 , n201198 );
or ( n33935 , n33933 , n33934 );
buf ( n201213 , n33935 );
buf ( n201214 , n201213 );
not ( n33938 , n201214 );
buf ( n201216 , n33938 );
or ( n33940 , n33897 , n201216 );
nand ( n33941 , n33896 , n33940 );
and ( n33942 , n33785 , n33941 );
and ( n33943 , n33709 , n33784 );
or ( n33944 , n33942 , n33943 );
buf ( n201222 , n33944 );
xor ( n33946 , n200975 , n201222 );
xor ( n33947 , n191801 , n24581 );
xor ( n33948 , n33947 , n24635 );
not ( n33949 , n33948 );
xor ( n33950 , n192048 , n192111 );
xor ( n33951 , n33950 , n192116 );
buf ( n201229 , n33951 );
not ( n33953 , n201229 );
or ( n33954 , n33949 , n33953 );
or ( n33955 , n201229 , n33948 );
buf ( n201233 , n191834 );
not ( n33957 , n201233 );
buf ( n201235 , n24534 );
not ( n33959 , n201235 );
or ( n33960 , n33957 , n33959 );
buf ( n201238 , n191814 );
buf ( n201239 , n191831 );
nand ( n33963 , n201238 , n201239 );
buf ( n201241 , n33963 );
buf ( n201242 , n201241 );
nand ( n33966 , n33960 , n201242 );
buf ( n201244 , n33966 );
not ( n33968 , n191852 );
and ( n33969 , n201244 , n33968 );
not ( n33970 , n201244 );
and ( n33971 , n33970 , n191852 );
nor ( n33972 , n33969 , n33971 );
not ( n33973 , n33972 );
not ( n33974 , n33973 );
xor ( n33975 , n192011 , n192028 );
xor ( n33976 , n33975 , n192043 );
buf ( n201254 , n33976 );
not ( n33978 , n201254 );
or ( n33979 , n33974 , n33978 );
not ( n33980 , n33972 );
buf ( n201258 , n201254 );
not ( n33982 , n201258 );
buf ( n201260 , n33982 );
not ( n33984 , n201260 );
or ( n33985 , n33980 , n33984 );
xor ( n33986 , n192082 , n192064 );
xor ( n33987 , n33986 , n192104 );
nand ( n33988 , n33985 , n33987 );
nand ( n33989 , n33979 , n33988 );
nand ( n33990 , n33955 , n33989 );
nand ( n33991 , n33954 , n33990 );
buf ( n201269 , n33991 );
and ( n33993 , n33946 , n201269 );
and ( n33994 , n200975 , n201222 );
or ( n33995 , n33993 , n33994 );
buf ( n201273 , n33995 );
buf ( n201274 , n201273 );
and ( n33998 , n33695 , n201274 );
and ( n33999 , n200967 , n200971 );
or ( n34000 , n33998 , n33999 );
buf ( n201278 , n34000 );
buf ( n201279 , n201278 );
xor ( n34003 , n200963 , n201279 );
xor ( n34004 , n191763 , n191767 );
xor ( n34005 , n34004 , n192141 );
buf ( n201283 , n34005 );
buf ( n201284 , n201283 );
and ( n34008 , n34003 , n201284 );
and ( n34009 , n200963 , n201279 );
or ( n34010 , n34008 , n34009 );
buf ( n201288 , n34010 );
and ( n34012 , n192164 , n201288 );
nand ( n34013 , n33682 , n34012 );
xor ( n34014 , n200943 , n200949 );
and ( n34015 , n34014 , n200954 );
and ( n34016 , n200943 , n200949 );
or ( n34017 , n34015 , n34016 );
buf ( n201295 , n34017 );
nand ( n34019 , n190324 , n201295 );
nand ( n34020 , n194823 , n200956 );
nand ( n34021 , n34019 , n34020 );
not ( n34022 , n34021 );
buf ( n201300 , n188497 );
buf ( n201301 , n189427 );
xor ( n34025 , n201300 , n201301 );
buf ( n201303 , n189823 );
xor ( n34027 , n34025 , n201303 );
buf ( n201305 , n34027 );
xor ( n34029 , n189854 , n189858 );
and ( n34030 , n34029 , n190322 );
and ( n34031 , n189854 , n189858 );
or ( n34032 , n34030 , n34031 );
buf ( n201310 , n34032 );
nand ( n34034 , n201305 , n201310 );
nand ( n34035 , n34013 , n34022 , n34034 );
nor ( n34036 , n33649 , n34035 );
xor ( n34037 , n190711 , n23716 );
and ( n34038 , n34037 , n191051 );
and ( n34039 , n190711 , n23716 );
or ( n34040 , n34038 , n34039 );
buf ( n201318 , n34040 );
xor ( n34042 , n191098 , n191313 );
and ( n34043 , n34042 , n191336 );
and ( n34044 , n191098 , n191313 );
or ( n34045 , n34043 , n34044 );
buf ( n201323 , n34045 );
xor ( n34047 , n201318 , n201323 );
xor ( n34048 , n200811 , n200815 );
xor ( n34049 , n34048 , n200820 );
buf ( n201327 , n34049 );
buf ( n201328 , n201327 );
and ( n34052 , n34047 , n201328 );
and ( n34053 , n201318 , n201323 );
or ( n34054 , n34052 , n34053 );
buf ( n201332 , n34054 );
not ( n34056 , n201332 );
not ( n34057 , n34056 );
xor ( n34058 , n200805 , n200825 );
xor ( n34059 , n34058 , n200830 );
buf ( n201337 , n34059 );
not ( n34061 , n201337 );
not ( n34062 , n34061 );
or ( n34063 , n34057 , n34062 );
xor ( n34064 , n201318 , n201323 );
xor ( n34065 , n34064 , n201328 );
buf ( n201343 , n34065 );
or ( n34067 , n201343 , n24107 );
nand ( n34068 , n34063 , n34067 );
not ( n34069 , n34068 );
not ( n34070 , n34069 );
or ( n34071 , n34036 , n34070 );
not ( n34072 , n34056 );
nor ( n34073 , n34072 , n201337 );
nand ( n34074 , n201343 , n24107 );
or ( n34075 , n34073 , n34074 );
not ( n34076 , n34056 );
buf ( n34077 , n201337 );
nand ( n34078 , n34076 , n34077 );
nand ( n34079 , n34075 , n34078 );
not ( n34080 , n34079 );
nand ( n34081 , n34071 , n34080 );
not ( n34082 , n33649 );
not ( n34083 , n33636 );
nand ( n34084 , n34083 , n33632 );
not ( n34085 , n200923 );
not ( n34086 , n189835 );
nand ( n34087 , n34085 , n34086 );
nand ( n34088 , n34084 , n34087 );
not ( n34089 , n34088 );
nor ( n34090 , n201305 , n201310 );
nor ( n34091 , n190324 , n201295 );
or ( n34092 , n34090 , n34091 );
nand ( n34093 , n34092 , n34034 );
nand ( n34094 , n34089 , n34093 );
nand ( n34095 , n34082 , n34094 , n34080 );
nand ( n34096 , n33509 , n33558 );
nand ( n34097 , n34096 , n33568 );
nor ( n34098 , n33461 , n34097 );
nand ( n34099 , n34098 , n33428 );
not ( n34100 , n34099 );
nand ( n34101 , n34081 , n34095 , n34100 );
nand ( n34102 , n33605 , n34101 );
not ( n34103 , n34102 );
or ( n34104 , n32873 , n34103 );
not ( n34105 , n200956 );
not ( n34106 , n194823 );
and ( n34107 , n34105 , n34106 );
nor ( n34108 , n192164 , n201288 );
nor ( n34109 , n34107 , n34108 );
not ( n34110 , n34109 );
not ( n34111 , n201305 );
not ( n34112 , n201310 );
nand ( n34113 , n34111 , n34112 );
not ( n34114 , n190324 );
not ( n34115 , n201295 );
nand ( n34116 , n34114 , n34115 );
nand ( n34117 , n34113 , n34116 );
nor ( n34118 , n34110 , n34117 );
not ( n34119 , n34086 );
not ( n34120 , n34085 );
or ( n34121 , n34119 , n34120 );
nand ( n34122 , n34121 , n34084 );
nor ( n34123 , n34068 , n34122 );
nand ( n34124 , n34118 , n34123 );
nor ( n34125 , n34124 , n34099 );
not ( n34126 , n34125 );
not ( n34127 , n34126 );
and ( n34128 , n34127 , n32872 );
buf ( n201406 , n842 );
buf ( n201407 , n890 );
xor ( n34131 , n201406 , n201407 );
buf ( n201409 , n34131 );
buf ( n201410 , n201409 );
not ( n34134 , n201410 );
buf ( n201412 , n188751 );
not ( n34136 , n201412 );
or ( n34137 , n34134 , n34136 );
buf ( n201415 , n20902 );
buf ( n201416 , n192052 );
nand ( n34140 , n201415 , n201416 );
buf ( n201418 , n34140 );
buf ( n201419 , n201418 );
nand ( n34143 , n34137 , n201419 );
buf ( n201421 , n34143 );
not ( n34145 , n201421 );
buf ( n201423 , n850 );
buf ( n201424 , n882 );
xor ( n34148 , n201423 , n201424 );
buf ( n201426 , n34148 );
buf ( n201427 , n201426 );
not ( n34151 , n201427 );
buf ( n201429 , n19613 );
not ( n34153 , n201429 );
or ( n34154 , n34151 , n34153 );
buf ( n201432 , n26571 );
buf ( n201433 , n200990 );
nand ( n34157 , n201432 , n201433 );
buf ( n201435 , n34157 );
buf ( n201436 , n201435 );
nand ( n34160 , n34154 , n201436 );
buf ( n201438 , n34160 );
not ( n34162 , n201438 );
nand ( n34163 , n34145 , n34162 );
not ( n34164 , n34163 );
buf ( n201442 , n863 );
buf ( n201443 , n871 );
or ( n34167 , n201442 , n201443 );
buf ( n201445 , n872 );
nand ( n34169 , n34167 , n201445 );
buf ( n201447 , n34169 );
buf ( n201448 , n201447 );
buf ( n201449 , n863 );
buf ( n201450 , n871 );
nand ( n34174 , n201449 , n201450 );
buf ( n201452 , n34174 );
buf ( n201453 , n201452 );
buf ( n201454 , n870 );
nand ( n34178 , n201448 , n201453 , n201454 );
buf ( n201456 , n34178 );
not ( n34180 , n201456 );
buf ( n201458 , n841 );
buf ( n201459 , n892 );
xor ( n34183 , n201458 , n201459 );
buf ( n201461 , n34183 );
buf ( n201462 , n201461 );
not ( n34186 , n201462 );
buf ( n201464 , n190485 );
not ( n34188 , n201464 );
or ( n34189 , n34186 , n34188 );
buf ( n201467 , n190128 );
buf ( n201468 , n33763 );
nand ( n34192 , n201467 , n201468 );
buf ( n201470 , n34192 );
buf ( n201471 , n201470 );
nand ( n34195 , n34189 , n201471 );
buf ( n201473 , n34195 );
nand ( n34197 , n34180 , n201473 );
not ( n34198 , n34197 );
not ( n34199 , n34198 );
or ( n34200 , n34164 , n34199 );
nand ( n34201 , n201438 , n201421 );
nand ( n34202 , n34200 , n34201 );
xor ( n34203 , n191875 , n191892 );
buf ( n201481 , n34203 );
buf ( n201482 , n191910 );
xnor ( n34206 , n201481 , n201482 );
buf ( n201484 , n34206 );
xor ( n34208 , n34202 , n201484 );
and ( n34209 , n33732 , n201002 );
not ( n34210 , n33732 );
and ( n34211 , n34210 , n201014 );
nor ( n34212 , n34209 , n34211 );
buf ( n34213 , n201057 );
and ( n34214 , n34212 , n34213 );
not ( n34215 , n34212 );
not ( n34216 , n34213 );
and ( n34217 , n34215 , n34216 );
nor ( n34218 , n34214 , n34217 );
xor ( n34219 , n34208 , n34218 );
buf ( n34220 , n34219 );
buf ( n201498 , n34220 );
not ( n34222 , n201498 );
xor ( n34223 , n201132 , n201149 );
xor ( n34224 , n34223 , n201167 );
buf ( n201502 , n34224 );
buf ( n201503 , n201502 );
xor ( n34227 , n201078 , n201094 );
and ( n34228 , n34227 , n201111 );
not ( n34229 , n34227 );
buf ( n201507 , n201111 );
not ( n34231 , n201507 );
buf ( n201509 , n34231 );
and ( n34233 , n34229 , n201509 );
nor ( n34234 , n34228 , n34233 );
buf ( n201512 , n34234 );
xor ( n34236 , n201503 , n201512 );
xor ( n34237 , n201421 , n34162 );
xor ( n34238 , n34237 , n34197 );
buf ( n201516 , n34238 );
and ( n34240 , n34236 , n201516 );
and ( n34241 , n201503 , n201512 );
or ( n34242 , n34240 , n34241 );
buf ( n201520 , n34242 );
buf ( n201521 , n201520 );
not ( n34245 , n201521 );
not ( n34246 , n33973 );
and ( n34247 , n33987 , n34246 );
not ( n34248 , n33987 );
and ( n34249 , n34248 , n33973 );
nor ( n34250 , n34247 , n34249 );
buf ( n201528 , n34250 );
buf ( n201529 , n201254 );
and ( n34253 , n201528 , n201529 );
not ( n34254 , n201528 );
buf ( n34255 , n201260 );
buf ( n201533 , n34255 );
and ( n34257 , n34254 , n201533 );
nor ( n34258 , n34253 , n34257 );
buf ( n201536 , n34258 );
buf ( n201537 , n201536 );
not ( n34261 , n201537 );
and ( n34262 , n34245 , n34261 );
buf ( n201540 , n201520 );
buf ( n201541 , n201536 );
and ( n34265 , n201540 , n201541 );
nor ( n34266 , n34262 , n34265 );
buf ( n201544 , n34266 );
buf ( n201545 , n201544 );
not ( n34269 , n201545 );
or ( n34270 , n34222 , n34269 );
buf ( n201548 , n201544 );
buf ( n201549 , n34220 );
or ( n34273 , n201548 , n201549 );
nand ( n34274 , n34270 , n34273 );
buf ( n201552 , n34274 );
buf ( n201553 , n201552 );
buf ( n201554 , n852 );
buf ( n201555 , n882 );
xor ( n34279 , n201554 , n201555 );
buf ( n201557 , n34279 );
buf ( n201558 , n201557 );
not ( n34282 , n201558 );
buf ( n201560 , n26567 );
not ( n34284 , n201560 );
or ( n34285 , n34282 , n34284 );
buf ( n201563 , n26571 );
buf ( n201564 , n851 );
buf ( n201565 , n882 );
xor ( n34289 , n201564 , n201565 );
buf ( n201567 , n34289 );
buf ( n201568 , n201567 );
nand ( n34292 , n201563 , n201568 );
buf ( n201570 , n34292 );
buf ( n201571 , n201570 );
nand ( n34295 , n34285 , n201571 );
buf ( n201573 , n34295 );
buf ( n201574 , n201573 );
buf ( n201575 , n197086 );
not ( n34299 , n201575 );
buf ( n201577 , n20632 );
not ( n34301 , n201577 );
or ( n34302 , n34299 , n34301 );
buf ( n201580 , n190491 );
buf ( n201581 , n842 );
buf ( n201582 , n892 );
xor ( n34306 , n201581 , n201582 );
buf ( n201584 , n34306 );
buf ( n201585 , n201584 );
nand ( n34309 , n201580 , n201585 );
buf ( n201587 , n34309 );
buf ( n201588 , n201587 );
nand ( n34312 , n34302 , n201588 );
buf ( n201590 , n34312 );
buf ( n201591 , n201590 );
not ( n34315 , n201591 );
buf ( n201593 , n863 );
buf ( n201594 , n873 );
or ( n34318 , n201593 , n201594 );
buf ( n201596 , n874 );
nand ( n34320 , n34318 , n201596 );
buf ( n201598 , n34320 );
buf ( n201599 , n201598 );
buf ( n201600 , n863 );
buf ( n201601 , n873 );
nand ( n34325 , n201600 , n201601 );
buf ( n201603 , n34325 );
buf ( n201604 , n201603 );
buf ( n201605 , n872 );
nand ( n34329 , n201599 , n201604 , n201605 );
buf ( n201607 , n34329 );
buf ( n201608 , n201607 );
nor ( n34332 , n34315 , n201608 );
buf ( n201610 , n34332 );
buf ( n201611 , n201610 );
xor ( n34335 , n201574 , n201611 );
buf ( n201613 , n197123 );
not ( n34337 , n201613 );
buf ( n201615 , n19098 );
not ( n34339 , n201615 );
or ( n34340 , n34337 , n34339 );
buf ( n201618 , n20279 );
buf ( n201619 , n858 );
buf ( n201620 , n876 );
xor ( n34344 , n201619 , n201620 );
buf ( n201622 , n34344 );
buf ( n201623 , n201622 );
nand ( n34347 , n201618 , n201623 );
buf ( n201625 , n34347 );
buf ( n201626 , n201625 );
nand ( n34350 , n34340 , n201626 );
buf ( n201628 , n34350 );
buf ( n201629 , n201628 );
buf ( n201630 , n197141 );
not ( n34354 , n201630 );
buf ( n201632 , n18992 );
not ( n34356 , n201632 );
or ( n34357 , n34354 , n34356 );
buf ( n201635 , n188823 );
buf ( n201636 , n860 );
buf ( n201637 , n874 );
xor ( n34361 , n201636 , n201637 );
buf ( n201639 , n34361 );
buf ( n201640 , n201639 );
nand ( n34364 , n201635 , n201640 );
buf ( n201642 , n34364 );
buf ( n201643 , n201642 );
nand ( n34367 , n34357 , n201643 );
buf ( n201645 , n34367 );
buf ( n201646 , n201645 );
xor ( n34370 , n201629 , n201646 );
not ( n34371 , n23353 );
buf ( n201649 , n848 );
buf ( n201650 , n886 );
xor ( n34374 , n201649 , n201650 );
buf ( n201652 , n34374 );
not ( n34376 , n201652 );
or ( n34377 , n34371 , n34376 );
buf ( n201655 , n197016 );
not ( n34379 , n201655 );
buf ( n201657 , n34379 );
or ( n34381 , n190334 , n201657 );
nand ( n34382 , n34377 , n34381 );
buf ( n201660 , n34382 );
and ( n34384 , n34370 , n201660 );
and ( n34385 , n201629 , n201646 );
or ( n34386 , n34384 , n34385 );
buf ( n201664 , n34386 );
buf ( n201665 , n201664 );
and ( n34389 , n34335 , n201665 );
and ( n34390 , n201574 , n201611 );
or ( n34391 , n34389 , n34390 );
buf ( n201669 , n34391 );
buf ( n201670 , n201669 );
buf ( n201671 , n186441 );
buf ( n201672 , n863 );
and ( n34396 , n201671 , n201672 );
buf ( n201674 , n34396 );
buf ( n201675 , n201674 );
not ( n34399 , n201675 );
buf ( n201677 , n846 );
buf ( n201678 , n888 );
xor ( n34402 , n201677 , n201678 );
buf ( n201680 , n34402 );
buf ( n201681 , n201680 );
not ( n34405 , n201681 );
buf ( n201683 , n22336 );
not ( n34407 , n201683 );
or ( n34408 , n34405 , n34407 );
buf ( n201686 , n20396 );
buf ( n201687 , n845 );
buf ( n201688 , n888 );
xor ( n34412 , n201687 , n201688 );
buf ( n201690 , n34412 );
buf ( n201691 , n201690 );
nand ( n34415 , n201686 , n201691 );
buf ( n201693 , n34415 );
buf ( n201694 , n201693 );
nand ( n34418 , n34408 , n201694 );
buf ( n201696 , n34418 );
buf ( n201697 , n201696 );
not ( n34421 , n201697 );
or ( n34422 , n34399 , n34421 );
buf ( n201700 , n201696 );
buf ( n201701 , n201674 );
or ( n34425 , n201700 , n201701 );
buf ( n201703 , n201584 );
not ( n34427 , n201703 );
buf ( n201705 , n190485 );
not ( n34429 , n201705 );
or ( n34430 , n34427 , n34429 );
buf ( n201708 , n190128 );
buf ( n201709 , n201461 );
nand ( n34433 , n201708 , n201709 );
buf ( n201711 , n34433 );
buf ( n201712 , n201711 );
nand ( n34436 , n34430 , n201712 );
buf ( n201714 , n34436 );
buf ( n201715 , n201714 );
nand ( n34439 , n34425 , n201715 );
buf ( n201717 , n34439 );
buf ( n201718 , n201717 );
nand ( n34442 , n34422 , n201718 );
buf ( n201720 , n34442 );
buf ( n201721 , n201720 );
buf ( n201722 , n862 );
buf ( n201723 , n872 );
xor ( n34447 , n201722 , n201723 );
buf ( n201725 , n34447 );
buf ( n201726 , n201725 );
not ( n34450 , n201726 );
buf ( n201728 , n25318 );
not ( n34452 , n201728 );
or ( n34453 , n34450 , n34452 );
buf ( n201731 , n19264 );
buf ( n201732 , n861 );
buf ( n201733 , n872 );
xor ( n34457 , n201732 , n201733 );
buf ( n201735 , n34457 );
buf ( n201736 , n201735 );
nand ( n34460 , n201731 , n201736 );
buf ( n201738 , n34460 );
buf ( n201739 , n201738 );
nand ( n34463 , n34453 , n201739 );
buf ( n201741 , n34463 );
buf ( n201742 , n201741 );
not ( n34466 , n201742 );
buf ( n201744 , n844 );
buf ( n201745 , n890 );
xor ( n34469 , n201744 , n201745 );
buf ( n201747 , n34469 );
buf ( n201748 , n201747 );
not ( n34472 , n201748 );
buf ( n201750 , n188751 );
not ( n34474 , n201750 );
or ( n34475 , n34472 , n34474 );
buf ( n201753 , n20902 );
buf ( n201754 , n843 );
buf ( n201755 , n890 );
xor ( n34479 , n201754 , n201755 );
buf ( n201757 , n34479 );
buf ( n201758 , n201757 );
nand ( n34482 , n201753 , n201758 );
buf ( n201760 , n34482 );
buf ( n201761 , n201760 );
nand ( n34485 , n34475 , n201761 );
buf ( n201763 , n34485 );
buf ( n201764 , n201763 );
not ( n34488 , n201764 );
or ( n34489 , n34466 , n34488 );
buf ( n201767 , n201763 );
buf ( n201768 , n201741 );
or ( n34492 , n201767 , n201768 );
buf ( n201770 , n850 );
buf ( n201771 , n884 );
xor ( n34495 , n201770 , n201771 );
buf ( n201773 , n34495 );
buf ( n201774 , n201773 );
not ( n34498 , n201774 );
buf ( n201776 , n20727 );
not ( n34500 , n201776 );
or ( n34501 , n34498 , n34500 );
buf ( n201779 , n192573 );
buf ( n201780 , n849 );
buf ( n201781 , n884 );
xor ( n34505 , n201780 , n201781 );
buf ( n201783 , n34505 );
buf ( n201784 , n201783 );
nand ( n34508 , n201779 , n201784 );
buf ( n201786 , n34508 );
buf ( n201787 , n201786 );
nand ( n34511 , n34501 , n201787 );
buf ( n201789 , n34511 );
buf ( n201790 , n201789 );
nand ( n34514 , n34492 , n201790 );
buf ( n201792 , n34514 );
buf ( n201793 , n201792 );
nand ( n34517 , n34489 , n201793 );
buf ( n201795 , n34517 );
buf ( n201796 , n201795 );
xor ( n34520 , n201721 , n201796 );
buf ( n201798 , n201567 );
not ( n34522 , n201798 );
buf ( n201800 , n19613 );
not ( n34524 , n201800 );
or ( n34525 , n34522 , n34524 );
buf ( n201803 , n19942 );
buf ( n201804 , n201426 );
nand ( n34528 , n201803 , n201804 );
buf ( n201806 , n34528 );
buf ( n201807 , n201806 );
nand ( n34531 , n34525 , n201807 );
buf ( n201809 , n34531 );
buf ( n201810 , n201809 );
buf ( n201811 , n863 );
buf ( n201812 , n870 );
xor ( n34536 , n201811 , n201812 );
buf ( n201814 , n34536 );
buf ( n201815 , n201814 );
not ( n34539 , n201815 );
buf ( n201817 , n186432 );
not ( n34541 , n201817 );
or ( n34542 , n34539 , n34541 );
buf ( n201820 , n186441 );
buf ( n201821 , n201154 );
nand ( n34545 , n201820 , n201821 );
buf ( n201823 , n34545 );
buf ( n201824 , n201823 );
nand ( n34548 , n34542 , n201824 );
buf ( n201826 , n34548 );
buf ( n201827 , n201826 );
xor ( n34551 , n201810 , n201827 );
buf ( n201829 , n201757 );
not ( n34553 , n201829 );
buf ( n201831 , n188751 );
not ( n34555 , n201831 );
or ( n34556 , n34553 , n34555 );
buf ( n201834 , n20902 );
buf ( n201835 , n201409 );
nand ( n34559 , n201834 , n201835 );
buf ( n201837 , n34559 );
buf ( n201838 , n201837 );
nand ( n34562 , n34556 , n201838 );
buf ( n201840 , n34562 );
buf ( n201841 , n201840 );
xor ( n34565 , n34551 , n201841 );
buf ( n201843 , n34565 );
buf ( n201844 , n201843 );
xor ( n34568 , n34520 , n201844 );
buf ( n201846 , n34568 );
buf ( n201847 , n201846 );
xor ( n34571 , n201670 , n201847 );
buf ( n201849 , n201714 );
buf ( n201850 , n189037 );
buf ( n201851 , n863 );
and ( n34575 , n201850 , n201851 );
buf ( n201853 , n34575 );
buf ( n201854 , n201853 );
and ( n34578 , n201849 , n201854 );
not ( n34579 , n201849 );
buf ( n201857 , n201853 );
not ( n34581 , n201857 );
buf ( n201859 , n34581 );
buf ( n201860 , n201859 );
and ( n34584 , n34579 , n201860 );
nor ( n34585 , n34578 , n34584 );
buf ( n201863 , n34585 );
buf ( n201864 , n201863 );
buf ( n201865 , n201696 );
and ( n34589 , n201864 , n201865 );
not ( n34590 , n201864 );
buf ( n201868 , n201696 );
not ( n34592 , n201868 );
buf ( n201870 , n34592 );
buf ( n201871 , n201870 );
and ( n34595 , n34590 , n201871 );
nor ( n34596 , n34589 , n34595 );
buf ( n201874 , n34596 );
buf ( n201875 , n201874 );
not ( n34599 , n201875 );
not ( n34600 , n201652 );
not ( n34601 , n20554 );
or ( n34602 , n34600 , n34601 );
buf ( n201880 , n20558 );
buf ( n201881 , n847 );
buf ( n201882 , n886 );
xor ( n34606 , n201881 , n201882 );
buf ( n201884 , n34606 );
buf ( n201885 , n201884 );
nand ( n34609 , n201880 , n201885 );
buf ( n201887 , n34609 );
nand ( n34611 , n34602 , n201887 );
buf ( n201889 , n854 );
buf ( n201890 , n880 );
xor ( n34614 , n201889 , n201890 );
buf ( n201892 , n34614 );
not ( n34616 , n201892 );
not ( n34617 , n18862 );
or ( n34618 , n34616 , n34617 );
buf ( n201896 , n20358 );
buf ( n201897 , n853 );
buf ( n201898 , n880 );
xor ( n34622 , n201897 , n201898 );
buf ( n201900 , n34622 );
buf ( n201901 , n201900 );
nand ( n34625 , n201896 , n201901 );
buf ( n201903 , n34625 );
nand ( n34627 , n34618 , n201903 );
xor ( n34628 , n34611 , n34627 );
buf ( n201906 , n856 );
buf ( n201907 , n878 );
xor ( n34631 , n201906 , n201907 );
buf ( n201909 , n34631 );
not ( n34633 , n201909 );
not ( n34634 , n186569 );
or ( n34635 , n34633 , n34634 );
buf ( n201913 , n186575 );
buf ( n201914 , n855 );
buf ( n201915 , n878 );
xor ( n34639 , n201914 , n201915 );
buf ( n201917 , n34639 );
buf ( n201918 , n201917 );
nand ( n34642 , n201913 , n201918 );
buf ( n201920 , n34642 );
nand ( n34644 , n34635 , n201920 );
xor ( n34645 , n34628 , n34644 );
buf ( n201923 , n34645 );
not ( n34647 , n201923 );
or ( n34648 , n34599 , n34647 );
buf ( n201926 , n34645 );
buf ( n201927 , n201874 );
or ( n34651 , n201926 , n201927 );
buf ( n201929 , n840 );
buf ( n201930 , n894 );
xor ( n34654 , n201929 , n201930 );
buf ( n201932 , n34654 );
buf ( n201933 , n201932 );
not ( n34657 , n201933 );
buf ( n201935 , n21330 );
not ( n34659 , n201935 );
or ( n34660 , n34657 , n34659 );
buf ( n201938 , n839 );
buf ( n201939 , n894 );
xor ( n34663 , n201938 , n201939 );
buf ( n201941 , n34663 );
buf ( n201942 , n201941 );
buf ( n201943 , n895 );
nand ( n34667 , n201942 , n201943 );
buf ( n201945 , n34667 );
buf ( n201946 , n201945 );
nand ( n34670 , n34660 , n201946 );
buf ( n201948 , n34670 );
buf ( n201949 , n201948 );
buf ( n201950 , n201622 );
not ( n34674 , n201950 );
buf ( n201952 , n19098 );
not ( n34676 , n201952 );
or ( n34677 , n34674 , n34676 );
buf ( n201955 , n19103 );
buf ( n201956 , n857 );
buf ( n201957 , n876 );
xor ( n34681 , n201956 , n201957 );
buf ( n201959 , n34681 );
buf ( n201960 , n201959 );
nand ( n34684 , n201955 , n201960 );
buf ( n201962 , n34684 );
buf ( n201963 , n201962 );
nand ( n34687 , n34677 , n201963 );
buf ( n201965 , n34687 );
buf ( n201966 , n201965 );
xor ( n34690 , n201949 , n201966 );
buf ( n201968 , n201639 );
not ( n34692 , n201968 );
buf ( n201970 , n186287 );
not ( n34694 , n201970 );
or ( n34695 , n34692 , n34694 );
buf ( n201973 , n186297 );
xor ( n34697 , n874 , n859 );
buf ( n201975 , n34697 );
nand ( n34699 , n201973 , n201975 );
buf ( n201977 , n34699 );
buf ( n201978 , n201977 );
nand ( n34702 , n34695 , n201978 );
buf ( n201980 , n34702 );
buf ( n201981 , n201980 );
xor ( n34705 , n34690 , n201981 );
buf ( n201983 , n34705 );
buf ( n201984 , n201983 );
nand ( n34708 , n34651 , n201984 );
buf ( n201986 , n34708 );
buf ( n201987 , n201986 );
nand ( n34711 , n34648 , n201987 );
buf ( n201989 , n34711 );
buf ( n201990 , n201989 );
and ( n34714 , n34571 , n201990 );
and ( n34715 , n201670 , n201847 );
or ( n34716 , n34714 , n34715 );
buf ( n201994 , n34716 );
buf ( n201995 , n201994 );
not ( n34719 , n23321 );
not ( n34720 , n197105 );
or ( n34721 , n34719 , n34720 );
buf ( n201999 , n201932 );
buf ( n202000 , n895 );
nand ( n34724 , n201999 , n202000 );
buf ( n202002 , n34724 );
nand ( n34726 , n34721 , n202002 );
not ( n34727 , n196960 );
not ( n34728 , n188751 );
or ( n34729 , n34727 , n34728 );
buf ( n202007 , n20902 );
buf ( n202008 , n201747 );
nand ( n34732 , n202007 , n202008 );
buf ( n202010 , n34732 );
nand ( n34734 , n34729 , n202010 );
xor ( n34735 , n34726 , n34734 );
not ( n34736 , n19265 );
not ( n34737 , n201725 );
or ( n34738 , n34736 , n34737 );
buf ( n202016 , n863 );
buf ( n202017 , n872 );
xor ( n34741 , n202016 , n202017 );
buf ( n202019 , n34741 );
nand ( n34743 , n19260 , n202019 );
nand ( n34744 , n34738 , n34743 );
and ( n34745 , n34735 , n34744 );
and ( n34746 , n34726 , n34734 );
or ( n34747 , n34745 , n34746 );
buf ( n202025 , n34747 );
xor ( n34749 , n201741 , n201763 );
xor ( n34750 , n34749 , n201789 );
buf ( n202028 , n34750 );
xor ( n34752 , n202025 , n202028 );
not ( n34753 , n197067 );
not ( n34754 , n190454 );
or ( n34755 , n34753 , n34754 );
buf ( n202033 , n20396 );
buf ( n202034 , n201680 );
nand ( n34758 , n202033 , n202034 );
buf ( n202036 , n34758 );
nand ( n34760 , n34755 , n202036 );
not ( n34761 , n34760 );
not ( n34762 , n34761 );
buf ( n202040 , n197045 );
not ( n34764 , n202040 );
buf ( n202042 , n186569 );
not ( n34766 , n202042 );
or ( n34767 , n34764 , n34766 );
buf ( n202045 , n186575 );
buf ( n202046 , n201909 );
nand ( n34770 , n202045 , n202046 );
buf ( n202048 , n34770 );
buf ( n202049 , n202048 );
nand ( n34773 , n34767 , n202049 );
buf ( n202051 , n34773 );
not ( n34775 , n202051 );
not ( n34776 , n34775 );
or ( n34777 , n34762 , n34776 );
buf ( n202055 , n197030 );
not ( n34779 , n202055 );
buf ( n202057 , n186924 );
not ( n34781 , n202057 );
or ( n34782 , n34779 , n34781 );
buf ( n202060 , n22304 );
buf ( n202061 , n201892 );
nand ( n34785 , n202060 , n202061 );
buf ( n202063 , n34785 );
buf ( n202064 , n202063 );
nand ( n34788 , n34782 , n202064 );
buf ( n202066 , n34788 );
nand ( n34790 , n34777 , n202066 );
nand ( n34791 , n202051 , n34760 );
nand ( n34792 , n34790 , n34791 );
buf ( n202070 , n34792 );
and ( n34794 , n34752 , n202070 );
and ( n34795 , n202025 , n202028 );
or ( n34796 , n34794 , n34795 );
buf ( n202074 , n34796 );
buf ( n202075 , n202074 );
not ( n34799 , n202075 );
or ( n34800 , n34627 , n34611 );
nand ( n34801 , n34800 , n34644 );
nand ( n34802 , n34627 , n34611 );
nand ( n34803 , n34801 , n34802 );
not ( n34804 , n201456 );
not ( n34805 , n34804 );
not ( n34806 , n201473 );
or ( n34807 , n34805 , n34806 );
or ( n34808 , n201473 , n34804 );
nand ( n34809 , n34807 , n34808 );
xor ( n34810 , n34803 , n34809 );
xor ( n34811 , n201949 , n201966 );
and ( n34812 , n34811 , n201981 );
and ( n34813 , n201949 , n201966 );
or ( n34814 , n34812 , n34813 );
buf ( n202092 , n34814 );
xor ( n34816 , n34810 , n202092 );
buf ( n202094 , n34816 );
not ( n34818 , n202094 );
buf ( n202096 , n34818 );
buf ( n202097 , n202096 );
not ( n34821 , n202097 );
or ( n34822 , n34799 , n34821 );
buf ( n202100 , n34816 );
not ( n34824 , n202100 );
buf ( n202102 , n202074 );
not ( n34826 , n202102 );
buf ( n202104 , n34826 );
buf ( n202105 , n202104 );
not ( n34829 , n202105 );
or ( n34830 , n34824 , n34829 );
buf ( n202108 , n201941 );
not ( n34832 , n202108 );
buf ( n202110 , n20165 );
not ( n34834 , n202110 );
or ( n34835 , n34832 , n34834 );
buf ( n202113 , n201178 );
buf ( n202114 , n895 );
nand ( n34838 , n202113 , n202114 );
buf ( n202116 , n34838 );
buf ( n202117 , n202116 );
nand ( n34841 , n34835 , n202117 );
buf ( n202119 , n34841 );
buf ( n202120 , n202119 );
buf ( n202121 , n201783 );
not ( n34845 , n202121 );
buf ( n202123 , n20727 );
not ( n34847 , n202123 );
or ( n34848 , n34845 , n34847 );
buf ( n202126 , n188010 );
buf ( n202127 , n201136 );
nand ( n34851 , n202126 , n202127 );
buf ( n202129 , n34851 );
buf ( n202130 , n202129 );
nand ( n34854 , n34848 , n202130 );
buf ( n202132 , n34854 );
buf ( n202133 , n202132 );
xor ( n34857 , n202120 , n202133 );
buf ( n202135 , n201735 );
not ( n34859 , n202135 );
buf ( n202137 , n25318 );
not ( n34861 , n202137 );
or ( n34862 , n34859 , n34861 );
buf ( n202140 , n19265 );
buf ( n202141 , n33842 );
nand ( n34865 , n202140 , n202141 );
buf ( n202143 , n34865 );
buf ( n202144 , n202143 );
nand ( n34868 , n34862 , n202144 );
buf ( n202146 , n34868 );
buf ( n202147 , n202146 );
xor ( n34871 , n34857 , n202147 );
buf ( n202149 , n34871 );
buf ( n202150 , n202149 );
buf ( n202151 , n201900 );
not ( n34875 , n202151 );
buf ( n202153 , n18862 );
not ( n34877 , n202153 );
or ( n34878 , n34875 , n34877 );
buf ( n202156 , n18875 );
buf ( n202157 , n201066 );
nand ( n34881 , n202156 , n202157 );
buf ( n202159 , n34881 );
buf ( n202160 , n202159 );
nand ( n34884 , n34878 , n202160 );
buf ( n202162 , n34884 );
buf ( n202163 , n201690 );
not ( n34887 , n202163 );
buf ( n202165 , n22336 );
not ( n34889 , n202165 );
or ( n34890 , n34887 , n34889 );
buf ( n202168 , n20396 );
buf ( n202169 , n33748 );
nand ( n34893 , n202168 , n202169 );
buf ( n202171 , n34893 );
buf ( n202172 , n202171 );
nand ( n34896 , n34890 , n202172 );
buf ( n202174 , n34896 );
xor ( n34898 , n202162 , n202174 );
buf ( n202176 , n201917 );
not ( n34900 , n202176 );
buf ( n202178 , n186569 );
not ( n34902 , n202178 );
or ( n34903 , n34900 , n34902 );
buf ( n202181 , n186575 );
buf ( n202182 , n201099 );
nand ( n34906 , n202181 , n202182 );
buf ( n202184 , n34906 );
buf ( n202185 , n202184 );
nand ( n34909 , n34903 , n202185 );
buf ( n202187 , n34909 );
xor ( n34911 , n34898 , n202187 );
buf ( n202189 , n34911 );
xor ( n34913 , n202150 , n202189 );
buf ( n202191 , n201959 );
not ( n34915 , n202191 );
buf ( n202193 , n19177 );
not ( n34917 , n202193 );
or ( n34918 , n34915 , n34917 );
buf ( n202196 , n19103 );
buf ( n202197 , n201203 );
nand ( n34921 , n202196 , n202197 );
buf ( n202199 , n34921 );
buf ( n202200 , n202199 );
nand ( n34924 , n34918 , n202200 );
buf ( n202202 , n34924 );
buf ( n202203 , n201884 );
not ( n34927 , n202203 );
buf ( n202205 , n21850 );
not ( n34929 , n202205 );
or ( n34930 , n34927 , n34929 );
buf ( n202208 , n20558 );
buf ( n202209 , n201082 );
nand ( n34933 , n202208 , n202209 );
buf ( n202211 , n34933 );
buf ( n202212 , n202211 );
nand ( n34936 , n34930 , n202212 );
buf ( n202214 , n34936 );
xor ( n34938 , n202202 , n202214 );
buf ( n202216 , n186287 );
buf ( n202217 , n34697 );
and ( n34941 , n202216 , n202217 );
buf ( n202219 , n187865 );
buf ( n202220 , n33915 );
and ( n34944 , n202219 , n202220 );
nor ( n34945 , n34941 , n34944 );
buf ( n202223 , n34945 );
xnor ( n34947 , n34938 , n202223 );
buf ( n202225 , n34947 );
xor ( n34949 , n34913 , n202225 );
buf ( n202227 , n34949 );
buf ( n202228 , n202227 );
nand ( n34952 , n34830 , n202228 );
buf ( n202230 , n34952 );
buf ( n202231 , n202230 );
nand ( n34955 , n34822 , n202231 );
buf ( n202233 , n34955 );
buf ( n202234 , n202233 );
xor ( n34958 , n201995 , n202234 );
buf ( n202236 , n34809 );
not ( n34960 , n202236 );
buf ( n202238 , n34803 );
not ( n34962 , n202238 );
buf ( n202240 , n34962 );
buf ( n202241 , n202240 );
not ( n34965 , n202241 );
or ( n34966 , n34960 , n34965 );
buf ( n202244 , n202092 );
nand ( n34968 , n34966 , n202244 );
buf ( n202246 , n34968 );
buf ( n202247 , n202246 );
not ( n34971 , n34802 );
not ( n34972 , n34801 );
or ( n34973 , n34971 , n34972 );
not ( n34974 , n34809 );
nand ( n34975 , n34973 , n34974 );
buf ( n202253 , n34975 );
nand ( n34977 , n202247 , n202253 );
buf ( n202255 , n34977 );
buf ( n202256 , n202255 );
xor ( n34980 , n201721 , n201796 );
and ( n34981 , n34980 , n201844 );
and ( n34982 , n201721 , n201796 );
or ( n34983 , n34981 , n34982 );
buf ( n202261 , n34983 );
buf ( n202262 , n202261 );
xor ( n34986 , n202256 , n202262 );
xor ( n34987 , n202150 , n202189 );
and ( n34988 , n34987 , n202225 );
and ( n34989 , n202150 , n202189 );
or ( n34990 , n34988 , n34989 );
buf ( n202268 , n34990 );
buf ( n202269 , n202268 );
xor ( n34993 , n34986 , n202269 );
buf ( n202271 , n34993 );
buf ( n202272 , n202271 );
and ( n34996 , n34958 , n202272 );
and ( n34997 , n201995 , n202234 );
or ( n34998 , n34996 , n34997 );
buf ( n202276 , n34998 );
buf ( n202277 , n202276 );
xor ( n35001 , n201553 , n202277 );
xor ( n35002 , n202256 , n202262 );
and ( n35003 , n35002 , n202269 );
and ( n35004 , n202256 , n202262 );
or ( n35005 , n35003 , n35004 );
buf ( n202283 , n35005 );
buf ( n202284 , n202283 );
buf ( n202285 , n202162 );
not ( n35009 , n202285 );
buf ( n202287 , n202174 );
not ( n35011 , n202287 );
or ( n35012 , n35009 , n35011 );
buf ( n202290 , n202174 );
buf ( n202291 , n202162 );
or ( n35015 , n202290 , n202291 );
buf ( n202293 , n202187 );
nand ( n35017 , n35015 , n202293 );
buf ( n202295 , n35017 );
buf ( n202296 , n202295 );
nand ( n35020 , n35012 , n202296 );
buf ( n202298 , n35020 );
not ( n35022 , n202298 );
xor ( n35023 , n202120 , n202133 );
and ( n35024 , n35023 , n202147 );
and ( n35025 , n202120 , n202133 );
or ( n35026 , n35024 , n35025 );
buf ( n202304 , n35026 );
buf ( n202305 , n202304 );
not ( n35029 , n202305 );
buf ( n202307 , n35029 );
nand ( n35031 , n35022 , n202307 );
not ( n35032 , n35031 );
not ( n35033 , n202214 );
not ( n35034 , n202202 );
or ( n35035 , n35033 , n35034 );
buf ( n202313 , n202214 );
buf ( n202314 , n202202 );
nor ( n35038 , n202313 , n202314 );
buf ( n202316 , n35038 );
or ( n35040 , n202316 , n202223 );
nand ( n35041 , n35035 , n35040 );
not ( n35042 , n35041 );
or ( n35043 , n35032 , n35042 );
buf ( n202321 , n202298 );
buf ( n202322 , n202304 );
nand ( n35046 , n202321 , n202322 );
buf ( n202324 , n35046 );
nand ( n35048 , n35043 , n202324 );
buf ( n202326 , n35048 );
xor ( n35050 , n201024 , n201038 );
xor ( n35051 , n35050 , n201053 );
buf ( n202329 , n35051 );
not ( n35053 , n202329 );
xor ( n35054 , n201810 , n201827 );
and ( n35055 , n35054 , n201841 );
and ( n35056 , n201810 , n201827 );
or ( n35057 , n35055 , n35056 );
buf ( n202335 , n35057 );
not ( n35059 , n202335 );
or ( n35060 , n35053 , n35059 );
or ( n35061 , n202329 , n202335 );
xor ( n35062 , n201191 , n201198 );
xor ( n35063 , n35062 , n201209 );
buf ( n202341 , n35063 );
nand ( n35065 , n35061 , n202341 );
nand ( n35066 , n35060 , n35065 );
buf ( n202344 , n35066 );
xor ( n35068 , n202326 , n202344 );
and ( n35069 , n33840 , n201216 );
not ( n35070 , n33840 );
and ( n35071 , n35070 , n201213 );
nor ( n35072 , n35069 , n35071 );
buf ( n202350 , n35072 );
buf ( n202351 , n201171 );
not ( n35075 , n202351 );
buf ( n202353 , n35075 );
buf ( n202354 , n202353 );
and ( n35078 , n202350 , n202354 );
not ( n35079 , n202350 );
buf ( n202357 , n201171 );
and ( n35081 , n35079 , n202357 );
nor ( n35082 , n35078 , n35081 );
buf ( n202360 , n35082 );
buf ( n202361 , n202360 );
xor ( n35085 , n35068 , n202361 );
buf ( n202363 , n35085 );
buf ( n202364 , n202363 );
xor ( n35088 , n202284 , n202364 );
xor ( n35089 , n201503 , n201512 );
xor ( n35090 , n35089 , n201516 );
buf ( n202368 , n35090 );
buf ( n202369 , n202368 );
buf ( n202370 , n202298 );
not ( n35094 , n202370 );
buf ( n202372 , n35041 );
not ( n35096 , n202372 );
buf ( n202374 , n35096 );
buf ( n202375 , n202374 );
not ( n35099 , n202375 );
or ( n35100 , n35094 , n35099 );
buf ( n202378 , n202374 );
buf ( n202379 , n202298 );
or ( n35103 , n202378 , n202379 );
nand ( n35104 , n35100 , n35103 );
buf ( n202382 , n35104 );
buf ( n202383 , n202382 );
buf ( n202384 , n202307 );
and ( n35108 , n202383 , n202384 );
not ( n35109 , n202383 );
buf ( n202387 , n202304 );
and ( n35111 , n35109 , n202387 );
nor ( n35112 , n35108 , n35111 );
buf ( n202390 , n35112 );
buf ( n202391 , n202390 );
not ( n35115 , n202391 );
buf ( n202393 , n35115 );
buf ( n202394 , n202393 );
or ( n35118 , n202369 , n202394 );
xor ( n35119 , n202335 , n202329 );
xor ( n35120 , n35119 , n202341 );
buf ( n202398 , n35120 );
nand ( n35122 , n35118 , n202398 );
buf ( n202400 , n35122 );
buf ( n202401 , n202400 );
buf ( n202402 , n202393 );
buf ( n202403 , n202368 );
nand ( n35127 , n202402 , n202403 );
buf ( n202405 , n35127 );
buf ( n202406 , n202405 );
nand ( n35130 , n202401 , n202406 );
buf ( n202408 , n35130 );
buf ( n202409 , n202408 );
xor ( n35133 , n35088 , n202409 );
buf ( n202411 , n35133 );
buf ( n202412 , n202411 );
and ( n35136 , n35001 , n202412 );
and ( n35137 , n201553 , n202277 );
or ( n35138 , n35136 , n35137 );
buf ( n202416 , n35138 );
not ( n35140 , n202416 );
xor ( n35141 , n34202 , n201484 );
and ( n35142 , n35141 , n34218 );
and ( n35143 , n34202 , n201484 );
or ( n35144 , n35142 , n35143 );
buf ( n202422 , n35144 );
buf ( n202423 , n24662 );
not ( n35147 , n202423 );
buf ( n202425 , n191948 );
not ( n35149 , n202425 );
or ( n35150 , n35147 , n35149 );
buf ( n202428 , n24662 );
buf ( n202429 , n191948 );
or ( n35153 , n202428 , n202429 );
nand ( n35154 , n35150 , n35153 );
buf ( n202432 , n35154 );
buf ( n202433 , n202432 );
buf ( n202434 , n191957 );
and ( n35158 , n202433 , n202434 );
not ( n35159 , n202433 );
buf ( n35160 , n191927 );
buf ( n202438 , n35160 );
and ( n35162 , n35159 , n202438 );
nor ( n35163 , n35158 , n35162 );
buf ( n202441 , n35163 );
buf ( n202442 , n202441 );
xor ( n35166 , n202422 , n202442 );
xor ( n35167 , n202326 , n202344 );
and ( n35168 , n35167 , n202361 );
and ( n35169 , n202326 , n202344 );
or ( n35170 , n35168 , n35169 );
buf ( n202448 , n35170 );
buf ( n202449 , n202448 );
xor ( n35173 , n35166 , n202449 );
buf ( n202451 , n35173 );
buf ( n202452 , n202451 );
xor ( n35176 , n202284 , n202364 );
and ( n35177 , n35176 , n202409 );
and ( n35178 , n202284 , n202364 );
or ( n35179 , n35177 , n35178 );
buf ( n202457 , n35179 );
buf ( n202458 , n202457 );
xor ( n35182 , n202452 , n202458 );
xor ( n35183 , n33709 , n33784 );
xor ( n35184 , n35183 , n33941 );
buf ( n202462 , n35184 );
buf ( n202463 , n33989 );
not ( n35187 , n202463 );
buf ( n202465 , n33948 );
not ( n35189 , n202465 );
buf ( n202467 , n35189 );
buf ( n202468 , n202467 );
not ( n35192 , n202468 );
or ( n35193 , n35187 , n35192 );
not ( n35194 , n33989 );
nand ( n35195 , n35194 , n33948 );
buf ( n202473 , n35195 );
nand ( n35197 , n35193 , n202473 );
buf ( n202475 , n35197 );
buf ( n202476 , n202475 );
buf ( n202477 , n201229 );
buf ( n35201 , n202477 );
buf ( n202479 , n35201 );
buf ( n202480 , n202479 );
xor ( n35204 , n202476 , n202480 );
buf ( n202482 , n35204 );
buf ( n202483 , n202482 );
xor ( n35207 , n202462 , n202483 );
not ( n35208 , n201520 );
not ( n35209 , n34219 );
or ( n35210 , n35208 , n35209 );
buf ( n202488 , n34219 );
buf ( n202489 , n201520 );
or ( n35213 , n202488 , n202489 );
buf ( n202491 , n201536 );
not ( n35215 , n202491 );
buf ( n202493 , n35215 );
buf ( n202494 , n202493 );
nand ( n35218 , n35213 , n202494 );
buf ( n202496 , n35218 );
nand ( n35220 , n35210 , n202496 );
buf ( n202498 , n35220 );
xor ( n35222 , n35207 , n202498 );
buf ( n202500 , n35222 );
buf ( n202501 , n202500 );
xor ( n35225 , n35182 , n202501 );
buf ( n202503 , n35225 );
not ( n35227 , n202503 );
nand ( n35228 , n35140 , n35227 );
xor ( n35229 , n202422 , n202442 );
and ( n35230 , n35229 , n202449 );
and ( n35231 , n202422 , n202442 );
or ( n35232 , n35230 , n35231 );
buf ( n202510 , n35232 );
buf ( n202511 , n202510 );
xor ( n35235 , n202462 , n202483 );
and ( n35236 , n35235 , n202498 );
and ( n35237 , n202462 , n202483 );
or ( n35238 , n35236 , n35237 );
buf ( n202516 , n35238 );
buf ( n202517 , n202516 );
xor ( n35241 , n202511 , n202517 );
xor ( n35242 , n191774 , n191916 );
xor ( n35243 , n35242 , n191964 );
buf ( n202521 , n35243 );
buf ( n202522 , n202521 );
buf ( n202523 , n24706 );
not ( n35247 , n202523 );
buf ( n202525 , n192120 );
not ( n35249 , n202525 );
and ( n35250 , n35247 , n35249 );
buf ( n202528 , n24706 );
buf ( n202529 , n192120 );
and ( n35253 , n202528 , n202529 );
nor ( n35254 , n35250 , n35253 );
buf ( n202532 , n35254 );
buf ( n202533 , n202532 );
buf ( n202534 , n191991 );
and ( n35258 , n202533 , n202534 );
not ( n35259 , n202533 );
buf ( n202537 , n192129 );
and ( n35261 , n35259 , n202537 );
nor ( n35262 , n35258 , n35261 );
buf ( n202540 , n35262 );
buf ( n202541 , n202540 );
xor ( n35265 , n202522 , n202541 );
xor ( n35266 , n200975 , n201222 );
xor ( n35267 , n35266 , n201269 );
buf ( n202545 , n35267 );
buf ( n202546 , n202545 );
xor ( n35270 , n35265 , n202546 );
buf ( n202548 , n35270 );
buf ( n202549 , n202548 );
xor ( n35273 , n35241 , n202549 );
buf ( n202551 , n35273 );
not ( n35275 , n202551 );
xor ( n35276 , n202452 , n202458 );
and ( n35277 , n35276 , n202501 );
and ( n35278 , n202452 , n202458 );
or ( n35279 , n35277 , n35278 );
buf ( n202557 , n35279 );
not ( n35281 , n202557 );
nand ( n35282 , n35275 , n35281 );
nand ( n35283 , n35228 , n35282 );
not ( n35284 , n35283 );
xor ( n35285 , n202511 , n202517 );
and ( n35286 , n35285 , n202549 );
and ( n35287 , n202511 , n202517 );
or ( n35288 , n35286 , n35287 );
buf ( n202566 , n35288 );
xor ( n35290 , n191771 , n191969 );
xor ( n35291 , n35290 , n192136 );
buf ( n202569 , n35291 );
buf ( n202570 , n202569 );
xor ( n35294 , n200967 , n200971 );
xor ( n35295 , n35294 , n201274 );
buf ( n202573 , n35295 );
buf ( n202574 , n202573 );
xor ( n35298 , n202570 , n202574 );
xor ( n35299 , n202522 , n202541 );
and ( n35300 , n35299 , n202546 );
and ( n35301 , n202522 , n202541 );
or ( n35302 , n35300 , n35301 );
buf ( n202580 , n35302 );
buf ( n202581 , n202580 );
xor ( n35305 , n35298 , n202581 );
buf ( n202583 , n35305 );
nor ( n35307 , n202566 , n202583 );
xor ( n35308 , n200963 , n201279 );
xor ( n35309 , n35308 , n201284 );
buf ( n202587 , n35309 );
xor ( n35311 , n202570 , n202574 );
and ( n35312 , n35311 , n202581 );
and ( n35313 , n202570 , n202574 );
or ( n35314 , n35312 , n35313 );
buf ( n202592 , n35314 );
nor ( n35316 , n202587 , n202592 );
nor ( n35317 , n35307 , n35316 );
nand ( n35318 , n35284 , n35317 );
not ( n35319 , n35318 );
xor ( n35320 , n201553 , n202277 );
xor ( n35321 , n35320 , n202412 );
buf ( n202599 , n35321 );
xor ( n35323 , n202390 , n202368 );
xnor ( n35324 , n35323 , n35120 );
buf ( n202602 , n35324 );
buf ( n202603 , n196977 );
not ( n35327 , n202603 );
buf ( n202605 , n192332 );
not ( n35329 , n202605 );
or ( n35330 , n35327 , n35329 );
buf ( n202608 , n192573 );
buf ( n202609 , n201773 );
nand ( n35333 , n202608 , n202609 );
buf ( n202611 , n35333 );
buf ( n202612 , n202611 );
nand ( n35336 , n35330 , n202612 );
buf ( n202614 , n35336 );
buf ( n202615 , n202614 );
buf ( n202616 , n196995 );
not ( n35340 , n202616 );
buf ( n202618 , n19613 );
not ( n35342 , n202618 );
or ( n35343 , n35340 , n35342 );
buf ( n202621 , n26571 );
buf ( n202622 , n201557 );
nand ( n35346 , n202621 , n202622 );
buf ( n202624 , n35346 );
buf ( n202625 , n202624 );
nand ( n35349 , n35343 , n202625 );
buf ( n202627 , n35349 );
buf ( n202628 , n202627 );
xor ( n35352 , n202615 , n202628 );
buf ( n202630 , n201590 );
not ( n35354 , n202630 );
buf ( n202632 , n201607 );
not ( n35356 , n202632 );
or ( n35357 , n35354 , n35356 );
buf ( n202635 , n201590 );
buf ( n202636 , n201607 );
or ( n35360 , n202635 , n202636 );
nand ( n35361 , n35357 , n35360 );
buf ( n202639 , n35361 );
buf ( n202640 , n202639 );
and ( n35364 , n35352 , n202640 );
and ( n35365 , n202615 , n202628 );
or ( n35366 , n35364 , n35365 );
buf ( n202644 , n35366 );
buf ( n202645 , n202644 );
xor ( n35369 , n201574 , n201611 );
xor ( n35370 , n35369 , n201665 );
buf ( n202648 , n35370 );
buf ( n202649 , n202648 );
xor ( n35373 , n202645 , n202649 );
xor ( n35374 , n197058 , n197075 );
and ( n35375 , n35374 , n197093 );
and ( n35376 , n197058 , n197075 );
or ( n35377 , n35375 , n35376 );
buf ( n202655 , n35377 );
buf ( n202656 , n202655 );
xor ( n35380 , n197113 , n197130 );
and ( n35381 , n35380 , n197148 );
and ( n35382 , n197113 , n197130 );
or ( n35383 , n35381 , n35382 );
buf ( n202661 , n35383 );
buf ( n202662 , n202661 );
xor ( n35386 , n202656 , n202662 );
xor ( n35387 , n196967 , n196984 );
and ( n35388 , n35387 , n197002 );
and ( n35389 , n196967 , n196984 );
or ( n35390 , n35388 , n35389 );
buf ( n202668 , n35390 );
buf ( n202669 , n202668 );
and ( n35393 , n35386 , n202669 );
and ( n35394 , n202656 , n202662 );
or ( n35395 , n35393 , n35394 );
buf ( n202673 , n35395 );
buf ( n202674 , n202673 );
and ( n35398 , n35373 , n202674 );
and ( n35399 , n202645 , n202649 );
or ( n35400 , n35398 , n35399 );
buf ( n202678 , n35400 );
buf ( n202679 , n202678 );
xor ( n35403 , n201670 , n201847 );
xor ( n35404 , n35403 , n201990 );
buf ( n202682 , n35404 );
buf ( n202683 , n202682 );
xor ( n35407 , n202679 , n202683 );
buf ( n202685 , n29757 );
buf ( n202686 , n197022 );
or ( n35410 , n202685 , n202686 );
buf ( n202688 , n197051 );
nand ( n35412 , n35410 , n202688 );
buf ( n202690 , n35412 );
buf ( n202691 , n202690 );
buf ( n202692 , n29757 );
buf ( n202693 , n197022 );
nand ( n35417 , n202692 , n202693 );
buf ( n202695 , n35417 );
buf ( n202696 , n202695 );
nand ( n35420 , n202691 , n202696 );
buf ( n202698 , n35420 );
buf ( n202699 , n202698 );
xor ( n35423 , n34726 , n34734 );
xor ( n35424 , n35423 , n34744 );
buf ( n202702 , n35424 );
xor ( n35426 , n202699 , n202702 );
xor ( n35427 , n201629 , n201646 );
xor ( n35428 , n35427 , n201660 );
buf ( n202706 , n35428 );
buf ( n202707 , n202706 );
and ( n35431 , n35426 , n202707 );
and ( n35432 , n202699 , n202702 );
or ( n35433 , n35431 , n35432 );
buf ( n202711 , n35433 );
buf ( n202712 , n202711 );
not ( n35436 , n202712 );
buf ( n202714 , n35436 );
buf ( n202715 , n202714 );
not ( n35439 , n202715 );
xor ( n35440 , n202025 , n202028 );
xor ( n35441 , n35440 , n202070 );
buf ( n202719 , n35441 );
buf ( n202720 , n202719 );
not ( n35444 , n202720 );
buf ( n202722 , n35444 );
buf ( n202723 , n202722 );
not ( n35447 , n202723 );
or ( n35448 , n35439 , n35447 );
xor ( n35449 , n201983 , n201874 );
xor ( n35450 , n35449 , n34645 );
buf ( n202728 , n35450 );
nand ( n35452 , n35448 , n202728 );
buf ( n202730 , n35452 );
buf ( n202731 , n202730 );
buf ( n202732 , n202719 );
buf ( n202733 , n202711 );
nand ( n35457 , n202732 , n202733 );
buf ( n202735 , n35457 );
buf ( n202736 , n202735 );
nand ( n35460 , n202731 , n202736 );
buf ( n202738 , n35460 );
buf ( n202739 , n202738 );
and ( n35463 , n35407 , n202739 );
and ( n35464 , n202679 , n202683 );
or ( n35465 , n35463 , n35464 );
buf ( n202743 , n35465 );
buf ( n202744 , n202743 );
xor ( n35468 , n202602 , n202744 );
xor ( n35469 , n201995 , n202234 );
xor ( n35470 , n35469 , n202272 );
buf ( n202748 , n35470 );
buf ( n202749 , n202748 );
and ( n35473 , n35468 , n202749 );
and ( n35474 , n202602 , n202744 );
or ( n35475 , n35473 , n35474 );
buf ( n202753 , n35475 );
nor ( n35477 , n202599 , n202753 );
xor ( n35478 , n202602 , n202744 );
xor ( n35479 , n35478 , n202749 );
buf ( n202757 , n35479 );
xor ( n35481 , n202104 , n202096 );
not ( n35482 , n202227 );
xor ( n35483 , n35481 , n35482 );
xor ( n35484 , n34760 , n34775 );
not ( n35485 , n202066 );
xor ( n35486 , n35484 , n35485 );
buf ( n202764 , n35486 );
xor ( n35488 , n202615 , n202628 );
xor ( n35489 , n35488 , n202640 );
buf ( n202767 , n35489 );
buf ( n202768 , n202767 );
xor ( n35492 , n202764 , n202768 );
xor ( n35493 , n196884 , n196904 );
and ( n35494 , n35493 , n196911 );
and ( n35495 , n196884 , n196904 );
or ( n35496 , n35494 , n35495 );
buf ( n202774 , n35496 );
buf ( n202775 , n202774 );
and ( n35499 , n35492 , n202775 );
and ( n35500 , n202764 , n202768 );
or ( n35501 , n35499 , n35500 );
buf ( n202779 , n35501 );
buf ( n202780 , n202779 );
xor ( n35504 , n202645 , n202649 );
xor ( n35505 , n35504 , n202674 );
buf ( n202783 , n35505 );
buf ( n202784 , n202783 );
xor ( n35508 , n202780 , n202784 );
xor ( n35509 , n202656 , n202662 );
xor ( n35510 , n35509 , n202669 );
buf ( n202788 , n35510 );
buf ( n202789 , n202788 );
xor ( n35513 , n196950 , n197005 );
and ( n35514 , n35513 , n197053 );
and ( n35515 , n196950 , n197005 );
or ( n35516 , n35514 , n35515 );
buf ( n202794 , n35516 );
buf ( n202795 , n202794 );
xor ( n35519 , n202789 , n202795 );
xor ( n35520 , n202699 , n202702 );
xor ( n35521 , n35520 , n202707 );
buf ( n202799 , n35521 );
buf ( n202800 , n202799 );
and ( n35524 , n35519 , n202800 );
and ( n35525 , n202789 , n202795 );
or ( n35526 , n35524 , n35525 );
buf ( n202804 , n35526 );
buf ( n202805 , n202804 );
and ( n35529 , n35508 , n202805 );
and ( n35530 , n202780 , n202784 );
or ( n35531 , n35529 , n35530 );
buf ( n202809 , n35531 );
xor ( n35533 , n35483 , n202809 );
xor ( n35534 , n202679 , n202683 );
xor ( n35535 , n35534 , n202739 );
buf ( n202813 , n35535 );
and ( n35537 , n35533 , n202813 );
and ( n35538 , n35483 , n202809 );
or ( n35539 , n35537 , n35538 );
nor ( n35540 , n202757 , n35539 );
nor ( n35541 , n35477 , n35540 );
xor ( n35542 , n35483 , n202809 );
xor ( n35543 , n35542 , n202813 );
xor ( n35544 , n202714 , n202719 );
xnor ( n35545 , n35544 , n35450 );
buf ( n202823 , n35545 );
xor ( n35547 , n197096 , n197151 );
and ( n35548 , n35547 , n197158 );
and ( n35549 , n197096 , n197151 );
or ( n35550 , n35548 , n35549 );
buf ( n202828 , n35550 );
xor ( n35552 , n202764 , n202768 );
xor ( n35553 , n35552 , n202775 );
buf ( n202831 , n35553 );
xor ( n35555 , n202828 , n202831 );
xor ( n35556 , n202789 , n202795 );
xor ( n35557 , n35556 , n202800 );
buf ( n202835 , n35557 );
and ( n35559 , n35555 , n202835 );
and ( n35560 , n202828 , n202831 );
or ( n35561 , n35559 , n35560 );
buf ( n202839 , n35561 );
xor ( n35563 , n202823 , n202839 );
xor ( n35564 , n202780 , n202784 );
xor ( n35565 , n35564 , n202805 );
buf ( n202843 , n35565 );
buf ( n202844 , n202843 );
and ( n35568 , n35563 , n202844 );
and ( n35569 , n202823 , n202839 );
or ( n35570 , n35568 , n35569 );
buf ( n202848 , n35570 );
nor ( n35572 , n35543 , n202848 );
xor ( n35573 , n202823 , n202839 );
xor ( n35574 , n35573 , n202844 );
buf ( n202852 , n35574 );
xor ( n35576 , n196914 , n196920 );
and ( n35577 , n35576 , n196927 );
and ( n35578 , n196914 , n196920 );
or ( n35579 , n35577 , n35578 );
buf ( n202857 , n35579 );
buf ( n35581 , n202857 );
not ( n35582 , n35581 );
not ( n35583 , n35582 );
xor ( n35584 , n197056 , n197161 );
and ( n35585 , n35584 , n197168 );
and ( n35586 , n197056 , n197161 );
or ( n35587 , n35585 , n35586 );
buf ( n202865 , n35587 );
not ( n35589 , n202865 );
not ( n35590 , n35589 );
or ( n35591 , n35583 , n35590 );
xor ( n35592 , n202828 , n202831 );
xor ( n35593 , n35592 , n202835 );
nand ( n35594 , n35591 , n35593 );
nand ( n35595 , n202865 , n35581 );
nand ( n35596 , n35594 , n35595 );
nor ( n35597 , n202852 , n35596 );
nor ( n35598 , n35572 , n35597 );
and ( n35599 , n35541 , n35598 );
nand ( n35600 , n35319 , n35599 );
xor ( n35601 , n195314 , n195591 );
xor ( n35602 , n35601 , n195873 );
buf ( n202880 , n35602 );
not ( n35604 , n202880 );
xor ( n35605 , n196015 , n196185 );
and ( n35606 , n35605 , n196207 );
and ( n35607 , n196015 , n196185 );
or ( n35608 , n35606 , n35607 );
buf ( n202886 , n35608 );
not ( n35610 , n202886 );
nand ( n35611 , n35604 , n35610 );
or ( n35612 , n196209 , n196298 );
nand ( n35613 , n35611 , n35612 );
not ( n35614 , n197182 );
not ( n35615 , n35614 );
xor ( n35616 , n202857 , n202865 );
xnor ( n35617 , n35616 , n35593 );
not ( n35618 , n35617 );
or ( n35619 , n35615 , n35618 );
xor ( n35620 , n196930 , n197171 );
xor ( n35621 , n35620 , n197178 );
buf ( n202899 , n35621 );
not ( n35623 , n202899 );
not ( n35624 , n195877 );
nand ( n35625 , n35623 , n35624 );
nand ( n35626 , n35619 , n35625 );
nor ( n35627 , n35613 , n35626 );
not ( n35628 , n35627 );
xor ( n35629 , n28988 , n28995 );
xnor ( n35630 , n35629 , n28983 );
buf ( n202908 , n35630 );
xor ( n35632 , n194192 , n194303 );
and ( n35633 , n35632 , n194358 );
and ( n35634 , n194192 , n194303 );
or ( n35635 , n35633 , n35634 );
buf ( n202913 , n35635 );
buf ( n202914 , n202913 );
xor ( n35638 , n202908 , n202914 );
xor ( n35639 , n194195 , n194243 );
and ( n35640 , n35639 , n194300 );
and ( n35641 , n194195 , n194243 );
or ( n35642 , n35640 , n35641 );
buf ( n202920 , n35642 );
buf ( n202921 , n202920 );
xor ( n35645 , n28944 , n28948 );
xor ( n35646 , n35645 , n196240 );
buf ( n202924 , n35646 );
xor ( n35648 , n202921 , n202924 );
not ( n35649 , n26587 );
not ( n35650 , n26473 );
or ( n35651 , n35649 , n35650 );
nand ( n35652 , n26519 , n26583 );
nand ( n35653 , n35651 , n35652 );
buf ( n202931 , n35653 );
xor ( n35655 , n35648 , n202931 );
buf ( n202933 , n35655 );
buf ( n202934 , n202933 );
and ( n35658 , n35638 , n202934 );
and ( n35659 , n202908 , n202914 );
or ( n35660 , n35658 , n35659 );
buf ( n202938 , n35660 );
xor ( n35662 , n196056 , n196060 );
xor ( n35663 , n35662 , n196076 );
buf ( n202941 , n35663 );
buf ( n202942 , n202941 );
xor ( n35666 , n202921 , n202924 );
and ( n35667 , n35666 , n202931 );
and ( n35668 , n202921 , n202924 );
or ( n35669 , n35667 , n35668 );
buf ( n202947 , n35669 );
buf ( n202948 , n202947 );
xor ( n35672 , n202942 , n202948 );
xor ( n35673 , n196244 , n196248 );
xor ( n35674 , n35673 , n196279 );
buf ( n202952 , n35674 );
buf ( n202953 , n202952 );
xor ( n35677 , n35672 , n202953 );
buf ( n202955 , n35677 );
nor ( n35679 , n202938 , n202955 );
xor ( n35680 , n196214 , n196284 );
xor ( n35681 , n35680 , n196294 );
buf ( n202959 , n35681 );
xor ( n35683 , n202942 , n202948 );
and ( n35684 , n35683 , n202953 );
and ( n35685 , n202942 , n202948 );
or ( n35686 , n35684 , n35685 );
buf ( n202964 , n35686 );
nor ( n35688 , n202959 , n202964 );
nor ( n35689 , n35679 , n35688 );
not ( n35690 , n35689 );
xor ( n35691 , n194368 , n194485 );
and ( n35692 , n35691 , n194490 );
and ( n35693 , n194368 , n194485 );
or ( n35694 , n35692 , n35693 );
buf ( n202972 , n35694 );
nand ( n35696 , n194363 , n202972 );
not ( n35697 , n35696 );
xor ( n35698 , n202908 , n202914 );
xor ( n35699 , n35698 , n202934 );
buf ( n202977 , n35699 );
xor ( n35701 , n193873 , n194185 );
and ( n35702 , n35701 , n194361 );
and ( n35703 , n193873 , n194185 );
or ( n35704 , n35702 , n35703 );
buf ( n202982 , n35704 );
nand ( n35706 , n202977 , n202982 );
not ( n35707 , n35706 );
or ( n35708 , n35697 , n35707 );
not ( n35709 , n202977 );
not ( n35710 , n202982 );
nand ( n35711 , n35709 , n35710 );
nand ( n35712 , n35708 , n35711 );
not ( n35713 , n35712 );
not ( n35714 , n35713 );
or ( n35715 , n35690 , n35714 );
not ( n35716 , n35688 );
nand ( n35717 , n202938 , n202955 );
not ( n35718 , n35717 );
and ( n35719 , n35716 , n35718 );
and ( n35720 , n202959 , n202964 );
nor ( n35721 , n35719 , n35720 );
nand ( n35722 , n35715 , n35721 );
not ( n35723 , n35722 );
or ( n35724 , n35628 , n35723 );
xor ( n35725 , n202857 , n202865 );
xor ( n35726 , n35725 , n35593 );
not ( n35727 , n35726 );
and ( n35728 , n35727 , n35614 );
nor ( n35729 , n202899 , n195877 );
nor ( n35730 , n35728 , n35729 );
not ( n35731 , n35730 );
not ( n35732 , n35611 );
and ( n35733 , n196209 , n196298 );
not ( n35734 , n35733 );
or ( n35735 , n35732 , n35734 );
not ( n35736 , n35604 );
not ( n35737 , n35610 );
nand ( n35738 , n35736 , n35737 );
nand ( n35739 , n35735 , n35738 );
not ( n35740 , n35739 );
or ( n35741 , n35731 , n35740 );
and ( n35742 , n202899 , n195877 );
nand ( n35743 , n35617 , n35614 );
and ( n35744 , n35742 , n35743 );
nand ( n35745 , n35726 , n197182 );
not ( n35746 , n35745 );
nor ( n35747 , n35744 , n35746 );
nand ( n35748 , n35741 , n35747 );
not ( n35749 , n35748 );
nand ( n35750 , n35724 , n35749 );
not ( n35751 , n35688 );
not ( n35752 , n202977 );
not ( n35753 , n202982 );
and ( n35754 , n35752 , n35753 );
nor ( n35755 , n194363 , n202972 );
nor ( n35756 , n35754 , n35755 );
not ( n35757 , n35679 );
and ( n35758 , n35751 , n35756 , n35757 );
not ( n35759 , n35613 );
xor ( n35760 , n194054 , n194122 );
xor ( n35761 , n35760 , n194175 );
buf ( n203039 , n35761 );
buf ( n203040 , n203039 );
xor ( n35764 , n194869 , n194873 );
and ( n35765 , n35764 , n194906 );
and ( n35766 , n194869 , n194873 );
or ( n35767 , n35765 , n35766 );
buf ( n203045 , n35767 );
buf ( n203046 , n203045 );
xor ( n35770 , n203040 , n203046 );
xor ( n35771 , n194372 , n194376 );
xor ( n35772 , n35771 , n194480 );
buf ( n203050 , n35772 );
buf ( n203051 , n203050 );
xor ( n35775 , n35770 , n203051 );
buf ( n203053 , n35775 );
not ( n35777 , n203053 );
xor ( n35778 , n194828 , n194855 );
and ( n35779 , n35778 , n194909 );
and ( n35780 , n194828 , n194855 );
or ( n35781 , n35779 , n35780 );
buf ( n203059 , n35781 );
not ( n35783 , n203059 );
and ( n35784 , n35777 , n35783 );
xor ( n35785 , n194888 , n194894 );
xor ( n35786 , n35785 , n194901 );
buf ( n203064 , n35786 );
buf ( n203065 , n203064 );
xor ( n35789 , n194568 , n194583 );
and ( n35790 , n35789 , n194627 );
and ( n35791 , n194568 , n194583 );
or ( n35792 , n35790 , n35791 );
buf ( n203070 , n35792 );
buf ( n203071 , n203070 );
xor ( n35795 , n203065 , n203071 );
xor ( n35796 , n194832 , n194836 );
xor ( n35797 , n35796 , n194850 );
buf ( n203075 , n35797 );
buf ( n203076 , n203075 );
and ( n35800 , n35795 , n203076 );
and ( n35801 , n203065 , n203071 );
or ( n35802 , n35800 , n35801 );
buf ( n203080 , n35802 );
not ( n35804 , n203080 );
not ( n35805 , n35804 );
not ( n35806 , n194911 );
not ( n35807 , n35806 );
or ( n35808 , n35805 , n35807 );
xor ( n35809 , n203065 , n203071 );
xor ( n35810 , n35809 , n203076 );
buf ( n203088 , n35810 );
xor ( n35812 , n194562 , n194630 );
and ( n35813 , n35812 , n194637 );
and ( n35814 , n194562 , n194630 );
or ( n35815 , n35813 , n35814 );
buf ( n203093 , n35815 );
or ( n35817 , n203088 , n203093 );
nand ( n35818 , n35808 , n35817 );
nor ( n35819 , n35784 , n35818 );
not ( n35820 , n194639 );
xor ( n35821 , n190394 , n190533 );
and ( n35822 , n35821 , n190646 );
and ( n35823 , n190394 , n190533 );
or ( n35824 , n35822 , n35823 );
buf ( n203102 , n35824 );
not ( n35826 , n203102 );
nand ( n35827 , n35820 , n35826 );
buf ( n35828 , n35827 );
buf ( n203106 , n20902 );
buf ( n203107 , n863 );
and ( n35831 , n203106 , n203107 );
buf ( n203109 , n35831 );
buf ( n203110 , n203109 );
buf ( n203111 , n194807 );
not ( n35835 , n203111 );
buf ( n203113 , n21330 );
not ( n35837 , n203113 );
or ( n35838 , n35835 , n35837 );
buf ( n203116 , n859 );
buf ( n203117 , n894 );
xor ( n35841 , n203116 , n203117 );
buf ( n203119 , n35841 );
buf ( n203120 , n203119 );
buf ( n203121 , n895 );
nand ( n35845 , n203120 , n203121 );
buf ( n203123 , n35845 );
buf ( n203124 , n203123 );
nand ( n35848 , n35838 , n203124 );
buf ( n203126 , n35848 );
buf ( n203127 , n203126 );
xor ( n35851 , n203110 , n203127 );
buf ( n203129 , n862 );
buf ( n203130 , n892 );
xor ( n35854 , n203129 , n203130 );
buf ( n203132 , n35854 );
buf ( n203133 , n203132 );
not ( n35857 , n203133 );
buf ( n203135 , n190485 );
not ( n35859 , n203135 );
or ( n35860 , n35857 , n35859 );
buf ( n203138 , n190491 );
buf ( n203139 , n861 );
buf ( n203140 , n892 );
xor ( n35864 , n203139 , n203140 );
buf ( n203142 , n35864 );
buf ( n203143 , n203142 );
nand ( n35867 , n203138 , n203143 );
buf ( n203145 , n35867 );
buf ( n203146 , n203145 );
nand ( n35870 , n35860 , n203146 );
buf ( n203148 , n35870 );
buf ( n203149 , n203148 );
xor ( n35873 , n35851 , n203149 );
buf ( n203151 , n35873 );
and ( n35875 , n194794 , n194815 );
buf ( n203153 , n35875 );
nand ( n35877 , n203151 , n203153 );
not ( n35878 , n35877 );
not ( n35879 , n35878 );
buf ( n203157 , n203142 );
not ( n35881 , n203157 );
buf ( n203159 , n190485 );
not ( n35883 , n203159 );
or ( n35884 , n35881 , n35883 );
buf ( n203162 , n190491 );
buf ( n203163 , n860 );
buf ( n203164 , n892 );
xor ( n35888 , n203163 , n203164 );
buf ( n203166 , n35888 );
buf ( n203167 , n203166 );
nand ( n35891 , n203162 , n203167 );
buf ( n203169 , n35891 );
buf ( n203170 , n203169 );
nand ( n35894 , n35884 , n203170 );
buf ( n203172 , n35894 );
buf ( n203173 , n203172 );
buf ( n203174 , n863 );
buf ( n203175 , n890 );
xor ( n35899 , n203174 , n203175 );
buf ( n203177 , n35899 );
buf ( n203178 , n203177 );
not ( n35902 , n203178 );
buf ( n203180 , n188751 );
not ( n35904 , n203180 );
or ( n35905 , n35902 , n35904 );
buf ( n203183 , n20902 );
buf ( n203184 , n862 );
buf ( n203185 , n890 );
xor ( n35909 , n203184 , n203185 );
buf ( n203187 , n35909 );
buf ( n203188 , n203187 );
nand ( n35912 , n203183 , n203188 );
buf ( n203190 , n35912 );
buf ( n203191 , n203190 );
nand ( n35915 , n35905 , n203191 );
buf ( n203193 , n35915 );
buf ( n203194 , n203193 );
xor ( n35918 , n203173 , n203194 );
not ( n35919 , n203119 );
not ( n35920 , n21330 );
or ( n35921 , n35919 , n35920 );
buf ( n203199 , n858 );
buf ( n203200 , n894 );
xor ( n35924 , n203199 , n203200 );
buf ( n203202 , n35924 );
buf ( n203203 , n203202 );
buf ( n203204 , n895 );
nand ( n35928 , n203203 , n203204 );
buf ( n203206 , n35928 );
nand ( n35930 , n35921 , n203206 );
buf ( n203208 , n863 );
buf ( n203209 , n891 );
or ( n35933 , n203208 , n203209 );
buf ( n203211 , n892 );
nand ( n35935 , n35933 , n203211 );
buf ( n203213 , n35935 );
buf ( n203214 , n863 );
buf ( n203215 , n891 );
nand ( n35939 , n203214 , n203215 );
buf ( n203217 , n35939 );
nand ( n35941 , n203213 , n203217 , n890 );
not ( n35942 , n35941 );
and ( n35943 , n35930 , n35942 );
not ( n35944 , n35930 );
and ( n35945 , n35944 , n35941 );
nor ( n35946 , n35943 , n35945 );
buf ( n203224 , n35946 );
xor ( n35948 , n35918 , n203224 );
buf ( n203226 , n35948 );
not ( n35950 , n203226 );
xor ( n35951 , n203110 , n203127 );
and ( n35952 , n35951 , n203149 );
and ( n35953 , n203110 , n203127 );
or ( n35954 , n35952 , n35953 );
buf ( n203232 , n35954 );
not ( n35956 , n203232 );
nand ( n35957 , n35950 , n35956 );
not ( n35958 , n35957 );
or ( n35959 , n35879 , n35958 );
nand ( n35960 , n203226 , n203232 );
nand ( n35961 , n35959 , n35960 );
not ( n35962 , n203226 );
nand ( n35963 , n35962 , n35956 );
buf ( n203241 , n863 );
buf ( n203242 , n892 );
xor ( n35966 , n203241 , n203242 );
buf ( n203244 , n35966 );
buf ( n203245 , n203244 );
not ( n35969 , n203245 );
buf ( n203247 , n20632 );
not ( n35971 , n203247 );
or ( n35972 , n35969 , n35971 );
buf ( n203250 , n190491 );
buf ( n203251 , n203132 );
nand ( n35975 , n203250 , n203251 );
buf ( n203253 , n35975 );
buf ( n203254 , n203253 );
nand ( n35978 , n35972 , n203254 );
buf ( n203256 , n35978 );
nand ( n35980 , n194817 , n203256 );
buf ( n203258 , n196308 );
not ( n35982 , n203258 );
buf ( n203260 , n22809 );
not ( n35984 , n203260 );
or ( n35985 , n35982 , n35984 );
buf ( n203263 , n194798 );
buf ( n203264 , n895 );
nand ( n35988 , n203263 , n203264 );
buf ( n203266 , n35988 );
buf ( n203267 , n203266 );
nand ( n35991 , n35985 , n203267 );
buf ( n203269 , n35991 );
buf ( n203270 , n190491 );
buf ( n203271 , n863 );
and ( n35995 , n203270 , n203271 );
buf ( n203273 , n35995 );
nor ( n35997 , n203269 , n203273 );
buf ( n203275 , n863 );
buf ( n203276 , n895 );
nand ( n36000 , n203275 , n203276 );
buf ( n203278 , n36000 );
buf ( n203279 , n203278 );
buf ( n203280 , n894 );
and ( n36004 , n203279 , n203280 );
buf ( n203282 , n36004 );
nand ( n36006 , n203282 , n196315 );
nor ( n36007 , n35997 , n36006 );
and ( n36008 , n203269 , n203273 );
or ( n36009 , n36007 , n36008 );
or ( n36010 , n203256 , n194817 );
nand ( n36011 , n36009 , n36010 );
nand ( n36012 , n35980 , n36011 );
or ( n36013 , n203151 , n203153 );
nand ( n36014 , n35963 , n36012 , n36013 );
not ( n36015 , n36014 );
or ( n36016 , n35961 , n36015 );
buf ( n203294 , n863 );
buf ( n203295 , n20396 );
nand ( n36019 , n203294 , n203295 );
buf ( n203297 , n36019 );
buf ( n203298 , n203297 );
not ( n36022 , n203298 );
buf ( n203300 , n36022 );
buf ( n203301 , n203300 );
not ( n36025 , n203301 );
buf ( n203303 , n203202 );
not ( n36027 , n203303 );
buf ( n203305 , n23321 );
not ( n36029 , n203305 );
or ( n36030 , n36027 , n36029 );
buf ( n203308 , n194734 );
buf ( n203309 , n895 );
nand ( n36033 , n203308 , n203309 );
buf ( n203311 , n36033 );
buf ( n203312 , n203311 );
nand ( n36036 , n36030 , n203312 );
buf ( n203314 , n36036 );
buf ( n203315 , n203314 );
not ( n36039 , n203315 );
or ( n36040 , n36025 , n36039 );
buf ( n203318 , n203314 );
not ( n36042 , n203318 );
buf ( n203320 , n36042 );
buf ( n203321 , n203320 );
not ( n36045 , n203321 );
buf ( n203323 , n203297 );
not ( n36047 , n203323 );
or ( n36048 , n36045 , n36047 );
buf ( n203326 , n203166 );
not ( n36050 , n203326 );
buf ( n203328 , n190485 );
not ( n36052 , n203328 );
or ( n36053 , n36050 , n36052 );
buf ( n203331 , n190491 );
buf ( n203332 , n194644 );
nand ( n36056 , n203331 , n203332 );
buf ( n203334 , n36056 );
buf ( n203335 , n203334 );
nand ( n36059 , n36053 , n203335 );
buf ( n203337 , n36059 );
buf ( n203338 , n203337 );
nand ( n36062 , n36048 , n203338 );
buf ( n203340 , n36062 );
buf ( n203341 , n203340 );
nand ( n36065 , n36040 , n203341 );
buf ( n203343 , n36065 );
buf ( n203344 , n203343 );
not ( n36068 , n203344 );
buf ( n203346 , n194746 );
buf ( n203347 , n194762 );
and ( n36071 , n203346 , n203347 );
not ( n36072 , n203346 );
buf ( n203350 , n194765 );
and ( n36074 , n36072 , n203350 );
nor ( n36075 , n36071 , n36074 );
buf ( n203353 , n36075 );
buf ( n203354 , n203353 );
not ( n36078 , n203354 );
and ( n36079 , n36068 , n36078 );
buf ( n203357 , n203343 );
buf ( n203358 , n203353 );
and ( n36082 , n203357 , n203358 );
nor ( n36083 , n36079 , n36082 );
buf ( n203361 , n36083 );
xor ( n36085 , n27379 , n27395 );
xor ( n36086 , n36085 , n27409 );
xnor ( n36087 , n203361 , n36086 );
not ( n36088 , n36087 );
buf ( n203366 , n203187 );
not ( n36090 , n203366 );
buf ( n203368 , n188751 );
not ( n36092 , n203368 );
or ( n36093 , n36090 , n36092 );
buf ( n203371 , n20902 );
buf ( n203372 , n194660 );
nand ( n36096 , n203371 , n203372 );
buf ( n203374 , n36096 );
buf ( n203375 , n203374 );
nand ( n36099 , n36093 , n203375 );
buf ( n203377 , n36099 );
buf ( n203378 , n203377 );
not ( n36102 , n203378 );
buf ( n203380 , n36102 );
nand ( n36104 , n35930 , n35942 );
nand ( n36105 , n203380 , n36104 );
buf ( n203383 , n36105 );
not ( n36107 , n203383 );
xor ( n36108 , n203300 , n203320 );
xor ( n36109 , n36108 , n203337 );
buf ( n203387 , n36109 );
not ( n36111 , n203387 );
buf ( n203389 , n36111 );
buf ( n203390 , n203389 );
not ( n36114 , n203390 );
or ( n36115 , n36107 , n36114 );
not ( n36116 , n36104 );
nand ( n36117 , n36116 , n203377 );
buf ( n203395 , n36117 );
nand ( n36119 , n36115 , n203395 );
buf ( n203397 , n36119 );
not ( n36121 , n203397 );
nand ( n36122 , n36088 , n36121 );
and ( n36123 , n36104 , n203380 );
not ( n36124 , n36104 );
and ( n36125 , n36124 , n203377 );
nor ( n36126 , n36123 , n36125 );
buf ( n203404 , n36126 );
not ( n36128 , n203404 );
buf ( n203406 , n36128 );
buf ( n203407 , n203406 );
not ( n36131 , n203407 );
buf ( n203409 , n203389 );
not ( n36133 , n203409 );
or ( n36134 , n36131 , n36133 );
buf ( n203412 , n36109 );
buf ( n203413 , n36126 );
nand ( n36137 , n203412 , n203413 );
buf ( n203415 , n36137 );
buf ( n203416 , n203415 );
nand ( n36140 , n36134 , n203416 );
buf ( n203418 , n36140 );
not ( n36142 , n203418 );
xor ( n36143 , n203173 , n203194 );
and ( n36144 , n36143 , n203224 );
and ( n36145 , n203173 , n203194 );
or ( n36146 , n36144 , n36145 );
buf ( n203424 , n36146 );
not ( n36148 , n203424 );
nand ( n36149 , n36142 , n36148 );
nand ( n36150 , n36016 , n36122 , n36149 );
nand ( n36151 , n203418 , n203424 );
not ( n36152 , n36151 );
or ( n36153 , n36087 , n203397 );
and ( n36154 , n36152 , n36153 );
nand ( n36155 , n36087 , n203397 );
not ( n36156 , n36155 );
nor ( n36157 , n36154 , n36156 );
nand ( n36158 , n36150 , n36157 );
buf ( n203436 , n194717 );
buf ( n203437 , n194771 );
or ( n36161 , n203436 , n203437 );
buf ( n203439 , n194729 );
nand ( n36163 , n36161 , n203439 );
buf ( n203441 , n36163 );
buf ( n203442 , n203441 );
buf ( n203443 , n194717 );
buf ( n203444 , n194771 );
nand ( n36168 , n203443 , n203444 );
buf ( n203446 , n36168 );
buf ( n203447 , n203446 );
nand ( n36171 , n203442 , n203447 );
buf ( n203449 , n36171 );
buf ( n203450 , n203449 );
xor ( n36174 , n190609 , n190622 );
xor ( n36175 , n36174 , n190638 );
buf ( n203453 , n36175 );
buf ( n203454 , n203453 );
xor ( n36178 , n203450 , n203454 );
xor ( n36179 , n190412 , n190475 );
xor ( n36180 , n36179 , n190528 );
buf ( n203458 , n36180 );
buf ( n203459 , n203458 );
and ( n36183 , n36178 , n203459 );
and ( n36184 , n203450 , n203454 );
or ( n36185 , n36183 , n36184 );
buf ( n203463 , n36185 );
not ( n36187 , n203463 );
not ( n36188 , n190648 );
nand ( n36189 , n36187 , n36188 );
xor ( n36190 , n203450 , n203454 );
xor ( n36191 , n36190 , n203459 );
buf ( n203469 , n36191 );
not ( n36193 , n27427 );
not ( n36194 , n27498 );
or ( n36195 , n36193 , n36194 );
nand ( n36196 , n36195 , n27412 );
or ( n36197 , n27498 , n27427 );
nand ( n36198 , n36196 , n36197 );
nor ( n36199 , n203469 , n36198 );
buf ( n203477 , n203343 );
not ( n36201 , n203477 );
buf ( n203479 , n203353 );
nand ( n36203 , n36201 , n203479 );
buf ( n203481 , n36203 );
buf ( n203482 , n203481 );
not ( n36206 , n203482 );
buf ( n203484 , n36086 );
not ( n36208 , n203484 );
or ( n36209 , n36206 , n36208 );
buf ( n203487 , n203353 );
not ( n36211 , n203487 );
buf ( n203489 , n203343 );
nand ( n36213 , n36211 , n203489 );
buf ( n203491 , n36213 );
buf ( n203492 , n203491 );
nand ( n36216 , n36209 , n203492 );
buf ( n203494 , n36216 );
nor ( n36218 , n27500 , n203494 );
nor ( n36219 , n36199 , n36218 );
and ( n36220 , n35828 , n36158 , n36189 , n36219 );
xor ( n36221 , n203040 , n203046 );
and ( n36222 , n36221 , n203051 );
and ( n36223 , n203040 , n203046 );
or ( n36224 , n36222 , n36223 );
buf ( n203502 , n36224 );
or ( n36226 , n194492 , n203502 );
nand ( n36227 , n35819 , n36220 , n36226 );
nor ( n36228 , n194492 , n203502 );
nor ( n36229 , n203053 , n203059 );
nor ( n36230 , n36228 , n36229 );
nand ( n36231 , n203088 , n203093 );
not ( n36232 , n36231 );
not ( n36233 , n36232 );
nand ( n36234 , n35806 , n35804 );
not ( n36235 , n36234 );
or ( n36236 , n36233 , n36235 );
nand ( n36237 , n194911 , n203080 );
nand ( n36238 , n36236 , n36237 );
and ( n36239 , n36230 , n36238 );
nand ( n36240 , n203053 , n203059 );
or ( n36241 , n36228 , n36240 );
nand ( n36242 , n194492 , n203502 );
nand ( n36243 , n36241 , n36242 );
nor ( n36244 , n36239 , n36243 );
nand ( n36245 , n27500 , n203494 );
nor ( n36246 , n203469 , n36198 );
or ( n36247 , n36245 , n36246 );
nand ( n36248 , n203469 , n36198 );
nand ( n36249 , n36247 , n36248 );
not ( n36250 , n36249 );
not ( n36251 , n203463 );
nand ( n36252 , n36251 , n36188 );
and ( n36253 , n35827 , n36252 );
not ( n36254 , n36253 );
or ( n36255 , n36250 , n36254 );
nand ( n36256 , n190648 , n203463 );
not ( n36257 , n36256 );
not ( n36258 , n36257 );
not ( n36259 , n35827 );
or ( n36260 , n36258 , n36259 );
not ( n36261 , n35820 );
nand ( n36262 , n36261 , n203102 );
nand ( n36263 , n36260 , n36262 );
not ( n36264 , n36263 );
nand ( n36265 , n36255 , n36264 );
not ( n36266 , n35818 );
nand ( n36267 , n36265 , n36230 , n36266 );
nand ( n36268 , n36227 , n36244 , n36267 );
and ( n36269 , n35758 , n35759 , n36268 , n35730 );
nor ( n36270 , n35750 , n36269 );
or ( n36271 , n35600 , n36270 );
nand ( n36272 , n202852 , n35596 );
nand ( n36273 , n35543 , n202848 );
nand ( n36274 , n36272 , n36273 );
not ( n36275 , n35539 );
not ( n36276 , n202757 );
nand ( n36277 , n36275 , n36276 );
nand ( n36278 , n36274 , n36277 );
not ( n36279 , n36278 );
not ( n36280 , n36279 );
nor ( n36281 , n35477 , n35572 );
not ( n36282 , n36281 );
or ( n36283 , n36280 , n36282 );
nand ( n36284 , n202757 , n35539 );
not ( n36285 , n36284 );
not ( n36286 , n36285 );
not ( n36287 , n202599 );
not ( n36288 , n202753 );
nand ( n36289 , n36287 , n36288 );
not ( n36290 , n36289 );
or ( n36291 , n36286 , n36290 );
nand ( n36292 , n202599 , n202753 );
nand ( n36293 , n36291 , n36292 );
not ( n36294 , n36293 );
nand ( n36295 , n36283 , n36294 );
and ( n36296 , n35319 , n36295 );
not ( n36297 , n35317 );
not ( n36298 , n202416 );
nor ( n36299 , n36298 , n35227 );
not ( n36300 , n36299 );
not ( n36301 , n35282 );
or ( n36302 , n36300 , n36301 );
not ( n36303 , n35281 );
buf ( n36304 , n202551 );
nand ( n36305 , n36303 , n36304 );
nand ( n36306 , n36302 , n36305 );
not ( n36307 , n36306 );
or ( n36308 , n36297 , n36307 );
and ( n36309 , n202583 , n202566 );
not ( n36310 , n202587 );
not ( n36311 , n202592 );
nand ( n36312 , n36310 , n36311 );
and ( n36313 , n36309 , n36312 );
and ( n36314 , n202587 , n202592 );
nor ( n36315 , n36313 , n36314 );
nand ( n36316 , n36308 , n36315 );
nor ( n36317 , n36296 , n36316 );
nand ( n36318 , n36271 , n36317 );
buf ( n36319 , n36318 );
buf ( n36320 , n36319 );
and ( n36321 , n34128 , n36320 );
not ( n36322 , n32871 );
not ( n36323 , n36322 );
not ( n36324 , n32806 );
not ( n36325 , n36324 );
nand ( n36326 , n32538 , n187405 );
nor ( n36327 , n199823 , n193688 );
or ( n36328 , n36326 , n36327 );
nand ( n36329 , n199823 , n193688 );
nand ( n36330 , n36328 , n36329 );
not ( n36331 , n36330 );
or ( n36332 , n36325 , n36331 );
and ( n36333 , n199832 , n199998 );
and ( n36334 , n32805 , n36333 );
not ( n36335 , n200074 );
nor ( n36336 , n36335 , n32804 );
nor ( n36337 , n36334 , n36336 );
nand ( n36338 , n36332 , n36337 );
not ( n36339 , n36338 );
not ( n36340 , n36339 );
not ( n36341 , n36340 );
or ( n36342 , n36323 , n36341 );
nand ( n36343 , n200141 , n200146 );
not ( n36344 , n36343 );
not ( n36345 , n36344 );
not ( n36346 , n32861 );
or ( n36347 , n36345 , n36346 );
nand ( n36348 , n200120 , n200137 );
nand ( n36349 , n36347 , n36348 );
not ( n36350 , n36349 );
nand ( n36351 , n36342 , n36350 );
nor ( n36352 , n36321 , n36351 );
nand ( n36353 , n34104 , n36352 );
not ( n36354 , n196880 );
xor ( n36355 , n200124 , n200128 );
and ( n36356 , n36355 , n200135 );
and ( n36357 , n200124 , n200128 );
or ( n36358 , n36356 , n36357 );
buf ( n203636 , n36358 );
not ( n36360 , n203636 );
nand ( n36361 , n36354 , n36360 );
not ( n36362 , n196880 );
nor ( n36363 , n36362 , n36360 );
not ( n36364 , n36363 );
nand ( n36365 , n36361 , n36364 );
not ( n36366 , n36365 );
and ( n36367 , n36353 , n36366 );
not ( n36368 , n36353 );
and ( n36369 , n36368 , n36365 );
nor ( n36370 , n36367 , n36369 );
not ( n36371 , n34126 );
not ( n36372 , n32808 );
and ( n36373 , n36371 , n36372 );
buf ( n36374 , n36319 );
and ( n36375 , n36373 , n36374 );
nor ( n36376 , n36375 , n36340 );
not ( n36377 , n32808 );
not ( n36378 , n33604 );
nand ( n36379 , n34081 , n34095 , n34100 );
nand ( n36380 , n36378 , n36379 );
nand ( n36381 , n36377 , n36380 );
nand ( n36382 , n36376 , n36381 );
not ( n36383 , n32870 );
or ( n36384 , n36344 , n36383 );
not ( n36385 , n36384 );
and ( n36386 , n36382 , n36385 );
not ( n36387 , n36382 );
and ( n36388 , n36387 , n36384 );
nor ( n36389 , n36386 , n36388 );
not ( n36390 , n34109 );
nor ( n36391 , n36390 , n34091 );
not ( n36392 , n36391 );
not ( n36393 , n36319 );
or ( n36394 , n36392 , n36393 );
buf ( n36395 , n34116 );
not ( n36396 , n36395 );
not ( n36397 , n34020 );
not ( n36398 , n36397 );
nand ( n36399 , n34013 , n36398 );
not ( n36400 , n36399 );
or ( n36401 , n36396 , n36400 );
buf ( n36402 , n34019 );
nand ( n36403 , n36401 , n36402 );
not ( n36404 , n36403 );
nand ( n36405 , n36394 , n36404 );
buf ( n36406 , n34034 );
nand ( n36407 , n34113 , n36406 );
nand ( n36408 , n36405 , n36407 );
nor ( n36409 , n32808 , n36383 );
not ( n36410 , n36409 );
not ( n36411 , n36380 );
or ( n36412 , n36410 , n36411 );
not ( n36413 , n36319 );
buf ( n36414 , n34125 );
nand ( n36415 , n36414 , n36409 );
nor ( n36416 , n36413 , n36415 );
not ( n36417 , n32870 );
not ( n36418 , n36338 );
or ( n36419 , n36417 , n36418 );
nand ( n36420 , n36419 , n36343 );
nor ( n36421 , n36416 , n36420 );
nand ( n36422 , n36412 , n36421 );
xor ( n36423 , n196500 , n196690 );
and ( n36424 , n36423 , n196878 );
and ( n36425 , n196500 , n196690 );
or ( n36426 , n36424 , n36425 );
buf ( n203704 , n36426 );
xor ( n36428 , n196383 , n196440 );
and ( n36429 , n36428 , n196497 );
and ( n36430 , n196383 , n196440 );
or ( n36431 , n36429 , n36430 );
buf ( n203709 , n36431 );
buf ( n203710 , n203709 );
xor ( n36434 , n196503 , n196520 );
and ( n36435 , n36434 , n196541 );
and ( n36436 , n196503 , n196520 );
or ( n36437 , n36435 , n36436 );
buf ( n203715 , n36437 );
buf ( n203716 , n203715 );
buf ( n203717 , n196457 );
not ( n36441 , n203717 );
buf ( n203719 , n196449 );
not ( n36443 , n203719 );
or ( n36444 , n36441 , n36443 );
buf ( n203722 , n186254 );
xor ( n36446 , n866 , n836 );
buf ( n203724 , n36446 );
nand ( n36448 , n203722 , n203724 );
buf ( n203726 , n36448 );
buf ( n203727 , n203726 );
nand ( n36451 , n36444 , n203727 );
buf ( n203729 , n36451 );
buf ( n203730 , n203729 );
not ( n36454 , n186539 );
buf ( n203732 , n19265 );
not ( n36456 , n203732 );
buf ( n203734 , n36456 );
not ( n36458 , n203734 );
or ( n36459 , n36454 , n36458 );
nand ( n36460 , n36459 , n872 );
buf ( n203738 , n36460 );
xor ( n36462 , n203730 , n203738 );
buf ( n203740 , n196531 );
not ( n36464 , n203740 );
buf ( n203742 , n186435 );
not ( n36466 , n203742 );
or ( n36467 , n36464 , n36466 );
buf ( n203745 , n186444 );
buf ( n203746 , n832 );
buf ( n203747 , n870 );
xor ( n36471 , n203746 , n203747 );
buf ( n203749 , n36471 );
buf ( n203750 , n203749 );
nand ( n36474 , n203745 , n203750 );
buf ( n203752 , n36474 );
buf ( n203753 , n203752 );
nand ( n36477 , n36467 , n203753 );
buf ( n203755 , n36477 );
buf ( n203756 , n203755 );
xor ( n36480 , n36462 , n203756 );
buf ( n203758 , n36480 );
buf ( n203759 , n203758 );
xor ( n36483 , n203716 , n203759 );
buf ( n203761 , n196537 );
buf ( n203762 , n196493 );
buf ( n203763 , n196463 );
or ( n36487 , n203762 , n203763 );
buf ( n203765 , n196475 );
nand ( n36489 , n36487 , n203765 );
buf ( n203767 , n36489 );
buf ( n203768 , n203767 );
buf ( n203769 , n196493 );
buf ( n203770 , n196463 );
nand ( n36494 , n203769 , n203770 );
buf ( n203772 , n36494 );
buf ( n203773 , n203772 );
nand ( n36497 , n203768 , n203773 );
buf ( n203775 , n36497 );
buf ( n203776 , n203775 );
xor ( n36500 , n203761 , n203776 );
and ( n36501 , n196368 , n196369 );
buf ( n203779 , n36501 );
buf ( n203780 , n203779 );
buf ( n203781 , n196487 );
not ( n36505 , n203781 );
buf ( n203783 , n186640 );
not ( n36507 , n203783 );
or ( n36508 , n36505 , n36507 );
buf ( n203786 , n186340 );
buf ( n203787 , n864 );
buf ( n203788 , n838 );
xor ( n36512 , n203787 , n203788 );
buf ( n203790 , n36512 );
buf ( n203791 , n203790 );
nand ( n36515 , n203786 , n203791 );
buf ( n203793 , n36515 );
buf ( n203794 , n203793 );
nand ( n36518 , n36508 , n203794 );
buf ( n203796 , n36518 );
buf ( n203797 , n203796 );
xor ( n36521 , n203780 , n203797 );
buf ( n203799 , n196513 );
not ( n36523 , n203799 );
buf ( n203801 , n186197 );
not ( n36525 , n203801 );
or ( n36526 , n36523 , n36525 );
buf ( n203804 , n186208 );
buf ( n203805 , n834 );
buf ( n203806 , n868 );
xor ( n36530 , n203805 , n203806 );
buf ( n203808 , n36530 );
buf ( n203809 , n203808 );
nand ( n36533 , n203804 , n203809 );
buf ( n203811 , n36533 );
buf ( n203812 , n203811 );
nand ( n36536 , n36526 , n203812 );
buf ( n203814 , n36536 );
buf ( n203815 , n203814 );
xor ( n36539 , n36521 , n203815 );
buf ( n203817 , n36539 );
buf ( n203818 , n203817 );
xor ( n36542 , n36500 , n203818 );
buf ( n203820 , n36542 );
buf ( n203821 , n203820 );
xor ( n36545 , n36483 , n203821 );
buf ( n203823 , n36545 );
buf ( n203824 , n203823 );
xor ( n36548 , n203710 , n203824 );
xor ( n36549 , n196544 , n196629 );
and ( n36550 , n36549 , n196687 );
and ( n36551 , n196544 , n196629 );
or ( n36552 , n36550 , n36551 );
buf ( n203830 , n36552 );
buf ( n203831 , n203830 );
xor ( n36555 , n36548 , n203831 );
buf ( n203833 , n36555 );
or ( n36557 , n203704 , n203833 );
nand ( n36558 , n36361 , n36557 );
nor ( n36559 , n32871 , n36558 );
and ( n36560 , n32807 , n36559 );
buf ( n36561 , n36560 );
not ( n36562 , n36561 );
not ( n36563 , n34102 );
or ( n36564 , n36562 , n36563 );
nand ( n36565 , n36414 , n36560 );
nor ( n36566 , n36565 , n36413 );
not ( n36567 , n36559 );
not ( n36568 , n36338 );
or ( n36569 , n36567 , n36568 );
not ( n36570 , n36558 );
not ( n36571 , n36570 );
not ( n36572 , n36349 );
or ( n36573 , n36571 , n36572 );
and ( n36574 , n36363 , n36557 );
and ( n36575 , n203704 , n203833 );
nor ( n36576 , n36574 , n36575 );
nand ( n36577 , n36573 , n36576 );
not ( n36578 , n36577 );
nand ( n36579 , n36569 , n36578 );
buf ( n36580 , n36579 );
nor ( n36581 , n36566 , n36580 );
nand ( n36582 , n36564 , n36581 );
buf ( n36583 , n34108 );
not ( n36584 , n36583 );
not ( n36585 , n36584 );
not ( n36586 , n36319 );
or ( n36587 , n36585 , n36586 );
not ( n36588 , n34012 );
nand ( n36589 , n36587 , n36588 );
and ( n36590 , n34098 , n33347 );
not ( n36591 , n36590 );
not ( n36592 , n34124 );
not ( n36593 , n36592 );
nor ( n36594 , n36591 , n36593 );
not ( n36595 , n36594 );
not ( n36596 , n36319 );
or ( n36597 , n36595 , n36596 );
not ( n36598 , n36590 );
buf ( n36599 , n34123 );
not ( n36600 , n36599 );
and ( n36601 , n34035 , n34093 );
not ( n36602 , n36601 );
or ( n36603 , n36600 , n36602 );
not ( n36604 , n33649 );
not ( n36605 , n34069 );
or ( n36606 , n36604 , n36605 );
nand ( n36607 , n36606 , n34080 );
not ( n36608 , n36607 );
nand ( n36609 , n36603 , n36608 );
not ( n36610 , n36609 );
or ( n36611 , n36598 , n36610 );
buf ( n36612 , n33585 );
not ( n36613 , n200567 );
buf ( n36614 , n33346 );
nand ( n36615 , n36613 , n36614 );
and ( n36616 , n36612 , n36615 );
buf ( n36617 , n33592 );
not ( n36618 , n36617 );
nor ( n36619 , n36616 , n36618 );
nand ( n36620 , n36611 , n36619 );
not ( n36621 , n36620 );
nand ( n36622 , n36597 , n36621 );
buf ( n36623 , n34097 );
nor ( n36624 , n36593 , n36623 );
not ( n36625 , n36624 );
not ( n36626 , n36374 );
or ( n36627 , n36625 , n36626 );
not ( n36628 , n36623 );
not ( n36629 , n36628 );
not ( n36630 , n36599 );
not ( n36631 , n36601 );
or ( n36632 , n36630 , n36631 );
nand ( n36633 , n36632 , n36608 );
not ( n36634 , n36633 );
or ( n36635 , n36629 , n36634 );
buf ( n36636 , n33574 );
not ( n36637 , n36636 );
nand ( n36638 , n36635 , n36637 );
not ( n36639 , n36638 );
nand ( n36640 , n36627 , n36639 );
not ( n36641 , n36405 );
not ( n36642 , n36281 );
not ( n36643 , n36279 );
or ( n36644 , n36642 , n36643 );
nand ( n36645 , n36644 , n36294 );
not ( n36646 , n36645 );
not ( n36647 , n35750 );
not ( n36648 , n36647 );
not ( n36649 , n35599 );
not ( n36650 , n36649 );
nand ( n36651 , n36648 , n36650 );
not ( n36652 , n35758 );
not ( n36653 , n36652 );
not ( n36654 , n35759 );
not ( n36655 , n36654 );
buf ( n36656 , n35730 );
nand ( n36657 , n36653 , n36655 , n36656 );
not ( n36658 , n36657 );
buf ( n36659 , n36268 );
buf ( n36660 , n36659 );
nand ( n36661 , n36658 , n36650 , n36660 );
nand ( n36662 , n36646 , n36651 , n36661 );
buf ( n36663 , n35228 );
not ( n36664 , n36299 );
nand ( n36665 , n36663 , n36664 );
not ( n36666 , n36665 );
and ( n36667 , n36662 , n36666 );
not ( n36668 , n36662 );
and ( n36669 , n36668 , n36665 );
nor ( n36670 , n36667 , n36669 );
buf ( n36671 , n33389 );
not ( n36672 , n36671 );
buf ( n36673 , n34098 );
nand ( n36674 , n36672 , n36673 );
nor ( n36675 , n36593 , n36674 );
not ( n36676 , n36675 );
not ( n36677 , n36374 );
or ( n36678 , n36676 , n36677 );
not ( n36679 , n36633 );
not ( n36680 , n36674 );
not ( n36681 , n36680 );
or ( n36682 , n36679 , n36681 );
and ( n36683 , n36672 , n36612 );
buf ( n36684 , n33596 );
nor ( n36685 , n36683 , n36684 );
nand ( n36686 , n36682 , n36685 );
not ( n36687 , n36686 );
nand ( n36688 , n36678 , n36687 );
buf ( n36689 , n33460 );
not ( n36690 , n36689 );
nor ( n36691 , n36690 , n36623 );
not ( n36692 , n36691 );
nor ( n36693 , n36692 , n36593 );
not ( n36694 , n36693 );
not ( n36695 , n36319 );
or ( n36696 , n36694 , n36695 );
not ( n36697 , n36691 );
not ( n36698 , n36609 );
or ( n36699 , n36697 , n36698 );
not ( n36700 , n36689 );
not ( n36701 , n36636 );
or ( n36702 , n36700 , n36701 );
buf ( n36703 , n33579 );
nand ( n36704 , n36702 , n36703 );
not ( n36705 , n36704 );
nand ( n36706 , n36699 , n36705 );
not ( n36707 , n36706 );
nand ( n36708 , n36696 , n36707 );
not ( n36709 , n36269 );
not ( n36710 , n36709 );
or ( n36711 , n36710 , n36648 );
buf ( n36712 , n35283 );
not ( n36713 , n36712 );
not ( n36714 , n35307 );
nand ( n36715 , n36713 , n36714 );
nor ( n36716 , n36715 , n36649 );
nand ( n36717 , n36711 , n36716 );
not ( n36718 , n36715 );
and ( n36719 , n36718 , n36645 );
not ( n36720 , n36714 );
buf ( n36721 , n36306 );
not ( n36722 , n36721 );
or ( n36723 , n36720 , n36722 );
buf ( n36724 , n36309 );
not ( n36725 , n36724 );
nand ( n36726 , n36723 , n36725 );
nor ( n36727 , n36719 , n36726 );
nand ( n36728 , n36717 , n36727 );
not ( n36729 , n36728 );
not ( n36730 , n36414 );
and ( n36731 , n32807 , n36559 );
buf ( n204009 , n36446 );
not ( n36733 , n204009 );
buf ( n204011 , n196449 );
not ( n36735 , n204011 );
or ( n36736 , n36733 , n36735 );
buf ( n204014 , n186254 );
buf ( n204015 , n835 );
buf ( n204016 , n866 );
xor ( n36740 , n204015 , n204016 );
buf ( n204018 , n36740 );
buf ( n204019 , n204018 );
nand ( n36743 , n204014 , n204019 );
buf ( n204021 , n36743 );
buf ( n204022 , n204021 );
nand ( n36746 , n36736 , n204022 );
buf ( n204024 , n36746 );
buf ( n204025 , n204024 );
buf ( n204026 , n203808 );
not ( n36750 , n204026 );
buf ( n204028 , n186197 );
not ( n36752 , n204028 );
or ( n36753 , n36750 , n36752 );
buf ( n204031 , n833 );
buf ( n204032 , n868 );
xnor ( n36756 , n204031 , n204032 );
buf ( n204034 , n36756 );
buf ( n204035 , n204034 );
not ( n36759 , n204035 );
buf ( n204037 , n186208 );
nand ( n36761 , n36759 , n204037 );
buf ( n204039 , n36761 );
buf ( n204040 , n204039 );
nand ( n36764 , n36753 , n204040 );
buf ( n204042 , n36764 );
buf ( n204043 , n204042 );
not ( n36767 , n204043 );
buf ( n204045 , n36767 );
buf ( n204046 , n204045 );
xor ( n36770 , n204025 , n204046 );
xor ( n36771 , n203780 , n203797 );
and ( n36772 , n36771 , n203815 );
and ( n36773 , n203780 , n203797 );
or ( n36774 , n36772 , n36773 );
buf ( n204052 , n36774 );
buf ( n204053 , n204052 );
and ( n36777 , n36770 , n204053 );
and ( n36778 , n204025 , n204046 );
or ( n36779 , n36777 , n36778 );
buf ( n204057 , n36779 );
buf ( n204058 , n204057 );
and ( n36782 , n196484 , n196485 );
buf ( n204060 , n36782 );
buf ( n204061 , n204060 );
buf ( n204062 , n203790 );
not ( n36786 , n204062 );
buf ( n204064 , n186640 );
not ( n36788 , n204064 );
or ( n36789 , n36786 , n36788 );
buf ( n204067 , n186340 );
buf ( n204068 , n864 );
buf ( n204069 , n837 );
xor ( n36793 , n204068 , n204069 );
buf ( n204071 , n36793 );
buf ( n204072 , n204071 );
nand ( n36796 , n204067 , n204072 );
buf ( n204074 , n36796 );
buf ( n204075 , n204074 );
nand ( n36799 , n36789 , n204075 );
buf ( n204077 , n36799 );
buf ( n204078 , n204077 );
xor ( n36802 , n204061 , n204078 );
buf ( n204080 , n203749 );
not ( n36804 , n204080 );
buf ( n204082 , n186435 );
not ( n36806 , n204082 );
or ( n36807 , n36804 , n36806 );
buf ( n204085 , n186444 );
buf ( n204086 , n870 );
nand ( n36810 , n204085 , n204086 );
buf ( n204088 , n36810 );
buf ( n204089 , n204088 );
nand ( n36813 , n36807 , n204089 );
buf ( n204091 , n36813 );
buf ( n204092 , n204091 );
xor ( n36816 , n36802 , n204092 );
buf ( n204094 , n36816 );
buf ( n204095 , n204094 );
xor ( n36819 , n203730 , n203738 );
and ( n36820 , n36819 , n203756 );
and ( n36821 , n203730 , n203738 );
or ( n36822 , n36820 , n36821 );
buf ( n204100 , n36822 );
buf ( n204101 , n204100 );
xor ( n36825 , n204095 , n204101 );
xor ( n36826 , n204025 , n204046 );
xor ( n36827 , n36826 , n204053 );
buf ( n204105 , n36827 );
buf ( n204106 , n204105 );
and ( n36830 , n36825 , n204106 );
and ( n36831 , n204095 , n204101 );
or ( n36832 , n36830 , n36831 );
buf ( n204110 , n36832 );
buf ( n204111 , n204110 );
xor ( n36835 , n204058 , n204111 );
xor ( n36836 , n204061 , n204078 );
and ( n36837 , n36836 , n204092 );
and ( n36838 , n204061 , n204078 );
or ( n36839 , n36837 , n36838 );
buf ( n204117 , n36839 );
buf ( n204118 , n204117 );
and ( n36842 , n203787 , n203788 );
buf ( n204120 , n36842 );
buf ( n204121 , n204120 );
buf ( n204122 , n204018 );
not ( n36846 , n204122 );
buf ( n204124 , n196449 );
not ( n36848 , n204124 );
or ( n36849 , n36846 , n36848 );
buf ( n204127 , n834 );
buf ( n204128 , n866 );
xnor ( n36852 , n204127 , n204128 );
buf ( n204130 , n36852 );
buf ( n204131 , n204130 );
not ( n36855 , n204131 );
buf ( n204133 , n186254 );
nand ( n36857 , n36855 , n204133 );
buf ( n204135 , n36857 );
buf ( n204136 , n204135 );
nand ( n36860 , n36849 , n204136 );
buf ( n204138 , n36860 );
buf ( n204139 , n204138 );
xor ( n36863 , n204121 , n204139 );
buf ( n204141 , n204042 );
xor ( n36865 , n36863 , n204141 );
buf ( n204143 , n36865 );
buf ( n204144 , n204143 );
xor ( n36868 , n204118 , n204144 );
buf ( n204146 , n204071 );
not ( n36870 , n204146 );
buf ( n204148 , n186640 );
not ( n36872 , n204148 );
or ( n36873 , n36870 , n36872 );
buf ( n204151 , n186340 );
buf ( n204152 , n864 );
buf ( n204153 , n836 );
xor ( n36877 , n204152 , n204153 );
buf ( n204155 , n36877 );
buf ( n204156 , n204155 );
nand ( n36880 , n204151 , n204156 );
buf ( n204158 , n36880 );
buf ( n204159 , n204158 );
nand ( n36883 , n36873 , n204159 );
buf ( n204161 , n36883 );
buf ( n204162 , n204161 );
buf ( n204163 , n186444 );
buf ( n204164 , n186435 );
or ( n36888 , n204163 , n204164 );
buf ( n204166 , n870 );
nand ( n36890 , n36888 , n204166 );
buf ( n204168 , n36890 );
buf ( n204169 , n204168 );
xor ( n36893 , n204162 , n204169 );
buf ( n204171 , n186197 );
not ( n36895 , n204171 );
buf ( n204173 , n36895 );
buf ( n204174 , n204173 );
buf ( n204175 , n204034 );
or ( n36899 , n204174 , n204175 );
buf ( n204177 , n186205 );
buf ( n204178 , n868 );
buf ( n204179 , n832 );
not ( n36903 , n204179 );
buf ( n204181 , n36903 );
buf ( n204182 , n204181 );
and ( n36906 , n204178 , n204182 );
not ( n36907 , n204178 );
buf ( n204185 , n832 );
and ( n36909 , n36907 , n204185 );
nor ( n36910 , n36906 , n36909 );
buf ( n204188 , n36910 );
buf ( n204189 , n204188 );
or ( n36913 , n204177 , n204189 );
nand ( n36914 , n36899 , n36913 );
buf ( n204192 , n36914 );
buf ( n204193 , n204192 );
xor ( n36917 , n36893 , n204193 );
buf ( n204195 , n36917 );
buf ( n204196 , n204195 );
xor ( n36920 , n36868 , n204196 );
buf ( n204198 , n36920 );
buf ( n204199 , n204198 );
xor ( n36923 , n36835 , n204199 );
buf ( n204201 , n36923 );
xor ( n36925 , n203761 , n203776 );
and ( n36926 , n36925 , n203818 );
and ( n36927 , n203761 , n203776 );
or ( n36928 , n36926 , n36927 );
buf ( n204206 , n36928 );
buf ( n204207 , n204206 );
xor ( n36931 , n204095 , n204101 );
xor ( n36932 , n36931 , n204106 );
buf ( n204210 , n36932 );
buf ( n204211 , n204210 );
xor ( n36935 , n204207 , n204211 );
xor ( n36936 , n203716 , n203759 );
and ( n36937 , n36936 , n203821 );
and ( n36938 , n203716 , n203759 );
or ( n36939 , n36937 , n36938 );
buf ( n204217 , n36939 );
buf ( n204218 , n204217 );
and ( n36942 , n36935 , n204218 );
and ( n36943 , n204207 , n204211 );
or ( n36944 , n36942 , n36943 );
buf ( n204222 , n36944 );
or ( n36946 , n204201 , n204222 );
xor ( n36947 , n203710 , n203824 );
and ( n36948 , n36947 , n203831 );
and ( n36949 , n203710 , n203824 );
or ( n36950 , n36948 , n36949 );
buf ( n204228 , n36950 );
xor ( n36952 , n204207 , n204211 );
xor ( n36953 , n36952 , n204218 );
buf ( n204231 , n36953 );
or ( n36955 , n204228 , n204231 );
nand ( n36956 , n36946 , n36955 );
not ( n36957 , n36956 );
nand ( n36958 , n36731 , n36957 );
nor ( n36959 , n36730 , n36958 );
nand ( n36960 , n36959 , n36374 );
not ( n36961 , n35756 );
not ( n36962 , n36659 );
or ( n36963 , n36961 , n36962 );
buf ( n36964 , n35712 );
nand ( n36965 , n36963 , n36964 );
nand ( n36966 , n35757 , n35717 );
not ( n36967 , n36966 );
and ( n36968 , n36965 , n36967 );
not ( n36969 , n36965 );
and ( n36970 , n36969 , n36966 );
nor ( n36971 , n36968 , n36970 );
nor ( n36972 , n36654 , n35729 );
nand ( n36973 , n36972 , n36659 , n36653 );
buf ( n36974 , n35722 );
nand ( n36975 , n36972 , n36974 );
not ( n36976 , n35625 );
buf ( n36977 , n35739 );
not ( n36978 , n36977 );
or ( n36979 , n36976 , n36978 );
not ( n36980 , n35742 );
nand ( n36981 , n36979 , n36980 );
not ( n36982 , n36981 );
nand ( n36983 , n36973 , n36975 , n36982 );
nand ( n36984 , n35743 , n35745 );
nand ( n36985 , n36983 , n36984 );
not ( n36986 , n36647 );
and ( n36987 , n35598 , n36277 );
nand ( n36988 , n36986 , n36987 );
nand ( n36989 , n36658 , n36987 , n36660 );
not ( n36990 , n202848 );
not ( n36991 , n35543 );
nand ( n36992 , n36990 , n36991 );
and ( n36993 , n36992 , n36274 );
not ( n36994 , n35540 );
and ( n36995 , n36993 , n36994 );
nor ( n36996 , n36995 , n36285 );
nand ( n36997 , n36988 , n36989 , n36996 );
nand ( n36998 , n36709 , n36647 );
buf ( n36999 , n36998 );
nor ( n37000 , n36649 , n36712 );
nand ( n37001 , n36710 , n37000 );
not ( n37002 , n36663 );
nor ( n37003 , n37002 , n36649 );
nand ( n37004 , n37003 , n36710 );
buf ( n37005 , n35612 );
not ( n37006 , n37005 );
nor ( n37007 , n36652 , n37006 );
not ( n37008 , n37007 );
not ( n37009 , n36659 );
or ( n37010 , n37008 , n37009 );
not ( n37011 , n37005 );
not ( n37012 , n35722 );
or ( n37013 , n37011 , n37012 );
not ( n37014 , n35733 );
nand ( n37015 , n37013 , n37014 );
not ( n37016 , n37015 );
nand ( n37017 , n37010 , n37016 );
not ( n37018 , n36983 );
not ( n37019 , n36659 );
buf ( n37020 , n35597 );
nor ( n37021 , n37019 , n37020 );
nand ( n37022 , n36658 , n37021 );
not ( n37023 , n36249 );
not ( n37024 , n36253 );
or ( n37025 , n37023 , n37024 );
nand ( n37026 , n37025 , n36264 );
nand ( n37027 , n37026 , n35817 );
and ( n37028 , n36253 , n36219 );
not ( n37029 , n36158 );
not ( n37030 , n37029 );
nand ( n37031 , n37028 , n37030 , n35817 );
buf ( n37032 , n36231 );
nand ( n37033 , n37027 , n37031 , n37032 );
and ( n37034 , n36234 , n36237 );
and ( n37035 , n37033 , n37034 );
not ( n37036 , n37033 );
not ( n37037 , n37034 );
and ( n37038 , n37036 , n37037 );
nor ( n37039 , n37035 , n37038 );
not ( n37040 , n35755 );
nand ( n37041 , n37040 , n35696 );
not ( n37042 , n37041 );
not ( n37043 , n36659 );
or ( n37044 , n37042 , n37043 );
or ( n37045 , n36659 , n37041 );
nand ( n37046 , n37044 , n37045 );
and ( n37047 , n35756 , n35757 );
not ( n37048 , n37047 );
not ( n37049 , n36659 );
or ( n37050 , n37048 , n37049 );
not ( n37051 , n36964 );
and ( n37052 , n37051 , n35757 );
not ( n37053 , n35717 );
nor ( n37054 , n37052 , n37053 );
nand ( n37055 , n37050 , n37054 );
not ( n37056 , n36653 );
not ( n37057 , n36659 );
or ( n37058 , n37056 , n37057 );
not ( n37059 , n36974 );
nand ( n37060 , n37058 , n37059 );
not ( n37061 , n36238 );
nand ( n37062 , n37028 , n36266 , n37030 );
nand ( n37063 , n37026 , n36266 );
nand ( n37064 , n37061 , n37062 , n37063 );
nand ( n37065 , n35777 , n35783 );
buf ( n37066 , n36240 );
nand ( n37067 , n37065 , n37066 );
not ( n37068 , n37067 );
and ( n37069 , n37064 , n37068 );
not ( n37070 , n37064 );
and ( n37071 , n37070 , n37067 );
nor ( n37072 , n37069 , n37071 );
not ( n37073 , n36219 );
not ( n37074 , n36158 );
or ( n37075 , n37073 , n37074 );
not ( n37076 , n36249 );
nand ( n37077 , n37075 , n37076 );
buf ( n37078 , n36256 );
nand ( n37079 , n36189 , n37078 );
not ( n37080 , n37079 );
and ( n37081 , n37077 , n37080 );
not ( n37082 , n37077 );
and ( n37083 , n37082 , n37079 );
nor ( n37084 , n37081 , n37083 );
not ( n37085 , n36218 );
not ( n37086 , n37085 );
not ( n37087 , n36158 );
or ( n37088 , n37086 , n37087 );
nand ( n37089 , n37088 , n36245 );
not ( n37090 , n36199 );
nand ( n37091 , n37090 , n36248 );
not ( n37092 , n37091 );
and ( n37093 , n37089 , n37092 );
not ( n37094 , n37089 );
and ( n37095 , n37094 , n37091 );
nor ( n37096 , n37093 , n37095 );
nand ( n37097 , n36955 , n36560 );
not ( n37098 , n37097 );
nand ( n37099 , n36380 , n37098 );
buf ( n37100 , n34102 );
xor ( n37101 , n204121 , n204139 );
and ( n37102 , n37101 , n204141 );
and ( n37103 , n204121 , n204139 );
or ( n37104 , n37102 , n37103 );
buf ( n204382 , n37104 );
buf ( n204383 , n204382 );
xor ( n37107 , n204118 , n204144 );
and ( n37108 , n37107 , n204196 );
and ( n37109 , n204118 , n204144 );
or ( n37110 , n37108 , n37109 );
buf ( n204388 , n37110 );
buf ( n204389 , n204388 );
xor ( n37113 , n204383 , n204389 );
buf ( n204391 , n204188 );
not ( n37115 , n204391 );
buf ( n204393 , n37115 );
buf ( n204394 , n204393 );
not ( n37118 , n204394 );
buf ( n204396 , n186197 );
not ( n37120 , n204396 );
or ( n37121 , n37118 , n37120 );
buf ( n204399 , n186208 );
buf ( n204400 , n868 );
nand ( n37124 , n204399 , n204400 );
buf ( n204402 , n37124 );
buf ( n204403 , n204402 );
nand ( n37127 , n37121 , n204403 );
buf ( n204405 , n37127 );
buf ( n204406 , n204405 );
not ( n37130 , n204406 );
buf ( n204408 , n37130 );
buf ( n204409 , n204408 );
xor ( n37133 , n204162 , n204169 );
and ( n37134 , n37133 , n204193 );
and ( n37135 , n204162 , n204169 );
or ( n37136 , n37134 , n37135 );
buf ( n204414 , n37136 );
buf ( n204415 , n204414 );
xor ( n37139 , n204409 , n204415 );
and ( n37140 , n204068 , n204069 );
buf ( n204418 , n37140 );
buf ( n204419 , n204418 );
buf ( n204420 , n204155 );
not ( n37144 , n204420 );
buf ( n204422 , n186640 );
not ( n37146 , n204422 );
or ( n37147 , n37144 , n37146 );
buf ( n204425 , n864 );
buf ( n204426 , n835 );
xnor ( n37150 , n204425 , n204426 );
buf ( n204428 , n37150 );
buf ( n204429 , n204428 );
not ( n37153 , n204429 );
buf ( n204431 , n186340 );
nand ( n37155 , n37153 , n204431 );
buf ( n204433 , n37155 );
buf ( n204434 , n204433 );
nand ( n37158 , n37147 , n204434 );
buf ( n204436 , n37158 );
buf ( n204437 , n204436 );
xor ( n37161 , n204419 , n204437 );
buf ( n204439 , n196446 );
buf ( n204440 , n204130 );
or ( n37164 , n204439 , n204440 );
buf ( n204442 , n186251 );
buf ( n204443 , n866 );
buf ( n204444 , n833 );
not ( n37168 , n204444 );
buf ( n204446 , n37168 );
buf ( n204447 , n204446 );
and ( n37171 , n204443 , n204447 );
not ( n37172 , n204443 );
buf ( n204450 , n833 );
and ( n37174 , n37172 , n204450 );
nor ( n37175 , n37171 , n37174 );
buf ( n204453 , n37175 );
buf ( n204454 , n204453 );
or ( n37178 , n204442 , n204454 );
nand ( n37179 , n37164 , n37178 );
buf ( n204457 , n37179 );
buf ( n204458 , n204457 );
xor ( n37182 , n37161 , n204458 );
buf ( n204460 , n37182 );
buf ( n204461 , n204460 );
xor ( n37185 , n37139 , n204461 );
buf ( n204463 , n37185 );
buf ( n204464 , n204463 );
and ( n37188 , n37113 , n204464 );
and ( n37189 , n204383 , n204389 );
or ( n37190 , n37188 , n37189 );
buf ( n204468 , n37190 );
and ( n37192 , n204152 , n204153 );
buf ( n204470 , n37192 );
buf ( n204471 , n204470 );
buf ( n204472 , n186205 );
not ( n37196 , n204472 );
buf ( n204474 , n204173 );
not ( n37198 , n204474 );
or ( n37199 , n37196 , n37198 );
buf ( n204477 , n868 );
nand ( n37201 , n37199 , n204477 );
buf ( n204479 , n37201 );
buf ( n204480 , n204479 );
xor ( n37204 , n204471 , n204480 );
buf ( n204482 , n196446 );
buf ( n204483 , n204453 );
or ( n37207 , n204482 , n204483 );
buf ( n204485 , n186251 );
buf ( n204486 , n832 );
buf ( n204487 , n866 );
xnor ( n37211 , n204486 , n204487 );
buf ( n204489 , n37211 );
buf ( n204490 , n204489 );
or ( n37214 , n204485 , n204490 );
nand ( n37215 , n37207 , n37214 );
buf ( n204493 , n37215 );
buf ( n204494 , n204493 );
xor ( n37218 , n37204 , n204494 );
buf ( n204496 , n37218 );
buf ( n204497 , n204496 );
buf ( n204498 , n204405 );
buf ( n204499 , n186326 );
buf ( n204500 , n204428 );
or ( n37224 , n204499 , n204500 );
buf ( n204502 , n186343 );
buf ( n204503 , n864 );
buf ( n204504 , n834 );
xnor ( n37228 , n204503 , n204504 );
buf ( n204506 , n37228 );
buf ( n204507 , n204506 );
or ( n37231 , n204502 , n204507 );
nand ( n37232 , n37224 , n37231 );
buf ( n204510 , n37232 );
buf ( n204511 , n204510 );
xor ( n37235 , n204498 , n204511 );
xor ( n37236 , n204419 , n204437 );
and ( n37237 , n37236 , n204458 );
and ( n37238 , n204419 , n204437 );
or ( n37239 , n37237 , n37238 );
buf ( n204517 , n37239 );
buf ( n204518 , n204517 );
xor ( n37242 , n37235 , n204518 );
buf ( n204520 , n37242 );
buf ( n204521 , n204520 );
xor ( n37245 , n204497 , n204521 );
xor ( n37246 , n204409 , n204415 );
and ( n37247 , n37246 , n204461 );
and ( n37248 , n204409 , n204415 );
or ( n37249 , n37247 , n37248 );
buf ( n204527 , n37249 );
buf ( n204528 , n204527 );
xor ( n37252 , n37245 , n204528 );
buf ( n204530 , n37252 );
nor ( n37254 , n204468 , n204530 );
not ( n37255 , n37254 );
xor ( n37256 , n204058 , n204111 );
and ( n37257 , n37256 , n204199 );
and ( n37258 , n204058 , n204111 );
or ( n37259 , n37257 , n37258 );
buf ( n204537 , n37259 );
xor ( n37261 , n204383 , n204389 );
xor ( n37262 , n37261 , n204464 );
buf ( n204540 , n37262 );
or ( n37264 , n204537 , n204540 );
nand ( n37265 , n37255 , n37264 );
nor ( n37266 , n36956 , n37265 );
xor ( n37267 , n204497 , n204521 );
and ( n37268 , n37267 , n204528 );
and ( n37269 , n204497 , n204521 );
or ( n37270 , n37268 , n37269 );
buf ( n204548 , n37270 );
xor ( n37272 , n204471 , n204480 );
and ( n37273 , n37272 , n204494 );
and ( n37274 , n204471 , n204480 );
or ( n37275 , n37273 , n37274 );
buf ( n204553 , n37275 );
buf ( n204554 , n204553 );
buf ( n204555 , n835 );
buf ( n204556 , n864 );
and ( n37280 , n204555 , n204556 );
buf ( n204558 , n37280 );
buf ( n204559 , n204558 );
buf ( n204560 , n204489 );
not ( n37284 , n204560 );
buf ( n204562 , n196449 );
nand ( n37286 , n37284 , n204562 );
buf ( n204564 , n37286 );
buf ( n204565 , n204564 );
buf ( n204566 , n186254 );
buf ( n204567 , n866 );
nand ( n37291 , n204566 , n204567 );
buf ( n204569 , n37291 );
buf ( n204570 , n204569 );
and ( n37294 , n204565 , n204570 );
buf ( n204572 , n37294 );
buf ( n204573 , n204572 );
xor ( n37297 , n204559 , n204573 );
buf ( n204575 , n186326 );
buf ( n204576 , n204506 );
or ( n37300 , n204575 , n204576 );
buf ( n204578 , n186343 );
buf ( n204579 , n864 );
buf ( n204580 , n204446 );
and ( n37304 , n204579 , n204580 );
not ( n37305 , n204579 );
buf ( n204583 , n833 );
and ( n37307 , n37305 , n204583 );
nor ( n37308 , n37304 , n37307 );
buf ( n204586 , n37308 );
buf ( n204587 , n204586 );
or ( n37311 , n204578 , n204587 );
nand ( n37312 , n37300 , n37311 );
buf ( n204590 , n37312 );
buf ( n204591 , n204590 );
xor ( n37315 , n37297 , n204591 );
buf ( n204593 , n37315 );
buf ( n204594 , n204593 );
xor ( n37318 , n204554 , n204594 );
xor ( n37319 , n204498 , n204511 );
and ( n37320 , n37319 , n204518 );
and ( n37321 , n204498 , n204511 );
or ( n37322 , n37320 , n37321 );
buf ( n204600 , n37322 );
buf ( n204601 , n204600 );
xor ( n37325 , n37318 , n204601 );
buf ( n204603 , n37325 );
nor ( n37327 , n204548 , n204603 );
xor ( n37328 , n204554 , n204594 );
and ( n37329 , n37328 , n204601 );
and ( n37330 , n204554 , n204594 );
or ( n37331 , n37329 , n37330 );
buf ( n204609 , n37331 );
buf ( n204610 , n204572 );
not ( n37334 , n204610 );
buf ( n204612 , n37334 );
buf ( n204613 , n204612 );
xor ( n37337 , n204559 , n204573 );
and ( n37338 , n37337 , n204591 );
and ( n37339 , n204559 , n204573 );
or ( n37340 , n37338 , n37339 );
buf ( n204618 , n37340 );
buf ( n204619 , n204618 );
xor ( n37343 , n204613 , n204619 );
buf ( n204621 , n196449 );
buf ( n204622 , n186254 );
or ( n37346 , n204621 , n204622 );
buf ( n204624 , n866 );
nand ( n37348 , n37346 , n204624 );
buf ( n204626 , n37348 );
buf ( n204627 , n204626 );
buf ( n204628 , n834 );
buf ( n204629 , n864 );
and ( n37353 , n204628 , n204629 );
buf ( n204631 , n37353 );
buf ( n204632 , n204631 );
xor ( n37356 , n204627 , n204632 );
buf ( n204634 , n186326 );
buf ( n204635 , n204586 );
or ( n37359 , n204634 , n204635 );
buf ( n204637 , n186343 );
buf ( n204638 , n864 );
buf ( n204639 , n204181 );
and ( n37363 , n204638 , n204639 );
not ( n37364 , n204638 );
buf ( n204642 , n832 );
and ( n37366 , n37364 , n204642 );
nor ( n37367 , n37363 , n37366 );
buf ( n204645 , n37367 );
buf ( n204646 , n204645 );
or ( n37370 , n204637 , n204646 );
nand ( n37371 , n37359 , n37370 );
buf ( n204649 , n37371 );
buf ( n204650 , n204649 );
xor ( n37374 , n37356 , n204650 );
buf ( n204652 , n37374 );
buf ( n204653 , n204652 );
xor ( n37377 , n37343 , n204653 );
buf ( n204655 , n37377 );
nor ( n37379 , n204609 , n204655 );
nor ( n37380 , n37327 , n37379 );
xor ( n37381 , n204613 , n204619 );
and ( n37382 , n37381 , n204653 );
and ( n37383 , n204613 , n204619 );
or ( n37384 , n37382 , n37383 );
buf ( n204662 , n37384 );
buf ( n204663 , n833 );
buf ( n204664 , n864 );
nand ( n37388 , n204663 , n204664 );
buf ( n204666 , n37388 );
buf ( n204667 , n204666 );
buf ( n204668 , n186326 );
buf ( n204669 , n204645 );
or ( n37393 , n204668 , n204669 );
buf ( n204671 , n186343 );
buf ( n204672 , n864 );
not ( n37396 , n204672 );
buf ( n204674 , n37396 );
buf ( n204675 , n204674 );
or ( n37399 , n204671 , n204675 );
nand ( n37400 , n37393 , n37399 );
buf ( n204678 , n37400 );
buf ( n204679 , n204678 );
xor ( n37403 , n204667 , n204679 );
xor ( n37404 , n204627 , n204632 );
and ( n37405 , n37404 , n204650 );
and ( n37406 , n204627 , n204632 );
or ( n37407 , n37405 , n37406 );
buf ( n204685 , n37407 );
buf ( n204686 , n204685 );
xor ( n37410 , n37403 , n204686 );
buf ( n204688 , n37410 );
or ( n37412 , n204662 , n204688 );
and ( n37413 , n37380 , n37412 );
and ( n37414 , n37266 , n37413 );
and ( n37415 , n36561 , n37414 );
nand ( n37416 , n37100 , n37415 );
and ( n37417 , n36252 , n36219 );
not ( n37418 , n37417 );
not ( n37419 , n36158 );
or ( n37420 , n37418 , n37419 );
not ( n37421 , n36189 );
not ( n37422 , n36249 );
or ( n37423 , n37421 , n37422 );
nand ( n37424 , n37423 , n37078 );
not ( n37425 , n37424 );
nand ( n37426 , n37420 , n37425 );
not ( n37427 , n36380 );
not ( n37428 , n36673 );
not ( n37429 , n36609 );
or ( n37430 , n37428 , n37429 );
not ( n37431 , n36612 );
nand ( n37432 , n37430 , n37431 );
not ( n37433 , n37432 );
not ( n37434 , n36957 );
not ( n37435 , n36579 );
or ( n37436 , n37434 , n37435 );
not ( n37437 , n36946 );
and ( n37438 , n204231 , n204228 );
not ( n37439 , n37438 );
or ( n37440 , n37437 , n37439 );
nand ( n37441 , n204201 , n204222 );
nand ( n37442 , n37440 , n37441 );
not ( n37443 , n37442 );
nand ( n37444 , n37436 , n37443 );
not ( n37445 , n37444 );
not ( n37446 , n36955 );
not ( n37447 , n36579 );
or ( n37448 , n37446 , n37447 );
not ( n37449 , n37438 );
nand ( n37450 , n37448 , n37449 );
not ( n37451 , n37450 );
buf ( n37452 , n34096 );
not ( n37453 , n37452 );
not ( n37454 , n36633 );
or ( n37455 , n37453 , n37454 );
not ( n37456 , n33559 );
nand ( n37457 , n37455 , n37456 );
not ( n37458 , n37457 );
buf ( n37459 , n33417 );
not ( n37460 , n37459 );
nor ( n37461 , n37460 , n36671 );
nand ( n37462 , n37461 , n36673 );
not ( n37463 , n37462 );
not ( n37464 , n37463 );
not ( n37465 , n36633 );
or ( n37466 , n37464 , n37465 );
not ( n37467 , n37461 );
not ( n37468 , n36612 );
or ( n37469 , n37467 , n37468 );
and ( n37470 , n36684 , n37459 );
not ( n37471 , n33599 );
nor ( n37472 , n37470 , n37471 );
nand ( n37473 , n37469 , n37472 );
not ( n37474 , n37473 );
nand ( n37475 , n37466 , n37474 );
not ( n37476 , n37475 );
not ( n37477 , n37264 );
nor ( n37478 , n37477 , n36956 );
not ( n37479 , n37478 );
not ( n37480 , n36579 );
or ( n37481 , n37479 , n37480 );
not ( n37482 , n37264 );
not ( n37483 , n37442 );
or ( n37484 , n37482 , n37483 );
nand ( n37485 , n204537 , n204540 );
nand ( n37486 , n37484 , n37485 );
not ( n37487 , n37486 );
nand ( n37488 , n37481 , n37487 );
nand ( n37489 , n37000 , n36648 );
not ( n37490 , n35597 );
nand ( n37491 , n36648 , n37490 );
nand ( n37492 , n37003 , n36648 );
not ( n37493 , n36012 );
not ( n37494 , n36013 );
or ( n37495 , n37493 , n37494 );
nand ( n37496 , n37495 , n35877 );
not ( n37497 , n36663 );
not ( n37498 , n36645 );
or ( n37499 , n37497 , n37498 );
nand ( n37500 , n37499 , n36664 );
nand ( n37501 , n36013 , n35877 );
buf ( n37502 , n36012 );
nand ( n37503 , n37501 , n37502 );
not ( n37504 , n36712 );
not ( n37505 , n37504 );
not ( n37506 , n36645 );
or ( n37507 , n37505 , n37506 );
not ( n37508 , n36721 );
nand ( n37509 , n37507 , n37508 );
not ( n37510 , n37380 );
not ( n37511 , n37265 );
not ( n37512 , n37511 );
not ( n37513 , n37442 );
or ( n37514 , n37512 , n37513 );
not ( n37515 , n37485 );
not ( n37516 , n37254 );
and ( n37517 , n37515 , n37516 );
and ( n37518 , n204468 , n204530 );
nor ( n37519 , n37517 , n37518 );
nand ( n37520 , n37514 , n37519 );
not ( n37521 , n37520 );
or ( n37522 , n37510 , n37521 );
nand ( n37523 , n204548 , n204603 );
or ( n37524 , n37523 , n37379 );
nand ( n37525 , n204609 , n204655 );
nand ( n37526 , n37524 , n37525 );
not ( n37527 , n37526 );
nand ( n37528 , n37522 , n37527 );
not ( n37529 , n37327 );
not ( n37530 , n37529 );
not ( n37531 , n37520 );
or ( n37532 , n37530 , n37531 );
nand ( n37533 , n37532 , n37523 );
not ( n37534 , n37533 );
not ( n37535 , n36609 );
not ( n37536 , n37413 );
not ( n37537 , n37520 );
or ( n37538 , n37536 , n37537 );
and ( n37539 , n37526 , n37412 );
and ( n37540 , n204662 , n204688 );
nor ( n37541 , n37539 , n37540 );
nand ( n37542 , n37538 , n37541 );
buf ( n37543 , n201343 );
or ( n37544 , n37543 , n24107 );
not ( n37545 , n34088 );
nand ( n37546 , n37544 , n37545 );
not ( n37547 , n37546 );
buf ( n37548 , n36601 );
and ( n37549 , n37547 , n37548 );
not ( n37550 , n37544 );
not ( n37551 , n34082 );
not ( n37552 , n37551 );
or ( n37553 , n37550 , n37552 );
nand ( n37554 , n37553 , n34074 );
nor ( n37555 , n37549 , n37554 );
not ( n37556 , n36414 );
nor ( n37557 , n37556 , n37097 );
not ( n37558 , n34127 );
and ( n37559 , n36322 , n36361 );
nand ( n37560 , n36372 , n37559 );
nor ( n37561 , n37558 , n37560 );
not ( n37562 , n32723 );
buf ( n37563 , n32550 );
nor ( n37564 , n37562 , n37563 );
and ( n37565 , n36371 , n37564 );
nand ( n37566 , n36010 , n35980 );
not ( n37567 , n36007 );
not ( n37568 , n36008 );
nand ( n37569 , n37567 , n37568 );
nand ( n37570 , n37566 , n37569 );
not ( n37571 , n37548 );
nor ( n37572 , n36593 , n37462 );
and ( n37573 , n37266 , n37380 );
nand ( n37574 , n36561 , n37573 );
nand ( n37575 , n36561 , n37266 );
and ( n37576 , n37266 , n37529 );
nand ( n37577 , n36561 , n37576 );
not ( n37578 , n32723 );
not ( n37579 , n36330 );
or ( n37580 , n37578 , n37579 );
not ( n37581 , n36333 );
nand ( n37582 , n37580 , n37581 );
buf ( n37583 , n34118 );
not ( n37584 , n37583 );
nor ( n37585 , n37584 , n34088 );
not ( n37586 , n36399 );
and ( n37587 , n35957 , n35878 );
not ( n37588 , n35960 );
nor ( n37589 , n37587 , n37588 );
nand ( n37590 , n33637 , n33633 );
and ( n37591 , n37590 , n34084 );
not ( n37592 , n37591 );
nand ( n37593 , n35711 , n35706 );
not ( n37594 , n37593 );
nand ( n37595 , n37459 , n33599 );
not ( n37596 , n37595 );
nand ( n37597 , n36689 , n36703 );
not ( n37598 , n37597 );
nand ( n37599 , n36714 , n36725 );
not ( n37600 , n37599 );
not ( n37601 , n36390 );
nand ( n37602 , n36955 , n37449 );
nand ( n37603 , n37264 , n37485 );
nand ( n37604 , n37005 , n37014 );
nand ( n37605 , n32861 , n36348 );
not ( n37606 , n35828 );
not ( n37607 , n37606 );
nand ( n37608 , n37607 , n36262 );
nand ( n37609 , n37452 , n37456 );
nand ( n37610 , n35957 , n35960 );
not ( n37611 , n36314 );
nand ( n37612 , n37611 , n36312 );
not ( n37613 , n37612 );
nand ( n37614 , n35817 , n36231 );
not ( n37615 , n37614 );
not ( n37616 , n36984 );
buf ( n37617 , n37254 );
nor ( n37618 , n37518 , n37617 );
not ( n37619 , n37618 );
not ( n37620 , n35751 );
nor ( n37621 , n37620 , n35720 );
not ( n37622 , n37621 );
not ( n37623 , n36407 );
not ( n37624 , n36088 );
not ( n37625 , n36121 );
or ( n37626 , n37624 , n37625 );
nand ( n37627 , n37626 , n36155 );
not ( n37628 , n37627 );
not ( n37629 , n37563 );
nand ( n37630 , n36584 , n36588 );
buf ( n204908 , n204666 );
not ( n37632 , n204908 );
buf ( n204910 , n832 );
buf ( n204911 , n864 );
nand ( n37635 , n204910 , n204911 );
buf ( n204913 , n37635 );
buf ( n204914 , n204913 );
not ( n37638 , n204914 );
buf ( n204916 , n186640 );
buf ( n204917 , n186340 );
or ( n37641 , n204916 , n204917 );
buf ( n204919 , n864 );
nand ( n37643 , n37641 , n204919 );
buf ( n204921 , n37643 );
buf ( n204922 , n204921 );
not ( n37646 , n204922 );
or ( n37647 , n37638 , n37646 );
buf ( n204925 , n204921 );
buf ( n204926 , n204913 );
or ( n37650 , n204925 , n204926 );
nand ( n37651 , n37647 , n37650 );
buf ( n204929 , n37651 );
buf ( n204930 , n204929 );
not ( n37654 , n204930 );
or ( n37655 , n37632 , n37654 );
buf ( n204933 , n204929 );
buf ( n204934 , n204666 );
or ( n37658 , n204933 , n204934 );
nand ( n37659 , n37655 , n37658 );
buf ( n204937 , n37659 );
not ( n37661 , n204937 );
xor ( n37662 , n204667 , n204679 );
and ( n37663 , n37662 , n204686 );
and ( n37664 , n204667 , n204679 );
or ( n37665 , n37663 , n37664 );
buf ( n204943 , n37665 );
not ( n37667 , n204943 );
or ( n37668 , n37661 , n37667 );
or ( n37669 , n204943 , n204937 );
nand ( n37670 , n37668 , n37669 );
not ( n37671 , n37379 );
nand ( n37672 , n37671 , n37525 );
nand ( n37673 , n36992 , n36273 );
nand ( n37674 , n37085 , n36245 );
not ( n37675 , n203418 );
nand ( n37676 , n37675 , n36148 );
and ( n37677 , n37266 , n36580 );
nor ( n37678 , n37677 , n37520 );
and ( n37679 , n37414 , n36580 );
nor ( n37680 , n37679 , n37542 );
and ( n37681 , n35759 , n36974 );
nor ( n37682 , n37681 , n36977 );
or ( n37683 , n203282 , n196315 );
and ( n37684 , n36006 , n37683 );
not ( n37685 , n37509 );
nand ( n37686 , n37685 , n37489 , n37001 );
nand ( n37687 , n36731 , n37478 );
not ( n37688 , n37687 );
nand ( n37689 , n37688 , n36380 );
not ( n37690 , n36958 );
nand ( n37691 , n37690 , n34102 );
not ( n37692 , n37575 );
nand ( n37693 , n37692 , n37100 );
not ( n37694 , n37560 );
nand ( n37695 , n37694 , n34102 );
not ( n37696 , n35997 );
nand ( n37697 , n37696 , n37568 );
xor ( n37698 , n37697 , n36006 );
not ( n37699 , n36266 );
nor ( n37700 , n37699 , n36229 );
not ( n37701 , n33589 );
nand ( n37702 , n37701 , n33595 );
not ( n37703 , n37452 );
nor ( n37704 , n37703 , n36593 );
not ( n37705 , n36285 );
nand ( n37706 , n37705 , n36277 );
and ( n37707 , n31829 , n198286 );
xor ( n37708 , n183994 , n183988 );
not ( n37709 , n37708 );
buf ( n204987 , n183526 );
buf ( n204988 , n183266 );
and ( n37712 , n204987 , n204988 );
buf ( n204990 , n37712 );
not ( n37714 , n204990 );
and ( n37715 , n37709 , n37714 );
and ( n37716 , n183259 , n182960 );
buf ( n204994 , n37716 );
xor ( n37718 , n183266 , n183526 );
buf ( n204996 , n37718 );
nor ( n37720 , n204994 , n204996 );
buf ( n204998 , n37720 );
nor ( n37722 , n37715 , n204998 );
nand ( n37723 , n37707 , n37722 );
buf ( n205001 , n37723 );
not ( n37725 , n205001 );
buf ( n205003 , n37725 );
not ( n37727 , n31792 );
and ( n37728 , n205003 , n37727 );
nor ( n37729 , n204990 , n37708 );
nor ( n37730 , n37729 , n204998 );
not ( n37731 , n37730 );
not ( n37732 , n31799 );
or ( n37733 , n31826 , n199105 );
not ( n37734 , n37733 );
or ( n37735 , n37732 , n37734 );
nand ( n37736 , n37735 , n31831 );
not ( n37737 , n37736 );
or ( n37738 , n37731 , n37737 );
not ( n37739 , n37729 );
buf ( n205017 , n37716 );
buf ( n205018 , n37718 );
nand ( n37742 , n205017 , n205018 );
buf ( n205020 , n37742 );
not ( n37744 , n205020 );
and ( n37745 , n37739 , n37744 );
nand ( n37746 , n37708 , n204990 );
not ( n37747 , n37746 );
nor ( n37748 , n37745 , n37747 );
nand ( n37749 , n37738 , n37748 );
nor ( n37750 , n37728 , n37749 );
buf ( n205028 , n37750 );
buf ( n205029 , n199058 );
buf ( n205030 , n37723 );
or ( n37754 , n205029 , n205030 );
buf ( n205032 , n37754 );
buf ( n205033 , n205032 );
not ( n37757 , n31065 );
nand ( n37758 , n37757 , n205003 );
buf ( n205036 , n37758 );
nand ( n37760 , n205028 , n205033 , n205036 );
buf ( n205038 , n37760 );
buf ( n205039 , n205038 );
buf ( n205040 , n31749 );
not ( n37764 , n37730 );
not ( n37765 , n37736 );
or ( n37766 , n37764 , n37765 );
nand ( n37767 , n37766 , n37748 );
buf ( n205045 , n37767 );
not ( n37769 , n205045 );
buf ( n205047 , n37769 );
buf ( n205048 , n205047 );
and ( n37772 , n205040 , n205048 );
buf ( n205050 , n37772 );
buf ( n205051 , n205050 );
buf ( n205052 , n199058 );
buf ( n205053 , n199003 );
buf ( n205054 , n31791 );
nor ( n37778 , n205053 , n205054 );
buf ( n205056 , n37778 );
buf ( n205057 , n205056 );
and ( n37781 , n205052 , n205057 );
buf ( n205059 , n37781 );
buf ( n205060 , n205059 );
buf ( n205061 , n198980 );
nand ( n37785 , n205051 , n205060 , n205061 );
buf ( n205063 , n37785 );
buf ( n205064 , n205063 );
nand ( n37788 , n205039 , n205064 );
buf ( n205066 , n37788 );
buf ( n205067 , n205066 );
buf ( n37791 , n205067 );
buf ( n205069 , n37791 );
buf ( n205070 , n205069 );
not ( n37794 , n205070 );
buf ( n205072 , n37794 );
not ( n37796 , n205072 );
buf ( n205074 , n184771 );
buf ( n205075 , n184900 );
xor ( n37799 , n205074 , n205075 );
buf ( n205077 , n37799 );
buf ( n205078 , n205077 );
buf ( n205079 , n184910 );
buf ( n205080 , n184946 );
and ( n37804 , n205079 , n205080 );
buf ( n205082 , n37804 );
buf ( n205083 , n205082 );
nor ( n37807 , n205078 , n205083 );
buf ( n205085 , n37807 );
buf ( n205086 , n205085 );
buf ( n205087 , n184982 );
xor ( n37811 , n205079 , n205080 );
buf ( n205089 , n37811 );
buf ( n205090 , n205089 );
nor ( n37814 , n205087 , n205090 );
buf ( n205092 , n37814 );
buf ( n205093 , n205092 );
nor ( n37817 , n205086 , n205093 );
buf ( n205095 , n37817 );
buf ( n205096 , n205095 );
buf ( n205097 , n183988 );
buf ( n205098 , n183994 );
and ( n37822 , n205097 , n205098 );
buf ( n205100 , n37822 );
buf ( n205101 , n205100 );
xor ( n37825 , n185001 , n185004 );
buf ( n205103 , n37825 );
nor ( n37827 , n205101 , n205103 );
buf ( n205105 , n37827 );
buf ( n205106 , n205105 );
buf ( n205107 , n185004 );
buf ( n205108 , n185001 );
and ( n37832 , n205107 , n205108 );
buf ( n205110 , n37832 );
buf ( n205111 , n205110 );
buf ( n205112 , n185033 );
nor ( n37836 , n205111 , n205112 );
buf ( n205114 , n37836 );
buf ( n205115 , n205114 );
nor ( n37839 , n205106 , n205115 );
buf ( n205117 , n37839 );
buf ( n205118 , n205117 );
nand ( n37842 , n205096 , n205118 );
buf ( n205120 , n37842 );
buf ( n205121 , n205120 );
and ( n37845 , n205074 , n205075 );
buf ( n205123 , n37845 );
buf ( n205124 , n205123 );
not ( n37848 , n205124 );
buf ( n205126 , n185231 );
buf ( n205127 , n185058 );
xor ( n37851 , n205126 , n205127 );
buf ( n205129 , n37851 );
buf ( n205130 , n205129 );
not ( n37854 , n205130 );
buf ( n205132 , n37854 );
buf ( n205133 , n205132 );
nand ( n37857 , n37848 , n205133 );
buf ( n205135 , n37857 );
buf ( n205136 , n205135 );
xor ( n37860 , n185399 , n185393 );
buf ( n205138 , n37860 );
and ( n37862 , n205126 , n205127 );
buf ( n205140 , n37862 );
buf ( n205141 , n205140 );
or ( n37865 , n205138 , n205141 );
buf ( n205143 , n37865 );
buf ( n205144 , n205143 );
and ( n37868 , n205136 , n205144 );
buf ( n205146 , n37868 );
buf ( n205147 , n205146 );
and ( n37871 , n185399 , n185393 );
buf ( n205149 , n37871 );
buf ( n205150 , n185661 );
buf ( n205151 , n185667 );
xor ( n37875 , n205150 , n205151 );
buf ( n205153 , n37875 );
buf ( n205154 , n205153 );
nor ( n37878 , n205149 , n205154 );
buf ( n205156 , n37878 );
buf ( n205157 , n205156 );
and ( n37881 , n205150 , n205151 );
buf ( n205159 , n37881 );
buf ( n205160 , n205159 );
xor ( n37884 , n185538 , n185544 );
and ( n37885 , n37884 , n185592 );
and ( n37886 , n185538 , n185544 );
or ( n37887 , n37885 , n37886 );
buf ( n205165 , n37887 );
buf ( n205166 , n205165 );
xor ( n37890 , n185598 , n185615 );
and ( n37891 , n37890 , n185633 );
and ( n37892 , n185598 , n185615 );
or ( n37893 , n37891 , n37892 );
buf ( n205171 , n37893 );
buf ( n205172 , n205171 );
or ( n37896 , n170019 , n2554 );
nand ( n37897 , n37896 , n808 );
buf ( n205175 , n37897 );
buf ( n205176 , n18313 );
not ( n37900 , n205176 );
buf ( n205178 , n181588 );
not ( n37902 , n205178 );
or ( n37903 , n37900 , n37902 );
buf ( n205181 , n181594 );
buf ( n205182 , n806 );
buf ( n205183 , n768 );
and ( n37907 , n205182 , n205183 );
not ( n37908 , n205182 );
buf ( n205186 , n768 );
not ( n37910 , n205186 );
buf ( n205188 , n37910 );
buf ( n205189 , n205188 );
and ( n37913 , n37908 , n205189 );
nor ( n37914 , n37907 , n37913 );
buf ( n205192 , n37914 );
buf ( n205193 , n205192 );
nand ( n37917 , n205181 , n205193 );
buf ( n205195 , n37917 );
buf ( n205196 , n205195 );
nand ( n37920 , n37903 , n205196 );
buf ( n205198 , n37920 );
buf ( n205199 , n205198 );
xor ( n37923 , n205175 , n205199 );
buf ( n205201 , n185584 );
not ( n37925 , n205201 );
buf ( n205203 , n170419 );
not ( n37927 , n205203 );
or ( n37928 , n37925 , n37927 );
buf ( n205206 , n168870 );
buf ( n205207 , n772 );
buf ( n205208 , n802 );
xor ( n37932 , n205207 , n205208 );
buf ( n205210 , n37932 );
buf ( n205211 , n205210 );
nand ( n37935 , n205206 , n205211 );
buf ( n205213 , n37935 );
buf ( n205214 , n205213 );
nand ( n37938 , n37928 , n205214 );
buf ( n205216 , n37938 );
buf ( n205217 , n205216 );
xor ( n37941 , n37923 , n205217 );
buf ( n205219 , n37941 );
buf ( n205220 , n205219 );
xor ( n37944 , n205172 , n205220 );
buf ( n205222 , n185629 );
xor ( n37946 , n185561 , n185573 );
and ( n37947 , n37946 , n185590 );
and ( n37948 , n185561 , n185573 );
or ( n37949 , n37947 , n37948 );
buf ( n205227 , n37949 );
xor ( n37951 , n205222 , n205227 );
and ( n37952 , n185303 , n185304 );
buf ( n205230 , n37952 );
buf ( n205231 , n205230 );
buf ( n205232 , n185555 );
not ( n37956 , n205232 );
buf ( n205234 , n177819 );
not ( n37958 , n205234 );
or ( n37959 , n37956 , n37958 );
buf ( n205237 , n170972 );
buf ( n205238 , n774 );
buf ( n205239 , n800 );
xor ( n37963 , n205238 , n205239 );
buf ( n205241 , n37963 );
buf ( n205242 , n205241 );
nand ( n37966 , n205237 , n205242 );
buf ( n205244 , n37966 );
buf ( n205245 , n205244 );
nand ( n37969 , n37959 , n205245 );
buf ( n205247 , n37969 );
buf ( n205248 , n205247 );
xor ( n37972 , n205231 , n205248 );
buf ( n205250 , n185608 );
not ( n37974 , n205250 );
buf ( n205252 , n183183 );
not ( n37976 , n205252 );
or ( n37977 , n37974 , n37976 );
buf ( n205255 , n178447 );
buf ( n205256 , n770 );
buf ( n205257 , n804 );
xor ( n37981 , n205256 , n205257 );
buf ( n205259 , n37981 );
buf ( n205260 , n205259 );
nand ( n37984 , n205255 , n205260 );
buf ( n205262 , n37984 );
buf ( n205263 , n205262 );
nand ( n37987 , n37977 , n205263 );
buf ( n205265 , n37987 );
buf ( n205266 , n205265 );
xor ( n37990 , n37972 , n205266 );
buf ( n205268 , n37990 );
buf ( n205269 , n205268 );
xor ( n37993 , n37951 , n205269 );
buf ( n205271 , n37993 );
buf ( n205272 , n205271 );
xor ( n37996 , n37944 , n205272 );
buf ( n205274 , n37996 );
buf ( n205275 , n205274 );
xor ( n37999 , n205166 , n205275 );
xor ( n38000 , n185636 , n185642 );
and ( n38001 , n38000 , n185649 );
and ( n38002 , n185636 , n185642 );
or ( n38003 , n38001 , n38002 );
buf ( n205281 , n38003 );
buf ( n205282 , n205281 );
xor ( n38006 , n37999 , n205282 );
buf ( n205284 , n38006 );
buf ( n205285 , n205284 );
xor ( n38009 , n185595 , n185652 );
and ( n38010 , n38009 , n185659 );
and ( n38011 , n185595 , n185652 );
or ( n38012 , n38010 , n38011 );
buf ( n205290 , n38012 );
buf ( n205291 , n205290 );
xor ( n38015 , n205285 , n205291 );
buf ( n205293 , n38015 );
buf ( n205294 , n205293 );
nor ( n38018 , n205160 , n205294 );
buf ( n205296 , n38018 );
buf ( n205297 , n205296 );
nor ( n38021 , n205157 , n205297 );
buf ( n205299 , n38021 );
buf ( n205300 , n205299 );
nand ( n38024 , n205147 , n205300 );
buf ( n205302 , n38024 );
buf ( n205303 , n205302 );
nor ( n38027 , n205121 , n205303 );
buf ( n205305 , n38027 );
buf ( n205306 , n205305 );
and ( n38030 , n205285 , n205291 );
buf ( n205308 , n38030 );
buf ( n205309 , n205308 );
xor ( n38033 , n205222 , n205227 );
and ( n38034 , n38033 , n205269 );
and ( n38035 , n205222 , n205227 );
or ( n38036 , n38034 , n38035 );
buf ( n205314 , n38036 );
buf ( n205315 , n205314 );
and ( n38039 , n185552 , n185553 );
buf ( n205317 , n38039 );
buf ( n205318 , n205317 );
buf ( n205319 , n205241 );
not ( n38043 , n205319 );
buf ( n205321 , n177819 );
not ( n38045 , n205321 );
or ( n38046 , n38043 , n38045 );
buf ( n205324 , n800 );
buf ( n205325 , n773 );
xnor ( n38049 , n205324 , n205325 );
buf ( n205327 , n38049 );
buf ( n205328 , n205327 );
not ( n38052 , n205328 );
buf ( n205330 , n170972 );
nand ( n38054 , n38052 , n205330 );
buf ( n205332 , n38054 );
buf ( n205333 , n205332 );
nand ( n38057 , n38046 , n205333 );
buf ( n205335 , n38057 );
buf ( n205336 , n205335 );
xor ( n38060 , n205318 , n205336 );
buf ( n205338 , n205192 );
not ( n38062 , n205338 );
buf ( n205340 , n181588 );
not ( n38064 , n205340 );
or ( n38065 , n38062 , n38064 );
buf ( n205343 , n181594 );
buf ( n205344 , n806 );
nand ( n38068 , n205343 , n205344 );
buf ( n205346 , n38068 );
buf ( n205347 , n205346 );
nand ( n38071 , n38065 , n205347 );
buf ( n205349 , n38071 );
buf ( n205350 , n205349 );
xor ( n38074 , n38060 , n205350 );
buf ( n205352 , n38074 );
buf ( n205353 , n205352 );
xor ( n38077 , n205175 , n205199 );
and ( n38078 , n38077 , n205217 );
and ( n38079 , n205175 , n205199 );
or ( n38080 , n38078 , n38079 );
buf ( n205358 , n38080 );
buf ( n205359 , n205358 );
xor ( n38083 , n205353 , n205359 );
buf ( n205361 , n205259 );
not ( n38085 , n205361 );
buf ( n205363 , n183183 );
not ( n38087 , n205363 );
or ( n38088 , n38085 , n38087 );
buf ( n205366 , n178447 );
buf ( n205367 , n769 );
buf ( n205368 , n804 );
xor ( n38092 , n205367 , n205368 );
buf ( n205370 , n38092 );
buf ( n205371 , n205370 );
nand ( n38095 , n205366 , n205371 );
buf ( n205373 , n38095 );
buf ( n205374 , n205373 );
nand ( n38098 , n38088 , n205374 );
buf ( n205376 , n38098 );
buf ( n205377 , n205376 );
not ( n38101 , n205377 );
buf ( n205379 , n38101 );
buf ( n205380 , n205379 );
buf ( n205381 , n205210 );
not ( n38105 , n205381 );
buf ( n205383 , n170419 );
not ( n38107 , n205383 );
or ( n38108 , n38105 , n38107 );
buf ( n205386 , n168870 );
buf ( n205387 , n771 );
buf ( n205388 , n802 );
xor ( n38112 , n205387 , n205388 );
buf ( n205390 , n38112 );
buf ( n205391 , n205390 );
nand ( n38115 , n205386 , n205391 );
buf ( n205393 , n38115 );
buf ( n205394 , n205393 );
nand ( n38118 , n38108 , n205394 );
buf ( n205396 , n38118 );
buf ( n205397 , n205396 );
xor ( n38121 , n205380 , n205397 );
xor ( n38122 , n205231 , n205248 );
and ( n38123 , n38122 , n205266 );
and ( n38124 , n205231 , n205248 );
or ( n38125 , n38123 , n38124 );
buf ( n205403 , n38125 );
buf ( n205404 , n205403 );
xor ( n38128 , n38121 , n205404 );
buf ( n205406 , n38128 );
buf ( n205407 , n205406 );
xor ( n38131 , n38083 , n205407 );
buf ( n205409 , n38131 );
buf ( n205410 , n205409 );
xor ( n38134 , n205315 , n205410 );
xor ( n38135 , n205172 , n205220 );
and ( n38136 , n38135 , n205272 );
and ( n38137 , n205172 , n205220 );
or ( n38138 , n38136 , n38137 );
buf ( n205416 , n38138 );
buf ( n205417 , n205416 );
xor ( n38141 , n38134 , n205417 );
buf ( n205419 , n38141 );
buf ( n205420 , n205419 );
xor ( n38144 , n205166 , n205275 );
and ( n38145 , n38144 , n205282 );
and ( n38146 , n205166 , n205275 );
or ( n38147 , n38145 , n38146 );
buf ( n205425 , n38147 );
buf ( n205426 , n205425 );
xor ( n38150 , n205420 , n205426 );
buf ( n205428 , n38150 );
buf ( n205429 , n205428 );
nor ( n38153 , n205309 , n205429 );
buf ( n205431 , n38153 );
buf ( n205432 , n205431 );
not ( n38156 , n205432 );
buf ( n205434 , n38156 );
buf ( n205435 , n205434 );
and ( n38159 , n205306 , n205435 );
buf ( n205437 , n38159 );
not ( n38161 , n205437 );
or ( n38162 , n37796 , n38161 );
not ( n38163 , n31065 );
and ( n38164 , n31748 , n31146 );
and ( n38165 , n32173 , n37707 , n37722 );
not ( n38166 , n31200 );
and ( n38167 , n31113 , n38166 );
nand ( n38168 , n38163 , n38164 , n38165 , n38167 );
not ( n38169 , n38168 );
buf ( n205447 , n38169 );
buf ( n205448 , n205437 );
and ( n38172 , n205447 , n205448 );
buf ( n205450 , n38172 );
and ( n38174 , n199278 , n205450 );
buf ( n205452 , n205434 );
not ( n38176 , n205452 );
buf ( n205454 , n205302 );
not ( n38178 , n205454 );
buf ( n205456 , n38178 );
buf ( n205457 , n205456 );
not ( n38181 , n205457 );
buf ( n205459 , n205095 );
not ( n38183 , n205459 );
not ( n38184 , n205110 );
not ( n38185 , n185033 );
or ( n38186 , n38184 , n38185 );
not ( n38187 , n205114 );
nand ( n38188 , n38187 , n37825 , n205100 );
nand ( n38189 , n38186 , n38188 );
buf ( n205467 , n38189 );
not ( n38191 , n205467 );
or ( n38192 , n38183 , n38191 );
buf ( n205470 , n205085 );
not ( n38194 , n205470 );
buf ( n205472 , n38194 );
buf ( n205473 , n205472 );
buf ( n205474 , n184982 );
buf ( n205475 , n205089 );
and ( n38199 , n205474 , n205475 );
buf ( n205477 , n38199 );
buf ( n205478 , n205477 );
and ( n38202 , n205473 , n205478 );
buf ( n205480 , n205077 );
buf ( n205481 , n205082 );
and ( n38205 , n205480 , n205481 );
buf ( n205483 , n38205 );
buf ( n205484 , n205483 );
nor ( n38208 , n38202 , n205484 );
buf ( n205486 , n38208 );
buf ( n205487 , n205486 );
nand ( n38211 , n38192 , n205487 );
buf ( n205489 , n38211 );
buf ( n205490 , n205489 );
not ( n38214 , n205490 );
or ( n38215 , n38181 , n38214 );
buf ( n205493 , n205299 );
not ( n38217 , n205493 );
buf ( n205495 , n205143 );
not ( n38219 , n205495 );
buf ( n205497 , n205132 );
not ( n38221 , n205497 );
buf ( n205499 , n205123 );
nand ( n38223 , n38221 , n205499 );
buf ( n205501 , n38223 );
buf ( n205502 , n205501 );
not ( n38226 , n205502 );
buf ( n205504 , n38226 );
buf ( n205505 , n205504 );
not ( n38229 , n205505 );
or ( n38230 , n38219 , n38229 );
nand ( n38231 , n205140 , n37860 );
buf ( n205509 , n38231 );
nand ( n38233 , n38230 , n205509 );
buf ( n205511 , n38233 );
buf ( n205512 , n205511 );
not ( n38236 , n205512 );
or ( n38237 , n38217 , n38236 );
buf ( n205515 , n37871 );
buf ( n205516 , n205153 );
and ( n38240 , n205515 , n205516 );
buf ( n205518 , n38240 );
buf ( n205519 , n205518 );
buf ( n205520 , n205296 );
not ( n38244 , n205520 );
buf ( n205522 , n38244 );
buf ( n205523 , n205522 );
and ( n38247 , n205519 , n205523 );
buf ( n205525 , n205159 );
buf ( n205526 , n205293 );
and ( n38250 , n205525 , n205526 );
buf ( n205528 , n38250 );
buf ( n205529 , n205528 );
nor ( n38253 , n38247 , n205529 );
buf ( n205531 , n38253 );
buf ( n205532 , n205531 );
nand ( n38256 , n38237 , n205532 );
buf ( n205534 , n38256 );
buf ( n205535 , n205534 );
not ( n38259 , n205535 );
buf ( n205537 , n38259 );
buf ( n205538 , n205537 );
nand ( n38262 , n38215 , n205538 );
buf ( n205540 , n38262 );
buf ( n205541 , n205540 );
not ( n38265 , n205541 );
or ( n38266 , n38176 , n38265 );
buf ( n205544 , n205308 );
buf ( n205545 , n205428 );
and ( n38269 , n205544 , n205545 );
buf ( n205547 , n38269 );
buf ( n205548 , n205547 );
not ( n38272 , n205548 );
buf ( n205550 , n38272 );
buf ( n205551 , n205550 );
nand ( n38275 , n38266 , n205551 );
buf ( n205553 , n38275 );
nor ( n38277 , n38174 , n205553 );
nand ( n38278 , n38162 , n38277 );
not ( n38279 , n38278 );
and ( n38280 , n205420 , n205426 );
buf ( n205558 , n38280 );
buf ( n205559 , n205558 );
xor ( n38283 , n205315 , n205410 );
and ( n38284 , n38283 , n205417 );
and ( n38285 , n205315 , n205410 );
or ( n38286 , n38284 , n38285 );
buf ( n205564 , n38286 );
buf ( n205565 , n205564 );
xor ( n38289 , n205380 , n205397 );
and ( n38290 , n38289 , n205404 );
and ( n38291 , n205380 , n205397 );
or ( n38292 , n38290 , n38291 );
buf ( n205570 , n38292 );
buf ( n205571 , n205570 );
xor ( n38295 , n205353 , n205359 );
and ( n38296 , n38295 , n205407 );
and ( n38297 , n205353 , n205359 );
or ( n38298 , n38296 , n38297 );
buf ( n205576 , n38298 );
buf ( n205577 , n205576 );
xor ( n38301 , n205571 , n205577 );
xor ( n38302 , n205318 , n205336 );
and ( n38303 , n38302 , n205350 );
and ( n38304 , n205318 , n205336 );
or ( n38305 , n38303 , n38304 );
buf ( n205583 , n38305 );
buf ( n205584 , n205583 );
and ( n38308 , n205238 , n205239 );
buf ( n205586 , n38308 );
buf ( n205587 , n205586 );
buf ( n205588 , n205376 );
xor ( n38312 , n205587 , n205588 );
buf ( n205590 , n802 );
buf ( n205591 , n770 );
and ( n38315 , n205590 , n205591 );
not ( n38316 , n205590 );
buf ( n205594 , n770 );
not ( n38318 , n205594 );
buf ( n205596 , n38318 );
buf ( n205597 , n205596 );
and ( n38321 , n38316 , n205597 );
nor ( n38322 , n38315 , n38321 );
buf ( n205600 , n38322 );
buf ( n205601 , n205600 );
not ( n38325 , n205601 );
buf ( n205603 , n168870 );
not ( n38327 , n205603 );
or ( n38328 , n38325 , n38327 );
buf ( n205606 , n170419 );
buf ( n205607 , n205390 );
nand ( n38331 , n205606 , n205607 );
buf ( n205609 , n38331 );
buf ( n205610 , n205609 );
nand ( n38334 , n38328 , n205610 );
buf ( n205612 , n38334 );
buf ( n205613 , n205612 );
xor ( n38337 , n38312 , n205613 );
buf ( n205615 , n38337 );
buf ( n205616 , n205615 );
xor ( n38340 , n205584 , n205616 );
buf ( n205618 , n205370 );
not ( n38342 , n205618 );
buf ( n205620 , n183183 );
not ( n38344 , n205620 );
or ( n38345 , n38342 , n38344 );
buf ( n205623 , n804 );
buf ( n205624 , n768 );
xnor ( n38348 , n205623 , n205624 );
buf ( n205626 , n38348 );
buf ( n205627 , n205626 );
not ( n38351 , n205627 );
buf ( n205629 , n178447 );
nand ( n38353 , n38351 , n205629 );
buf ( n205631 , n38353 );
buf ( n205632 , n205631 );
nand ( n38356 , n38345 , n205632 );
buf ( n205634 , n38356 );
buf ( n205635 , n205634 );
buf ( n205636 , n181594 );
buf ( n205637 , n181588 );
or ( n38361 , n205636 , n205637 );
buf ( n205639 , n806 );
nand ( n38363 , n38361 , n205639 );
buf ( n205641 , n38363 );
buf ( n205642 , n205641 );
xor ( n38366 , n205635 , n205642 );
buf ( n205644 , n177819 );
not ( n38368 , n205644 );
buf ( n205646 , n38368 );
buf ( n205647 , n205646 );
buf ( n205648 , n205327 );
or ( n38372 , n205647 , n205648 );
buf ( n205650 , n170972 );
not ( n38374 , n205650 );
buf ( n205652 , n38374 );
buf ( n205653 , n205652 );
buf ( n205654 , n800 );
buf ( n205655 , n772 );
xor ( n38379 , n205654 , n205655 );
buf ( n205657 , n38379 );
buf ( n205658 , n205657 );
not ( n38382 , n205658 );
buf ( n205660 , n38382 );
buf ( n205661 , n205660 );
or ( n38385 , n205653 , n205661 );
nand ( n38386 , n38372 , n38385 );
buf ( n205664 , n38386 );
buf ( n205665 , n205664 );
xor ( n38389 , n38366 , n205665 );
buf ( n205667 , n38389 );
buf ( n205668 , n205667 );
xor ( n38392 , n38340 , n205668 );
buf ( n205670 , n38392 );
buf ( n205671 , n205670 );
xor ( n38395 , n38301 , n205671 );
buf ( n205673 , n38395 );
buf ( n205674 , n205673 );
xor ( n38398 , n205565 , n205674 );
buf ( n205676 , n38398 );
buf ( n205677 , n205676 );
nor ( n38401 , n205559 , n205677 );
buf ( n205679 , n38401 );
buf ( n205680 , n205679 );
not ( n38404 , n205680 );
buf ( n205682 , n38404 );
buf ( n205683 , n205682 );
buf ( n205684 , n205558 );
buf ( n205685 , n205676 );
nand ( n38409 , n205684 , n205685 );
buf ( n205687 , n38409 );
buf ( n205688 , n205687 );
nand ( n38412 , n205683 , n205688 );
buf ( n205690 , n38412 );
not ( n38414 , n205690 );
nor ( n38415 , n38414 , n831 );
nand ( n38416 , n38279 , n38415 );
buf ( n205694 , n205284 );
buf ( n205695 , n205290 );
and ( n38419 , n205694 , n205695 );
buf ( n205697 , n38419 );
buf ( n205698 , n205697 );
buf ( n205699 , n205419 );
buf ( n205700 , n205425 );
xor ( n38424 , n205699 , n205700 );
buf ( n205702 , n38424 );
buf ( n205703 , n205702 );
nor ( n38427 , n205698 , n205703 );
buf ( n205705 , n38427 );
buf ( n205706 , n205705 );
not ( n38430 , n205706 );
buf ( n205708 , n38430 );
not ( n38432 , n205708 );
buf ( n205710 , n185406 );
buf ( n205711 , n185673 );
xor ( n38435 , n205290 , n205284 );
buf ( n205713 , n38435 );
and ( n38437 , n185662 , n185668 );
buf ( n205715 , n38437 );
buf ( n205716 , n205715 );
nor ( n38440 , n205713 , n205716 );
buf ( n205718 , n38440 );
buf ( n205719 , n205718 );
nor ( n38443 , n205711 , n205719 );
buf ( n205721 , n38443 );
buf ( n205722 , n205721 );
nand ( n38446 , n205710 , n205722 );
buf ( n205724 , n38446 );
buf ( n205725 , n205724 );
not ( n38449 , n205725 );
buf ( n205727 , n38449 );
not ( n38451 , n205727 );
not ( n38452 , n185491 );
or ( n38453 , n38451 , n38452 );
buf ( n205731 , n205721 );
not ( n38455 , n205731 );
buf ( n205733 , n185519 );
not ( n38457 , n205733 );
or ( n38458 , n38455 , n38457 );
buf ( n205736 , n185680 );
buf ( n205737 , n205718 );
nor ( n38461 , n205736 , n205737 );
buf ( n205739 , n38461 );
buf ( n205740 , n205739 );
buf ( n205741 , n205715 );
buf ( n205742 , n38435 );
and ( n38466 , n205741 , n205742 );
buf ( n205744 , n38466 );
buf ( n205745 , n205744 );
nor ( n38469 , n205740 , n205745 );
buf ( n205747 , n38469 );
buf ( n205748 , n205747 );
nand ( n38472 , n38458 , n205748 );
buf ( n205750 , n38472 );
buf ( n205751 , n205750 );
not ( n38475 , n205751 );
buf ( n205753 , n38475 );
nand ( n38477 , n38453 , n205753 );
not ( n38478 , n38477 );
or ( n38479 , n38432 , n38478 );
buf ( n205757 , n205697 );
buf ( n205758 , n205702 );
nand ( n38482 , n205757 , n205758 );
buf ( n205760 , n38482 );
nand ( n38484 , n38479 , n205760 );
not ( n38485 , n38484 );
buf ( n205763 , n184143 );
buf ( n205764 , n185042 );
buf ( n205765 , n205724 );
nor ( n38489 , n205764 , n205765 );
buf ( n205767 , n38489 );
buf ( n205768 , n205767 );
buf ( n205769 , n205708 );
and ( n38493 , n205768 , n205769 );
buf ( n205771 , n38493 );
buf ( n205772 , n205771 );
nand ( n38496 , n205763 , n205772 );
buf ( n205774 , n38496 );
nand ( n38498 , n177727 , n185881 , n205771 );
nand ( n38499 , n38485 , n205774 , n38498 );
not ( n38500 , n38499 );
and ( n38501 , n205699 , n205700 );
buf ( n205779 , n38501 );
buf ( n205780 , n205779 );
buf ( n205781 , n205564 );
buf ( n205782 , n205673 );
xor ( n38506 , n205781 , n205782 );
buf ( n205784 , n38506 );
buf ( n205785 , n205784 );
nor ( n38509 , n205780 , n205785 );
buf ( n205787 , n38509 );
buf ( n205788 , n205787 );
not ( n38512 , n205788 );
buf ( n205790 , n38512 );
buf ( n205791 , n205790 );
buf ( n205792 , n205779 );
buf ( n205793 , n205784 );
nand ( n38517 , n205792 , n205793 );
buf ( n205795 , n38517 );
buf ( n205796 , n205795 );
nand ( n38520 , n205791 , n205796 );
buf ( n205798 , n38520 );
and ( n38522 , n205798 , n831 );
nand ( n38523 , n38500 , n38522 );
buf ( n205801 , n205798 );
not ( n38525 , n205801 );
buf ( n205803 , n38525 );
nand ( n38527 , n38499 , n205803 , n831 );
nor ( n38528 , n205690 , n831 );
nand ( n38529 , n38278 , n38528 );
nand ( n38530 , n38416 , n38523 , n38527 , n38529 );
not ( n38531 , n38530 );
buf ( n38532 , n38531 );
buf ( n38533 , n38532 );
buf ( n205811 , n170419 );
not ( n38535 , n205811 );
buf ( n205813 , n38535 );
buf ( n205814 , n205813 );
buf ( n205815 , n768 );
buf ( n205816 , n802 );
xnor ( n38540 , n205815 , n205816 );
buf ( n205818 , n38540 );
buf ( n205819 , n205818 );
or ( n38543 , n205814 , n205819 );
buf ( n205821 , n168870 );
not ( n38545 , n205821 );
buf ( n205823 , n38545 );
buf ( n205824 , n205823 );
buf ( n205825 , n802 );
not ( n38549 , n205825 );
buf ( n205827 , n38549 );
buf ( n205828 , n205827 );
or ( n38552 , n205824 , n205828 );
nand ( n38553 , n38543 , n38552 );
buf ( n205831 , n38553 );
buf ( n205832 , n205831 );
buf ( n205833 , n770 );
buf ( n205834 , n800 );
and ( n38558 , n205833 , n205834 );
buf ( n205836 , n38558 );
buf ( n205837 , n205836 );
buf ( n205838 , n205646 );
buf ( n205839 , n800 );
not ( n38563 , n205839 );
buf ( n205841 , n38563 );
buf ( n205842 , n205841 );
buf ( n205843 , n769 );
and ( n38567 , n205842 , n205843 );
buf ( n205845 , n178502 );
buf ( n205846 , n800 );
and ( n38570 , n205845 , n205846 );
nor ( n38571 , n38567 , n38570 );
buf ( n205849 , n38571 );
buf ( n205850 , n205849 );
or ( n38574 , n205838 , n205850 );
buf ( n205852 , n205652 );
buf ( n205853 , n205841 );
buf ( n205854 , n768 );
and ( n38578 , n205853 , n205854 );
buf ( n205856 , n205188 );
buf ( n205857 , n800 );
and ( n38581 , n205856 , n205857 );
nor ( n38582 , n38578 , n38581 );
buf ( n205860 , n38582 );
buf ( n205861 , n205860 );
or ( n38585 , n205852 , n205861 );
nand ( n38586 , n38574 , n38585 );
buf ( n205864 , n38586 );
buf ( n205865 , n205864 );
xor ( n38589 , n205837 , n205865 );
buf ( n205867 , n170419 );
buf ( n205868 , n168870 );
or ( n38592 , n205867 , n205868 );
buf ( n205870 , n802 );
nand ( n38594 , n38592 , n205870 );
buf ( n205872 , n38594 );
buf ( n205873 , n205872 );
xor ( n38597 , n38589 , n205873 );
buf ( n205875 , n38597 );
buf ( n205876 , n205875 );
xor ( n38600 , n205832 , n205876 );
buf ( n205878 , n771 );
buf ( n205879 , n800 );
and ( n38603 , n205878 , n205879 );
buf ( n205881 , n38603 );
buf ( n205882 , n205881 );
buf ( n205883 , n205646 );
buf ( n205884 , n205841 );
buf ( n205885 , n770 );
and ( n38609 , n205884 , n205885 );
buf ( n205887 , n205596 );
buf ( n205888 , n800 );
and ( n38612 , n205887 , n205888 );
nor ( n38613 , n38609 , n38612 );
buf ( n205891 , n38613 );
buf ( n205892 , n205891 );
or ( n38616 , n205883 , n205892 );
buf ( n205894 , n205652 );
buf ( n205895 , n205849 );
or ( n38619 , n205894 , n205895 );
nand ( n38620 , n38616 , n38619 );
buf ( n205898 , n38620 );
buf ( n205899 , n205898 );
xor ( n38623 , n205882 , n205899 );
buf ( n205901 , n205831 );
not ( n38625 , n205901 );
buf ( n205903 , n38625 );
buf ( n205904 , n205903 );
and ( n38628 , n38623 , n205904 );
and ( n38629 , n205882 , n205899 );
or ( n38630 , n38628 , n38629 );
buf ( n205908 , n38630 );
buf ( n205909 , n205908 );
xor ( n38633 , n38600 , n205909 );
buf ( n205911 , n38633 );
buf ( n205912 , n205911 );
and ( n38636 , n205654 , n205655 );
buf ( n205914 , n38636 );
buf ( n205915 , n205914 );
buf ( n205916 , n178447 );
not ( n38640 , n205916 );
buf ( n205918 , n38640 );
buf ( n205919 , n205918 );
not ( n38643 , n205919 );
buf ( n205921 , n183183 );
not ( n38645 , n205921 );
buf ( n205923 , n38645 );
buf ( n205924 , n205923 );
not ( n38648 , n205924 );
or ( n38649 , n38643 , n38648 );
buf ( n205927 , n804 );
nand ( n38651 , n38649 , n205927 );
buf ( n205929 , n38651 );
buf ( n205930 , n205929 );
xor ( n38654 , n205915 , n205930 );
buf ( n205932 , n205813 );
buf ( n205933 , n769 );
buf ( n205934 , n802 );
xnor ( n38658 , n205933 , n205934 );
buf ( n205936 , n38658 );
buf ( n205937 , n205936 );
or ( n38661 , n205932 , n205937 );
buf ( n205939 , n205823 );
buf ( n205940 , n205818 );
or ( n38664 , n205939 , n205940 );
nand ( n38665 , n38661 , n38664 );
buf ( n205943 , n38665 );
buf ( n205944 , n205943 );
and ( n38668 , n38654 , n205944 );
and ( n38669 , n205915 , n205930 );
or ( n38670 , n38668 , n38669 );
buf ( n205948 , n38670 );
buf ( n205949 , n205948 );
xor ( n38673 , n205882 , n205899 );
xor ( n38674 , n38673 , n205904 );
buf ( n205952 , n38674 );
buf ( n205953 , n205952 );
xor ( n38677 , n205949 , n205953 );
buf ( n205955 , n205923 );
buf ( n205956 , n205626 );
or ( n38680 , n205955 , n205956 );
buf ( n205958 , n205918 );
buf ( n205959 , n804 );
not ( n38683 , n205959 );
buf ( n205961 , n38683 );
buf ( n205962 , n205961 );
or ( n38686 , n205958 , n205962 );
nand ( n38687 , n38680 , n38686 );
buf ( n205965 , n38687 );
buf ( n205966 , n205965 );
buf ( n205967 , n205646 );
buf ( n205968 , n800 );
buf ( n205969 , n771 );
xnor ( n38693 , n205968 , n205969 );
buf ( n205971 , n38693 );
buf ( n205972 , n205971 );
or ( n38696 , n205967 , n205972 );
buf ( n205974 , n205652 );
buf ( n205975 , n205891 );
or ( n38699 , n205974 , n205975 );
nand ( n38700 , n38696 , n38699 );
buf ( n205978 , n38700 );
buf ( n205979 , n205978 );
xor ( n38703 , n205966 , n205979 );
buf ( n205981 , n773 );
buf ( n205982 , n800 );
and ( n38706 , n205981 , n205982 );
buf ( n205984 , n38706 );
buf ( n205985 , n205984 );
buf ( n205986 , n205657 );
not ( n38710 , n205986 );
buf ( n205988 , n177819 );
not ( n38712 , n205988 );
or ( n38713 , n38710 , n38712 );
buf ( n205991 , n205971 );
not ( n38715 , n205991 );
buf ( n205993 , n170972 );
nand ( n38717 , n38715 , n205993 );
buf ( n205995 , n38717 );
buf ( n205996 , n205995 );
nand ( n38720 , n38713 , n205996 );
buf ( n205998 , n38720 );
buf ( n205999 , n205998 );
xor ( n38723 , n205985 , n205999 );
buf ( n206001 , n205600 );
not ( n38725 , n206001 );
buf ( n206003 , n170419 );
not ( n38727 , n206003 );
or ( n38728 , n38725 , n38727 );
buf ( n206006 , n205936 );
not ( n38730 , n206006 );
buf ( n206008 , n168870 );
nand ( n38732 , n38730 , n206008 );
buf ( n206010 , n38732 );
buf ( n206011 , n206010 );
nand ( n38735 , n38728 , n206011 );
buf ( n206013 , n38735 );
buf ( n206014 , n206013 );
and ( n38738 , n38723 , n206014 );
and ( n38739 , n205985 , n205999 );
or ( n38740 , n38738 , n38739 );
buf ( n206018 , n38740 );
buf ( n206019 , n206018 );
and ( n38743 , n38703 , n206019 );
and ( n38744 , n205966 , n205979 );
or ( n38745 , n38743 , n38744 );
buf ( n206023 , n38745 );
buf ( n206024 , n206023 );
and ( n38748 , n38677 , n206024 );
and ( n38749 , n205949 , n205953 );
or ( n38750 , n38748 , n38749 );
buf ( n206028 , n38750 );
buf ( n206029 , n206028 );
and ( n38753 , n205912 , n206029 );
buf ( n206031 , n38753 );
buf ( n206032 , n206031 );
buf ( n206033 , n769 );
buf ( n206034 , n800 );
nand ( n38758 , n206033 , n206034 );
buf ( n206036 , n38758 );
buf ( n206037 , n206036 );
buf ( n206038 , n205646 );
buf ( n206039 , n205860 );
or ( n38763 , n206038 , n206039 );
buf ( n206041 , n205652 );
buf ( n206042 , n205841 );
or ( n38766 , n206041 , n206042 );
nand ( n38767 , n38763 , n38766 );
buf ( n206045 , n38767 );
buf ( n206046 , n206045 );
xor ( n38770 , n206037 , n206046 );
xor ( n38771 , n205837 , n205865 );
and ( n38772 , n38771 , n205873 );
and ( n38773 , n205837 , n205865 );
or ( n38774 , n38772 , n38773 );
buf ( n206052 , n38774 );
buf ( n206053 , n206052 );
xor ( n38777 , n38770 , n206053 );
buf ( n206055 , n38777 );
buf ( n206056 , n206055 );
xor ( n38780 , n205832 , n205876 );
and ( n38781 , n38780 , n205909 );
and ( n38782 , n205832 , n205876 );
or ( n38783 , n38781 , n38782 );
buf ( n206061 , n38783 );
buf ( n206062 , n206061 );
xor ( n38786 , n206056 , n206062 );
buf ( n206064 , n38786 );
buf ( n206065 , n206064 );
and ( n38789 , n206032 , n206065 );
buf ( n206067 , n38789 );
buf ( n206068 , n206067 );
not ( n38792 , n206068 );
buf ( n206070 , n206031 );
buf ( n206071 , n206064 );
or ( n38795 , n206070 , n206071 );
buf ( n206073 , n38795 );
buf ( n206074 , n206073 );
nand ( n38798 , n38792 , n206074 );
buf ( n206076 , n38798 );
not ( n38800 , n206076 );
buf ( n206078 , n177727 );
buf ( n38802 , n206078 );
buf ( n206080 , n38802 );
buf ( n206081 , n206080 );
buf ( n206082 , n185446 );
buf ( n206083 , n205767 );
buf ( n38807 , n206083 );
buf ( n206085 , n38807 );
buf ( n206086 , n206085 );
xor ( n38810 , n205915 , n205930 );
xor ( n38811 , n38810 , n205944 );
buf ( n206089 , n38811 );
buf ( n206090 , n206089 );
xor ( n38814 , n205966 , n205979 );
xor ( n38815 , n38814 , n206019 );
buf ( n206093 , n38815 );
buf ( n206094 , n206093 );
xor ( n38818 , n206090 , n206094 );
buf ( n206096 , n205965 );
not ( n38820 , n206096 );
buf ( n206098 , n38820 );
buf ( n206099 , n206098 );
xor ( n38823 , n205985 , n205999 );
xor ( n38824 , n38823 , n206014 );
buf ( n206102 , n38824 );
buf ( n206103 , n206102 );
xor ( n38827 , n206099 , n206103 );
xor ( n38828 , n205635 , n205642 );
and ( n38829 , n38828 , n205665 );
and ( n38830 , n205635 , n205642 );
or ( n38831 , n38829 , n38830 );
buf ( n206109 , n38831 );
buf ( n206110 , n206109 );
and ( n38834 , n38827 , n206110 );
and ( n38835 , n206099 , n206103 );
or ( n38836 , n38834 , n38835 );
buf ( n206114 , n38836 );
buf ( n206115 , n206114 );
xor ( n38839 , n38818 , n206115 );
buf ( n206117 , n38839 );
buf ( n206118 , n206117 );
xor ( n38842 , n205587 , n205588 );
and ( n38843 , n38842 , n205613 );
and ( n38844 , n205587 , n205588 );
or ( n38845 , n38843 , n38844 );
buf ( n206123 , n38845 );
buf ( n206124 , n206123 );
xor ( n38848 , n206099 , n206103 );
xor ( n38849 , n38848 , n206110 );
buf ( n206127 , n38849 );
buf ( n206128 , n206127 );
xor ( n38852 , n206124 , n206128 );
xor ( n38853 , n205584 , n205616 );
and ( n38854 , n38853 , n205668 );
and ( n38855 , n205584 , n205616 );
or ( n38856 , n38854 , n38855 );
buf ( n206134 , n38856 );
buf ( n206135 , n206134 );
and ( n38859 , n38852 , n206135 );
and ( n38860 , n206124 , n206128 );
or ( n38861 , n38859 , n38860 );
buf ( n206139 , n38861 );
buf ( n206140 , n206139 );
and ( n38864 , n206118 , n206140 );
buf ( n206142 , n38864 );
buf ( n206143 , n206142 );
xor ( n38867 , n205949 , n205953 );
xor ( n38868 , n38867 , n206024 );
buf ( n206146 , n38868 );
buf ( n206147 , n206146 );
xor ( n38871 , n206090 , n206094 );
and ( n38872 , n38871 , n206115 );
and ( n38873 , n206090 , n206094 );
or ( n38874 , n38872 , n38873 );
buf ( n206152 , n38874 );
buf ( n206153 , n206152 );
xor ( n38877 , n206147 , n206153 );
buf ( n206155 , n38877 );
buf ( n206156 , n206155 );
nor ( n38880 , n206143 , n206156 );
buf ( n206158 , n38880 );
buf ( n206159 , n206158 );
and ( n38883 , n206147 , n206153 );
buf ( n206161 , n38883 );
buf ( n206162 , n206161 );
xor ( n38886 , n205912 , n206029 );
buf ( n206164 , n38886 );
buf ( n206165 , n206164 );
nor ( n38889 , n206162 , n206165 );
buf ( n206167 , n38889 );
buf ( n206168 , n206167 );
nor ( n38892 , n206159 , n206168 );
buf ( n206170 , n38892 );
buf ( n206171 , n206170 );
not ( n38895 , n206171 );
xor ( n38896 , n206124 , n206128 );
xor ( n38897 , n38896 , n206135 );
buf ( n206175 , n38897 );
buf ( n206176 , n206175 );
xor ( n38900 , n205571 , n205577 );
and ( n38901 , n38900 , n205671 );
and ( n38902 , n205571 , n205577 );
or ( n38903 , n38901 , n38902 );
buf ( n206181 , n38903 );
buf ( n206182 , n206181 );
xor ( n38906 , n206176 , n206182 );
buf ( n206184 , n38906 );
buf ( n206185 , n206184 );
and ( n38909 , n205781 , n205782 );
buf ( n206187 , n38909 );
buf ( n206188 , n206187 );
nor ( n38912 , n206185 , n206188 );
buf ( n206190 , n38912 );
buf ( n206191 , n206190 );
and ( n38915 , n206176 , n206182 );
buf ( n206193 , n38915 );
buf ( n206194 , n206193 );
xor ( n38918 , n206118 , n206140 );
buf ( n206196 , n38918 );
buf ( n206197 , n206196 );
nor ( n38921 , n206194 , n206197 );
buf ( n206199 , n38921 );
buf ( n206200 , n206199 );
nor ( n38924 , n206191 , n206200 );
buf ( n206202 , n38924 );
buf ( n206203 , n205787 );
buf ( n206204 , n205705 );
nor ( n38928 , n206203 , n206204 );
buf ( n206206 , n38928 );
nand ( n38930 , n206202 , n206206 );
buf ( n206208 , n38930 );
nor ( n38932 , n38895 , n206208 );
buf ( n206210 , n38932 );
buf ( n206211 , n206210 );
nand ( n38935 , n206086 , n206211 );
buf ( n206213 , n38935 );
buf ( n206214 , n206213 );
nor ( n38938 , n206082 , n206214 );
buf ( n206216 , n38938 );
buf ( n206217 , n206216 );
nand ( n38941 , n206081 , n206217 );
buf ( n206219 , n38941 );
not ( n38943 , n206213 );
nand ( n38944 , n38943 , n185895 );
buf ( n206222 , n206210 );
not ( n38946 , n206222 );
buf ( n206224 , n38477 );
not ( n38948 , n206224 );
or ( n38949 , n38946 , n38948 );
not ( n38950 , n206202 );
buf ( n206228 , n205790 );
not ( n38952 , n206228 );
buf ( n206230 , n205760 );
not ( n38954 , n206230 );
buf ( n206232 , n38954 );
buf ( n206233 , n206232 );
not ( n38957 , n206233 );
or ( n38958 , n38952 , n38957 );
buf ( n206236 , n205795 );
nand ( n38960 , n38958 , n206236 );
buf ( n206238 , n38960 );
not ( n38962 , n206238 );
or ( n38963 , n38950 , n38962 );
buf ( n206241 , n206184 );
buf ( n206242 , n206187 );
and ( n38966 , n206241 , n206242 );
buf ( n206244 , n38966 );
buf ( n206245 , n206244 );
buf ( n206246 , n206199 );
not ( n38970 , n206246 );
buf ( n206248 , n38970 );
buf ( n206249 , n206248 );
and ( n38973 , n206245 , n206249 );
buf ( n206251 , n206193 );
buf ( n206252 , n206196 );
nand ( n38976 , n206251 , n206252 );
buf ( n206254 , n38976 );
buf ( n206255 , n206254 );
not ( n38979 , n206255 );
buf ( n206257 , n38979 );
buf ( n206258 , n206257 );
nor ( n38982 , n38973 , n206258 );
buf ( n206260 , n38982 );
nand ( n38984 , n38963 , n206260 );
and ( n38985 , n206170 , n38984 );
buf ( n206263 , n206142 );
buf ( n206264 , n206155 );
nand ( n38988 , n206263 , n206264 );
buf ( n206266 , n38988 );
buf ( n206267 , n206266 );
buf ( n206268 , n206167 );
or ( n38992 , n206267 , n206268 );
buf ( n206270 , n206161 );
buf ( n206271 , n206164 );
nand ( n38995 , n206270 , n206271 );
buf ( n206273 , n38995 );
buf ( n206274 , n206273 );
nand ( n38998 , n38992 , n206274 );
buf ( n206276 , n38998 );
nor ( n39000 , n38985 , n206276 );
buf ( n206278 , n39000 );
nand ( n39002 , n38949 , n206278 );
buf ( n206280 , n39002 );
buf ( n206281 , n206280 );
not ( n39005 , n206281 );
buf ( n206283 , n39005 );
nand ( n39007 , n206219 , n38944 , n206283 );
not ( n39008 , n39007 );
or ( n39009 , n38800 , n39008 );
not ( n39010 , n206076 );
and ( n39011 , n206283 , n39010 );
nand ( n39012 , n39011 , n206219 , n38944 );
nand ( n39013 , n39009 , n39012 );
nor ( n39014 , n38533 , n39013 );
buf ( n206292 , n38477 );
buf ( n39016 , n206292 );
buf ( n206294 , n39016 );
not ( n39018 , n206294 );
buf ( n206296 , n185881 );
buf ( n206297 , n206085 );
and ( n39021 , n206296 , n206297 );
buf ( n206299 , n39021 );
nand ( n39023 , n177740 , n206299 );
buf ( n206301 , n185895 );
buf ( n206302 , n206085 );
nand ( n39026 , n206301 , n206302 );
buf ( n206304 , n39026 );
nand ( n39028 , n39018 , n39023 , n206304 );
buf ( n206306 , n205708 );
buf ( n206307 , n205760 );
nand ( n39031 , n206306 , n206307 );
buf ( n206309 , n39031 );
buf ( n206310 , n206309 );
not ( n39034 , n206310 );
buf ( n206312 , n39034 );
and ( n39036 , n206312 , n831 );
and ( n39037 , n39028 , n39036 );
not ( n39038 , n39028 );
and ( n39039 , n206309 , n831 );
and ( n39040 , n39038 , n39039 );
nor ( n39041 , n39037 , n39040 );
buf ( n206319 , n205069 );
not ( n39043 , n206319 );
buf ( n206321 , n39043 );
buf ( n206322 , n206321 );
buf ( n206323 , n205305 );
buf ( n39047 , n206323 );
buf ( n206325 , n39047 );
buf ( n206326 , n206325 );
nand ( n39050 , n206322 , n206326 );
buf ( n206328 , n39050 );
not ( n39052 , n206328 );
buf ( n206330 , n205434 );
buf ( n206331 , n205550 );
nand ( n39055 , n206330 , n206331 );
buf ( n206333 , n39055 );
nand ( n39057 , n39052 , n206333 );
buf ( n206335 , n199278 );
buf ( n206336 , n38169 );
buf ( n206337 , n206325 );
and ( n39061 , n206336 , n206337 );
buf ( n206339 , n39061 );
buf ( n206340 , n206339 );
nand ( n39064 , n206335 , n206340 );
buf ( n206342 , n39064 );
not ( n39066 , n206342 );
nand ( n39067 , n39066 , n206333 );
buf ( n206345 , n205456 );
not ( n39069 , n206345 );
buf ( n206347 , n205489 );
not ( n39071 , n206347 );
or ( n39072 , n39069 , n39071 );
buf ( n206350 , n205537 );
nand ( n39074 , n39072 , n206350 );
buf ( n206352 , n39074 );
buf ( n206353 , n206352 );
not ( n39077 , n206353 );
buf ( n206355 , n39077 );
buf ( n206356 , n206333 );
not ( n39080 , n206356 );
buf ( n206358 , n39080 );
and ( n39082 , n206355 , n206358 );
nand ( n39083 , n206328 , n206342 , n39082 );
or ( n39084 , n206355 , n206358 );
and ( n39085 , n39084 , n2047 );
nand ( n39086 , n39057 , n39067 , n39083 , n39085 );
nand ( n39087 , n39041 , n39086 );
not ( n39088 , n39087 );
buf ( n39089 , n39088 );
buf ( n206367 , n185446 );
buf ( n206368 , n206085 );
buf ( n206369 , n38930 );
buf ( n206370 , n206158 );
nor ( n39094 , n206369 , n206370 );
buf ( n206372 , n39094 );
buf ( n206373 , n206372 );
nand ( n39097 , n206368 , n206373 );
buf ( n206375 , n39097 );
buf ( n206376 , n206375 );
nor ( n39100 , n206367 , n206376 );
buf ( n206378 , n39100 );
nand ( n39102 , n206378 , n206080 );
buf ( n206380 , n206375 );
not ( n39104 , n206380 );
buf ( n206382 , n185895 );
nand ( n39106 , n39104 , n206382 );
buf ( n206384 , n39106 );
buf ( n206385 , n206372 );
buf ( n206386 , n38477 );
and ( n39110 , n206385 , n206386 );
buf ( n206388 , n206158 );
not ( n39112 , n206388 );
buf ( n206390 , n39112 );
buf ( n206391 , n206390 );
not ( n39115 , n206391 );
buf ( n206393 , n38984 );
not ( n39117 , n206393 );
or ( n39118 , n39115 , n39117 );
buf ( n206396 , n206266 );
nand ( n39120 , n39118 , n206396 );
buf ( n206398 , n39120 );
buf ( n206399 , n206398 );
nor ( n39123 , n39110 , n206399 );
buf ( n206401 , n39123 );
nand ( n39125 , n39102 , n206384 , n206401 );
not ( n39126 , n206167 );
nand ( n39127 , n39126 , n206273 );
not ( n39128 , n39127 );
and ( n39129 , n39125 , n39128 );
not ( n39130 , n39125 );
and ( n39131 , n39130 , n39127 );
nor ( n39132 , n39129 , n39131 );
nor ( n39133 , n39089 , n39132 );
nor ( n39134 , n39014 , n39133 );
not ( n39135 , n39134 );
not ( n39136 , n831 );
buf ( n206414 , n205767 );
buf ( n206415 , n206206 );
not ( n39139 , n206415 );
buf ( n206417 , n39139 );
buf ( n206418 , n206417 );
buf ( n206419 , n206190 );
nor ( n39143 , n206418 , n206419 );
buf ( n206421 , n39143 );
buf ( n206422 , n206421 );
and ( n39146 , n206414 , n206422 );
buf ( n206424 , n39146 );
nand ( n39148 , n177727 , n185881 , n206424 );
buf ( n206426 , n39148 );
buf ( n206427 , n185895 );
buf ( n206428 , n206424 );
nand ( n39152 , n206427 , n206428 );
buf ( n206430 , n39152 );
buf ( n206431 , n206430 );
buf ( n206432 , n206421 );
not ( n39156 , n206432 );
buf ( n206434 , n38477 );
not ( n39158 , n206434 );
or ( n39159 , n39156 , n39158 );
buf ( n206437 , n206238 );
buf ( n206438 , n206190 );
not ( n39162 , n206438 );
buf ( n206440 , n39162 );
buf ( n206441 , n206440 );
and ( n39165 , n206437 , n206441 );
buf ( n206443 , n206244 );
nor ( n39167 , n39165 , n206443 );
buf ( n206445 , n39167 );
buf ( n206446 , n206445 );
nand ( n39170 , n39159 , n206446 );
buf ( n206448 , n39170 );
buf ( n206449 , n206448 );
not ( n39173 , n206449 );
buf ( n206451 , n39173 );
buf ( n206452 , n206451 );
nand ( n39176 , n206426 , n206431 , n206452 );
buf ( n206454 , n39176 );
buf ( n206455 , n206248 );
buf ( n206456 , n206254 );
nand ( n39180 , n206455 , n206456 );
buf ( n206458 , n39180 );
buf ( n206459 , n206458 );
not ( n39183 , n206459 );
buf ( n206461 , n39183 );
and ( n39185 , n206454 , n206461 );
not ( n39186 , n206454 );
and ( n39187 , n39186 , n206458 );
nor ( n39188 , n39185 , n39187 );
not ( n39189 , n39188 );
or ( n39190 , n39136 , n39189 );
buf ( n206468 , n206175 );
buf ( n206469 , n206181 );
and ( n39193 , n206468 , n206469 );
buf ( n206471 , n39193 );
buf ( n206472 , n206471 );
buf ( n206473 , n206117 );
buf ( n206474 , n206139 );
xor ( n39198 , n206473 , n206474 );
buf ( n206476 , n39198 );
buf ( n206477 , n206476 );
nor ( n39201 , n206472 , n206477 );
buf ( n206479 , n39201 );
buf ( n206480 , n206479 );
not ( n39204 , n206480 );
buf ( n206482 , n39204 );
buf ( n206483 , n206482 );
buf ( n206484 , n206471 );
buf ( n206485 , n206476 );
nand ( n39209 , n206484 , n206485 );
buf ( n206487 , n39209 );
buf ( n206488 , n206487 );
nand ( n39212 , n206483 , n206488 );
buf ( n206490 , n39212 );
not ( n39214 , n206490 );
buf ( n206492 , n205679 );
buf ( n206493 , n205431 );
nor ( n39217 , n206492 , n206493 );
buf ( n206495 , n39217 );
buf ( n206496 , n206495 );
not ( n39220 , n206496 );
buf ( n206498 , n39220 );
buf ( n206499 , n206498 );
xor ( n39223 , n206468 , n206469 );
buf ( n206501 , n39223 );
buf ( n206502 , n206501 );
and ( n39226 , n205565 , n205674 );
buf ( n206504 , n39226 );
buf ( n206505 , n206504 );
nor ( n39229 , n206502 , n206505 );
buf ( n206507 , n39229 );
buf ( n206508 , n206507 );
nor ( n39232 , n206499 , n206508 );
buf ( n206510 , n39232 );
buf ( n206511 , n206510 );
not ( n39235 , n206511 );
buf ( n206513 , n205540 );
not ( n39237 , n206513 );
or ( n39238 , n39235 , n39237 );
buf ( n206516 , n205682 );
not ( n39240 , n206516 );
buf ( n206518 , n205547 );
not ( n39242 , n206518 );
or ( n39243 , n39240 , n39242 );
buf ( n206521 , n205687 );
nand ( n39245 , n39243 , n206521 );
buf ( n206523 , n39245 );
buf ( n206524 , n206523 );
buf ( n206525 , n206507 );
not ( n39249 , n206525 );
buf ( n206527 , n39249 );
buf ( n206528 , n206527 );
and ( n39252 , n206524 , n206528 );
buf ( n206530 , n206501 );
buf ( n206531 , n206504 );
and ( n39255 , n206530 , n206531 );
buf ( n206533 , n39255 );
buf ( n206534 , n206533 );
nor ( n39258 , n39252 , n206534 );
buf ( n206536 , n39258 );
buf ( n206537 , n206536 );
nand ( n39261 , n39238 , n206537 );
buf ( n206539 , n39261 );
not ( n39263 , n206539 );
buf ( n206541 , n205069 );
not ( n39265 , n206541 );
buf ( n206543 , n39265 );
buf ( n206544 , n206543 );
buf ( n206545 , n205305 );
buf ( n206546 , n206510 );
and ( n39270 , n206545 , n206546 );
buf ( n206548 , n39270 );
buf ( n206549 , n206548 );
nand ( n39273 , n206544 , n206549 );
buf ( n206551 , n39273 );
not ( n39275 , n38168 );
nand ( n39276 , n199278 , n39275 , n206548 );
nand ( n39277 , n39263 , n206551 , n39276 );
not ( n39278 , n39277 );
or ( n39279 , n39214 , n39278 );
not ( n39280 , n206539 );
not ( n39281 , n206490 );
nand ( n39282 , n206551 , n39280 , n39276 , n39281 );
nand ( n39283 , n39279 , n39282 );
nand ( n39284 , n39283 , n168462 );
nand ( n39285 , n39190 , n39284 );
buf ( n39286 , n39285 );
not ( n39287 , n39286 );
not ( n39288 , n39287 );
buf ( n206566 , n184143 );
buf ( n206567 , n206417 );
not ( n39291 , n206567 );
buf ( n206569 , n206085 );
nand ( n39293 , n39291 , n206569 );
buf ( n206571 , n39293 );
buf ( n206572 , n206571 );
not ( n39296 , n206572 );
buf ( n206574 , n39296 );
buf ( n206575 , n206574 );
nand ( n39299 , n206566 , n206575 );
buf ( n206577 , n39299 );
buf ( n206578 , n177727 );
buf ( n206579 , n185446 );
buf ( n206580 , n206571 );
nor ( n39304 , n206579 , n206580 );
buf ( n206582 , n39304 );
buf ( n206583 , n206582 );
nand ( n39307 , n206578 , n206583 );
buf ( n206585 , n39307 );
and ( n39309 , n206206 , n38477 );
nor ( n39310 , n39309 , n206238 );
nand ( n39311 , n206577 , n206585 , n39310 );
buf ( n206589 , n206244 );
buf ( n206590 , n206190 );
nor ( n39314 , n206589 , n206590 );
buf ( n206592 , n39314 );
xor ( n39316 , n39311 , n206592 );
not ( n39317 , n831 );
or ( n39318 , n39316 , n39317 );
buf ( n206596 , n206495 );
not ( n39320 , n206596 );
buf ( n206598 , n206352 );
not ( n39322 , n206598 );
or ( n39323 , n39320 , n39322 );
buf ( n206601 , n206523 );
not ( n39325 , n206601 );
buf ( n206603 , n39325 );
buf ( n206604 , n206603 );
nand ( n39328 , n39323 , n206604 );
buf ( n206606 , n39328 );
buf ( n206607 , n206606 );
not ( n39331 , n206607 );
buf ( n206609 , n39331 );
nor ( n39333 , n206533 , n206507 );
not ( n39334 , n39333 );
nand ( n39335 , n39334 , n39317 );
and ( n39336 , n206609 , n39335 );
buf ( n206614 , n206498 );
not ( n39338 , n206614 );
buf ( n206616 , n206325 );
nand ( n39340 , n39338 , n206616 );
buf ( n206618 , n39340 );
not ( n39342 , n206618 );
nand ( n39343 , n39342 , n206321 );
buf ( n206621 , n199278 );
buf ( n206622 , n39275 );
not ( n39346 , n206622 );
buf ( n206624 , n206618 );
nor ( n39348 , n39346 , n206624 );
buf ( n206626 , n39348 );
buf ( n206627 , n206626 );
nand ( n39351 , n206621 , n206627 );
buf ( n206629 , n39351 );
nand ( n39353 , n39336 , n39343 , n206629 );
not ( n39354 , n39343 );
nand ( n39355 , n39333 , n39317 );
nand ( n39356 , n39354 , n39355 );
not ( n39357 , n206609 );
not ( n39358 , n206629 );
or ( n39359 , n39357 , n39358 );
nand ( n39360 , n39359 , n39355 );
nand ( n39361 , n39353 , n39356 , n39360 );
nand ( n39362 , n39318 , n39361 );
not ( n39363 , n39362 );
not ( n39364 , n39363 );
not ( n39365 , n39364 );
not ( n39366 , n39365 );
buf ( n39367 , n39366 );
not ( n39368 , n39367 );
and ( n39369 , n206056 , n206062 );
buf ( n206647 , n39369 );
buf ( n206648 , n206647 );
not ( n39372 , n206648 );
xor ( n39373 , n206037 , n206046 );
and ( n39374 , n39373 , n206053 );
and ( n39375 , n206037 , n206046 );
or ( n39376 , n39374 , n39375 );
buf ( n206654 , n39376 );
buf ( n206655 , n206654 );
buf ( n206656 , n206036 );
not ( n39380 , n206656 );
buf ( n206658 , n768 );
buf ( n206659 , n800 );
nand ( n39383 , n206658 , n206659 );
buf ( n206661 , n39383 );
buf ( n206662 , n206661 );
not ( n39386 , n206662 );
buf ( n206664 , n177819 );
buf ( n206665 , n170972 );
or ( n39389 , n206664 , n206665 );
buf ( n206667 , n800 );
nand ( n39391 , n39389 , n206667 );
buf ( n206669 , n39391 );
buf ( n206670 , n206669 );
not ( n39394 , n206670 );
or ( n39395 , n39386 , n39394 );
buf ( n206673 , n206669 );
buf ( n206674 , n206661 );
or ( n39398 , n206673 , n206674 );
nand ( n39399 , n39395 , n39398 );
buf ( n206677 , n39399 );
buf ( n206678 , n206677 );
not ( n39402 , n206678 );
or ( n39403 , n39380 , n39402 );
buf ( n206681 , n206677 );
buf ( n206682 , n206036 );
or ( n39406 , n206681 , n206682 );
nand ( n39407 , n39403 , n39406 );
buf ( n206685 , n39407 );
buf ( n206686 , n206685 );
xor ( n39410 , n206655 , n206686 );
buf ( n206688 , n39410 );
buf ( n206689 , n206688 );
not ( n39413 , n206689 );
and ( n39414 , n39372 , n39413 );
buf ( n206692 , n206647 );
buf ( n206693 , n206688 );
and ( n39417 , n206692 , n206693 );
nor ( n39418 , n39414 , n39417 );
buf ( n206696 , n39418 );
not ( n39420 , n206696 );
not ( n39421 , n39420 );
buf ( n206699 , n206080 );
buf ( n206700 , n185446 );
buf ( n206701 , n206085 );
buf ( n206702 , n38930 );
buf ( n206703 , n206170 );
buf ( n206704 , n206073 );
nand ( n39428 , n206703 , n206704 );
buf ( n206706 , n39428 );
buf ( n206707 , n206706 );
nor ( n39431 , n206702 , n206707 );
buf ( n206709 , n39431 );
buf ( n206710 , n206709 );
nand ( n39434 , n206701 , n206710 );
buf ( n206712 , n39434 );
buf ( n206713 , n206712 );
nor ( n39437 , n206700 , n206713 );
buf ( n206715 , n39437 );
buf ( n206716 , n206715 );
nand ( n39440 , n206699 , n206716 );
buf ( n206718 , n39440 );
buf ( n206719 , n206709 );
not ( n39443 , n206719 );
buf ( n206721 , n206294 );
not ( n39445 , n206721 );
or ( n39446 , n39443 , n39445 );
buf ( n206724 , n206706 );
not ( n39448 , n206724 );
buf ( n206726 , n39448 );
and ( n39450 , n206726 , n38984 );
and ( n39451 , n206276 , n206073 );
nor ( n39452 , n39450 , n39451 , n206067 );
buf ( n206730 , n39452 );
nand ( n39454 , n39446 , n206730 );
buf ( n206732 , n39454 );
buf ( n206733 , n206732 );
not ( n39457 , n206733 );
buf ( n206735 , n39457 );
not ( n39459 , n206712 );
nand ( n39460 , n39459 , n184143 );
nand ( n39461 , n206718 , n206735 , n39460 );
not ( n39462 , n39461 );
or ( n39463 , n39421 , n39462 );
nand ( n39464 , n206718 , n206735 , n39460 , n206696 );
nand ( n39465 , n39463 , n39464 );
buf ( n39466 , n39465 );
or ( n39467 , n39368 , n39466 );
nand ( n39468 , n39288 , n39467 );
nor ( n39469 , n39135 , n39468 );
not ( n39470 , n39469 );
buf ( n206748 , n38169 );
not ( n39472 , n206748 );
buf ( n206750 , n39472 );
buf ( n206751 , n206750 );
buf ( n206752 , n205120 );
buf ( n39476 , n206752 );
buf ( n206754 , n39476 );
buf ( n206755 , n206754 );
not ( n39479 , n206755 );
buf ( n206757 , n39479 );
buf ( n206758 , n206757 );
buf ( n206759 , n205146 );
not ( n39483 , n206759 );
buf ( n206761 , n205156 );
nor ( n39485 , n39483 , n206761 );
buf ( n206763 , n39485 );
buf ( n206764 , n206763 );
nand ( n39488 , n206758 , n206764 );
buf ( n206766 , n39488 );
buf ( n206767 , n206766 );
nor ( n39491 , n206751 , n206767 );
buf ( n206769 , n39491 );
buf ( n206770 , n206769 );
not ( n39494 , n206770 );
buf ( n206772 , n199278 );
not ( n39496 , n206772 );
or ( n39497 , n39494 , n39496 );
buf ( n206775 , n206763 );
not ( n39499 , n206775 );
buf ( n206777 , n205489 );
buf ( n39501 , n206777 );
buf ( n206779 , n39501 );
buf ( n206780 , n206779 );
not ( n39504 , n206780 );
or ( n39505 , n39499 , n39504 );
buf ( n206783 , n205511 );
buf ( n206784 , n205156 );
not ( n39508 , n206784 );
buf ( n206786 , n39508 );
buf ( n206787 , n206786 );
and ( n39511 , n206783 , n206787 );
buf ( n206789 , n205518 );
nor ( n39513 , n39511 , n206789 );
buf ( n206791 , n39513 );
buf ( n206792 , n206791 );
nand ( n39516 , n39505 , n206792 );
buf ( n206794 , n39516 );
buf ( n206795 , n206794 );
not ( n39519 , n206795 );
buf ( n206797 , n39519 );
buf ( n206798 , n206797 );
nand ( n39522 , n39497 , n206798 );
buf ( n206800 , n39522 );
not ( n39524 , n206800 );
buf ( n206802 , n205528 );
not ( n39526 , n206802 );
buf ( n206804 , n205522 );
nand ( n39528 , n39526 , n206804 );
buf ( n206806 , n39528 );
buf ( n39530 , n168462 );
and ( n39531 , n206806 , n39530 );
nor ( n39532 , n205069 , n206766 );
nor ( n39533 , n39531 , n39532 );
nand ( n39534 , n39524 , n39533 );
not ( n39535 , n39534 );
or ( n39536 , n206800 , n39532 );
not ( n39537 , n206806 );
nand ( n39538 , n39537 , n39530 );
nand ( n39539 , n39536 , n39538 );
not ( n39540 , n39539 );
or ( n39541 , n39535 , n39540 );
buf ( n206819 , n185045 );
buf ( n206820 , n185406 );
buf ( n206821 , n185676 );
nand ( n39545 , n206820 , n206821 );
buf ( n206823 , n39545 );
buf ( n206824 , n206823 );
nor ( n39548 , n206819 , n206824 );
buf ( n206826 , n39548 );
buf ( n206827 , n206826 );
not ( n39551 , n206827 );
buf ( n206829 , n185895 );
not ( n39553 , n206829 );
or ( n39554 , n39551 , n39553 );
buf ( n206832 , n177727 );
buf ( n206833 , n185881 );
buf ( n206834 , n206826 );
and ( n39558 , n206833 , n206834 );
buf ( n206836 , n39558 );
buf ( n206837 , n206836 );
and ( n39561 , n206832 , n206837 );
buf ( n206839 , n206823 );
not ( n39563 , n206839 );
buf ( n206841 , n39563 );
buf ( n206842 , n206841 );
not ( n39566 , n206842 );
buf ( n206844 , n185494 );
not ( n39568 , n206844 );
or ( n39569 , n39566 , n39568 );
buf ( n206847 , n185676 );
not ( n39571 , n206847 );
buf ( n206849 , n185519 );
not ( n39573 , n206849 );
or ( n39574 , n39571 , n39573 );
buf ( n206852 , n185680 );
nand ( n39576 , n39574 , n206852 );
buf ( n206854 , n39576 );
buf ( n206855 , n206854 );
not ( n39579 , n206855 );
buf ( n206857 , n39579 );
buf ( n206858 , n206857 );
nand ( n39582 , n39569 , n206858 );
buf ( n206860 , n39582 );
buf ( n206861 , n206860 );
nor ( n39585 , n39561 , n206861 );
buf ( n206863 , n39585 );
buf ( n206864 , n206863 );
nand ( n39588 , n39554 , n206864 );
buf ( n206866 , n39588 );
buf ( n206867 , n205744 );
buf ( n206868 , n205718 );
nor ( n39592 , n206867 , n206868 );
buf ( n206870 , n39592 );
not ( n39594 , n206870 );
nor ( n39595 , n39594 , n39530 );
and ( n39596 , n206866 , n39595 );
not ( n39597 , n206866 );
buf ( n206875 , n206870 );
not ( n39599 , n206875 );
buf ( n206877 , n39599 );
not ( n39601 , n206877 );
nor ( n39602 , n39601 , n39530 );
and ( n39603 , n39597 , n39602 );
nor ( n39604 , n39596 , n39603 );
nand ( n39605 , n39541 , n39604 );
not ( n39606 , n39605 );
buf ( n39607 , n39606 );
buf ( n39608 , n39607 );
buf ( n206886 , n177740 );
buf ( n206887 , n185881 );
buf ( n206888 , n205767 );
not ( n39612 , n38930 );
buf ( n206890 , n39612 );
and ( n39614 , n206888 , n206890 );
buf ( n206892 , n39614 );
buf ( n206893 , n206892 );
and ( n39617 , n206887 , n206893 );
buf ( n206895 , n39617 );
buf ( n206896 , n206895 );
nand ( n39620 , n206886 , n206896 );
buf ( n206898 , n39620 );
and ( n39622 , n39612 , n38477 );
nor ( n39623 , n39622 , n38984 );
buf ( n206901 , n185895 );
buf ( n206902 , n206892 );
nand ( n39626 , n206901 , n206902 );
buf ( n206904 , n39626 );
nand ( n39628 , n206898 , n39623 , n206904 );
buf ( n206906 , n206390 );
buf ( n206907 , n206266 );
nand ( n39631 , n206906 , n206907 );
buf ( n206909 , n39631 );
xnor ( n39633 , n39628 , n206909 );
or ( n39634 , n39608 , n39633 );
buf ( n39635 , n39316 );
buf ( n39636 , n39635 );
not ( n39637 , n168462 );
buf ( n206915 , n205135 );
not ( n39639 , n206915 );
buf ( n206917 , n206779 );
not ( n39641 , n206917 );
or ( n39642 , n39639 , n39641 );
buf ( n206920 , n205501 );
nand ( n39644 , n39642 , n206920 );
buf ( n206922 , n39644 );
not ( n39646 , n206922 );
buf ( n206924 , n205072 );
not ( n39648 , n205135 );
nor ( n39649 , n39648 , n206754 );
buf ( n206927 , n39649 );
nand ( n39651 , n206924 , n206927 );
buf ( n206929 , n39651 );
nand ( n39653 , n199278 , n38169 , n39649 );
nand ( n39654 , n39646 , n206929 , n39653 );
buf ( n206932 , n39654 );
buf ( n206933 , n205143 );
buf ( n206934 , n38231 );
nand ( n39658 , n206933 , n206934 );
buf ( n206936 , n39658 );
buf ( n206937 , n206936 );
not ( n39661 , n206937 );
buf ( n206939 , n39661 );
buf ( n206940 , n206939 );
and ( n39664 , n206932 , n206940 );
not ( n39665 , n206932 );
buf ( n206943 , n206936 );
and ( n39667 , n39665 , n206943 );
nor ( n39668 , n39664 , n39667 );
buf ( n206946 , n39668 );
not ( n39670 , n206946 );
or ( n39671 , n39637 , n39670 );
buf ( n206949 , n185240 );
not ( n39673 , n206949 );
buf ( n206951 , n185494 );
not ( n39675 , n206951 );
or ( n39676 , n39673 , n39675 );
buf ( n206954 , n185506 );
nand ( n39678 , n39676 , n206954 );
buf ( n206956 , n39678 );
not ( n39680 , n206956 );
buf ( n206958 , n185443 );
buf ( n206959 , n185240 );
not ( n39683 , n206959 );
buf ( n206961 , n185045 );
nor ( n39685 , n39683 , n206961 );
buf ( n206963 , n39685 );
buf ( n206964 , n206963 );
and ( n39688 , n206958 , n206964 );
buf ( n206966 , n39688 );
buf ( n206967 , n206966 );
buf ( n206968 , n177727 );
nand ( n39692 , n206967 , n206968 );
buf ( n206970 , n39692 );
buf ( n206971 , n184143 );
buf ( n206972 , n206963 );
nand ( n39696 , n206971 , n206972 );
buf ( n206974 , n39696 );
nand ( n39698 , n39680 , n206970 , n206974 );
buf ( n206976 , n18087 );
buf ( n206977 , n185516 );
nand ( n39701 , n206976 , n206977 );
buf ( n206979 , n39701 );
buf ( n206980 , n206979 );
not ( n39704 , n206980 );
buf ( n206982 , n39704 );
and ( n39706 , n39698 , n206982 );
not ( n39707 , n39698 );
and ( n39708 , n39707 , n206979 );
nor ( n39709 , n39706 , n39708 );
nand ( n39710 , n39709 , n831 );
nand ( n39711 , n39671 , n39710 );
not ( n39712 , n39711 );
not ( n39713 , n39712 );
buf ( n39714 , n39713 );
or ( n39715 , n39636 , n39714 );
and ( n39716 , n831 , n18376 );
not ( n39717 , n831 );
buf ( n206995 , n206786 );
buf ( n206996 , n205518 );
not ( n39720 , n206996 );
and ( n39721 , n206995 , n39720 );
buf ( n206999 , n39721 );
not ( n39723 , n206999 );
not ( n39724 , n39723 );
buf ( n207002 , n206750 );
buf ( n207003 , n205146 );
buf ( n207004 , n206757 );
nand ( n39728 , n207003 , n207004 );
buf ( n207006 , n39728 );
buf ( n207007 , n207006 );
nor ( n39731 , n207002 , n207007 );
buf ( n207009 , n39731 );
nand ( n39733 , n207009 , n199278 );
not ( n39734 , n205069 );
not ( n39735 , n207006 );
nand ( n39736 , n39734 , n39735 );
and ( n39737 , n205146 , n206779 );
nor ( n39738 , n39737 , n205511 );
nand ( n39739 , n39733 , n39736 , n39738 );
not ( n39740 , n39739 );
or ( n39741 , n39724 , n39740 );
nand ( n39742 , n39733 , n39736 , n39738 , n206999 );
nand ( n39743 , n39741 , n39742 );
and ( n39744 , n39717 , n39743 );
nor ( n39745 , n39716 , n39744 );
not ( n39746 , n39745 );
buf ( n39747 , n39746 );
not ( n39748 , n39747 );
not ( n39749 , n39748 );
buf ( n39750 , n39188 );
or ( n39751 , n39749 , n39750 );
not ( n39752 , n831 );
buf ( n207030 , n185494 );
not ( n39754 , n207030 );
buf ( n207032 , n177740 );
buf ( n207033 , n185881 );
buf ( n207034 , n185048 );
and ( n39758 , n207033 , n207034 );
buf ( n207036 , n39758 );
buf ( n207037 , n207036 );
nand ( n39761 , n207032 , n207037 );
buf ( n207039 , n39761 );
buf ( n207040 , n207039 );
buf ( n207041 , n184143 );
buf ( n207042 , n185048 );
nand ( n39766 , n207041 , n207042 );
buf ( n207044 , n39766 );
buf ( n207045 , n207044 );
nand ( n39769 , n39754 , n207040 , n207045 );
buf ( n207047 , n39769 );
buf ( n207048 , n207047 );
buf ( n207049 , n185240 );
buf ( n207050 , n185506 );
nand ( n39774 , n207049 , n207050 );
buf ( n207052 , n39774 );
buf ( n207053 , n207052 );
not ( n39777 , n207053 );
buf ( n207055 , n39777 );
buf ( n207056 , n207055 );
and ( n39780 , n207048 , n207056 );
not ( n39781 , n207048 );
buf ( n207059 , n207052 );
and ( n39783 , n39781 , n207059 );
nor ( n39784 , n39780 , n39783 );
buf ( n207062 , n39784 );
not ( n39786 , n207062 );
or ( n39787 , n39752 , n39786 );
not ( n39788 , n206779 );
buf ( n207066 , n206543 );
buf ( n207067 , n206757 );
nand ( n39791 , n207066 , n207067 );
buf ( n207069 , n39791 );
nand ( n39793 , n199278 , n39275 , n206757 );
nand ( n39794 , n39788 , n207069 , n39793 );
buf ( n207072 , n39794 );
buf ( n207073 , n205135 );
buf ( n207074 , n205501 );
nand ( n39798 , n207073 , n207074 );
buf ( n207076 , n39798 );
buf ( n207077 , n207076 );
not ( n39801 , n207077 );
buf ( n207079 , n39801 );
buf ( n207080 , n207079 );
and ( n39804 , n207072 , n207080 );
not ( n39805 , n207072 );
buf ( n207083 , n207076 );
and ( n39807 , n39805 , n207083 );
nor ( n39808 , n39804 , n39807 );
buf ( n207086 , n39808 );
nand ( n39810 , n207086 , n168462 );
nand ( n39811 , n39787 , n39810 );
buf ( n39812 , n39811 );
buf ( n39813 , n38499 );
and ( n39814 , n39813 , n205803 );
not ( n39815 , n39813 );
and ( n39816 , n39815 , n205798 );
nor ( n39817 , n39814 , n39816 );
or ( n39818 , n39812 , n39817 );
and ( n39819 , n39634 , n39715 , n39751 , n39818 );
not ( n39820 , n39819 );
buf ( n207098 , n206543 );
buf ( n207099 , n205117 );
nand ( n39823 , n207098 , n207099 );
buf ( n207101 , n39823 );
buf ( n207102 , n207101 );
nand ( n39826 , n199278 , n39275 , n205117 );
buf ( n207104 , n39826 );
buf ( n207105 , n38189 );
buf ( n39829 , n207105 );
buf ( n207107 , n39829 );
buf ( n207108 , n207107 );
not ( n39832 , n207108 );
buf ( n207110 , n39832 );
buf ( n207111 , n207110 );
nand ( n39835 , n207102 , n207104 , n207111 );
buf ( n207113 , n39835 );
not ( n39837 , n207113 );
buf ( n207115 , n205477 );
buf ( n207116 , n205092 );
buf ( n39840 , n207116 );
buf ( n207118 , n39840 );
buf ( n207119 , n207118 );
nor ( n39843 , n207115 , n207119 );
buf ( n207121 , n39843 );
nor ( n39845 , n207121 , n831 );
nand ( n39846 , n39837 , n39845 );
not ( n39847 , n18155 );
buf ( n207125 , n177740 );
buf ( n207126 , n185881 );
buf ( n207127 , n185039 );
and ( n39851 , n207126 , n207127 );
buf ( n207129 , n39851 );
buf ( n207130 , n207129 );
nand ( n39854 , n207125 , n207130 );
buf ( n207132 , n39854 );
buf ( n207133 , n184143 );
buf ( n207134 , n185039 );
nand ( n39858 , n207133 , n207134 );
buf ( n207136 , n39858 );
nand ( n39860 , n39847 , n207132 , n207136 );
not ( n39861 , n39860 );
buf ( n207139 , n185868 );
buf ( n207140 , n185476 );
nand ( n39864 , n207139 , n207140 );
buf ( n207142 , n39864 );
and ( n39866 , n207142 , n831 );
nand ( n39867 , n39861 , n39866 );
not ( n39868 , n207121 );
nor ( n39869 , n39868 , n831 );
nand ( n39870 , n207113 , n39869 );
buf ( n207148 , n207142 );
not ( n39872 , n207148 );
buf ( n207150 , n39872 );
and ( n39874 , n207150 , n831 );
nand ( n39875 , n39860 , n39874 );
nand ( n39876 , n39846 , n39867 , n39870 , n39875 );
buf ( n39877 , n39876 );
not ( n39878 , n39877 );
not ( n39879 , n39878 );
not ( n39880 , n39879 );
buf ( n39881 , n206866 );
and ( n39882 , n39881 , n206870 );
not ( n39883 , n39881 );
and ( n39884 , n39883 , n206877 );
nor ( n39885 , n39882 , n39884 );
or ( n39886 , n39880 , n39885 );
buf ( n39887 , n168462 );
buf ( n207165 , n206543 );
not ( n39889 , n205117 );
nor ( n39890 , n39889 , n207118 );
buf ( n207168 , n39890 );
nand ( n39892 , n207165 , n207168 );
buf ( n207170 , n39892 );
buf ( n207171 , n207170 );
buf ( n207172 , n39275 );
buf ( n207173 , n39890 );
and ( n39897 , n207172 , n207173 );
buf ( n207175 , n39897 );
buf ( n207176 , n207175 );
buf ( n207177 , n199278 );
nand ( n39901 , n207176 , n207177 );
buf ( n207179 , n39901 );
buf ( n207180 , n207179 );
buf ( n207181 , n207107 );
buf ( n207182 , n207118 );
not ( n39906 , n207182 );
buf ( n207184 , n39906 );
buf ( n207185 , n207184 );
and ( n39909 , n207181 , n207185 );
buf ( n207187 , n205477 );
nor ( n39911 , n39909 , n207187 );
buf ( n207189 , n39911 );
buf ( n207190 , n207189 );
nand ( n39914 , n207171 , n207180 , n207190 );
buf ( n207192 , n39914 );
buf ( n207193 , n205472 );
not ( n39917 , n207193 );
buf ( n207195 , n205483 );
nor ( n39919 , n39917 , n207195 );
buf ( n207197 , n39919 );
xor ( n39921 , n207192 , n207197 );
and ( n39922 , n39887 , n39921 );
not ( n39923 , n39887 );
and ( n39924 , n39923 , n185916 );
nor ( n39925 , n39922 , n39924 );
buf ( n39926 , n39925 );
buf ( n39927 , n39926 );
buf ( n39928 , n39927 );
not ( n39929 , n39928 );
and ( n39930 , n39028 , n206312 );
not ( n39931 , n39028 );
and ( n39932 , n39931 , n206309 );
nor ( n39933 , n39930 , n39932 );
or ( n39934 , n39929 , n39933 );
nand ( n39935 , n39886 , n39934 );
buf ( n207213 , n37758 );
buf ( n207214 , n205105 );
nor ( n39938 , n207213 , n207214 );
buf ( n207216 , n39938 );
buf ( n207217 , n207216 );
not ( n39941 , n207217 );
buf ( n207219 , n32157 );
not ( n39943 , n207219 );
or ( n39944 , n39941 , n39943 );
buf ( n207222 , n205105 );
not ( n39946 , n207222 );
buf ( n207224 , n39946 );
buf ( n207225 , n207224 );
not ( n39949 , n207225 );
buf ( n207227 , n205003 );
not ( n39951 , n207227 );
buf ( n207229 , n199072 );
not ( n39953 , n207229 );
or ( n39954 , n39951 , n39953 );
buf ( n207232 , n205047 );
nand ( n39956 , n39954 , n207232 );
buf ( n207234 , n39956 );
buf ( n207235 , n207234 );
not ( n39959 , n207235 );
or ( n39960 , n39949 , n39959 );
buf ( n207238 , n37825 );
buf ( n207239 , n205100 );
nand ( n39963 , n207238 , n207239 );
buf ( n207241 , n39963 );
buf ( n207242 , n207241 );
nand ( n39966 , n39960 , n207242 );
buf ( n207244 , n39966 );
buf ( n207245 , n207244 );
not ( n39969 , n207245 );
buf ( n207247 , n39969 );
buf ( n207248 , n207247 );
nand ( n39972 , n39944 , n207248 );
buf ( n207250 , n39972 );
buf ( n207251 , n205114 );
not ( n39975 , n207251 );
buf ( n207253 , n205110 );
buf ( n39977 , n185033 );
buf ( n207255 , n39977 );
nand ( n39979 , n207253 , n207255 );
buf ( n207257 , n39979 );
buf ( n207258 , n207257 );
nand ( n39982 , n39975 , n207258 );
buf ( n207260 , n39982 );
buf ( n207261 , n207260 );
not ( n39985 , n207261 );
buf ( n207263 , n39985 );
and ( n39987 , n207250 , n207263 );
not ( n39988 , n207250 );
and ( n39989 , n39988 , n207260 );
nor ( n39990 , n39987 , n39989 );
not ( n39991 , n39990 );
not ( n39992 , n168462 );
or ( n39993 , n39991 , n39992 );
nand ( n39994 , n39993 , n32069 );
buf ( n39995 , n39994 );
not ( n39996 , n39995 );
not ( n39997 , n39996 );
nor ( n39998 , n39997 , n18377 );
not ( n39999 , n39998 );
buf ( n207277 , n39275 );
not ( n40001 , n207277 );
buf ( n207279 , n31665 );
not ( n40003 , n207279 );
or ( n40004 , n40001 , n40003 );
buf ( n207282 , n205069 );
nand ( n40006 , n40004 , n207282 );
buf ( n207284 , n40006 );
not ( n40008 , n207284 );
buf ( n207286 , n207224 );
buf ( n207287 , n207241 );
nand ( n40011 , n207286 , n207287 );
buf ( n207289 , n40011 );
not ( n40013 , n207289 );
nor ( n40014 , n40013 , n831 );
nand ( n40015 , n40008 , n40014 );
buf ( n207293 , n185443 );
not ( n40017 , n207293 );
buf ( n207295 , n177737 );
not ( n40019 , n207295 );
or ( n40020 , n40017 , n40019 );
buf ( n207298 , n16760 );
not ( n40022 , n207298 );
buf ( n207300 , n16787 );
not ( n40024 , n207300 );
or ( n40025 , n40022 , n40024 );
buf ( n207303 , n16805 );
nand ( n40027 , n40025 , n207303 );
buf ( n207305 , n40027 );
buf ( n207306 , n207305 );
nand ( n40030 , n40020 , n207306 );
buf ( n207308 , n40030 );
not ( n40032 , n207308 );
buf ( n207310 , n186097 );
buf ( n207311 , n185461 );
nand ( n40035 , n207310 , n207311 );
buf ( n207313 , n40035 );
nand ( n40037 , n40032 , n207313 , n831 );
not ( n40038 , n831 );
nor ( n40039 , n207313 , n40038 );
nand ( n40040 , n207308 , n40039 );
not ( n40041 , n207289 );
nand ( n40042 , n40041 , n207284 , n40038 );
nand ( n40043 , n40015 , n40037 , n40040 , n40042 );
not ( n40044 , n40043 );
buf ( n40045 , n40044 );
buf ( n40046 , n39698 );
and ( n40047 , n40046 , n206982 );
not ( n40048 , n40046 );
and ( n40049 , n40048 , n206979 );
nor ( n40050 , n40047 , n40049 );
or ( n40051 , n40045 , n40050 );
nand ( n40052 , n39999 , n40051 );
nor ( n40053 , n39935 , n40052 );
not ( n40054 , n40053 );
buf ( n207332 , n184023 );
buf ( n207333 , n14499 );
buf ( n40057 , n207333 );
buf ( n207335 , n40057 );
buf ( n207336 , n207335 );
buf ( n207337 , n182629 );
not ( n40061 , n207337 );
buf ( n207339 , n40061 );
buf ( n207340 , n207339 );
nand ( n40064 , n207336 , n207340 );
buf ( n207342 , n40064 );
buf ( n207343 , n207342 );
nor ( n40067 , n207332 , n207343 );
buf ( n207345 , n40067 );
buf ( n207346 , n207345 );
not ( n40070 , n207346 );
buf ( n207348 , n177727 );
not ( n40072 , n207348 );
or ( n40073 , n40070 , n40072 );
buf ( n207351 , n207342 );
not ( n40075 , n207351 );
buf ( n207353 , n40075 );
buf ( n207354 , n207353 );
not ( n40078 , n207354 );
buf ( n207356 , n16709 );
not ( n40080 , n207356 );
or ( n40081 , n40078 , n40080 );
buf ( n207359 , n207339 );
not ( n40083 , n207359 );
buf ( n40084 , n16303 );
buf ( n207362 , n40084 );
not ( n40086 , n207362 );
or ( n40087 , n40083 , n40086 );
buf ( n207365 , n183662 );
not ( n40089 , n207365 );
buf ( n207367 , n40089 );
buf ( n207368 , n207367 );
nand ( n40092 , n40087 , n207368 );
buf ( n207370 , n40092 );
buf ( n207371 , n207370 );
not ( n40095 , n207371 );
buf ( n207373 , n40095 );
buf ( n207374 , n207373 );
nand ( n40098 , n40081 , n207374 );
buf ( n207376 , n40098 );
buf ( n207377 , n207376 );
not ( n40101 , n207377 );
buf ( n207379 , n40101 );
buf ( n207380 , n207379 );
nand ( n40104 , n40073 , n207380 );
buf ( n207382 , n40104 );
buf ( n207383 , n182606 );
buf ( n207384 , n16329 );
and ( n40108 , n207383 , n207384 );
buf ( n207386 , n40108 );
and ( n40110 , n207382 , n207386 );
not ( n40111 , n207382 );
buf ( n207389 , n207386 );
not ( n40113 , n207389 );
buf ( n207391 , n40113 );
and ( n40115 , n40111 , n207391 );
nor ( n40116 , n40110 , n40115 );
and ( n40117 , n831 , n40116 );
not ( n40118 , n831 );
buf ( n207396 , n31215 );
not ( n40120 , n207396 );
buf ( n207398 , n40120 );
buf ( n207399 , n207398 );
buf ( n207400 , n31043 );
buf ( n40124 , n207400 );
buf ( n207402 , n40124 );
buf ( n207403 , n207402 );
buf ( n207404 , n198330 );
buf ( n40128 , n207404 );
buf ( n207406 , n40128 );
buf ( n207407 , n207406 );
nand ( n40131 , n207403 , n207407 );
buf ( n207409 , n40131 );
buf ( n207410 , n207409 );
nor ( n40134 , n207399 , n207410 );
buf ( n207412 , n40134 );
not ( n40136 , n207412 );
not ( n40137 , n31665 );
or ( n40138 , n40136 , n40137 );
buf ( n207416 , n207409 );
not ( n40140 , n207416 );
buf ( n207418 , n40140 );
buf ( n207419 , n207418 );
not ( n40143 , n207419 );
buf ( n207421 , n31754 );
not ( n40145 , n207421 );
or ( n40146 , n40143 , n40145 );
buf ( n207424 , n207406 );
not ( n40148 , n207424 );
buf ( n207426 , n199054 );
buf ( n40150 , n207426 );
buf ( n207428 , n40150 );
buf ( n207429 , n207428 );
not ( n40153 , n207429 );
or ( n40154 , n40148 , n40153 );
buf ( n207432 , n199064 );
not ( n40156 , n207432 );
buf ( n207434 , n40156 );
buf ( n207435 , n207434 );
nand ( n40159 , n40154 , n207435 );
buf ( n207437 , n40159 );
buf ( n207438 , n207437 );
not ( n40162 , n207438 );
buf ( n207440 , n40162 );
buf ( n207441 , n207440 );
nand ( n40165 , n40146 , n207441 );
buf ( n207443 , n40165 );
buf ( n207444 , n207443 );
not ( n40168 , n207444 );
buf ( n207446 , n40168 );
nand ( n40170 , n40138 , n207446 );
buf ( n40171 , n31790 );
nand ( n40172 , n40171 , n198339 );
not ( n40173 , n40172 );
and ( n40174 , n40170 , n40173 );
not ( n40175 , n40170 );
and ( n40176 , n40175 , n40172 );
nor ( n40177 , n40174 , n40176 );
and ( n40178 , n40118 , n40177 );
nor ( n40179 , n40117 , n40178 );
not ( n40180 , n40179 );
not ( n40181 , n40180 );
not ( n40182 , n40181 );
xnor ( n40183 , n207308 , n207313 );
or ( n40184 , n40182 , n40183 );
buf ( n207462 , n207398 );
buf ( n207463 , n198319 );
nor ( n40187 , n207462 , n207463 );
buf ( n207465 , n40187 );
buf ( n207466 , n207465 );
not ( n40190 , n207466 );
buf ( n207468 , n199278 );
not ( n40192 , n207468 );
or ( n40193 , n40190 , n40192 );
buf ( n207471 , n199438 );
not ( n40195 , n207471 );
buf ( n207473 , n31754 );
not ( n40197 , n207473 );
or ( n40198 , n40195 , n40197 );
buf ( n207476 , n199442 );
nand ( n40200 , n40198 , n207476 );
buf ( n207478 , n40200 );
buf ( n207479 , n207478 );
not ( n40203 , n207479 );
buf ( n207481 , n40203 );
buf ( n207482 , n207481 );
nand ( n40206 , n40193 , n207482 );
buf ( n207484 , n40206 );
not ( n40208 , n207484 );
buf ( n207486 , n31761 );
buf ( n207487 , n199051 );
and ( n40211 , n207486 , n207487 );
buf ( n207489 , n40211 );
nor ( n40213 , n207489 , n831 );
nand ( n40214 , n40208 , n40213 );
buf ( n207492 , n184023 );
buf ( n40216 , n181859 );
buf ( n207494 , n40216 );
nor ( n40218 , n207492 , n207494 );
buf ( n207496 , n40218 );
buf ( n207497 , n207496 );
not ( n40221 , n207497 );
buf ( n207499 , n177727 );
not ( n40223 , n207499 );
or ( n40224 , n40221 , n40223 );
buf ( n207502 , n40216 );
not ( n40226 , n207502 );
buf ( n207504 , n40226 );
buf ( n207505 , n207504 );
not ( n40229 , n207505 );
buf ( n207507 , n16709 );
not ( n40231 , n207507 );
or ( n40232 , n40229 , n40231 );
buf ( n40233 , n16298 );
buf ( n207511 , n40233 );
nand ( n40235 , n40232 , n207511 );
buf ( n207513 , n40235 );
buf ( n207514 , n207513 );
not ( n40238 , n207514 );
buf ( n207516 , n40238 );
buf ( n207517 , n207516 );
nand ( n40241 , n40224 , n207517 );
buf ( n207519 , n40241 );
not ( n40243 , n207519 );
buf ( n207521 , n183636 );
buf ( n207522 , n16302 );
and ( n40246 , n207521 , n207522 );
buf ( n207524 , n40246 );
buf ( n207525 , n207524 );
not ( n40249 , n207525 );
buf ( n207527 , n40249 );
and ( n40251 , n207527 , n831 );
nand ( n40252 , n40243 , n40251 );
nand ( n40253 , n207519 , n207524 , n831 );
not ( n40254 , n207489 );
nor ( n40255 , n40254 , n831 );
nand ( n40256 , n207484 , n40255 );
nand ( n40257 , n40214 , n40252 , n40253 , n40256 );
buf ( n40258 , n40257 );
not ( n40259 , n40258 );
buf ( n207537 , n177737 );
not ( n40261 , n207537 );
buf ( n207539 , n181081 );
buf ( n207540 , n182635 );
not ( n40264 , n207540 );
buf ( n207542 , n15909 );
nand ( n40266 , n40264 , n207542 );
buf ( n207544 , n40266 );
buf ( n207545 , n207544 );
nor ( n40269 , n207539 , n207545 );
buf ( n207547 , n40269 );
buf ( n207548 , n207547 );
not ( n40272 , n207548 );
or ( n40273 , n40261 , n40272 );
buf ( n207551 , n207544 );
not ( n40275 , n207551 );
buf ( n207553 , n40275 );
buf ( n207554 , n207553 );
not ( n40278 , n207554 );
buf ( n207556 , n16709 );
not ( n40280 , n207556 );
or ( n40281 , n40278 , n40280 );
buf ( n207559 , n15909 );
not ( n40283 , n207559 );
buf ( n207561 , n183678 );
not ( n40285 , n207561 );
or ( n40286 , n40283 , n40285 );
buf ( n207564 , n183704 );
not ( n40288 , n207564 );
buf ( n207566 , n40288 );
buf ( n207567 , n207566 );
nand ( n40291 , n40286 , n207567 );
buf ( n207569 , n40291 );
buf ( n207570 , n207569 );
not ( n40294 , n207570 );
buf ( n207572 , n40294 );
buf ( n207573 , n207572 );
nand ( n40297 , n40281 , n207573 );
buf ( n207575 , n40297 );
buf ( n207576 , n207575 );
not ( n40300 , n207576 );
buf ( n207578 , n40300 );
buf ( n207579 , n207578 );
nand ( n40303 , n40273 , n207579 );
buf ( n207581 , n40303 );
buf ( n207582 , n183533 );
buf ( n207583 , n183711 );
nand ( n40307 , n207582 , n207583 );
buf ( n207585 , n40307 );
buf ( n207586 , n207585 );
not ( n40310 , n207586 );
buf ( n207588 , n40310 );
and ( n40312 , n207581 , n207588 );
not ( n40313 , n207581 );
and ( n40314 , n40313 , n207585 );
nor ( n40315 , n40312 , n40314 );
or ( n40316 , n40259 , n40315 );
not ( n40317 , n831 );
buf ( n207595 , n181081 );
buf ( n207596 , n207335 );
not ( n40320 , n207596 );
buf ( n207598 , n40320 );
buf ( n207599 , n207598 );
nor ( n40323 , n207595 , n207599 );
buf ( n207601 , n40323 );
buf ( n207602 , n207601 );
not ( n40326 , n207602 );
buf ( n207604 , n177727 );
not ( n40328 , n207604 );
or ( n40329 , n40326 , n40328 );
buf ( n207607 , n207335 );
buf ( n207608 , n16283 );
and ( n40332 , n207607 , n207608 );
buf ( n207610 , n40084 );
nor ( n40334 , n40332 , n207610 );
buf ( n207612 , n40334 );
buf ( n207613 , n207612 );
nand ( n40337 , n40329 , n207613 );
buf ( n207615 , n40337 );
buf ( n207616 , n207339 );
buf ( n207617 , n207367 );
nand ( n40341 , n207616 , n207617 );
buf ( n207619 , n40341 );
buf ( n207620 , n207619 );
not ( n40344 , n207620 );
buf ( n207622 , n40344 );
and ( n40346 , n207615 , n207622 );
not ( n40347 , n207615 );
and ( n40348 , n40347 , n207619 );
nor ( n40349 , n40346 , n40348 );
not ( n40350 , n40349 );
or ( n40351 , n40317 , n40350 );
buf ( n207629 , n207402 );
not ( n40353 , n207629 );
buf ( n207631 , n207398 );
nor ( n40355 , n40353 , n207631 );
buf ( n207633 , n40355 );
buf ( n207634 , n207633 );
not ( n40358 , n207634 );
buf ( n207636 , n199278 );
not ( n40360 , n207636 );
or ( n40361 , n40358 , n40360 );
buf ( n207639 , n207402 );
not ( n40363 , n207639 );
buf ( n207641 , n31754 );
not ( n40365 , n207641 );
or ( n40366 , n40363 , n40365 );
buf ( n207644 , n207428 );
not ( n40368 , n207644 );
buf ( n207646 , n40368 );
buf ( n207647 , n207646 );
nand ( n40371 , n40366 , n207647 );
buf ( n207649 , n40371 );
buf ( n207650 , n207649 );
not ( n40374 , n207650 );
buf ( n207652 , n40374 );
buf ( n207653 , n207652 );
nand ( n40377 , n40361 , n207653 );
buf ( n207655 , n40377 );
buf ( n207656 , n207655 );
buf ( n207657 , n207406 );
buf ( n207658 , n207434 );
nand ( n40382 , n207657 , n207658 );
buf ( n207660 , n40382 );
buf ( n207661 , n207660 );
not ( n40385 , n207661 );
buf ( n207663 , n40385 );
buf ( n207664 , n207663 );
and ( n40388 , n207656 , n207664 );
not ( n40389 , n207656 );
buf ( n207667 , n207660 );
and ( n40391 , n40389 , n207667 );
nor ( n40392 , n40388 , n40391 );
buf ( n207670 , n40392 );
nand ( n40394 , n207670 , n168462 );
nand ( n40395 , n40351 , n40394 );
buf ( n40396 , n40395 );
buf ( n40397 , n40396 );
or ( n40398 , n40397 , n16683 );
nand ( n40399 , n207504 , n40233 );
not ( n40400 , n40399 );
and ( n40401 , n18785 , n40400 );
not ( n40402 , n18785 );
and ( n40403 , n40402 , n40399 );
nor ( n40404 , n40401 , n40403 );
not ( n40405 , n40404 );
not ( n40406 , n831 );
or ( n40407 , n40405 , n40406 );
nand ( n40408 , n40407 , n32172 );
buf ( n40409 , n40408 );
buf ( n40410 , n40409 );
or ( n40411 , n16750 , n40410 );
and ( n40412 , n40184 , n40316 , n40398 , n40411 );
not ( n40413 , n31848 );
buf ( n40414 , n40413 );
buf ( n40415 , n40414 );
and ( n40416 , n39860 , n207150 );
not ( n40417 , n39860 );
and ( n40418 , n40417 , n207142 );
nor ( n40419 , n40416 , n40418 );
or ( n40420 , n40415 , n40419 );
buf ( n40421 , n31880 );
buf ( n40422 , n40421 );
or ( n40423 , n40422 , n18814 );
nand ( n40424 , n40420 , n40423 );
and ( n40425 , n207581 , n207588 );
nor ( n40426 , n40425 , n40038 );
not ( n40427 , n40426 );
not ( n40428 , n207581 );
nand ( n40429 , n40428 , n207585 );
not ( n40430 , n40429 );
or ( n40431 , n40427 , n40430 );
buf ( n207709 , n198346 );
buf ( n207710 , n37707 );
not ( n40434 , n207710 );
buf ( n207712 , n40434 );
buf ( n207713 , n207712 );
nor ( n40437 , n207709 , n207713 );
buf ( n207715 , n40437 );
buf ( n207716 , n207715 );
buf ( n207717 , n31215 );
nand ( n40441 , n207716 , n207717 );
buf ( n207719 , n40441 );
buf ( n207720 , n207719 );
not ( n40444 , n207720 );
buf ( n207722 , n31664 );
not ( n40446 , n207722 );
and ( n40447 , n40444 , n40446 );
not ( n40448 , n207715 );
nand ( n40449 , n199030 , n198980 );
not ( n40450 , n40449 );
or ( n40451 , n40448 , n40450 );
buf ( n207729 , n199137 );
not ( n40453 , n207729 );
buf ( n207731 , n207712 );
not ( n40455 , n207731 );
and ( n40456 , n40453 , n40455 );
buf ( n207734 , n37736 );
nor ( n40458 , n40456 , n207734 );
buf ( n207736 , n40458 );
nand ( n40460 , n40451 , n207736 );
buf ( n207738 , n40460 );
nor ( n40462 , n40447 , n207738 );
buf ( n207740 , n40462 );
buf ( n207741 , n207740 );
buf ( n207742 , n204998 );
not ( n40466 , n207742 );
buf ( n207744 , n40466 );
buf ( n207745 , n207744 );
buf ( n207746 , n205020 );
nand ( n40470 , n207745 , n207746 );
buf ( n207748 , n40470 );
buf ( n207749 , n207748 );
and ( n40473 , n207741 , n207749 );
not ( n40474 , n207741 );
buf ( n207752 , n207748 );
not ( n40476 , n207752 );
buf ( n207754 , n40476 );
buf ( n207755 , n207754 );
and ( n40479 , n40474 , n207755 );
nor ( n40480 , n40473 , n40479 );
buf ( n207758 , n40480 );
nand ( n40482 , n207758 , n168462 );
nand ( n40483 , n40431 , n40482 );
buf ( n40484 , n40483 );
buf ( n40485 , n40484 );
or ( n40486 , n40485 , n18613 );
not ( n40487 , n31850 );
buf ( n207765 , n198346 );
buf ( n207766 , n37707 );
buf ( n207767 , n207744 );
nand ( n40491 , n207766 , n207767 );
buf ( n207769 , n40491 );
buf ( n207770 , n207769 );
nor ( n40494 , n207765 , n207770 );
buf ( n207772 , n40494 );
buf ( n207773 , n207772 );
buf ( n207774 , n31215 );
nand ( n40498 , n207773 , n207774 );
buf ( n207776 , n40498 );
nor ( n40500 , n40487 , n207776 );
not ( n40501 , n40500 );
not ( n40502 , n40501 );
buf ( n207780 , n37746 );
not ( n40504 , n207780 );
nor ( n40505 , n204990 , n37708 );
buf ( n207783 , n40505 );
nor ( n40507 , n40504 , n207783 );
buf ( n207785 , n40507 );
not ( n40509 , n207785 );
buf ( n207787 , n207772 );
not ( n40511 , n207787 );
buf ( n207789 , n31754 );
not ( n40513 , n207789 );
or ( n40514 , n40511 , n40513 );
buf ( n207792 , n199137 );
not ( n40516 , n207792 );
buf ( n207794 , n207769 );
not ( n40518 , n207794 );
and ( n40519 , n40516 , n40518 );
buf ( n207797 , n207744 );
not ( n40521 , n207797 );
buf ( n207799 , n37736 );
not ( n40523 , n207799 );
or ( n40524 , n40521 , n40523 );
buf ( n207802 , n205020 );
nand ( n40526 , n40524 , n207802 );
buf ( n207804 , n40526 );
buf ( n207805 , n207804 );
nor ( n40529 , n40519 , n207805 );
buf ( n207807 , n40529 );
buf ( n207808 , n207807 );
nand ( n40532 , n40514 , n207808 );
buf ( n207810 , n40532 );
nor ( n40534 , n40509 , n207810 );
not ( n40535 , n40534 );
or ( n40536 , n40502 , n40535 );
or ( n40537 , n40500 , n207810 );
not ( n40538 , n207785 );
nand ( n40539 , n40537 , n40538 );
nand ( n40540 , n40536 , n40539 );
not ( n40541 , n40540 );
not ( n40542 , n168462 );
or ( n40543 , n40541 , n40542 );
nand ( n40544 , n40543 , n32089 );
buf ( n40545 , n40544 );
not ( n40546 , n40545 );
not ( n40547 , n40546 );
buf ( n40548 , n40547 );
buf ( n40549 , n207062 );
or ( n40550 , n40548 , n40549 );
nand ( n40551 , n40486 , n40550 );
nor ( n40552 , n40424 , n40551 );
and ( n40553 , n40412 , n40552 );
not ( n40554 , n40553 );
not ( n40555 , n185979 );
not ( n40556 , n831 );
or ( n40557 , n40555 , n40556 );
nand ( n40558 , n40557 , n32040 );
buf ( n40559 , n40558 );
not ( n40560 , n40559 );
buf ( n40561 , n40560 );
not ( n40562 , n40561 );
and ( n40563 , n207519 , n207524 );
not ( n40564 , n207519 );
and ( n40565 , n40564 , n207527 );
nor ( n40566 , n40563 , n40565 );
or ( n40567 , n40562 , n40566 );
buf ( n40568 , n168462 );
nor ( n40569 , n31147 , n32023 );
buf ( n207847 , n40569 );
not ( n40571 , n207847 );
buf ( n207849 , n199278 );
not ( n40573 , n207849 );
or ( n40574 , n40571 , n40573 );
not ( n40575 , n32023 );
not ( n40576 , n40575 );
not ( n40577 , n32015 );
or ( n40578 , n40576 , n40577 );
nand ( n40579 , n40578 , n199305 );
buf ( n207857 , n40579 );
not ( n40581 , n207857 );
buf ( n207859 , n40581 );
buf ( n207860 , n207859 );
nand ( n40584 , n40574 , n207860 );
buf ( n207862 , n40584 );
buf ( n207863 , n207862 );
nand ( n40587 , n32173 , n199018 );
buf ( n207865 , n40587 );
not ( n40589 , n207865 );
buf ( n207867 , n40589 );
buf ( n207868 , n207867 );
and ( n40592 , n207863 , n207868 );
not ( n40593 , n207863 );
buf ( n207871 , n40587 );
and ( n40595 , n40593 , n207871 );
nor ( n40596 , n40592 , n40595 );
buf ( n207874 , n40596 );
and ( n40598 , n40568 , n207874 );
not ( n40599 , n40568 );
buf ( n207877 , n185794 );
buf ( n207878 , n12742 );
nor ( n40602 , n207877 , n207878 );
buf ( n207880 , n40602 );
not ( n40604 , n207880 );
not ( n40605 , n177727 );
or ( n40606 , n40604 , n40605 );
not ( n40607 , n18664 );
not ( n40608 , n18507 );
or ( n40609 , n40607 , n40608 );
nand ( n40610 , n40609 , n16225 );
buf ( n207888 , n40610 );
not ( n40612 , n207888 );
buf ( n207890 , n40612 );
nand ( n40614 , n40606 , n207890 );
nand ( n40615 , n185429 , n183588 );
not ( n40616 , n40615 );
and ( n40617 , n40614 , n40616 );
not ( n40618 , n40614 );
and ( n40619 , n40618 , n40615 );
nor ( n40620 , n40617 , n40619 );
and ( n40621 , n40599 , n40620 );
nor ( n40622 , n40598 , n40621 );
not ( n40623 , n40622 );
buf ( n40624 , n40623 );
buf ( n40625 , n40624 );
buf ( n40626 , n40349 );
or ( n40627 , n40625 , n40626 );
nand ( n40628 , n40567 , n40627 );
not ( n40629 , n168462 );
buf ( n207907 , n32175 );
not ( n40631 , n207907 );
buf ( n207909 , n31147 );
nor ( n40633 , n40631 , n207909 );
buf ( n207911 , n40633 );
buf ( n207912 , n207911 );
not ( n40636 , n207912 );
buf ( n207914 , n31850 );
not ( n40638 , n207914 );
or ( n207916 , n40636 , n40638 );
and ( n40640 , n32015 , n32175 );
nor ( n207918 , n40640 , n199479 );
buf ( n207919 , n207918 );
nand ( n207920 , n207916 , n207919 );
buf ( n207921 , n207920 );
buf ( n207922 , n199456 );
buf ( n207923 , n198988 );
nand ( n207924 , n207922 , n207923 );
buf ( n207925 , n207924 );
buf ( n207926 , n207925 );
not ( n40650 , n207926 );
buf ( n207928 , n40650 );
and ( n40652 , n207921 , n207928 );
not ( n207930 , n207921 );
and ( n40654 , n207930 , n207925 );
nor ( n207932 , n40652 , n40654 );
not ( n40656 , n207932 );
or ( n207934 , n40629 , n40656 );
nand ( n40658 , n207934 , n32090 );
buf ( n207936 , n40658 );
not ( n40660 , n207936 );
not ( n207938 , n40660 );
buf ( n40662 , n40116 );
or ( n207940 , n207938 , n40662 );
not ( n40664 , n831 );
not ( n207942 , n18545 );
or ( n40666 , n40664 , n207942 );
nand ( n207944 , n40666 , n32237 );
buf ( n40668 , n207944 );
buf ( n207946 , n40668 );
or ( n40670 , n207946 , n18425 );
nand ( n207948 , n207940 , n40670 );
nor ( n40672 , n40628 , n207948 );
not ( n207950 , n40672 );
not ( n40674 , n168462 );
buf ( n207952 , n198373 );
not ( n40676 , n207952 );
buf ( n207954 , n40676 );
buf ( n207955 , n207954 );
not ( n207956 , n207955 );
buf ( n207957 , n199278 );
not ( n207958 , n207957 );
or ( n40682 , n207956 , n207958 );
nand ( n207960 , n198357 , n198370 );
buf ( n207961 , n207960 );
buf ( n207962 , n207961 );
buf ( n207963 , n207962 );
buf ( n207964 , n207963 );
nand ( n40688 , n40682 , n207964 );
buf ( n207966 , n40688 );
buf ( n207967 , n207966 );
buf ( n207968 , n198389 );
not ( n40692 , n207968 );
buf ( n207970 , n31685 );
nand ( n40694 , n40692 , n207970 );
buf ( n207972 , n40694 );
buf ( n207973 , n207972 );
not ( n207974 , n207973 );
buf ( n207975 , n207974 );
buf ( n207976 , n207975 );
and ( n40700 , n207967 , n207976 );
not ( n207978 , n207967 );
buf ( n207979 , n207972 );
and ( n207980 , n207978 , n207979 );
nor ( n40704 , n40700 , n207980 );
buf ( n207982 , n40704 );
not ( n40706 , n207982 );
or ( n207984 , n40674 , n40706 );
nand ( n40708 , n185787 , n831 );
nand ( n207986 , n207984 , n40708 );
buf ( n40710 , n207986 );
or ( n207988 , n40710 , n18648 );
not ( n40712 , n207988 );
not ( n207990 , n831 );
not ( n40714 , n177745 );
or ( n207992 , n207990 , n40714 );
buf ( n207993 , n207954 );
buf ( n207994 , n207963 );
nand ( n40718 , n207993 , n207994 );
buf ( n207996 , n40718 );
not ( n40720 , n199278 );
xor ( n207998 , n207996 , n40720 );
nand ( n40722 , n207998 , n10010 );
nand ( n208000 , n207992 , n40722 );
buf ( n40724 , n208000 );
buf ( n208002 , n40724 );
buf ( n40726 , n40620 );
and ( n208004 , n208002 , n40726 );
not ( n40728 , n208004 );
or ( n208006 , n40712 , n40728 );
nand ( n40730 , n40710 , n18648 );
nand ( n208008 , n208006 , n40730 );
not ( n40732 , n31113 );
not ( n208010 , n31850 );
or ( n40734 , n40732 , n208010 );
buf ( n208012 , n31687 );
not ( n40736 , n208012 );
buf ( n208014 , n40736 );
nand ( n40738 , n40734 , n208014 );
nand ( n208016 , n198956 , n31688 );
buf ( n208017 , n208016 );
not ( n208018 , n208017 );
buf ( n208019 , n208018 );
and ( n208020 , n40738 , n208019 );
not ( n40744 , n40738 );
and ( n208022 , n40744 , n208016 );
nor ( n40746 , n208020 , n208022 );
not ( n208024 , n40746 );
not ( n40748 , n168462 );
or ( n208026 , n208024 , n40748 );
not ( n40750 , n18692 );
not ( n208028 , n185983 );
nand ( n40752 , n208028 , n177727 );
nand ( n208030 , n40750 , n40752 );
not ( n40754 , n185987 );
nand ( n208032 , n40754 , n185999 );
buf ( n208033 , n208032 );
not ( n208034 , n208033 );
buf ( n208035 , n208034 );
and ( n208036 , n208030 , n208035 );
not ( n40760 , n208030 );
and ( n208038 , n40760 , n208032 );
nor ( n40762 , n208036 , n208038 );
nand ( n208040 , n40762 , n831 );
nand ( n40764 , n208026 , n208040 );
not ( n208042 , n40764 );
buf ( n40766 , n208042 );
not ( n208044 , n40766 );
not ( n40768 , n208044 );
not ( n208046 , n40768 );
or ( n40770 , n208046 , n18546 );
and ( n208048 , n208008 , n40770 );
and ( n40772 , n208046 , n18546 );
nor ( n208050 , n208048 , n40772 );
not ( n40774 , n831 );
not ( n208052 , n18710 );
or ( n40776 , n40774 , n208052 );
and ( n208054 , n31113 , n31688 );
buf ( n208055 , n208054 );
not ( n208056 , n208055 );
buf ( n208057 , n31850 );
not ( n208058 , n208057 );
or ( n40782 , n208056 , n208058 );
and ( n208060 , n31689 , n198956 );
buf ( n208061 , n208060 );
nand ( n208062 , n40782 , n208061 );
buf ( n208063 , n208062 );
buf ( n208064 , n208063 );
or ( n40788 , n198974 , n32013 );
buf ( n208066 , n40788 );
not ( n40790 , n208066 );
buf ( n208068 , n40790 );
buf ( n208069 , n208068 );
and ( n208070 , n208064 , n208069 );
not ( n40794 , n208064 );
buf ( n208072 , n40788 );
and ( n40796 , n40794 , n208072 );
nor ( n208074 , n208070 , n40796 );
buf ( n208075 , n208074 );
nand ( n208076 , n208075 , n168462 );
nand ( n40800 , n40776 , n208076 );
buf ( n208078 , n40800 );
buf ( n40802 , n208078 );
buf ( n208080 , n40404 );
or ( n40804 , n40802 , n208080 );
not ( n208082 , n40804 );
or ( n40806 , n208050 , n208082 );
nand ( n208084 , n40802 , n208080 );
nand ( n40808 , n40806 , n208084 );
not ( n208086 , n40808 );
or ( n40810 , n207950 , n208086 );
not ( n208088 , n831 );
not ( n40812 , n208088 );
buf ( n208090 , n199401 );
not ( n40814 , n208090 );
buf ( n208092 , n40814 );
buf ( n208093 , n198706 );
not ( n208094 , n208093 );
buf ( n208095 , n31581 );
not ( n208096 , n208095 );
or ( n40820 , n208094 , n208096 );
buf ( n208098 , n199419 );
nand ( n40822 , n40820 , n208098 );
buf ( n208100 , n40822 );
buf ( n208101 , n208100 );
buf ( n208102 , n199411 );
nand ( n40826 , n208101 , n208102 );
buf ( n208104 , n40826 );
buf ( n208105 , n199411 );
buf ( n208106 , n198703 );
not ( n40830 , n208106 );
buf ( n208108 , n40830 );
buf ( n208109 , n208108 );
buf ( n208110 , n198592 );
and ( n40834 , n208109 , n208110 );
buf ( n208112 , n40834 );
buf ( n208113 , n208112 );
buf ( n208114 , n198630 );
nand ( n40838 , n208105 , n208113 , n208114 );
buf ( n208116 , n40838 );
nand ( n40840 , n208092 , n208104 , n208116 );
buf ( n208118 , n198888 );
not ( n40842 , n208118 );
buf ( n208120 , n40842 );
buf ( n208121 , n198907 );
buf ( n208122 , n208121 );
buf ( n208123 , n208122 );
nand ( n208124 , n208120 , n208123 );
and ( n40848 , n40840 , n208124 );
not ( n208126 , n40840 );
not ( n40850 , n208124 );
and ( n208128 , n208126 , n40850 );
nor ( n40852 , n40848 , n208128 );
not ( n208130 , n40852 );
or ( n40854 , n40812 , n208130 );
buf ( n208132 , n186063 );
not ( n40856 , n208132 );
buf ( n208134 , n186025 );
buf ( n208135 , n186034 );
nand ( n208136 , n208134 , n208135 );
buf ( n208137 , n208136 );
buf ( n208138 , n208137 );
buf ( n208139 , n186025 );
buf ( n208140 , n18738 );
not ( n40864 , n208140 );
buf ( n208142 , n40864 );
buf ( n208143 , n208142 );
buf ( n208144 , n198261 );
nand ( n40868 , n208139 , n208143 , n208144 );
buf ( n208146 , n40868 );
buf ( n208147 , n208146 );
nand ( n208148 , n40856 , n208138 , n208147 );
buf ( n208149 , n208148 );
not ( n208150 , n208149 );
buf ( n208151 , n5719 );
buf ( n208152 , n177679 );
not ( n40876 , n208152 );
buf ( n208154 , n40876 );
buf ( n208155 , n208154 );
nand ( n208156 , n208151 , n208155 );
buf ( n208157 , n208156 );
not ( n208158 , n208157 );
nand ( n40882 , n208150 , n208158 );
nand ( n208160 , n208149 , n208157 );
nand ( n40884 , n40882 , n208160 , n831 );
nand ( n208162 , n40854 , n40884 );
not ( n40886 , n208162 );
buf ( n208164 , n40886 );
not ( n40888 , n208164 );
not ( n208166 , n40888 );
nor ( n40890 , n18481 , n208166 );
not ( n208168 , n831 );
buf ( n208169 , n186022 );
buf ( n208170 , n5719 );
and ( n208171 , n208169 , n208170 );
buf ( n208172 , n208171 );
buf ( n208173 , n208172 );
buf ( n208174 , n186031 );
buf ( n208175 , n8688 );
nand ( n208176 , n208174 , n208175 );
buf ( n208177 , n208176 );
buf ( n208178 , n208177 );
nand ( n208179 , n208173 , n208178 );
buf ( n208180 , n208179 );
buf ( n208181 , n208180 );
buf ( n208182 , n208172 );
buf ( n208183 , n186042 );
nand ( n208184 , n208182 , n208183 );
buf ( n208185 , n208184 );
buf ( n208186 , n208185 );
buf ( n208187 , n5719 );
not ( n208188 , n208187 );
buf ( n208189 , n18759 );
not ( n208190 , n208189 );
or ( n208191 , n208188 , n208190 );
buf ( n208192 , n208154 );
nand ( n208193 , n208191 , n208192 );
buf ( n208194 , n208193 );
buf ( n208195 , n208194 );
not ( n208196 , n208195 );
buf ( n208197 , n208196 );
buf ( n208198 , n208197 );
nand ( n208199 , n208181 , n208186 , n208198 );
buf ( n208200 , n208199 );
buf ( n208201 , n172813 );
buf ( n208202 , n177688 );
nand ( n208203 , n208201 , n208202 );
buf ( n208204 , n208203 );
and ( n208205 , n208200 , n208204 );
not ( n208206 , n208200 );
not ( n208207 , n208204 );
and ( n208208 , n208206 , n208207 );
nor ( n208209 , n208205 , n208208 );
not ( n208210 , n208209 );
or ( n208211 , n208168 , n208210 );
buf ( n208212 , n199408 );
buf ( n208213 , n208120 );
and ( n208214 , n208212 , n208213 );
buf ( n208215 , n208214 );
buf ( n208216 , n208215 );
buf ( n208217 , n208100 );
nand ( n208218 , n208216 , n208217 );
buf ( n208219 , n208218 );
buf ( n208220 , n208219 );
buf ( n208221 , n208215 );
buf ( n208222 , n198703 );
buf ( n208223 , n198589 );
nor ( n208224 , n208222 , n208223 );
buf ( n208225 , n208224 );
buf ( n208226 , n208225 );
buf ( n208227 , n198146 );
and ( n208228 , n208226 , n208227 );
buf ( n208229 , n208228 );
buf ( n208230 , n208229 );
nand ( n208231 , n208221 , n208230 );
buf ( n208232 , n208231 );
buf ( n208233 , n208232 );
buf ( n208234 , n208120 );
not ( n208235 , n208234 );
buf ( n208236 , n199398 );
not ( n208237 , n208236 );
or ( n208238 , n208235 , n208237 );
buf ( n208239 , n208123 );
nand ( n208240 , n208238 , n208239 );
buf ( n208241 , n208240 );
buf ( n208242 , n208241 );
not ( n208243 , n208242 );
buf ( n208244 , n208243 );
buf ( n208245 , n208244 );
nand ( n208246 , n208220 , n208233 , n208245 );
buf ( n208247 , n208246 );
buf ( n208248 , n198884 );
not ( n208249 , n208248 );
buf ( n208250 , n198920 );
nand ( n208251 , n208249 , n208250 );
buf ( n208252 , n208251 );
nor ( n208253 , n208247 , n208252 );
not ( n208254 , n208253 );
nand ( n208255 , n208247 , n208252 );
not ( n208256 , n831 );
nand ( n208257 , n208254 , n208255 , n208256 );
nand ( n208258 , n208211 , n208257 );
not ( n208259 , n208258 );
buf ( n208260 , n208259 );
buf ( n208261 , n208260 );
buf ( n208262 , n208030 );
and ( n208263 , n208262 , n208035 );
not ( n208264 , n208262 );
and ( n208265 , n208264 , n208032 );
nor ( n208266 , n208263 , n208265 );
nor ( n208267 , n208261 , n208266 );
nor ( n208268 , n40890 , n208267 );
not ( n208269 , n198583 );
not ( n208270 , n199398 );
or ( n208271 , n208269 , n208270 );
buf ( n208272 , n198923 );
not ( n208273 , n208272 );
buf ( n208274 , n208273 );
nand ( n208275 , n208271 , n208274 );
not ( n208276 , n208275 );
buf ( n208277 , n198583 );
buf ( n208278 , n199408 );
and ( n208279 , n208277 , n208278 );
buf ( n208280 , n208279 );
buf ( n208281 , n208280 );
buf ( n208282 , n208229 );
nand ( n208283 , n208281 , n208282 );
buf ( n208284 , n208283 );
buf ( n208285 , n208280 );
buf ( n208286 , n208100 );
nand ( n208287 , n208285 , n208286 );
buf ( n208288 , n208287 );
nand ( n208289 , n208276 , n208284 , n208288 );
not ( n208290 , n208289 );
not ( n208291 , n2047 );
not ( n208292 , n31454 );
and ( n208293 , n208292 , n198929 );
nor ( n41017 , n208291 , n208293 );
nand ( n41018 , n208290 , n41017 );
buf ( n208296 , n173194 );
not ( n41020 , n208296 );
buf ( n208298 , n18759 );
not ( n41022 , n208298 );
or ( n41023 , n41020 , n41022 );
buf ( n208301 , n177691 );
not ( n41025 , n208301 );
buf ( n208303 , n41025 );
buf ( n208304 , n208303 );
nand ( n41028 , n41023 , n208304 );
buf ( n208306 , n41028 );
not ( n41030 , n208306 );
buf ( n208308 , n186022 );
buf ( n208309 , n173194 );
and ( n41033 , n208308 , n208309 );
buf ( n208311 , n41033 );
buf ( n208312 , n208311 );
buf ( n208313 , n186042 );
nand ( n41037 , n208312 , n208313 );
buf ( n208315 , n41037 );
buf ( n208316 , n208311 );
buf ( n208317 , n208177 );
nand ( n41041 , n208316 , n208317 );
buf ( n208319 , n41041 );
nand ( n41043 , n41030 , n208315 , n208319 );
not ( n41044 , n41043 );
buf ( n208322 , n172162 );
buf ( n208323 , n172483 );
nor ( n41047 , n208322 , n208323 );
buf ( n208325 , n41047 );
buf ( n208326 , n208325 );
not ( n41050 , n208326 );
buf ( n208328 , n41050 );
buf ( n208329 , n208328 );
buf ( n208330 , n177703 );
buf ( n41054 , n208330 );
buf ( n208332 , n41054 );
buf ( n208333 , n208332 );
nand ( n41057 , n208329 , n208333 );
buf ( n208335 , n41057 );
and ( n41059 , n208335 , n831 );
nand ( n41060 , n41044 , n41059 );
buf ( n208338 , n208335 );
not ( n41062 , n208338 );
buf ( n208340 , n41062 );
nand ( n41064 , n41043 , n208340 , n831 );
and ( n41065 , n208293 , n2047 );
nand ( n41066 , n208289 , n41065 );
nand ( n41067 , n41018 , n41060 , n41064 , n41066 );
not ( n41068 , n41067 );
buf ( n41069 , n41068 );
not ( n41070 , n41069 );
not ( n41071 , n41070 );
nor ( n41072 , n18711 , n41071 );
nand ( n41073 , n10299 , n177711 );
not ( n41074 , n41073 );
buf ( n208352 , n173191 );
buf ( n208353 , n208325 );
nor ( n41077 , n208352 , n208353 );
buf ( n208355 , n41077 );
buf ( n208356 , n208355 );
not ( n41080 , n208356 );
buf ( n208358 , n186063 );
not ( n41082 , n208358 );
or ( n41083 , n41080 , n41082 );
buf ( n208361 , n208328 );
not ( n41085 , n208361 );
buf ( n208363 , n177691 );
not ( n41087 , n208363 );
or ( n41088 , n41085 , n41087 );
buf ( n208366 , n208332 );
nand ( n41090 , n41088 , n208366 );
buf ( n208368 , n41090 );
buf ( n208369 , n208368 );
not ( n41093 , n208369 );
buf ( n208371 , n41093 );
buf ( n208372 , n208371 );
nand ( n41096 , n41083 , n208372 );
buf ( n208374 , n41096 );
buf ( n208375 , n208374 );
not ( n41099 , n208375 );
buf ( n208377 , n41099 );
buf ( n208378 , n186025 );
buf ( n208379 , n208355 );
and ( n41103 , n208378 , n208379 );
buf ( n208381 , n41103 );
buf ( n208382 , n208381 );
buf ( n41106 , n186042 );
buf ( n208384 , n41106 );
nand ( n41108 , n208382 , n208384 );
buf ( n208386 , n41108 );
buf ( n208387 , n208381 );
not ( n41111 , n186034 );
not ( n41112 , n41111 );
buf ( n208390 , n41112 );
nand ( n41114 , n208387 , n208390 );
buf ( n208392 , n41114 );
nand ( n41116 , n208377 , n208386 , n208392 );
not ( n41117 , n41116 );
or ( n41118 , n41074 , n41117 );
not ( n41119 , n41073 );
nand ( n41120 , n208377 , n208386 , n208392 , n41119 );
nand ( n41121 , n41118 , n41120 );
and ( n41122 , n831 , n41121 );
not ( n41123 , n831 );
buf ( n208401 , n198861 );
buf ( n208402 , n199419 );
nand ( n41126 , n208401 , n208402 );
buf ( n208404 , n41126 );
not ( n41128 , n208404 );
buf ( n208406 , n208229 );
not ( n41130 , n208406 );
buf ( n208408 , n41130 );
nand ( n41132 , n41128 , n208408 );
not ( n41133 , n41132 );
buf ( n208411 , n199411 );
and ( n41135 , n198583 , n208292 );
buf ( n208413 , n41135 );
and ( n41137 , n208411 , n208413 );
buf ( n208415 , n41137 );
not ( n41139 , n208415 );
or ( n41140 , n41133 , n41139 );
and ( n41141 , n41135 , n199401 );
not ( n41142 , n31469 );
not ( n41143 , n198923 );
or ( n41144 , n41142 , n41143 );
nand ( n41145 , n41144 , n198929 );
nor ( n41146 , n41141 , n41145 );
nand ( n41147 , n41140 , n41146 );
buf ( n208425 , n41147 );
not ( n41149 , n198739 );
and ( n41150 , n198935 , n198715 );
nor ( n41151 , n41149 , n41150 );
buf ( n208429 , n41151 );
and ( n41153 , n208425 , n208429 );
not ( n41154 , n208425 );
buf ( n208432 , n41151 );
not ( n41156 , n208432 );
buf ( n208434 , n41156 );
buf ( n208435 , n208434 );
and ( n41159 , n41154 , n208435 );
nor ( n41160 , n41153 , n41159 );
buf ( n208438 , n41160 );
and ( n41162 , n41123 , n208438 );
nor ( n41163 , n41122 , n41162 );
not ( n41164 , n41163 );
buf ( n41165 , n41164 );
nor ( n41166 , n18679 , n41165 );
nor ( n41167 , n41072 , n41166 );
and ( n41168 , n208268 , n41167 );
not ( n41169 , n41168 );
buf ( n208447 , n198621 );
not ( n41171 , n208447 );
buf ( n208449 , n41171 );
buf ( n208450 , n208449 );
not ( n41174 , n208450 );
buf ( n208452 , n198843 );
not ( n41176 , n208452 );
or ( n41177 , n41174 , n41176 );
buf ( n208455 , n198753 );
nand ( n41179 , n41177 , n208455 );
buf ( n208457 , n41179 );
not ( n41181 , n208457 );
buf ( n208459 , n198538 );
buf ( n208460 , n208449 );
and ( n41184 , n208459 , n208460 );
buf ( n208462 , n41184 );
nand ( n41186 , n208404 , n208462 );
buf ( n208464 , n208462 );
buf ( n208465 , n208112 );
buf ( n208466 , n199189 );
nand ( n41190 , n208464 , n208465 , n208466 );
buf ( n208468 , n41190 );
nand ( n41192 , n41181 , n41186 , n208468 );
buf ( n208470 , n41192 );
buf ( n208471 , n198745 );
buf ( n208472 , n198876 );
nand ( n41196 , n208471 , n208472 );
buf ( n208474 , n41196 );
buf ( n208475 , n208474 );
not ( n41199 , n208475 );
buf ( n208477 , n41199 );
buf ( n208478 , n208477 );
and ( n41202 , n208470 , n208478 );
not ( n41203 , n208470 );
buf ( n208481 , n208474 );
and ( n41205 , n41203 , n208481 );
nor ( n41206 , n41202 , n41205 );
buf ( n208484 , n41206 );
and ( n41208 , n168462 , n208484 );
not ( n41209 , n168462 );
buf ( n208487 , n174170 );
buf ( n208488 , n176171 );
not ( n41212 , n208488 );
buf ( n208490 , n41212 );
buf ( n208491 , n208490 );
and ( n41215 , n208487 , n208491 );
buf ( n208493 , n41215 );
not ( n41217 , n208493 );
not ( n41218 , n208142 );
not ( n41219 , n198255 );
or ( n41220 , n41218 , n41219 );
nand ( n41221 , n41220 , n41111 );
not ( n41222 , n41221 );
or ( n41223 , n41217 , n41222 );
and ( n41224 , n6181 , n173662 );
not ( n41225 , n41224 );
not ( n41226 , n208490 );
buf ( n41227 , n6725 );
not ( n41228 , n41227 );
or ( n41229 , n41226 , n41228 );
buf ( n208507 , n173636 );
buf ( n41231 , n208507 );
buf ( n208509 , n41231 );
nand ( n41233 , n41229 , n208509 );
nor ( n41234 , n41225 , n41233 );
nand ( n41235 , n41223 , n41234 );
and ( n41236 , n41227 , n208490 );
not ( n41237 , n208509 );
nor ( n41238 , n41236 , n41237 );
not ( n41239 , n41238 );
not ( n41240 , n41224 );
and ( n41241 , n41239 , n41240 );
not ( n41242 , n208493 );
nor ( n41243 , n41242 , n41224 );
and ( n41244 , n41221 , n41243 );
nor ( n41245 , n41241 , n41244 );
nand ( n41246 , n41235 , n41245 );
and ( n41247 , n41209 , n41246 );
nor ( n41248 , n41208 , n41247 );
buf ( n41249 , n41248 );
not ( n41250 , n41249 );
nor ( n41251 , n10346 , n41250 );
buf ( n208529 , n198538 );
not ( n41253 , n208529 );
buf ( n208531 , n208404 );
not ( n208532 , n208531 );
or ( n41256 , n41253 , n208532 );
not ( n208534 , n198538 );
buf ( n208535 , n198143 );
buf ( n208536 , n198090 );
buf ( n208537 , n197536 );
nand ( n208538 , n208536 , n208537 );
buf ( n208539 , n208538 );
buf ( n208540 , n208539 );
and ( n41264 , n208535 , n208540 );
buf ( n208542 , n41264 );
nor ( n208543 , n208534 , n208542 );
buf ( n208544 , n208543 );
buf ( n208545 , n208112 );
and ( n208546 , n208544 , n208545 );
buf ( n208547 , n198843 );
buf ( n41271 , n208547 );
buf ( n208549 , n41271 );
buf ( n208550 , n208549 );
nor ( n41274 , n208546 , n208550 );
buf ( n208552 , n41274 );
buf ( n208553 , n208552 );
nand ( n41277 , n41256 , n208553 );
buf ( n208555 , n41277 );
not ( n41279 , n208555 );
buf ( n208557 , n198753 );
buf ( n208558 , n208449 );
nand ( n41282 , n208557 , n208558 );
buf ( n208560 , n41282 );
not ( n208561 , n831 );
and ( n41285 , n208560 , n208561 );
nand ( n41286 , n41279 , n41285 );
not ( n208564 , n174170 );
not ( n41288 , n208177 );
or ( n41289 , n208564 , n41288 );
buf ( n208567 , n208142 );
buf ( n208568 , n174173 );
buf ( n208569 , n198252 );
nor ( n208570 , n208568 , n208569 );
buf ( n208571 , n208570 );
buf ( n208572 , n208571 );
and ( n208573 , n208567 , n208572 );
buf ( n208574 , n41227 );
nor ( n41298 , n208573 , n208574 );
buf ( n208576 , n41298 );
nand ( n41300 , n41289 , n208576 );
not ( n41301 , n41300 );
buf ( n208579 , n208490 );
buf ( n208580 , n208509 );
nand ( n41304 , n208579 , n208580 );
buf ( n208582 , n41304 );
and ( n41306 , n208582 , n831 );
nand ( n41307 , n41301 , n41306 );
buf ( n208585 , n208582 );
not ( n41309 , n208585 );
buf ( n208587 , n41309 );
not ( n208588 , n208587 );
nor ( n41312 , n208588 , n208561 );
nand ( n41313 , n41300 , n41312 );
nor ( n208591 , n208560 , n831 );
nand ( n41315 , n208555 , n208591 );
nand ( n41316 , n41286 , n41307 , n41313 , n41315 );
buf ( n208594 , n41316 );
buf ( n41318 , n208594 );
not ( n41319 , n41318 );
not ( n208597 , n41319 );
not ( n41321 , n208597 );
buf ( n41322 , n41121 );
buf ( n208600 , n41322 );
or ( n41324 , n41321 , n208600 );
buf ( n208602 , n208225 );
buf ( n208603 , n198146 );
buf ( n208604 , n198529 );
not ( n41328 , n208604 );
buf ( n208606 , n41328 );
buf ( n208607 , n208606 );
nand ( n41331 , n208602 , n208603 , n208607 );
buf ( n208609 , n41331 );
buf ( n208610 , n208609 );
buf ( n208611 , n198822 );
nand ( n208612 , n208610 , n208611 );
buf ( n208613 , n208612 );
buf ( n208614 , n208613 );
not ( n208615 , n208614 );
buf ( n208616 , n208100 );
buf ( n208617 , n208606 );
nand ( n208618 , n208616 , n208617 );
buf ( n208619 , n208618 );
buf ( n208620 , n208619 );
nand ( n208621 , n208615 , n208620 );
buf ( n208622 , n208621 );
buf ( n208623 , n198840 );
buf ( n208624 , n198830 );
nand ( n41348 , n208623 , n208624 );
buf ( n208626 , n41348 );
buf ( n208627 , n208626 );
not ( n41351 , n208627 );
buf ( n208629 , n41351 );
and ( n208630 , n208622 , n208629 );
not ( n41354 , n208622 );
and ( n41355 , n41354 , n208626 );
nor ( n208633 , n208630 , n41355 );
not ( n41357 , n208633 );
not ( n41358 , n168462 );
or ( n208636 , n41357 , n41358 );
buf ( n208637 , n208177 );
buf ( n208638 , n174164 );
not ( n208639 , n208638 );
buf ( n208640 , n208639 );
buf ( n208641 , n208640 );
nand ( n208642 , n208637 , n208641 );
buf ( n208643 , n208642 );
buf ( n208644 , n208643 );
buf ( n208645 , n208142 );
buf ( n208646 , n198261 );
buf ( n208647 , n208640 );
nand ( n208648 , n208645 , n208646 , n208647 );
buf ( n208649 , n208648 );
buf ( n208650 , n208649 );
buf ( n208651 , n174177 );
nand ( n41375 , n208644 , n208650 , n208651 );
buf ( n208653 , n41375 );
buf ( n208654 , n208653 );
buf ( n41378 , n174184 );
buf ( n208656 , n41378 );
buf ( n208657 , n174193 );
buf ( n208658 , n208657 );
and ( n41382 , n208656 , n208658 );
buf ( n208660 , n41382 );
buf ( n208661 , n208660 );
and ( n41385 , n208654 , n208661 );
not ( n208663 , n208654 );
buf ( n208664 , n208660 );
not ( n41388 , n208664 );
buf ( n208666 , n41388 );
buf ( n208667 , n208666 );
and ( n41391 , n208663 , n208667 );
nor ( n208669 , n41385 , n41391 );
buf ( n208670 , n208669 );
nand ( n41394 , n208670 , n831 );
nand ( n208672 , n208636 , n41394 );
buf ( n41396 , n208672 );
buf ( n41397 , n41396 );
and ( n208675 , n41043 , n208340 );
not ( n41399 , n41043 );
and ( n41400 , n41399 , n208335 );
nor ( n208678 , n208675 , n41400 );
or ( n41402 , n41397 , n208678 );
not ( n41403 , n168462 );
buf ( n208681 , n208404 );
not ( n41405 , n208681 );
buf ( n208683 , n208408 );
nand ( n208684 , n41405 , n208683 );
buf ( n208685 , n208684 );
buf ( n208686 , n208685 );
buf ( n208687 , n208606 );
buf ( n208688 , n198822 );
nand ( n41412 , n208687 , n208688 );
buf ( n208690 , n41412 );
buf ( n208691 , n208690 );
not ( n41415 , n208691 );
buf ( n208693 , n41415 );
buf ( n208694 , n208693 );
and ( n41418 , n208686 , n208694 );
not ( n208696 , n208686 );
buf ( n208697 , n208690 );
and ( n41421 , n208696 , n208697 );
nor ( n208699 , n41418 , n41421 );
buf ( n208700 , n208699 );
not ( n41424 , n208700 );
or ( n208702 , n41403 , n41424 );
not ( n41426 , n186048 );
buf ( n208704 , n208640 );
buf ( n208705 , n174177 );
nand ( n41429 , n208704 , n208705 );
buf ( n208707 , n41429 );
nor ( n208708 , n208707 , n208561 );
and ( n41432 , n41426 , n208708 );
buf ( n208710 , n208707 );
not ( n208711 , n208710 );
buf ( n208712 , n208711 );
nor ( n41436 , n208712 , n208561 );
and ( n208714 , n186048 , n41436 );
nor ( n41438 , n41432 , n208714 );
nand ( n208716 , n208702 , n41438 );
buf ( n208717 , n208716 );
not ( n208718 , n208717 );
buf ( n208719 , n208209 );
nand ( n208720 , n208718 , n208719 );
nand ( n208721 , n41324 , n41402 , n208720 );
nor ( n208722 , n41251 , n208721 );
not ( n208723 , n208722 );
buf ( n208724 , n208670 );
buf ( n208725 , n31944 );
not ( n208726 , n208725 );
not ( n208727 , n208726 );
nor ( n208728 , n208724 , n208727 );
buf ( n208729 , n208542 );
not ( n208730 , n208729 );
buf ( n208731 , n31422 );
buf ( n208732 , n198661 );
buf ( n208733 , n208732 );
buf ( n208734 , n208733 );
buf ( n208735 , n208734 );
nor ( n208736 , n208731 , n208735 );
buf ( n208737 , n208736 );
buf ( n208738 , n208737 );
buf ( n208739 , n198592 );
nand ( n208740 , n208738 , n208739 );
buf ( n208741 , n208740 );
buf ( n208742 , n208741 );
not ( n208743 , n208742 );
and ( n208744 , n208730 , n208743 );
buf ( n208745 , n208737 );
not ( n208746 , n208745 );
buf ( n208747 , n31581 );
not ( n208748 , n208747 );
or ( n208749 , n208746 , n208748 );
buf ( n208750 , n208734 );
not ( n208751 , n208750 );
buf ( n208752 , n208751 );
buf ( n208753 , n208752 );
not ( n208754 , n208753 );
buf ( n208755 , n198791 );
not ( n208756 , n208755 );
or ( n208757 , n208754 , n208756 );
buf ( n208758 , n198802 );
not ( n208759 , n208758 );
buf ( n208760 , n208759 );
buf ( n208761 , n208760 );
nand ( n208762 , n208757 , n208761 );
buf ( n208763 , n208762 );
buf ( n208764 , n208763 );
not ( n208765 , n208764 );
buf ( n208766 , n208765 );
buf ( n208767 , n208766 );
nand ( n208768 , n208749 , n208767 );
buf ( n208769 , n208768 );
buf ( n208770 , n208769 );
nor ( n208771 , n208744 , n208770 );
buf ( n208772 , n208771 );
not ( n208773 , n208772 );
buf ( n208774 , n198797 );
buf ( n208775 , n198808 );
nand ( n208776 , n208774 , n208775 );
buf ( n208777 , n208776 );
nor ( n208778 , n208777 , n831 );
nand ( n208779 , n208773 , n208778 );
buf ( n208780 , n176158 );
not ( n208781 , n208780 );
buf ( n208782 , n176144 );
nand ( n208783 , n208781 , n208782 );
buf ( n208784 , n208783 );
buf ( n208785 , n208784 );
not ( n208786 , n208785 );
buf ( n208787 , n208786 );
nor ( n208788 , n175034 , n18428 );
buf ( n208789 , n176116 );
not ( n208790 , n208789 );
buf ( n208791 , n208790 );
nand ( n208792 , n208788 , n208791 );
buf ( n208793 , n208792 );
buf ( n208794 , n176201 );
nor ( n208795 , n208793 , n208794 );
buf ( n208796 , n208795 );
buf ( n208797 , n208796 );
not ( n208798 , n208797 );
buf ( n208799 , n198255 );
not ( n208800 , n208799 );
or ( n208801 , n208798 , n208800 );
buf ( n208802 , n208792 );
not ( n208803 , n208802 );
buf ( n208804 , n208803 );
buf ( n208805 , n208804 );
buf ( n208806 , n31889 );
and ( n208807 , n208805 , n208806 );
buf ( n208808 , n208791 );
not ( n208809 , n208808 );
buf ( n208810 , n176123 );
not ( n208811 , n208810 );
buf ( n208812 , n8709 );
not ( n208813 , n208812 );
or ( n208814 , n208811 , n208813 );
buf ( n208815 , n8714 );
nand ( n208816 , n208814 , n208815 );
buf ( n208817 , n208816 );
buf ( n208818 , n208817 );
not ( n208819 , n208818 );
or ( n208820 , n208809 , n208819 );
buf ( n208821 , n176152 );
not ( n208822 , n208821 );
buf ( n208823 , n208822 );
buf ( n208824 , n208823 );
nand ( n208825 , n208820 , n208824 );
buf ( n208826 , n208825 );
buf ( n208827 , n208826 );
nor ( n208828 , n208807 , n208827 );
buf ( n208829 , n208828 );
buf ( n208830 , n208829 );
nand ( n208831 , n208801 , n208830 );
buf ( n208832 , n208831 );
nand ( n208833 , n208787 , n208832 , n831 );
not ( n208834 , n208832 );
not ( n208835 , n831 );
nor ( n208836 , n208787 , n208835 );
nand ( n208837 , n208834 , n208836 );
nand ( n208838 , n208772 , n208777 , n208835 );
nand ( n208839 , n208779 , n208833 , n208837 , n208838 );
buf ( n41563 , n208839 );
not ( n41564 , n41563 );
buf ( n41565 , n41564 );
buf ( n41566 , n40882 );
nand ( n41567 , n41566 , n208160 );
nor ( n41568 , n41565 , n41567 );
nor ( n41569 , n208728 , n41568 );
buf ( n208847 , n199202 );
not ( n41571 , n208847 );
buf ( n208849 , n31581 );
not ( n41573 , n208849 );
or ( n41574 , n41571 , n41573 );
buf ( n208852 , n199206 );
nand ( n41576 , n41574 , n208852 );
buf ( n208854 , n41576 );
buf ( n208855 , n208854 );
buf ( n208856 , n198592 );
buf ( n208857 , n199202 );
nand ( n41581 , n208856 , n208857 );
buf ( n208859 , n41581 );
buf ( n208860 , n208859 );
buf ( n208861 , n208542 );
nor ( n41585 , n208860 , n208861 );
buf ( n208863 , n41585 );
buf ( n208864 , n208863 );
nor ( n41588 , n208855 , n208864 );
buf ( n208866 , n41588 );
buf ( n208867 , n208866 );
buf ( n208868 , n31503 );
buf ( n208869 , n198788 );
and ( n41593 , n208868 , n208869 );
buf ( n208871 , n41593 );
buf ( n208872 , n208871 );
not ( n41596 , n208872 );
buf ( n208874 , n41596 );
buf ( n208875 , n208874 );
and ( n41599 , n208867 , n208875 );
not ( n41600 , n208867 );
buf ( n208878 , n208871 );
and ( n41602 , n41600 , n208878 );
nor ( n41603 , n41599 , n41602 );
buf ( n208881 , n41603 );
nand ( n41605 , n208881 , n168462 );
nand ( n41606 , n185766 , n831 );
nand ( n41607 , n41605 , n41606 );
buf ( n41608 , n41607 );
buf ( n41609 , n41608 );
and ( n41610 , n41301 , n208582 );
not ( n41611 , n41301 );
and ( n41612 , n41611 , n208587 );
nor ( n41613 , n41610 , n41612 );
nor ( n41614 , n41609 , n41613 );
buf ( n41615 , n41246 );
not ( n41616 , n831 );
buf ( n208894 , n177669 );
not ( n41618 , n208894 );
not ( n41619 , n208788 );
nor ( n41620 , n41619 , n176201 );
buf ( n208898 , n41620 );
not ( n41622 , n208898 );
or ( n41623 , n41618 , n41622 );
not ( n41624 , n208788 );
not ( n41625 , n8687 );
or ( n41626 , n41624 , n41625 );
buf ( n208904 , n208817 );
not ( n41628 , n208904 );
buf ( n208906 , n41628 );
nand ( n41630 , n41626 , n208906 );
buf ( n208908 , n41630 );
not ( n41632 , n208908 );
buf ( n208910 , n41632 );
buf ( n208911 , n208910 );
nand ( n41635 , n41623 , n208911 );
buf ( n208913 , n41635 );
buf ( n208914 , n208913 );
buf ( n208915 , n208791 );
buf ( n208916 , n208823 );
nand ( n41640 , n208915 , n208916 );
buf ( n208918 , n41640 );
buf ( n208919 , n208918 );
not ( n41643 , n208919 );
buf ( n208921 , n41643 );
buf ( n208922 , n208921 );
and ( n41646 , n208914 , n208922 );
not ( n41647 , n208914 );
buf ( n208925 , n208918 );
and ( n41649 , n41647 , n208925 );
nor ( n41650 , n41646 , n41649 );
buf ( n208928 , n41650 );
not ( n41652 , n208928 );
or ( n41653 , n41616 , n41652 );
buf ( n208931 , n198592 );
buf ( n208932 , n31422 );
not ( n41656 , n208932 );
buf ( n208934 , n41656 );
buf ( n208935 , n208934 );
nand ( n41659 , n208931 , n208935 );
buf ( n208937 , n41659 );
buf ( n208938 , n208937 );
not ( n41662 , n208938 );
buf ( n208940 , n208542 );
not ( n41664 , n208940 );
and ( n41665 , n41662 , n41664 );
buf ( n208943 , n208934 );
not ( n41667 , n208943 );
buf ( n208945 , n31581 );
not ( n41669 , n208945 );
or ( n41670 , n41667 , n41669 );
buf ( n208948 , n198791 );
not ( n41672 , n208948 );
buf ( n208950 , n41672 );
buf ( n208951 , n208950 );
nand ( n41675 , n41670 , n208951 );
buf ( n208953 , n41675 );
buf ( n208954 , n208953 );
nor ( n41678 , n41665 , n208954 );
buf ( n208956 , n41678 );
buf ( n208957 , n208956 );
buf ( n208958 , n208752 );
buf ( n41682 , n208958 );
buf ( n208960 , n41682 );
buf ( n208961 , n208960 );
buf ( n208962 , n208760 );
nand ( n41686 , n208961 , n208962 );
buf ( n208964 , n41686 );
buf ( n208965 , n208964 );
and ( n41689 , n208957 , n208965 );
not ( n41690 , n208957 );
buf ( n208968 , n208964 );
not ( n41692 , n208968 );
buf ( n208970 , n41692 );
buf ( n208971 , n208970 );
and ( n41695 , n41690 , n208971 );
nor ( n41696 , n41689 , n41695 );
buf ( n208974 , n41696 );
nand ( n41698 , n208974 , n168462 );
nand ( n41699 , n41653 , n41698 );
buf ( n41700 , n41699 );
buf ( n41701 , n41700 );
nor ( n41702 , n41615 , n41701 );
nor ( n41703 , n41614 , n41702 );
and ( n41704 , n41569 , n41703 );
not ( n41705 , n41704 );
and ( n41706 , n186048 , n208712 );
not ( n41707 , n186048 );
and ( n41708 , n41707 , n208707 );
nor ( n41709 , n41706 , n41708 );
or ( n41710 , n30962 , n41709 );
not ( n41711 , n41710 );
not ( n41712 , n831 );
not ( n41713 , n186143 );
or ( n41714 , n41712 , n41713 );
nand ( n41715 , n41714 , n32112 );
buf ( n41716 , n41715 );
and ( n41717 , n208832 , n208787 );
not ( n41718 , n208832 );
and ( n41719 , n41718 , n208784 );
nor ( n41720 , n41717 , n41719 );
or ( n41721 , n41716 , n41720 );
not ( n41722 , n41721 );
and ( n41723 , n30997 , n18460 );
not ( n41724 , n41723 );
buf ( n41725 , n31991 );
buf ( n41726 , n208928 );
or ( n41727 , n41725 , n41726 );
not ( n41728 , n41727 );
or ( n41729 , n41724 , n41728 );
nand ( n41730 , n41725 , n41726 );
nand ( n41731 , n41729 , n41730 );
not ( n41732 , n41731 );
or ( n41733 , n41722 , n41732 );
nand ( n41734 , n41716 , n41720 );
nand ( n41735 , n41733 , n41734 );
not ( n41736 , n41735 );
or ( n41737 , n41711 , n41736 );
nand ( n41738 , n30962 , n41709 );
nand ( n41739 , n41737 , n41738 );
not ( n41740 , n41739 );
or ( n41741 , n41705 , n41740 );
buf ( n41742 , n31901 );
buf ( n209020 , n9263 );
buf ( n209021 , n176446 );
not ( n41745 , n209021 );
buf ( n209023 , n41745 );
buf ( n209024 , n209023 );
and ( n41748 , n209020 , n209024 );
buf ( n209026 , n41748 );
buf ( n209027 , n209026 );
buf ( n209028 , n9748 );
buf ( n209029 , n177565 );
nand ( n41753 , n209027 , n209028 , n209029 );
buf ( n209031 , n41753 );
buf ( n209032 , n209031 );
buf ( n209033 , n209026 );
buf ( n209034 , n177613 );
nand ( n41758 , n209033 , n209034 );
buf ( n209036 , n41758 );
buf ( n209037 , n209036 );
buf ( n209038 , n209023 );
not ( n41762 , n209038 );
buf ( n209040 , n177638 );
not ( n41764 , n209040 );
or ( n41765 , n41762 , n41764 );
buf ( n209043 , n177645 );
not ( n41767 , n209043 );
buf ( n209045 , n41767 );
buf ( n209046 , n209045 );
nand ( n41770 , n41765 , n209046 );
buf ( n209048 , n41770 );
buf ( n209049 , n209048 );
not ( n41773 , n209049 );
buf ( n209051 , n41773 );
buf ( n209052 , n209051 );
nand ( n41776 , n209032 , n209037 , n209052 );
buf ( n209054 , n41776 );
buf ( n209055 , n177661 );
not ( n41779 , n209055 );
buf ( n209057 , n177654 );
nand ( n41781 , n41779 , n209057 );
buf ( n209059 , n41781 );
buf ( n209060 , n209059 );
not ( n41784 , n209060 );
buf ( n209062 , n41784 );
and ( n41786 , n209054 , n209062 );
not ( n41787 , n209054 );
and ( n41788 , n41787 , n209059 );
nor ( n41789 , n41786 , n41788 );
and ( n41790 , n831 , n41789 );
not ( n41791 , n831 );
buf ( n209069 , n198109 );
not ( n41793 , n209069 );
buf ( n209071 , n198087 );
not ( n41795 , n209071 );
or ( n41796 , n41793 , n41795 );
buf ( n209074 , n198127 );
not ( n41798 , n209074 );
buf ( n209076 , n41798 );
buf ( n209077 , n209076 );
nand ( n209078 , n41796 , n209077 );
buf ( n209079 , n209078 );
buf ( n209080 , n209079 );
not ( n41804 , n209080 );
buf ( n209082 , n198071 );
buf ( n209083 , n198087 );
and ( n209084 , n209082 , n209083 );
buf ( n209085 , n209084 );
buf ( n209086 , n209085 );
buf ( n209087 , n197481 );
buf ( n209088 , n197411 );
nand ( n209089 , n209086 , n209087 , n209088 );
buf ( n209090 , n209089 );
buf ( n209091 , n209090 );
buf ( n209092 , n209085 );
buf ( n209093 , n197533 );
not ( n41817 , n209093 );
buf ( n209095 , n41817 );
buf ( n209096 , n209095 );
nand ( n41820 , n209092 , n209096 );
buf ( n209098 , n41820 );
buf ( n209099 , n209098 );
nand ( n41823 , n41804 , n209091 , n209099 );
buf ( n209101 , n41823 );
buf ( n209102 , n198134 );
not ( n41826 , n209102 );
buf ( n209104 , n198051 );
nand ( n41828 , n41826 , n209104 );
buf ( n209106 , n41828 );
xnor ( n209107 , n209101 , n209106 );
and ( n41831 , n41791 , n209107 );
nor ( n41832 , n41790 , n41831 );
not ( n209110 , n41832 );
buf ( n41834 , n209110 );
buf ( n41835 , n41834 );
or ( n209113 , n41742 , n41835 );
not ( n41837 , n209113 );
buf ( n41838 , n197979 );
not ( n209116 , n831 );
buf ( n209117 , n177638 );
not ( n41841 , n209117 );
buf ( n209119 , n177613 );
buf ( n209120 , n9263 );
nand ( n41844 , n209119 , n209120 );
buf ( n209122 , n41844 );
buf ( n209123 , n209122 );
buf ( n209124 , n9748 );
buf ( n209125 , n9263 );
buf ( n209126 , n177565 );
nand ( n41850 , n209124 , n209125 , n209126 );
buf ( n209128 , n41850 );
buf ( n209129 , n209128 );
nand ( n41853 , n41841 , n209123 , n209129 );
buf ( n209131 , n41853 );
buf ( n209132 , n209131 );
buf ( n209133 , n209023 );
buf ( n209134 , n209045 );
nand ( n41858 , n209133 , n209134 );
buf ( n209136 , n41858 );
buf ( n209137 , n209136 );
not ( n41861 , n209137 );
buf ( n209139 , n41861 );
buf ( n209140 , n209139 );
and ( n41864 , n209132 , n209140 );
not ( n41865 , n209132 );
buf ( n209143 , n209136 );
and ( n41867 , n41865 , n209143 );
nor ( n41868 , n41864 , n41867 );
buf ( n209146 , n41868 );
not ( n41870 , n209146 );
or ( n41871 , n209116 , n41870 );
buf ( n209149 , n209095 );
buf ( n209150 , n198071 );
buf ( n41874 , n209150 );
buf ( n209152 , n41874 );
buf ( n209153 , n209152 );
nand ( n41877 , n209149 , n209153 );
buf ( n209155 , n41877 );
buf ( n209156 , n197481 );
buf ( n209157 , n209152 );
buf ( n209158 , n197411 );
nand ( n41882 , n209156 , n209157 , n209158 );
buf ( n209160 , n41882 );
not ( n209161 , n198109 );
nand ( n41885 , n209155 , n209160 , n209161 );
nand ( n41886 , n209076 , n198087 );
not ( n209164 , n41886 );
and ( n41888 , n41885 , n209164 );
not ( n41889 , n41885 );
and ( n209167 , n41889 , n41886 );
nor ( n41891 , n41888 , n209167 );
nand ( n41892 , n41891 , n168462 );
nand ( n209170 , n41871 , n41892 );
buf ( n41894 , n209170 );
nor ( n41895 , n41838 , n41894 );
not ( n209173 , n41895 );
not ( n41897 , n209173 );
nand ( n41898 , n199266 , n30292 );
not ( n209176 , n41898 );
not ( n41900 , n209176 );
buf ( n209178 , n177613 );
buf ( n209179 , n185854 );
nand ( n41903 , n209178 , n209179 );
buf ( n209181 , n41903 );
buf ( n209182 , n209181 );
buf ( n209183 , n9748 );
buf ( n209184 , n177565 );
buf ( n209185 , n185854 );
nand ( n41909 , n209183 , n209184 , n209185 );
buf ( n209187 , n41909 );
buf ( n209188 , n209187 );
buf ( n209189 , n177629 );
nand ( n41913 , n209182 , n209188 , n209189 );
buf ( n209191 , n41913 );
buf ( n209192 , n209191 );
buf ( n209193 , n177624 );
not ( n209194 , n209193 );
buf ( n209195 , n177635 );
nand ( n41919 , n209194 , n209195 );
buf ( n209197 , n41919 );
buf ( n209198 , n209197 );
not ( n41922 , n209198 );
buf ( n209200 , n41922 );
buf ( n209201 , n209200 );
and ( n41925 , n209192 , n209201 );
not ( n209203 , n209192 );
buf ( n209204 , n209197 );
and ( n41928 , n209203 , n209204 );
nor ( n209206 , n41925 , n41928 );
buf ( n209207 , n209206 );
and ( n41931 , n831 , n209207 );
not ( n209209 , n831 );
buf ( n209210 , n197533 );
not ( n41934 , n209210 );
buf ( n209212 , n197554 );
nand ( n41936 , n41934 , n209212 );
buf ( n209214 , n41936 );
buf ( n209215 , n209214 );
buf ( n209216 , n197481 );
buf ( n209217 , n197411 );
buf ( n209218 , n197554 );
nand ( n41942 , n209216 , n209217 , n209218 );
buf ( n209220 , n41942 );
buf ( n209221 , n209220 );
buf ( n209222 , n197562 );
nand ( n41946 , n209215 , n209221 , n209222 );
buf ( n209224 , n41946 );
buf ( n209225 , n209224 );
buf ( n209226 , n198099 );
not ( n209227 , n209226 );
buf ( n209228 , n198106 );
nand ( n41952 , n209227 , n209228 );
buf ( n209230 , n41952 );
buf ( n209231 , n209230 );
not ( n41955 , n209231 );
buf ( n209233 , n41955 );
buf ( n209234 , n209233 );
and ( n41958 , n209225 , n209234 );
not ( n209236 , n209225 );
buf ( n209237 , n209230 );
and ( n41961 , n209236 , n209237 );
nor ( n209239 , n41958 , n41961 );
buf ( n209240 , n209239 );
and ( n41964 , n209209 , n209240 );
nor ( n209242 , n41931 , n41964 );
not ( n41966 , n209242 );
nor ( n41967 , n18846 , n41966 );
not ( n209245 , n41967 );
not ( n41969 , n209245 );
or ( n41970 , n41900 , n41969 );
not ( n209248 , n41966 );
not ( n41972 , n209248 );
nand ( n41973 , n18846 , n41972 );
nand ( n209251 , n41970 , n41973 );
not ( n41975 , n209251 );
nor ( n41976 , n198266 , n30384 );
buf ( n209254 , n41789 );
not ( n41978 , n30558 );
buf ( n41979 , n41978 );
or ( n209257 , n209254 , n41979 );
buf ( n41981 , n30610 );
nor ( n41982 , n209146 , n41981 );
not ( n209260 , n41982 );
nand ( n41984 , n209257 , n209260 );
nor ( n209262 , n41976 , n41984 );
not ( n209263 , n209262 );
buf ( n209264 , n30498 );
xor ( n209265 , n209264 , n18560 );
buf ( n209266 , n30055 );
buf ( n209267 , n197381 );
not ( n209268 , n209267 );
buf ( n209269 , n209268 );
buf ( n209270 , n209269 );
nand ( n209271 , n209266 , n209270 );
buf ( n209272 , n209271 );
buf ( n209273 , n209272 );
buf ( n209274 , n197392 );
buf ( n209275 , n197758 );
nand ( n209276 , n209274 , n209275 );
buf ( n209277 , n209276 );
buf ( n209278 , n209277 );
not ( n209279 , n209278 );
buf ( n209280 , n209279 );
buf ( n209281 , n209280 );
and ( n209282 , n209273 , n209281 );
not ( n209283 , n209273 );
buf ( n209284 , n209277 );
and ( n209285 , n209283 , n209284 );
nor ( n209286 , n209282 , n209285 );
buf ( n209287 , n209286 );
and ( n209288 , n168462 , n209287 );
not ( n209289 , n168462 );
buf ( n209290 , n177552 );
not ( n209291 , n209290 );
buf ( n209292 , n209291 );
buf ( n209293 , n209292 );
buf ( n209294 , n177445 );
not ( n209295 , n209294 );
buf ( n209296 , n209295 );
buf ( n209297 , n209296 );
nand ( n209298 , n209293 , n209297 );
buf ( n209299 , n209298 );
buf ( n209300 , n209299 );
buf ( n209301 , n177453 );
buf ( n209302 , n177307 );
nand ( n209303 , n209301 , n209302 );
buf ( n209304 , n209303 );
buf ( n209305 , n209304 );
not ( n209306 , n209305 );
buf ( n209307 , n209306 );
buf ( n209308 , n209307 );
and ( n209309 , n209300 , n209308 );
not ( n209310 , n209300 );
buf ( n209311 , n209304 );
and ( n209312 , n209310 , n209311 );
nor ( n209313 , n209309 , n209312 );
buf ( n209314 , n209313 );
and ( n209315 , n209289 , n209314 );
or ( n209316 , n209288 , n209315 );
buf ( n209317 , n209316 );
or ( n209318 , n197658 , n209317 );
not ( n209319 , n209318 );
not ( n209320 , n168462 );
buf ( n209321 , n199350 );
not ( n209322 , n209321 );
buf ( n209323 , n30054 );
not ( n209324 , n209323 );
or ( n209325 , n209322 , n209324 );
buf ( n209326 , n197372 );
nand ( n209327 , n209325 , n209326 );
buf ( n209328 , n209327 );
buf ( n209329 , n209328 );
buf ( n209330 , n197367 );
not ( n209331 , n209330 );
buf ( n209332 , n197378 );
nand ( n209333 , n209331 , n209332 );
buf ( n209334 , n209333 );
buf ( n209335 , n209334 );
not ( n209336 , n209335 );
buf ( n209337 , n209336 );
buf ( n209338 , n209337 );
and ( n209339 , n209329 , n209338 );
not ( n209340 , n209329 );
buf ( n209341 , n209334 );
and ( n209342 , n209340 , n209341 );
nor ( n209343 , n209339 , n209342 );
buf ( n209344 , n209343 );
not ( n209345 , n209344 );
or ( n209346 , n209320 , n209345 );
nand ( n209347 , n209346 , n32068 );
buf ( n209348 , n209347 );
or ( n209349 , n197833 , n209348 );
not ( n209350 , n209349 );
not ( n209351 , n831 );
buf ( n209352 , n32041 );
buf ( n209353 , n177433 );
nand ( n209354 , n209352 , n209353 );
buf ( n209355 , n209354 );
xor ( n209356 , n197701 , n209355 );
not ( n209357 , n209356 );
or ( n209358 , n209351 , n209357 );
nand ( n209359 , n209358 , n32088 );
buf ( n209360 , n209359 );
or ( n209361 , n197885 , n209360 );
not ( n209362 , n209361 );
or ( n209363 , n197676 , n30643 );
not ( n209364 , n209363 );
not ( n209365 , n197728 );
not ( n209366 , n30666 );
nand ( n209367 , n209365 , n209366 );
not ( n209368 , n209367 );
nor ( n209369 , n209314 , n168523 );
not ( n209370 , n831 );
xor ( n209371 , n168493 , n863 );
not ( n209372 , n209371 );
or ( n209373 , n209370 , n209372 );
nand ( n209374 , n895 , n168462 );
nand ( n209375 , n209373 , n209374 );
nand ( n209376 , n199344 , n209375 );
or ( n209377 , n209369 , n209376 );
nand ( n209378 , n209314 , n168523 );
nand ( n209379 , n209377 , n209378 );
not ( n209380 , n209379 );
or ( n209381 , n209368 , n209380 );
nand ( n209382 , n30666 , n197728 );
nand ( n209383 , n209381 , n209382 );
not ( n209384 , n209383 );
or ( n209385 , n209364 , n209384 );
nand ( n209386 , n197676 , n30643 );
nand ( n209387 , n209385 , n209386 );
not ( n209388 , n209387 );
or ( n209389 , n209362 , n209388 );
nand ( n209390 , n197885 , n209360 );
nand ( n209391 , n209389 , n209390 );
not ( n209392 , n209391 );
or ( n209393 , n209350 , n209392 );
nand ( n209394 , n197833 , n209348 );
nand ( n209395 , n209393 , n209394 );
not ( n209396 , n209395 );
or ( n209397 , n209319 , n209396 );
nand ( n209398 , n197658 , n209317 );
nand ( n209399 , n209397 , n209398 );
and ( n209400 , n209265 , n209399 );
and ( n209401 , n209264 , n18560 );
or ( n209402 , n209400 , n209401 );
or ( n209403 , n209207 , n30412 );
and ( n209404 , n209402 , n209403 );
not ( n209405 , n209404 );
or ( n209406 , n209263 , n209405 );
not ( n209407 , n41976 );
nand ( n209408 , n209207 , n30412 );
or ( n209409 , n41982 , n209408 );
nand ( n209410 , n209146 , n41981 );
nand ( n209411 , n209409 , n209410 );
not ( n209412 , n209411 );
not ( n209413 , n209257 );
or ( n209414 , n209412 , n209413 );
nand ( n209415 , n209254 , n41979 );
nand ( n209416 , n209414 , n209415 );
and ( n209417 , n209407 , n209416 );
and ( n209418 , n198266 , n30384 );
nor ( n209419 , n209417 , n209418 );
nand ( n209420 , n209406 , n209419 );
nor ( n209421 , n199266 , n30292 );
nor ( n209422 , n41967 , n209421 );
nand ( n209423 , n209420 , n209422 );
nand ( n209424 , n41975 , n209423 );
not ( n209425 , n209424 );
or ( n209426 , n41897 , n209425 );
nand ( n209427 , n41838 , n41894 );
nand ( n209428 , n209426 , n209427 );
not ( n209429 , n209428 );
or ( n209430 , n41837 , n209429 );
nand ( n209431 , n41742 , n41835 );
nand ( n209432 , n209430 , n209431 );
or ( n209433 , n30997 , n18460 );
and ( n209434 , n41710 , n41721 , n41727 , n209433 );
and ( n209435 , n209432 , n209434 );
and ( n209436 , n209435 , n41704 );
not ( n209437 , n208726 );
nand ( n209438 , n208724 , n209437 );
or ( n209439 , n41614 , n209438 );
nand ( n209440 , n41609 , n41613 );
nand ( n209441 , n209439 , n209440 );
not ( n209442 , n41702 );
and ( n209443 , n209441 , n209442 );
nand ( n209444 , n41615 , n41701 );
not ( n209445 , n209444 );
nor ( n209446 , n209443 , n209445 );
or ( n209447 , n209446 , n41568 );
nand ( n209448 , n41567 , n41565 );
nand ( n209449 , n209447 , n209448 );
nor ( n209450 , n209436 , n209449 );
nand ( n209451 , n41741 , n209450 );
not ( n209452 , n209451 );
or ( n209453 , n208723 , n209452 );
not ( n209454 , n41324 );
not ( n209455 , n208717 );
nor ( n209456 , n209455 , n208719 );
not ( n209457 , n209456 );
not ( n209458 , n41402 );
or ( n209459 , n209457 , n209458 );
buf ( n209460 , n41397 );
nand ( n209461 , n209460 , n208678 );
nand ( n209462 , n209459 , n209461 );
not ( n209463 , n209462 );
or ( n209464 , n209454 , n209463 );
nand ( n209465 , n41321 , n208600 );
nand ( n209466 , n209464 , n209465 );
not ( n209467 , n41251 );
and ( n209468 , n209466 , n209467 );
and ( n209469 , n10346 , n41250 );
nor ( n209470 , n209468 , n209469 );
nand ( n209471 , n209453 , n209470 );
not ( n209472 , n209471 );
or ( n209473 , n41169 , n209472 );
nand ( n209474 , n18481 , n208166 );
or ( n209475 , n209474 , n208267 );
nand ( n209476 , n208261 , n208266 );
nand ( n209477 , n209475 , n209476 );
not ( n209478 , n209477 );
not ( n209479 , n41072 );
not ( n209480 , n209479 );
or ( n209481 , n209478 , n209480 );
nand ( n209482 , n18711 , n41071 );
nand ( n209483 , n209481 , n209482 );
not ( n209484 , n41166 );
and ( n209485 , n209483 , n209484 );
and ( n209486 , n18679 , n41165 );
nor ( n209487 , n209485 , n209486 );
nand ( n209488 , n209473 , n209487 );
or ( n209489 , n208002 , n40726 );
and ( n209490 , n40804 , n207988 , n40770 , n209489 );
and ( n209491 , n209488 , n209490 , n40672 );
not ( n209492 , n207940 );
and ( n209493 , n40562 , n40566 );
not ( n209494 , n209493 );
not ( n209495 , n40627 );
or ( n209496 , n209494 , n209495 );
nand ( n209497 , n40625 , n40626 );
nand ( n209498 , n209496 , n209497 );
not ( n209499 , n209498 );
or ( n209500 , n209492 , n209499 );
nand ( n209501 , n207938 , n40662 );
nand ( n209502 , n209500 , n209501 );
and ( n209503 , n209502 , n40670 );
and ( n209504 , n207946 , n18425 );
nor ( n209505 , n209503 , n209504 );
not ( n209506 , n209505 );
nor ( n209507 , n209491 , n209506 );
nand ( n209508 , n40810 , n209507 );
not ( n209509 , n209508 );
or ( n209510 , n40554 , n209509 );
not ( n209511 , n40184 );
not ( n209512 , n40398 );
nand ( n209513 , n16750 , n40410 );
not ( n209514 , n209513 );
not ( n209515 , n209514 );
not ( n209516 , n40316 );
or ( n209517 , n209515 , n209516 );
nand ( n209518 , n40259 , n40315 );
nand ( n209519 , n209517 , n209518 );
not ( n209520 , n209519 );
or ( n209521 , n209512 , n209520 );
nand ( n209522 , n40397 , n16683 );
nand ( n209523 , n209521 , n209522 );
not ( n209524 , n209523 );
or ( n209525 , n209511 , n209524 );
nand ( n209526 , n40182 , n40183 );
nand ( n209527 , n209525 , n209526 );
and ( n209528 , n209527 , n40552 );
not ( n209529 , n40420 );
and ( n209530 , n40422 , n18814 );
not ( n209531 , n209530 );
or ( n209532 , n209529 , n209531 );
nand ( n209533 , n40415 , n40419 );
nand ( n209534 , n209532 , n209533 );
and ( n209535 , n209534 , n40486 );
and ( n209536 , n40485 , n18613 );
nor ( n209537 , n209535 , n209536 );
not ( n209538 , n40550 );
or ( n209539 , n209537 , n209538 );
nand ( n209540 , n40548 , n40549 );
nand ( n209541 , n209539 , n209540 );
nor ( n209542 , n209528 , n209541 );
nand ( n209543 , n209510 , n209542 );
not ( n209544 , n209543 );
or ( n209545 , n40054 , n209544 );
not ( n209546 , n39886 );
nand ( n209547 , n40045 , n40050 );
or ( n209548 , n209547 , n39998 );
nand ( n209549 , n39997 , n18377 );
nand ( n209550 , n209548 , n209549 );
not ( n209551 , n209550 );
or ( n209552 , n209546 , n209551 );
nand ( n209553 , n39880 , n39885 );
nand ( n209554 , n209552 , n209553 );
and ( n209555 , n209554 , n39934 );
and ( n209556 , n39929 , n39933 );
nor ( n209557 , n209555 , n209556 );
nand ( n209558 , n209545 , n209557 );
not ( n209559 , n209558 );
or ( n209560 , n39820 , n209559 );
not ( n209561 , n39751 );
not ( n209562 , n39715 );
nand ( n209563 , n39817 , n39812 );
not ( n209564 , n209563 );
not ( n209565 , n209564 );
or ( n209566 , n209562 , n209565 );
nand ( n209567 , n39714 , n39636 );
nand ( n209568 , n209566 , n209567 );
not ( n209569 , n209568 );
or ( n209570 , n209561 , n209569 );
nand ( n209571 , n39749 , n39750 );
nand ( n209572 , n209570 , n209571 );
and ( n209573 , n209572 , n39634 );
and ( n209574 , n39608 , n39633 );
nor ( n209575 , n209573 , n209574 );
nand ( n209576 , n209560 , n209575 );
not ( n209577 , n209576 );
or ( n209578 , n39470 , n209577 );
not ( n209579 , n39287 );
nand ( n209580 , n39368 , n39466 );
not ( n209581 , n209580 );
and ( n209582 , n209579 , n209581 );
not ( n209583 , n39014 );
nand ( n209584 , n39089 , n39132 );
not ( n209585 , n209584 );
and ( n209586 , n209583 , n209585 );
and ( n209587 , n38533 , n39013 );
nor ( n209588 , n209586 , n209587 );
nor ( n209589 , n209588 , n39468 );
nor ( n209590 , n209582 , n209589 );
nand ( n209591 , n209578 , n209590 );
not ( n209592 , n168462 );
not ( n209593 , n199278 );
buf ( n209594 , n39275 );
not ( n209595 , n209594 );
buf ( n209596 , n209595 );
buf ( n209597 , n209596 );
buf ( n209598 , n206325 );
buf ( n209599 , n206495 );
buf ( n209600 , n206507 );
buf ( n209601 , n206479 );
nor ( n209602 , n209600 , n209601 );
buf ( n209603 , n209602 );
buf ( n209604 , n209603 );
and ( n209605 , n209599 , n209604 );
buf ( n209606 , n209605 );
buf ( n209607 , n209606 );
not ( n209608 , n209607 );
buf ( n209609 , n209608 );
buf ( n209610 , n209609 );
and ( n209611 , n206473 , n206474 );
buf ( n209612 , n209611 );
buf ( n209613 , n209612 );
buf ( n209614 , n206146 );
buf ( n209615 , n206152 );
xor ( n209616 , n209614 , n209615 );
buf ( n209617 , n209616 );
buf ( n209618 , n209617 );
nor ( n209619 , n209613 , n209618 );
buf ( n209620 , n209619 );
buf ( n209621 , n209620 );
nor ( n209622 , n209610 , n209621 );
buf ( n209623 , n209622 );
buf ( n209624 , n209623 );
nand ( n209625 , n209598 , n209624 );
buf ( n209626 , n209625 );
buf ( n209627 , n209626 );
nor ( n209628 , n209597 , n209627 );
buf ( n209629 , n209628 );
not ( n209630 , n209629 );
or ( n209631 , n209593 , n209630 );
buf ( n209632 , n209623 );
buf ( n209633 , n205540 );
and ( n209634 , n209632 , n209633 );
buf ( n209635 , n209620 );
not ( n209636 , n209635 );
buf ( n209637 , n209636 );
buf ( n209638 , n209637 );
not ( n209639 , n209638 );
buf ( n209640 , n209603 );
not ( n209641 , n209640 );
buf ( n209642 , n206523 );
not ( n209643 , n209642 );
or ( n209644 , n209641 , n209643 );
buf ( n209645 , n206533 );
buf ( n209646 , n206482 );
and ( n209647 , n209645 , n209646 );
buf ( n209648 , n206487 );
not ( n209649 , n209648 );
buf ( n209650 , n209649 );
buf ( n209651 , n209650 );
nor ( n209652 , n209647 , n209651 );
buf ( n209653 , n209652 );
buf ( n209654 , n209653 );
nand ( n209655 , n209644 , n209654 );
buf ( n209656 , n209655 );
buf ( n209657 , n209656 );
not ( n209658 , n209657 );
or ( n209659 , n209639 , n209658 );
buf ( n209660 , n209612 );
buf ( n209661 , n209617 );
nand ( n209662 , n209660 , n209661 );
buf ( n209663 , n209662 );
buf ( n209664 , n209663 );
nand ( n209665 , n209659 , n209664 );
buf ( n209666 , n209665 );
buf ( n209667 , n209666 );
nor ( n209668 , n209634 , n209667 );
buf ( n209669 , n209668 );
nand ( n209670 , n209631 , n209669 );
and ( n209671 , n209614 , n209615 );
buf ( n209672 , n209671 );
buf ( n209673 , n209672 );
buf ( n209674 , n205911 );
buf ( n209675 , n206028 );
xor ( n209676 , n209674 , n209675 );
buf ( n209677 , n209676 );
buf ( n209678 , n209677 );
nor ( n209679 , n209673 , n209678 );
buf ( n209680 , n209679 );
buf ( n209681 , n209680 );
not ( n209682 , n209681 );
buf ( n209683 , n209672 );
buf ( n209684 , n209677 );
nand ( n209685 , n209683 , n209684 );
buf ( n209686 , n209685 );
buf ( n209687 , n209686 );
nand ( n209688 , n209682 , n209687 );
buf ( n209689 , n209688 );
nor ( n209690 , n209670 , n209689 );
not ( n209691 , n209690 );
buf ( n209692 , n206321 );
not ( n209693 , n209692 );
buf ( n209694 , n209693 );
nor ( n209695 , n209626 , n209694 );
not ( n209696 , n209695 );
not ( n209697 , n209696 );
or ( n209698 , n209691 , n209697 );
or ( n209699 , n209695 , n209670 );
nand ( n209700 , n209699 , n209689 );
nand ( n209701 , n209698 , n209700 );
not ( n209702 , n209701 );
or ( n209703 , n209592 , n209702 );
nand ( n209704 , n39102 , n206384 , n206401 , n39127 );
nand ( n209705 , n39125 , n39128 );
nand ( n209706 , n209704 , n209705 , n831 );
nand ( n209707 , n209703 , n209706 );
not ( n209708 , n209707 );
buf ( n209709 , n209708 );
not ( n209710 , n209709 );
buf ( n209711 , n209710 );
not ( n209712 , n209711 );
buf ( n209713 , n209637 );
buf ( n209714 , n209663 );
nand ( n209715 , n209713 , n209714 );
buf ( n209716 , n209715 );
and ( n209717 , n168462 , n209716 );
not ( n209718 , n209717 );
not ( n209719 , n209718 );
buf ( n209720 , n205072 );
buf ( n209721 , n205305 );
buf ( n209722 , n206495 );
buf ( n209723 , n209603 );
and ( n209724 , n209722 , n209723 );
buf ( n209725 , n209724 );
buf ( n209726 , n209725 );
and ( n209727 , n209721 , n209726 );
buf ( n209728 , n209727 );
buf ( n209729 , n209728 );
nand ( n209730 , n209720 , n209729 );
buf ( n209731 , n209730 );
buf ( n209732 , n209725 );
not ( n209733 , n209732 );
buf ( n209734 , n205540 );
not ( n209735 , n209734 );
or ( n209736 , n209733 , n209735 );
buf ( n209737 , n209656 );
not ( n209738 , n209737 );
buf ( n209739 , n209738 );
buf ( n209740 , n209739 );
nand ( n209741 , n209736 , n209740 );
buf ( n209742 , n209741 );
buf ( n209743 , n209742 );
not ( n209744 , n209743 );
buf ( n209745 , n209744 );
buf ( n209746 , n38169 );
buf ( n209747 , n209728 );
and ( n209748 , n209746 , n209747 );
buf ( n209749 , n209748 );
buf ( n209750 , n209749 );
buf ( n209751 , n199278 );
nand ( n209752 , n209750 , n209751 );
buf ( n209753 , n209752 );
nand ( n209754 , n209731 , n209745 , n209753 );
not ( n209755 , n209754 );
or ( n209756 , n209719 , n209755 );
not ( n209757 , n168462 );
nor ( n209758 , n209757 , n209716 );
not ( n209759 , n209758 );
nand ( n209760 , n209759 , n209731 , n209745 , n209753 );
nand ( n209761 , n209756 , n209760 );
or ( n209762 , n39623 , n206909 );
nand ( n209763 , n209762 , n831 );
not ( n209764 , n209763 );
nand ( n209765 , n39623 , n206898 , n206904 , n206909 );
or ( n209766 , n206898 , n206909 );
or ( n209767 , n206904 , n206909 );
nand ( n209768 , n209764 , n209765 , n209766 , n209767 );
nand ( n209769 , n209761 , n209768 );
buf ( n209770 , n209769 );
not ( n209771 , n209770 );
nor ( n209772 , n209712 , n209771 );
nand ( n209773 , n209591 , n209772 );
and ( n209774 , n831 , n39013 );
not ( n209775 , n831 );
buf ( n209776 , n209694 );
not ( n209777 , n209776 );
buf ( n209778 , n206325 );
buf ( n209779 , n209620 );
buf ( n209780 , n209680 );
nor ( n209781 , n209779 , n209780 );
buf ( n209782 , n209781 );
buf ( n209783 , n209782 );
not ( n209784 , n209783 );
buf ( n209785 , n209609 );
nor ( n209786 , n209784 , n209785 );
buf ( n209787 , n209786 );
buf ( n209788 , n209787 );
nand ( n209789 , n209778 , n209788 );
buf ( n209790 , n209789 );
buf ( n209791 , n209790 );
not ( n209792 , n209791 );
and ( n209793 , n209777 , n209792 );
buf ( n209794 , n209596 );
buf ( n209795 , n209790 );
nor ( n209796 , n209794 , n209795 );
buf ( n209797 , n209796 );
buf ( n209798 , n209797 );
not ( n209799 , n209798 );
buf ( n209800 , n199278 );
not ( n209801 , n209800 );
or ( n209802 , n209799 , n209801 );
buf ( n209803 , n209787 );
buf ( n209804 , n206352 );
and ( n209805 , n209803 , n209804 );
buf ( n209806 , n209782 );
not ( n209807 , n209806 );
buf ( n209808 , n209656 );
not ( n209809 , n209808 );
or ( n209810 , n209807 , n209809 );
buf ( n209811 , n209663 );
buf ( n209812 , n209680 );
or ( n209813 , n209811 , n209812 );
buf ( n209814 , n209686 );
nand ( n209815 , n209813 , n209814 );
buf ( n209816 , n209815 );
buf ( n209817 , n209816 );
not ( n209818 , n209817 );
buf ( n209819 , n209818 );
buf ( n209820 , n209819 );
nand ( n209821 , n209810 , n209820 );
buf ( n209822 , n209821 );
buf ( n209823 , n209822 );
nor ( n209824 , n209805 , n209823 );
buf ( n209825 , n209824 );
buf ( n209826 , n209825 );
nand ( n209827 , n209802 , n209826 );
buf ( n209828 , n209827 );
buf ( n209829 , n209828 );
nor ( n209830 , n209793 , n209829 );
buf ( n209831 , n209830 );
buf ( n209832 , n209831 );
and ( n209833 , n209674 , n209675 );
buf ( n209834 , n209833 );
buf ( n209835 , n209834 );
buf ( n209836 , n206055 );
buf ( n209837 , n206061 );
xor ( n209838 , n209836 , n209837 );
buf ( n209839 , n209838 );
buf ( n209840 , n209839 );
and ( n209841 , n209835 , n209840 );
buf ( n209842 , n209841 );
buf ( n209843 , n209842 );
not ( n209844 , n209843 );
buf ( n209845 , n209834 );
buf ( n209846 , n209839 );
or ( n209847 , n209845 , n209846 );
buf ( n209848 , n209847 );
buf ( n209849 , n209848 );
nand ( n209850 , n209844 , n209849 );
buf ( n209851 , n209850 );
buf ( n209852 , n209851 );
and ( n209853 , n209832 , n209852 );
not ( n209854 , n209832 );
buf ( n209855 , n209851 );
not ( n209856 , n209855 );
buf ( n209857 , n209856 );
buf ( n209858 , n209857 );
and ( n209859 , n209854 , n209858 );
nor ( n209860 , n209853 , n209859 );
buf ( n209861 , n209860 );
and ( n209862 , n209775 , n209861 );
nor ( n209863 , n209774 , n209862 );
not ( n209864 , n209863 );
buf ( n209865 , n209864 );
buf ( n209866 , n209865 );
buf ( n209867 , n209866 );
not ( n209868 , n209867 );
nor ( n209869 , n209773 , n209868 );
not ( n209870 , n831 );
not ( n209871 , n39465 );
or ( n209872 , n209870 , n209871 );
not ( n209873 , n831 );
buf ( n209874 , n209694 );
not ( n209875 , n209874 );
buf ( n209876 , n206325 );
buf ( n209877 , n209609 );
buf ( n209878 , n209782 );
buf ( n209879 , n209848 );
nand ( n209880 , n209878 , n209879 );
buf ( n209881 , n209880 );
buf ( n209882 , n209881 );
nor ( n209883 , n209877 , n209882 );
buf ( n209884 , n209883 );
buf ( n209885 , n209884 );
nand ( n209886 , n209876 , n209885 );
buf ( n209887 , n209886 );
buf ( n209888 , n209887 );
not ( n209889 , n209888 );
and ( n209890 , n209875 , n209889 );
buf ( n209891 , n209596 );
buf ( n209892 , n209887 );
nor ( n209893 , n209891 , n209892 );
buf ( n209894 , n209893 );
buf ( n209895 , n209894 );
not ( n209896 , n209895 );
buf ( n209897 , n199278 );
not ( n209898 , n209897 );
or ( n209899 , n209896 , n209898 );
buf ( n209900 , n209884 );
not ( n209901 , n209900 );
buf ( n209902 , n206352 );
not ( n209903 , n209902 );
or ( n209904 , n209901 , n209903 );
buf ( n209905 , n209881 );
not ( n209906 , n209905 );
buf ( n209907 , n209906 );
buf ( n209908 , n209907 );
not ( n209909 , n209908 );
buf ( n209910 , n209656 );
not ( n209911 , n209910 );
or ( n209912 , n209909 , n209911 );
buf ( n209913 , n209816 );
buf ( n209914 , n209848 );
and ( n209915 , n209913 , n209914 );
buf ( n209916 , n209842 );
nor ( n209917 , n209915 , n209916 );
buf ( n209918 , n209917 );
buf ( n209919 , n209918 );
nand ( n209920 , n209912 , n209919 );
buf ( n209921 , n209920 );
buf ( n209922 , n209921 );
not ( n209923 , n209922 );
buf ( n209924 , n209923 );
buf ( n209925 , n209924 );
nand ( n209926 , n209904 , n209925 );
buf ( n209927 , n209926 );
buf ( n209928 , n209927 );
not ( n209929 , n209928 );
buf ( n209930 , n209929 );
buf ( n209931 , n209930 );
nand ( n209932 , n209899 , n209931 );
buf ( n209933 , n209932 );
buf ( n209934 , n209933 );
nor ( n209935 , n209890 , n209934 );
buf ( n209936 , n209935 );
buf ( n209937 , n209936 );
buf ( n209938 , n206688 );
not ( n209939 , n209938 );
and ( n209940 , n209836 , n209837 );
buf ( n209941 , n209940 );
buf ( n209942 , n209941 );
not ( n209943 , n209942 );
or ( n209944 , n209939 , n209943 );
buf ( n209945 , n209941 );
buf ( n209946 , n206688 );
or ( n209947 , n209945 , n209946 );
nand ( n209948 , n209944 , n209947 );
buf ( n209949 , n209948 );
buf ( n209950 , n209949 );
and ( n209951 , n209937 , n209950 );
not ( n209952 , n209937 );
buf ( n209953 , n209949 );
not ( n209954 , n209953 );
buf ( n209955 , n209954 );
buf ( n209956 , n209955 );
and ( n209957 , n209952 , n209956 );
nor ( n209958 , n209951 , n209957 );
buf ( n209959 , n209958 );
nand ( n209960 , n209873 , n209959 );
nand ( n209961 , n209872 , n209960 );
buf ( n209962 , n209961 );
not ( n209963 , n209962 );
not ( n209964 , n209963 );
not ( n209965 , n209964 );
not ( n209966 , n209965 );
buf ( n209967 , n209966 );
not ( n209968 , n209967 );
buf ( n209969 , n209968 );
buf ( n209970 , n209969 );
buf ( n209971 , n209970 );
buf ( n209972 , n209971 );
buf ( n209973 , n209972 );
buf ( n209974 , n209973 );
not ( n209975 , n209974 );
and ( n209976 , n209869 , n209975 );
not ( n209977 , n209869 );
and ( n209978 , n209977 , n209974 );
nor ( n209979 , n209976 , n209978 );
and ( n209980 , n209773 , n209868 );
not ( n209981 , n209773 );
and ( n209982 , n209981 , n209867 );
nor ( n209983 , n209980 , n209982 );
and ( n209984 , n209591 , n209770 );
not ( n209985 , n209591 );
and ( n209986 , n209985 , n209771 );
nor ( n209987 , n209984 , n209986 );
not ( n209988 , n39467 );
not ( n209989 , n39134 );
not ( n209990 , n209576 );
or ( n209991 , n209989 , n209990 );
nand ( n209992 , n209991 , n209588 );
not ( n209993 , n209992 );
or ( n209994 , n209988 , n209993 );
nand ( n209995 , n209994 , n209580 );
and ( n209996 , n209995 , n39288 );
not ( n209997 , n209995 );
and ( n209998 , n209997 , n39287 );
nor ( n209999 , n209996 , n209998 );
nand ( n210000 , n39467 , n209580 );
not ( n210001 , n210000 );
and ( n210002 , n209992 , n210001 );
not ( n210003 , n209992 );
and ( n210004 , n210003 , n210000 );
nor ( n210005 , n210002 , n210004 );
not ( n210006 , n39751 );
not ( n210007 , n209568 );
and ( n210008 , n39715 , n39818 );
nand ( n210009 , n209558 , n210008 );
nand ( n210010 , n210007 , n210009 );
not ( n210011 , n210010 );
or ( n210012 , n210006 , n210011 );
nand ( n210013 , n210012 , n209571 );
not ( n210014 , n209574 );
nand ( n210015 , n210014 , n39634 );
not ( n210016 , n210015 );
and ( n210017 , n210013 , n210016 );
not ( n210018 , n210013 );
and ( n210019 , n210018 , n210015 );
nor ( n210020 , n210017 , n210019 );
not ( n210021 , n39133 );
not ( n210022 , n210021 );
not ( n210023 , n209576 );
or ( n210024 , n210022 , n210023 );
nand ( n210025 , n210024 , n209584 );
not ( n210026 , n209576 );
nand ( n210027 , n210021 , n209584 );
and ( n210028 , n210026 , n210027 );
not ( n210029 , n210026 );
not ( n210030 , n210027 );
and ( n210031 , n210029 , n210030 );
nor ( n210032 , n210028 , n210031 );
nand ( n210033 , n209558 , n39818 );
nand ( n210034 , n210033 , n209563 );
not ( n210035 , n39886 );
not ( n210036 , n40052 );
not ( n210037 , n210036 );
not ( n210038 , n209543 );
or ( n210039 , n210037 , n210038 );
not ( n210040 , n209550 );
nand ( n210041 , n210039 , n210040 );
not ( n210042 , n210041 );
or ( n210043 , n210035 , n210042 );
nand ( n210044 , n210043 , n209553 );
not ( n210045 , n40486 );
not ( n210046 , n40424 );
not ( n210047 , n210046 );
not ( n210048 , n40412 );
not ( n210049 , n209508 );
or ( n210050 , n210048 , n210049 );
not ( n210051 , n209527 );
nand ( n210052 , n210050 , n210051 );
not ( n210053 , n210052 );
or ( n210054 , n210047 , n210053 );
not ( n210055 , n209534 );
nand ( n210056 , n210054 , n210055 );
not ( n210057 , n210056 );
or ( n210058 , n210045 , n210057 );
not ( n210059 , n209536 );
nand ( n210060 , n210058 , n210059 );
not ( n210061 , n40398 );
nand ( n210062 , n40411 , n209508 );
not ( n210063 , n40316 );
or ( n210064 , n210062 , n210063 );
not ( n210065 , n209519 );
nand ( n210066 , n210064 , n210065 );
not ( n210067 , n210066 );
or ( n210068 , n210061 , n210067 );
nand ( n210069 , n210068 , n209522 );
not ( n210070 , n40051 );
not ( n210071 , n209543 );
or ( n210072 , n210070 , n210071 );
nand ( n210073 , n210072 , n209547 );
not ( n210074 , n207940 );
not ( n210075 , n40628 );
not ( n210076 , n210075 );
not ( n210077 , n209490 );
not ( n210078 , n209488 );
or ( n210079 , n210077 , n210078 );
not ( n210080 , n40808 );
nand ( n210081 , n210079 , n210080 );
not ( n210082 , n210081 );
or ( n210083 , n210076 , n210082 );
not ( n210084 , n209498 );
nand ( n210085 , n210083 , n210084 );
not ( n210086 , n210085 );
or ( n210087 , n210074 , n210086 );
nand ( n210088 , n210087 , n209501 );
not ( n210089 , n40423 );
not ( n210090 , n210052 );
or ( n210091 , n210089 , n210090 );
not ( n210092 , n209530 );
nand ( n210093 , n210091 , n210092 );
not ( n210094 , n40567 );
not ( n210095 , n210081 );
or ( n210096 , n210094 , n210095 );
not ( n210097 , n209493 );
nand ( n210098 , n210096 , n210097 );
not ( n210099 , n210098 );
nand ( n210100 , n40627 , n209497 );
not ( n210101 , n210100 );
or ( n210102 , n210099 , n210101 );
or ( n210103 , n210100 , n210098 );
nand ( n210104 , n210102 , n210103 );
nand ( n210105 , n207940 , n209501 );
not ( n210106 , n210105 );
not ( n210107 , n210085 );
or ( n210108 , n210106 , n210107 );
or ( n210109 , n210105 , n210085 );
nand ( n210110 , n210108 , n210109 );
nand ( n210111 , n40051 , n209547 );
not ( n210112 , n210111 );
not ( n210113 , n209543 );
or ( n210114 , n210112 , n210113 );
or ( n210115 , n210111 , n209543 );
nand ( n210116 , n210114 , n210115 );
nand ( n210117 , n40423 , n210092 );
not ( n210118 , n210117 );
not ( n210119 , n210052 );
or ( n210120 , n210118 , n210119 );
or ( n210121 , n210117 , n210052 );
nand ( n210122 , n210120 , n210121 );
and ( n210123 , n209488 , n209489 );
and ( n210124 , n210123 , n207988 );
nor ( n210125 , n210124 , n208008 );
not ( n210126 , n40770 );
or ( n210127 , n210125 , n210126 );
not ( n210128 , n40772 );
nand ( n210129 , n210127 , n210128 );
not ( n210130 , n210125 );
nor ( n210131 , n210126 , n40772 );
not ( n210132 , n210131 );
or ( n210133 , n210130 , n210132 );
or ( n210134 , n210131 , n210125 );
nand ( n210135 , n210133 , n210134 );
not ( n210136 , n209508 );
nand ( n210137 , n40411 , n209513 );
not ( n210138 , n210137 );
or ( n210139 , n210136 , n210138 );
or ( n210140 , n210137 , n209508 );
nand ( n210141 , n210139 , n210140 );
not ( n210142 , n210081 );
nand ( n210143 , n40567 , n210097 );
not ( n210144 , n210143 );
or ( n210145 , n210142 , n210144 );
or ( n210146 , n210143 , n210081 );
nand ( n210147 , n210145 , n210146 );
nand ( n210148 , n207988 , n40730 );
not ( n210149 , n210148 );
not ( n210150 , n210123 );
not ( n210151 , n208004 );
nand ( n210152 , n210150 , n210151 );
not ( n210153 , n210152 );
or ( n210154 , n210149 , n210153 );
or ( n210155 , n210148 , n210152 );
nand ( n210156 , n210154 , n210155 );
and ( n210157 , n209471 , n208268 );
nor ( n210158 , n210157 , n209477 );
or ( n210159 , n210158 , n41072 );
nand ( n210160 , n210159 , n209482 );
not ( n210161 , n210160 );
not ( n210162 , n209486 );
nand ( n210163 , n210162 , n209484 );
not ( n210164 , n210163 );
or ( n210165 , n210161 , n210164 );
or ( n210166 , n210163 , n210160 );
nand ( n210167 , n210165 , n210166 );
nand ( n210168 , n209489 , n210151 );
not ( n210169 , n210168 );
not ( n210170 , n209488 );
or ( n210171 , n210169 , n210170 );
or ( n210172 , n210168 , n209488 );
nand ( n210173 , n210171 , n210172 );
not ( n210174 , n40890 );
not ( n210175 , n210174 );
not ( n210176 , n209471 );
or ( n210177 , n210175 , n210176 );
nand ( n210178 , n210177 , n209474 );
not ( n210179 , n210178 );
not ( n210180 , n208267 );
nand ( n210181 , n210180 , n209476 );
not ( n210182 , n210181 );
or ( n210183 , n210179 , n210182 );
or ( n210184 , n210181 , n210178 );
nand ( n210185 , n210183 , n210184 );
not ( n210186 , n41402 );
not ( n210187 , n209451 );
not ( n210188 , n208720 );
nor ( n210189 , n210187 , n210188 );
not ( n210190 , n210189 );
or ( n210191 , n210186 , n210190 );
not ( n210192 , n209462 );
nand ( n210193 , n210191 , n210192 );
nand ( n210194 , n41324 , n210193 );
nand ( n210195 , n210194 , n209465 );
not ( n210196 , n209471 );
nand ( n210197 , n210174 , n209474 );
not ( n210198 , n210197 );
or ( n210199 , n210196 , n210198 );
or ( n210200 , n210197 , n209471 );
nand ( n210201 , n210199 , n210200 );
or ( n210202 , n210189 , n209456 );
not ( n210203 , n210202 );
nand ( n210204 , n41402 , n209461 );
not ( n210205 , n210204 );
or ( n210206 , n210203 , n210205 );
or ( n210207 , n210204 , n210202 );
nand ( n210208 , n210206 , n210207 );
and ( n210209 , n209432 , n209433 );
and ( n210210 , n210209 , n41727 );
nor ( n210211 , n210210 , n41731 );
not ( n210212 , n41721 );
or ( n210213 , n210211 , n210212 );
nand ( n210214 , n210213 , n41734 );
not ( n210215 , n210214 );
nand ( n210216 , n41710 , n41738 );
not ( n210217 , n210216 );
or ( n210218 , n210215 , n210217 );
or ( n210219 , n210216 , n210214 );
nand ( n210220 , n210218 , n210219 );
not ( n210221 , n41614 );
nand ( n210222 , n210221 , n209440 );
not ( n210223 , n210222 );
or ( n210224 , n209435 , n41739 );
not ( n210225 , n210224 );
not ( n210226 , n208728 );
not ( n210227 , n210226 );
or ( n210228 , n210225 , n210227 );
nand ( n210229 , n210228 , n209438 );
not ( n210230 , n210229 );
or ( n210231 , n210223 , n210230 );
or ( n210232 , n210222 , n210229 );
nand ( n210233 , n210231 , n210232 );
nor ( n210234 , n210188 , n209456 );
not ( n210235 , n210234 );
not ( n210236 , n210187 );
or ( n210237 , n210235 , n210236 );
or ( n210238 , n210234 , n210187 );
nand ( n210239 , n210237 , n210238 );
not ( n210240 , n210211 );
and ( n210241 , n41721 , n41734 );
not ( n210242 , n210241 );
or ( n210243 , n210240 , n210242 );
or ( n210244 , n210241 , n210211 );
nand ( n210245 , n210243 , n210244 );
nand ( n210246 , n41727 , n41730 );
not ( n210247 , n210246 );
not ( n210248 , n210209 );
not ( n210249 , n41723 );
nand ( n210250 , n210248 , n210249 );
not ( n210251 , n210250 );
or ( n210252 , n210247 , n210251 );
or ( n210253 , n210246 , n210250 );
nand ( n210254 , n210252 , n210253 );
nand ( n210255 , n209433 , n210249 );
not ( n210256 , n210255 );
not ( n210257 , n209432 );
or ( n210258 , n210256 , n210257 );
or ( n210259 , n210255 , n209432 );
nand ( n210260 , n210258 , n210259 );
nand ( n210261 , n209113 , n209431 );
not ( n210262 , n210261 );
not ( n210263 , n209421 );
and ( n210264 , n209420 , n210263 );
and ( n210265 , n210264 , n209245 );
nor ( n210266 , n210265 , n209251 );
or ( n210267 , n210266 , n41895 );
nand ( n210268 , n210267 , n209427 );
not ( n210269 , n210268 );
or ( n210270 , n210262 , n210269 );
or ( n210271 , n210261 , n210268 );
nand ( n210272 , n210270 , n210271 );
not ( n210273 , n210266 );
and ( n210274 , n209173 , n209427 );
not ( n210275 , n210274 );
or ( n210276 , n210273 , n210275 );
or ( n210277 , n210274 , n210266 );
nand ( n210278 , n210276 , n210277 );
nand ( n210279 , n209245 , n41973 );
not ( n210280 , n210279 );
not ( n210281 , n210264 );
nand ( n210282 , n210281 , n41898 );
not ( n210283 , n210282 );
or ( n210284 , n210280 , n210283 );
or ( n210285 , n210279 , n210282 );
nand ( n210286 , n210284 , n210285 );
not ( n210287 , n209418 );
nand ( n210288 , n210287 , n209407 );
not ( n210289 , n210288 );
and ( n210290 , n209404 , n209260 );
nor ( n210291 , n210290 , n209411 );
not ( n210292 , n209257 );
or ( n210293 , n210291 , n210292 );
nand ( n210294 , n210293 , n209415 );
not ( n210295 , n210294 );
or ( n210296 , n210289 , n210295 );
or ( n210297 , n210288 , n210294 );
nand ( n210298 , n210296 , n210297 );
nand ( n210299 , n210263 , n41898 );
not ( n210300 , n210299 );
not ( n210301 , n209420 );
or ( n210302 , n210300 , n210301 );
or ( n210303 , n210299 , n209420 );
nand ( n210304 , n210302 , n210303 );
not ( n210305 , n210291 );
and ( n210306 , n209257 , n209415 );
not ( n210307 , n210306 );
or ( n210308 , n210305 , n210307 );
or ( n210309 , n210306 , n210291 );
nand ( n210310 , n210308 , n210309 );
nand ( n210311 , n209260 , n209410 );
not ( n210312 , n210311 );
not ( n210313 , n209404 );
nand ( n210314 , n210313 , n209408 );
not ( n210315 , n210314 );
or ( n210316 , n210312 , n210315 );
or ( n210317 , n210311 , n210314 );
nand ( n210318 , n210316 , n210317 );
nand ( n210319 , n209403 , n209408 );
not ( n210320 , n210319 );
not ( n210321 , n209402 );
or ( n210322 , n210320 , n210321 );
or ( n210323 , n210319 , n209402 );
nand ( n210324 , n210322 , n210323 );
xor ( n210325 , n209264 , n18560 );
xor ( n210326 , n210325 , n209399 );
nand ( n210327 , n209318 , n209398 );
not ( n210328 , n210327 );
not ( n210329 , n209395 );
or ( n210330 , n210328 , n210329 );
or ( n210331 , n210327 , n209395 );
nand ( n210332 , n210330 , n210331 );
nand ( n210333 , n209349 , n209394 );
not ( n210334 , n210333 );
not ( n210335 , n209391 );
or ( n210336 , n210334 , n210335 );
or ( n210337 , n210333 , n209391 );
nand ( n210338 , n210336 , n210337 );
nand ( n210339 , n209361 , n209390 );
not ( n210340 , n210339 );
not ( n210341 , n209387 );
or ( n210342 , n210340 , n210341 );
or ( n210343 , n210339 , n209387 );
nand ( n210344 , n210342 , n210343 );
not ( n210345 , n209379 );
nand ( n210346 , n209367 , n209382 );
not ( n210347 , n210346 );
or ( n210348 , n210345 , n210347 );
or ( n210349 , n209379 , n210346 );
nand ( n210350 , n210348 , n210349 );
not ( n210351 , n209378 );
nor ( n210352 , n210351 , n209369 );
not ( n210353 , n210352 );
not ( n210354 , n209376 );
or ( n210355 , n210353 , n210354 );
or ( n210356 , n209376 , n210352 );
nand ( n210357 , n210355 , n210356 );
nand ( n210358 , n40804 , n208084 );
and ( n210359 , n41324 , n209465 );
not ( n210360 , n209504 );
nand ( n210361 , n210360 , n40670 );
nand ( n210362 , n39886 , n209553 );
not ( n210363 , n39998 );
nand ( n210364 , n210363 , n209549 );
nand ( n210365 , n39751 , n209571 );
nand ( n210366 , n39715 , n209567 );
nand ( n210367 , n39818 , n209563 );
not ( n210368 , n209556 );
nand ( n210369 , n210368 , n39934 );
not ( n210370 , n209538 );
nand ( n210371 , n210370 , n209540 );
nand ( n210372 , n40486 , n210059 );
nand ( n210373 , n40420 , n209533 );
nor ( n210374 , n209445 , n41702 );
nor ( n210375 , n41251 , n209469 );
nand ( n210376 , n40184 , n209526 );
nand ( n210377 , n40398 , n209522 );
nor ( n210378 , n39014 , n209587 );
xnor ( n210379 , n210010 , n210365 );
xnor ( n210380 , n210129 , n210358 );
xnor ( n210381 , n210088 , n210361 );
xnor ( n210382 , n210041 , n210362 );
xnor ( n210383 , n210073 , n210364 );
xnor ( n210384 , n210034 , n210366 );
xnor ( n210385 , n209558 , n210367 );
xnor ( n210386 , n210044 , n210369 );
xnor ( n210387 , n210060 , n210371 );
xnor ( n210388 , n210056 , n210372 );
xnor ( n210389 , n210093 , n210373 );
xor ( n210390 , n210195 , n210375 );
xnor ( n210391 , n210069 , n210376 );
xnor ( n210392 , n210066 , n210377 );
xor ( n210393 , n210025 , n210378 );
buf ( n210394 , n204222 );
buf ( n210395 , n204201 );
buf ( n210396 , n209867 );
xor ( n210397 , n210394 , n210395 );
xor ( n210398 , n210397 , n210396 );
buf ( n210399 , n210398 );
xor ( n210400 , n210394 , n210395 );
and ( n210401 , n210400 , n210396 );
and ( n210402 , n210394 , n210395 );
or ( n210403 , n210401 , n210402 );
buf ( n210404 , n210403 );
buf ( n210405 , n204231 );
buf ( n210406 , n204228 );
buf ( n210407 , n209711 );
xor ( n210408 , n210405 , n210406 );
xor ( n210409 , n210408 , n210407 );
buf ( n210410 , n210409 );
xor ( n210411 , n210405 , n210406 );
and ( n210412 , n210411 , n210407 );
and ( n210413 , n210405 , n210406 );
or ( n210414 , n210412 , n210413 );
buf ( n210415 , n210414 );
buf ( n210416 , n203636 );
buf ( n210417 , n29604 );
buf ( n210418 , n39288 );
xor ( n210419 , n210416 , n210417 );
xor ( n210420 , n210419 , n210418 );
buf ( n210421 , n210420 );
xor ( n210422 , n210416 , n210417 );
and ( n210423 , n210422 , n210418 );
and ( n210424 , n210416 , n210417 );
or ( n210425 , n210423 , n210424 );
buf ( n210426 , n210425 );
buf ( n210427 , n204537 );
buf ( n210428 , n204540 );
not ( n210429 , n209972 );
buf ( n210430 , n210429 );
xor ( n210431 , n210427 , n210428 );
xor ( n210432 , n210431 , n210430 );
buf ( n210433 , n210432 );
xor ( n210434 , n210427 , n210428 );
and ( n210435 , n210434 , n210430 );
and ( n210436 , n210427 , n210428 );
or ( n210437 , n210435 , n210436 );
buf ( n210438 , n210437 );
buf ( n210439 , n203256 );
buf ( n210440 , n27541 );
buf ( n210441 , n30412 );
xor ( n210442 , n210439 , n210440 );
xor ( n210443 , n210442 , n210441 );
buf ( n210444 , n210443 );
xor ( n210445 , n210439 , n210440 );
and ( n210446 , n210445 , n210441 );
and ( n210447 , n210439 , n210440 );
or ( n210448 , n210446 , n210447 );
buf ( n210449 , n210448 );
buf ( n210450 , n203153 );
buf ( n210451 , n203151 );
buf ( n210452 , n41981 );
xor ( n210453 , n210450 , n210451 );
xor ( n210454 , n210453 , n210452 );
buf ( n210455 , n210454 );
xor ( n210456 , n210450 , n210451 );
and ( n210457 , n210456 , n210452 );
and ( n210458 , n210450 , n210451 );
or ( n210459 , n210457 , n210458 );
buf ( n210460 , n210459 );
buf ( n210461 , n203424 );
buf ( n210462 , n203418 );
buf ( n210463 , n30384 );
xor ( n210464 , n210461 , n210462 );
xor ( n210465 , n210464 , n210463 );
buf ( n210466 , n210465 );
xor ( n210467 , n210461 , n210462 );
and ( n210468 , n210467 , n210463 );
and ( n210469 , n210461 , n210462 );
or ( n210470 , n210468 , n210469 );
buf ( n210471 , n210470 );
buf ( n210472 , n36087 );
buf ( n210473 , n203397 );
buf ( n210474 , n30292 );
xor ( n210475 , n210472 , n210473 );
xor ( n210476 , n210475 , n210474 );
buf ( n210477 , n210476 );
xor ( n210478 , n210472 , n210473 );
and ( n210479 , n210478 , n210474 );
and ( n210480 , n210472 , n210473 );
or ( n210481 , n210479 , n210480 );
buf ( n210482 , n210481 );
buf ( n210483 , n23372 );
buf ( n210484 , n203463 );
buf ( n210485 , n41834 );
xor ( n210486 , n210483 , n210484 );
xor ( n210487 , n210486 , n210485 );
buf ( n210488 , n210487 );
xor ( n210489 , n210483 , n210484 );
and ( n210490 , n210489 , n210485 );
and ( n210491 , n210483 , n210484 );
or ( n210492 , n210490 , n210491 );
buf ( n210493 , n210492 );
buf ( n210494 , n203102 );
buf ( n210495 , n27363 );
buf ( n210496 , n30997 );
xor ( n210497 , n210494 , n210495 );
xor ( n210498 , n210497 , n210496 );
buf ( n210499 , n210498 );
xor ( n210500 , n210494 , n210495 );
and ( n210501 , n210500 , n210496 );
and ( n210502 , n210494 , n210495 );
or ( n210503 , n210501 , n210502 );
buf ( n210504 , n210503 );
buf ( n210505 , n203093 );
buf ( n210506 , n203088 );
buf ( n210507 , n41725 );
xor ( n210508 , n210505 , n210506 );
xor ( n210509 , n210508 , n210507 );
buf ( n210510 , n210509 );
xor ( n210511 , n210505 , n210506 );
and ( n210512 , n210511 , n210507 );
and ( n210513 , n210505 , n210506 );
or ( n210514 , n210512 , n210513 );
buf ( n210515 , n210514 );
buf ( n210516 , n203080 );
buf ( n210517 , n27635 );
buf ( n210518 , n41716 );
xor ( n210519 , n210516 , n210517 );
xor ( n210520 , n210519 , n210518 );
buf ( n210521 , n210520 );
xor ( n210522 , n210516 , n210517 );
and ( n210523 , n210522 , n210518 );
and ( n210524 , n210516 , n210517 );
or ( n210525 , n210523 , n210524 );
buf ( n210526 , n210525 );
buf ( n210527 , n203059 );
buf ( n210528 , n203053 );
buf ( n210529 , n30962 );
xor ( n210530 , n210527 , n210528 );
xor ( n210531 , n210530 , n210529 );
buf ( n210532 , n210531 );
xor ( n210533 , n210527 , n210528 );
and ( n210534 , n210533 , n210529 );
and ( n210535 , n210527 , n210528 );
or ( n210536 , n210534 , n210535 );
buf ( n210537 , n210536 );
buf ( n210538 , n202964 );
buf ( n210539 , n202959 );
buf ( n210540 , n208717 );
xor ( n210541 , n210538 , n210539 );
xor ( n210542 , n210541 , n210540 );
buf ( n210543 , n210542 );
xor ( n210544 , n210538 , n210539 );
and ( n210545 , n210544 , n210540 );
and ( n210546 , n210538 , n210539 );
or ( n210547 , n210545 , n210546 );
buf ( n210548 , n210547 );
buf ( n210549 , n28601 );
buf ( n210550 , n202899 );
buf ( n210551 , n41250 );
xor ( n210552 , n210549 , n210550 );
xor ( n210553 , n210552 , n210551 );
buf ( n210554 , n210553 );
xor ( n210555 , n210549 , n210550 );
and ( n210556 , n210555 , n210551 );
and ( n210557 , n210549 , n210550 );
or ( n210558 , n210556 , n210557 );
buf ( n210559 , n210558 );
buf ( n210560 , n202848 );
not ( n210561 , n36991 );
buf ( n210562 , n210561 );
buf ( n210563 , n41071 );
xor ( n210564 , n210560 , n210562 );
xor ( n210565 , n210564 , n210563 );
buf ( n210566 , n210565 );
xor ( n210567 , n210560 , n210562 );
and ( n210568 , n210567 , n210563 );
and ( n210569 , n210560 , n210562 );
or ( n210570 , n210568 , n210569 );
buf ( n210571 , n210570 );
buf ( n210572 , n35596 );
buf ( n210573 , n202852 );
buf ( n210574 , n208261 );
xor ( n210575 , n210572 , n210573 );
xor ( n210576 , n210575 , n210574 );
buf ( n210577 , n210576 );
xor ( n210578 , n210572 , n210573 );
and ( n210579 , n210578 , n210574 );
and ( n210580 , n210572 , n210573 );
or ( n210581 , n210579 , n210580 );
buf ( n210582 , n210581 );
buf ( n210583 , n202753 );
not ( n210584 , n36287 );
buf ( n210585 , n210584 );
buf ( n210586 , n208002 );
xor ( n210587 , n210583 , n210585 );
xor ( n210588 , n210587 , n210586 );
buf ( n210589 , n210588 );
xor ( n210590 , n210583 , n210585 );
and ( n210591 , n210590 , n210586 );
and ( n210592 , n210583 , n210585 );
or ( n210593 , n210591 , n210592 );
buf ( n210594 , n210593 );
buf ( n210595 , n40710 );
buf ( n210596 , n202503 );
buf ( n210597 , n210596 );
buf ( n210598 , n202416 );
xor ( n210599 , n210595 , n210597 );
xor ( n210600 , n210599 , n210598 );
buf ( n210601 , n210600 );
xor ( n210602 , n210595 , n210597 );
and ( n210603 , n210602 , n210598 );
and ( n210604 , n210595 , n210597 );
or ( n210605 , n210603 , n210604 );
buf ( n210606 , n210605 );
buf ( n210607 , n202566 );
buf ( n210608 , n202583 );
buf ( n210609 , n210608 );
buf ( n210610 , n210609 );
buf ( n210611 , n40802 );
xor ( n210612 , n210607 , n210610 );
xor ( n210613 , n210612 , n210611 );
buf ( n210614 , n210613 );
xor ( n210615 , n210607 , n210610 );
and ( n210616 , n210615 , n210611 );
and ( n210617 , n210607 , n210610 );
or ( n210618 , n210616 , n210617 );
buf ( n210619 , n210618 );
buf ( n210620 , n202592 );
buf ( n210621 , n210620 );
not ( n210622 , n36310 );
buf ( n210623 , n210622 );
buf ( n210624 , n40562 );
xor ( n210625 , n210621 , n210623 );
xor ( n210626 , n210625 , n210624 );
buf ( n210627 , n210626 );
xor ( n210628 , n210621 , n210623 );
and ( n210629 , n210628 , n210624 );
and ( n210630 , n210621 , n210623 );
or ( n210631 , n210629 , n210630 );
buf ( n210632 , n210631 );
not ( n210633 , n33680 );
buf ( n210634 , n210633 );
buf ( n210635 , n27547 );
buf ( n210636 , n207938 );
xor ( n210637 , n210634 , n210635 );
xor ( n210638 , n210637 , n210636 );
buf ( n210639 , n210638 );
xor ( n210640 , n210634 , n210635 );
and ( n210641 , n210640 , n210636 );
and ( n210642 , n210634 , n210635 );
or ( n210643 , n210641 , n210642 );
buf ( n210644 , n210643 );
buf ( n210645 , n22559 );
buf ( n210646 , n200923 );
buf ( n210647 , n210646 );
buf ( n210648 , n40259 );
xor ( n210649 , n210645 , n210647 );
xor ( n210650 , n210649 , n210648 );
buf ( n210651 , n210650 );
xor ( n210652 , n210645 , n210647 );
and ( n210653 , n210652 , n210648 );
and ( n210654 , n210645 , n210647 );
or ( n210655 , n210653 , n210654 );
buf ( n210656 , n210655 );
buf ( n210657 , n24108 );
buf ( n210658 , n37543 );
buf ( n210659 , n40182 );
xor ( n210660 , n210657 , n210658 );
xor ( n210661 , n210660 , n210659 );
buf ( n210662 , n210661 );
xor ( n210663 , n210657 , n210658 );
and ( n210664 , n210663 , n210659 );
and ( n210665 , n210657 , n210658 );
or ( n210666 , n210664 , n210665 );
buf ( n210667 , n210666 );
buf ( n210668 , n200834 );
not ( n210669 , n33509 );
buf ( n210670 , n210669 );
buf ( n210671 , n40414 );
xor ( n210672 , n210668 , n210670 );
xor ( n210673 , n210672 , n210671 );
buf ( n210674 , n210673 );
xor ( n210675 , n210668 , n210670 );
and ( n210676 , n210675 , n210671 );
and ( n210677 , n210668 , n210670 );
or ( n210678 , n210676 , n210677 );
buf ( n210679 , n210678 );
buf ( n210680 , n200137 );
buf ( n210681 , n200120 );
buf ( n210682 , n39368 );
xor ( n210683 , n210680 , n210681 );
xor ( n210684 , n210683 , n210682 );
buf ( n210685 , n210684 );
xor ( n210686 , n210680 , n210681 );
and ( n210687 , n210686 , n210682 );
and ( n210688 , n210680 , n210681 );
or ( n210689 , n210687 , n210688 );
buf ( n210690 , n210689 );
buf ( n210691 , n200567 );
buf ( n210692 , n200622 );
buf ( n210693 , n39997 );
xor ( n210694 , n210691 , n210692 );
xor ( n210695 , n210694 , n210693 );
buf ( n210696 , n210695 );
xor ( n210697 , n210691 , n210692 );
and ( n210698 , n210697 , n210693 );
and ( n210699 , n210691 , n210692 );
or ( n210700 , n210698 , n210699 );
buf ( n210701 , n210700 );
buf ( n210702 , n200663 );
buf ( n210703 , n200657 );
buf ( n210704 , n210703 );
buf ( n210705 , n39880 );
xor ( n210706 , n210702 , n210704 );
xor ( n210707 , n210706 , n210705 );
buf ( n210708 , n210707 );
xor ( n210709 , n210702 , n210704 );
and ( n210710 , n210709 , n210705 );
and ( n210711 , n210702 , n210704 );
or ( n210712 , n210710 , n210711 );
buf ( n210713 , n210712 );
buf ( n210714 , n33419 );
buf ( n210715 , n33424 );
buf ( n210716 , n39812 );
xor ( n210717 , n210714 , n210715 );
xor ( n210718 , n210717 , n210716 );
buf ( n210719 , n210718 );
xor ( n210720 , n210714 , n210715 );
and ( n210721 , n210720 , n210716 );
and ( n210722 , n210714 , n210715 );
or ( n210723 , n210721 , n210722 );
buf ( n210724 , n210723 );
buf ( n210725 , n203833 );
buf ( n210726 , n203704 );
buf ( n210727 , n209770 );
xor ( n210728 , n210725 , n210726 );
xor ( n210729 , n210728 , n210727 );
buf ( n210730 , n210729 );
xor ( n210731 , n210725 , n210726 );
and ( n210732 , n210731 , n210727 );
and ( n210733 , n210725 , n210726 );
or ( n210734 , n210732 , n210733 );
buf ( n210735 , n210734 );
buf ( n210736 , n200074 );
buf ( n210737 , n200080 );
buf ( n210738 , n39089 );
xor ( n210739 , n210736 , n210737 );
xor ( n210740 , n210739 , n210738 );
buf ( n210741 , n210740 );
xor ( n210742 , n210736 , n210737 );
and ( n210743 , n210742 , n210738 );
and ( n210744 , n210736 , n210737 );
or ( n210745 , n210743 , n210744 );
buf ( n210746 , n210745 );
buf ( n210747 , n204603 );
buf ( n210748 , n204548 );
xor ( n210749 , n210747 , n210748 );
buf ( n210750 , n210749 );
and ( n210751 , n210747 , n210748 );
buf ( n210752 , n210751 );
buf ( n210753 , n204530 );
buf ( n210754 , n204468 );
xor ( n210755 , n210753 , n210754 );
buf ( n210756 , n210755 );
and ( n210757 , n210753 , n210754 );
buf ( n210758 , n210757 );
buf ( n210759 , n204655 );
buf ( n210760 , n204609 );
xor ( n210761 , n210759 , n210760 );
buf ( n210762 , n210761 );
and ( n210763 , n210759 , n210760 );
buf ( n210764 , n210763 );
buf ( n210765 , n204688 );
buf ( n210766 , n204662 );
xor ( n210767 , n210765 , n210766 );
buf ( n210768 , n210767 );
and ( n210769 , n210765 , n210766 );
buf ( n210770 , n210769 );
buf ( n210771 , n204943 );
buf ( n210772 , n204937 );
xor ( n210773 , n210771 , n210772 );
buf ( n210774 , n210773 );
buf ( n210775 , n210768 );
buf ( n210776 , n210764 );
buf ( n210777 , n210758 );
buf ( n210778 , n210750 );
or ( n210779 , n210777 , n210778 );
buf ( n210780 , n210779 );
buf ( n210781 , n210780 );
not ( n210782 , n210781 );
buf ( n210783 , n210752 );
buf ( n210784 , n210762 );
nor ( n210785 , n210783 , n210784 );
buf ( n210786 , n210785 );
buf ( n210787 , n210786 );
nor ( n210788 , n210782 , n210787 );
buf ( n210789 , n210788 );
buf ( n210790 , n210789 );
not ( n210791 , n210790 );
buf ( n210792 , n199998 );
buf ( n210793 , n199832 );
xor ( n210794 , n210792 , n210793 );
buf ( n210795 , n39608 );
xor ( n210796 , n210794 , n210795 );
buf ( n210797 , n210796 );
buf ( n210798 , n210797 );
not ( n210799 , n210798 );
xor ( n210800 , n199823 , n26412 );
and ( n210801 , n210800 , n39749 );
and ( n210802 , n199823 , n26412 );
nor ( n210803 , n210801 , n210802 );
buf ( n210804 , n210803 );
nand ( n210805 , n210799 , n210804 );
buf ( n210806 , n210805 );
buf ( n210807 , n210806 );
xor ( n210808 , n210792 , n210793 );
and ( n210809 , n210808 , n210795 );
and ( n210810 , n210792 , n210793 );
or ( n210811 , n210809 , n210810 );
buf ( n210812 , n210811 );
buf ( n210813 , n210812 );
buf ( n210814 , n210741 );
or ( n210815 , n210813 , n210814 );
buf ( n210816 , n210815 );
buf ( n210817 , n210816 );
and ( n210818 , n210807 , n210817 );
buf ( n210819 , n210818 );
buf ( n210820 , n210819 );
buf ( n210821 , n210724 );
xnor ( n210822 , n20129 , n32538 );
not ( n210823 , n39714 );
and ( n210824 , n210822 , n210823 );
not ( n210825 , n210822 );
and ( n210826 , n210825 , n39714 );
nor ( n210827 , n210824 , n210826 );
buf ( n210828 , n210827 );
nor ( n210829 , n210821 , n210828 );
buf ( n210830 , n210829 );
buf ( n210831 , n210830 );
xor ( n210832 , n199823 , n26412 );
xor ( n210833 , n210832 , n39749 );
or ( n210834 , n20129 , n32538 );
not ( n210835 , n210834 );
not ( n210836 , n39714 );
or ( n210837 , n210835 , n210836 );
nand ( n210838 , n20129 , n32538 );
nand ( n210839 , n210837 , n210838 );
nor ( n210840 , n210833 , n210839 );
buf ( n210841 , n210840 );
nor ( n210842 , n210831 , n210841 );
buf ( n210843 , n210842 );
buf ( n210844 , n210843 );
nand ( n210845 , n210820 , n210844 );
buf ( n210846 , n210845 );
buf ( n210847 , n210846 );
buf ( n210848 , n210746 );
buf ( n210849 , n200146 );
buf ( n210850 , n210849 );
buf ( n210851 , n200141 );
buf ( n210852 , n210851 );
xor ( n210853 , n210850 , n210852 );
buf ( n210854 , n38533 );
xor ( n210855 , n210853 , n210854 );
buf ( n210856 , n210855 );
buf ( n210857 , n210856 );
nor ( n210858 , n210848 , n210857 );
buf ( n210859 , n210858 );
buf ( n210860 , n210859 );
buf ( n210861 , n210685 );
xor ( n210862 , n210850 , n210852 );
and ( n210863 , n210862 , n210854 );
and ( n210864 , n210850 , n210852 );
or ( n210865 , n210863 , n210864 );
buf ( n210866 , n210865 );
buf ( n210867 , n210866 );
nor ( n210868 , n210861 , n210867 );
buf ( n210869 , n210868 );
buf ( n210870 , n210869 );
nor ( n210871 , n210860 , n210870 );
buf ( n210872 , n210871 );
buf ( n210873 , n210872 );
buf ( n210874 , n210730 );
buf ( n210875 , n210426 );
nor ( n210876 , n210874 , n210875 );
buf ( n210877 , n210876 );
buf ( n210878 , n210877 );
buf ( n210879 , n210421 );
buf ( n210880 , n210690 );
nor ( n210881 , n210879 , n210880 );
buf ( n210882 , n210881 );
buf ( n210883 , n210882 );
nor ( n210884 , n210878 , n210883 );
buf ( n210885 , n210884 );
buf ( n210886 , n210885 );
nand ( n210887 , n210873 , n210886 );
buf ( n210888 , n210887 );
buf ( n210889 , n210888 );
nor ( n210890 , n210847 , n210889 );
buf ( n210891 , n210890 );
buf ( n210892 , n210891 );
not ( n210893 , n210892 );
buf ( n210894 , n210708 );
buf ( n210895 , n210701 );
nor ( n210896 , n210894 , n210895 );
buf ( n210897 , n210896 );
buf ( n210898 , n210897 );
buf ( n210899 , n200729 );
buf ( n210900 , n200709 );
buf ( n210901 , n210900 );
xor ( n210902 , n210899 , n210901 );
buf ( n210903 , n40045 );
and ( n210904 , n210902 , n210903 );
and ( n210905 , n210899 , n210901 );
or ( n210906 , n210904 , n210905 );
buf ( n210907 , n210906 );
buf ( n210908 , n210907 );
buf ( n210909 , n210696 );
nor ( n210910 , n210908 , n210909 );
buf ( n210911 , n210910 );
buf ( n210912 , n210911 );
nor ( n210913 , n210898 , n210912 );
buf ( n210914 , n210913 );
buf ( n210915 , n210914 );
buf ( n210916 , n210719 );
not ( n210917 , n210916 );
xor ( n210918 , n33415 , n200671 );
not ( n210919 , n39928 );
and ( n210920 , n210918 , n210919 );
and ( n210921 , n33415 , n200671 );
or ( n210922 , n210920 , n210921 );
buf ( n210923 , n210922 );
not ( n210924 , n210923 );
buf ( n210925 , n210924 );
buf ( n210926 , n210925 );
nand ( n210927 , n210917 , n210926 );
buf ( n210928 , n210927 );
buf ( n210929 , n210928 );
xor ( n210930 , n33415 , n200671 );
xor ( n210931 , n210930 , n210919 );
buf ( n210932 , n210931 );
not ( n210933 , n210932 );
buf ( n210934 , n210713 );
not ( n210935 , n210934 );
buf ( n210936 , n210935 );
buf ( n210937 , n210936 );
nand ( n210938 , n210933 , n210937 );
buf ( n210939 , n210938 );
buf ( n210940 , n210939 );
and ( n210941 , n210915 , n210929 , n210940 );
buf ( n210942 , n210941 );
buf ( n210943 , n210942 );
not ( n210944 , n210943 );
xor ( n210945 , n210899 , n210901 );
xor ( n210946 , n210945 , n210903 );
buf ( n210947 , n210946 );
buf ( n210948 , n210947 );
not ( n210949 , n210948 );
xor ( n210950 , n26418 , n40548 );
not ( n210951 , n33459 );
and ( n210952 , n210950 , n210951 );
and ( n210953 , n26418 , n40548 );
or ( n210954 , n210952 , n210953 );
not ( n210955 , n210954 );
buf ( n210956 , n210955 );
nand ( n210957 , n210949 , n210956 );
buf ( n210958 , n210957 );
buf ( n210959 , n210958 );
not ( n210960 , n210959 );
buf ( n210961 , n210674 );
buf ( n210962 , n34077 );
buf ( n210963 , n201332 );
xor ( n210964 , n210962 , n210963 );
buf ( n210965 , n40422 );
and ( n210966 , n210964 , n210965 );
and ( n210967 , n210962 , n210963 );
or ( n210968 , n210966 , n210967 );
buf ( n210969 , n210968 );
buf ( n210970 , n210969 );
nand ( n210971 , n210961 , n210970 );
buf ( n210972 , n210971 );
buf ( n210973 , n210679 );
buf ( n210974 , n200843 );
xor ( n210975 , n210974 , n26216 );
xor ( n210976 , n210975 , n40485 );
buf ( n210977 , n210976 );
nor ( n210978 , n210973 , n210977 );
buf ( n210979 , n210978 );
or ( n210980 , n210972 , n210979 );
buf ( n210981 , n210679 );
buf ( n210982 , n210976 );
nand ( n210983 , n210981 , n210982 );
buf ( n210984 , n210983 );
nand ( n210985 , n210980 , n210984 );
not ( n210986 , n210985 );
xor ( n210987 , n26418 , n40548 );
not ( n210988 , n33459 );
xor ( n210989 , n210987 , n210988 );
xor ( n210990 , n210974 , n26216 );
and ( n210991 , n210990 , n40485 );
and ( n210992 , n210974 , n26216 );
nor ( n210993 , n210991 , n210992 );
not ( n210994 , n210993 );
or ( n210995 , n210989 , n210994 );
not ( n210996 , n210995 );
or ( n210997 , n210986 , n210996 );
not ( n210998 , n210993 );
nand ( n210999 , n210998 , n210989 );
nand ( n211000 , n210997 , n210999 );
buf ( n211001 , n211000 );
not ( n211002 , n211001 );
or ( n211003 , n210960 , n211002 );
buf ( n211004 , n210955 );
not ( n211005 , n211004 );
buf ( n211006 , n210947 );
nand ( n211007 , n211005 , n211006 );
buf ( n211008 , n211007 );
buf ( n211009 , n211008 );
nand ( n211010 , n211003 , n211009 );
buf ( n211011 , n211010 );
buf ( n211012 , n211011 );
not ( n211013 , n211012 );
or ( n211014 , n210944 , n211013 );
buf ( n211015 , n210939 );
not ( n211016 , n211015 );
buf ( n211017 , n210907 );
buf ( n211018 , n210696 );
and ( n211019 , n211017 , n211018 );
buf ( n211020 , n211019 );
buf ( n211021 , n211020 );
not ( n211022 , n211021 );
buf ( n211023 , n210897 );
not ( n211024 , n211023 );
buf ( n211025 , n211024 );
buf ( n211026 , n211025 );
not ( n211027 , n211026 );
or ( n211028 , n211022 , n211027 );
buf ( n211029 , n210708 );
buf ( n211030 , n210701 );
nand ( n211031 , n211029 , n211030 );
buf ( n211032 , n211031 );
buf ( n211033 , n211032 );
nand ( n211034 , n211028 , n211033 );
buf ( n211035 , n211034 );
buf ( n211036 , n211035 );
not ( n211037 , n211036 );
or ( n211038 , n211016 , n211037 );
buf ( n211039 , n210936 );
not ( n211040 , n211039 );
buf ( n211041 , n210931 );
nand ( n211042 , n211040 , n211041 );
buf ( n211043 , n211042 );
buf ( n211044 , n211043 );
nand ( n211045 , n211038 , n211044 );
buf ( n211046 , n211045 );
buf ( n211047 , n211046 );
buf ( n211048 , n210928 );
and ( n211049 , n211047 , n211048 );
buf ( n211050 , n210925 );
not ( n211051 , n211050 );
buf ( n211052 , n210719 );
nand ( n211053 , n211051 , n211052 );
buf ( n211054 , n211053 );
buf ( n211055 , n211054 );
not ( n211056 , n211055 );
buf ( n211057 , n211056 );
buf ( n211058 , n211057 );
nor ( n211059 , n211049 , n211058 );
buf ( n211060 , n211059 );
buf ( n211061 , n211060 );
nand ( n211062 , n211014 , n211061 );
buf ( n211063 , n211062 );
buf ( n211064 , n211063 );
not ( n211065 , n211064 );
buf ( n211066 , n210942 );
buf ( n211067 , n210995 );
or ( n211068 , n210969 , n210674 );
buf ( n211069 , n211068 );
buf ( n211070 , n210958 );
buf ( n211071 , n210979 );
not ( n211072 , n211071 );
buf ( n211073 , n211072 );
buf ( n211074 , n211073 );
and ( n211075 , n211067 , n211069 , n211070 , n211074 );
buf ( n211076 , n211075 );
buf ( n211077 , n211076 );
and ( n211078 , n211066 , n211077 );
buf ( n211079 , n211078 );
buf ( n211080 , n211079 );
buf ( n211081 , n202886 );
buf ( n211082 , n202880 );
buf ( n211083 , n211082 );
xor ( n211084 , n211081 , n211083 );
buf ( n211085 , n41319 );
xor ( n211086 , n211084 , n211085 );
buf ( n211087 , n211086 );
buf ( n211088 , n211087 );
buf ( n211089 , n29022 );
buf ( n211090 , n28933 );
xor ( n211091 , n211089 , n211090 );
buf ( n211092 , n41397 );
and ( n211093 , n211091 , n211092 );
and ( n211094 , n211089 , n211090 );
or ( n211095 , n211093 , n211094 );
buf ( n211096 , n211095 );
buf ( n211097 , n211096 );
nor ( n211098 , n211088 , n211097 );
buf ( n211099 , n211098 );
buf ( n211100 , n211099 );
xor ( n211101 , n211089 , n211090 );
xor ( n211102 , n211101 , n211092 );
buf ( n211103 , n211102 );
buf ( n211104 , n211103 );
buf ( n211105 , n210548 );
nor ( n211106 , n211104 , n211105 );
buf ( n211107 , n211106 );
buf ( n211108 , n211107 );
nor ( n211109 , n211100 , n211108 );
buf ( n211110 , n211109 );
buf ( n211111 , n211110 );
xor ( n211112 , n211081 , n211083 );
and ( n211113 , n211112 , n211085 );
and ( n211114 , n211081 , n211083 );
or ( n211115 , n211113 , n211114 );
buf ( n211116 , n211115 );
or ( n211117 , n210554 , n211116 );
buf ( n211118 , n211117 );
buf ( n211119 , n29906 );
not ( n211120 , n35727 );
buf ( n211121 , n211120 );
xor ( n211122 , n211119 , n211121 );
buf ( n211123 , n208166 );
xor ( n211124 , n211122 , n211123 );
buf ( n211125 , n211124 );
buf ( n211126 , n211125 );
buf ( n211127 , n210559 );
or ( n211128 , n211126 , n211127 );
buf ( n211129 , n211128 );
buf ( n211130 , n211129 );
and ( n211131 , n211111 , n211118 , n211130 );
buf ( n211132 , n211131 );
buf ( n211133 , n211132 );
buf ( n211134 , n210526 );
buf ( n211135 , n210532 );
or ( n211136 , n211134 , n211135 );
buf ( n211137 , n211136 );
buf ( n211138 , n211137 );
not ( n211139 , n211138 );
buf ( n211140 , n210515 );
buf ( n211141 , n210521 );
nor ( n211142 , n211140 , n211141 );
buf ( n211143 , n211142 );
buf ( n211144 , n211143 );
buf ( n211145 , n210510 );
buf ( n211146 , n210504 );
nand ( n211147 , n211145 , n211146 );
buf ( n211148 , n211147 );
buf ( n211149 , n211148 );
or ( n211150 , n211144 , n211149 );
buf ( n211151 , n210515 );
buf ( n211152 , n210521 );
nand ( n211153 , n211151 , n211152 );
buf ( n211154 , n211153 );
buf ( n211155 , n211154 );
nand ( n211156 , n211150 , n211155 );
buf ( n211157 , n211156 );
buf ( n211158 , n211157 );
not ( n211159 , n211158 );
or ( n211160 , n211139 , n211159 );
buf ( n211161 , n210526 );
buf ( n211162 , n210532 );
nand ( n211163 , n211161 , n211162 );
buf ( n211164 , n211163 );
buf ( n211165 , n211164 );
nand ( n211166 , n211160 , n211165 );
buf ( n211167 , n211166 );
buf ( n211168 , n211167 );
not ( n211169 , n211168 );
buf ( n211170 , n203502 );
buf ( n211171 , n27216 );
xor ( n211172 , n211170 , n211171 );
buf ( n211173 , n209437 );
xor ( n211174 , n211172 , n211173 );
buf ( n211175 , n211174 );
buf ( n211176 , n211175 );
buf ( n211177 , n210537 );
nor ( n211178 , n211176 , n211177 );
buf ( n211179 , n211178 );
buf ( n211180 , n211179 );
not ( n211181 , n211180 );
buf ( n211182 , n211181 );
buf ( n211183 , n211182 );
not ( n211184 , n211183 );
or ( n211185 , n211169 , n211184 );
buf ( n211186 , n210537 );
buf ( n211187 , n211175 );
nand ( n211188 , n211186 , n211187 );
buf ( n211189 , n211188 );
buf ( n211190 , n211189 );
nand ( n211191 , n211185 , n211190 );
buf ( n211192 , n211191 );
buf ( n211193 , n211192 );
not ( n211194 , n211193 );
buf ( n211195 , n210488 );
buf ( n211196 , n36198 );
buf ( n211197 , n203469 );
xor ( n211198 , n211196 , n211197 );
buf ( n211199 , n209170 );
and ( n211200 , n211198 , n211199 );
and ( n211201 , n211196 , n211197 );
or ( n211202 , n211200 , n211201 );
buf ( n211203 , n211202 );
buf ( n211204 , n211203 );
or ( n211205 , n211195 , n211204 );
buf ( n211206 , n211205 );
buf ( n211207 , n211206 );
not ( n211208 , n211207 );
buf ( n211209 , n203494 );
buf ( n211210 , n27501 );
xor ( n211211 , n211209 , n211210 );
buf ( n211212 , n41966 );
and ( n211213 , n211211 , n211212 );
and ( n211214 , n211209 , n211210 );
or ( n211215 , n211213 , n211214 );
buf ( n211216 , n211215 );
buf ( n211217 , n211216 );
xor ( n211218 , n211196 , n211197 );
xor ( n211219 , n211218 , n211199 );
buf ( n211220 , n211219 );
buf ( n211221 , n211220 );
nor ( n211222 , n211217 , n211221 );
buf ( n211223 , n211222 );
buf ( n211224 , n211223 );
xor ( n211225 , n211209 , n211210 );
xor ( n211226 , n211225 , n211212 );
buf ( n211227 , n211226 );
buf ( n211228 , n211227 );
buf ( n211229 , n210482 );
nand ( n211230 , n211228 , n211229 );
buf ( n211231 , n211230 );
buf ( n211232 , n211231 );
or ( n211233 , n211224 , n211232 );
buf ( n211234 , n211216 );
buf ( n211235 , n211220 );
nand ( n211236 , n211234 , n211235 );
buf ( n211237 , n211236 );
buf ( n211238 , n211237 );
nand ( n211239 , n211233 , n211238 );
buf ( n211240 , n211239 );
buf ( n211241 , n211240 );
not ( n211242 , n211241 );
or ( n211243 , n211208 , n211242 );
buf ( n211244 , n210488 );
buf ( n211245 , n211203 );
nand ( n211246 , n211244 , n211245 );
buf ( n211247 , n211246 );
buf ( n211248 , n211247 );
nand ( n211249 , n211243 , n211248 );
buf ( n211250 , n211249 );
buf ( n211251 , n211250 );
not ( n211252 , n211251 );
buf ( n211253 , n210499 );
buf ( n211254 , n210493 );
or ( n211255 , n211253 , n211254 );
buf ( n211256 , n211255 );
buf ( n211257 , n211256 );
not ( n211258 , n211257 );
or ( n211259 , n211252 , n211258 );
buf ( n211260 , n210499 );
buf ( n211261 , n210493 );
nand ( n211262 , n211260 , n211261 );
buf ( n211263 , n211262 );
buf ( n211264 , n211263 );
nand ( n211265 , n211259 , n211264 );
buf ( n211266 , n211265 );
buf ( n211267 , n211266 );
not ( n211268 , n211267 );
buf ( n211269 , n210471 );
buf ( n211270 , n210477 );
xor ( n211271 , n211269 , n211270 );
buf ( n211272 , n210466 );
buf ( n211273 , n203226 );
buf ( n211274 , n203232 );
xor ( n211275 , n211273 , n211274 );
buf ( n211276 , n41979 );
and ( n211277 , n211275 , n211276 );
and ( n211278 , n211273 , n211274 );
or ( n211279 , n211277 , n211278 );
buf ( n211280 , n211279 );
buf ( n211281 , n211280 );
xor ( n211282 , n211272 , n211281 );
xor ( n211283 , n211273 , n211274 );
xor ( n211284 , n211283 , n211276 );
buf ( n211285 , n211284 );
buf ( n211286 , n211285 );
buf ( n211287 , n210460 );
xor ( n211288 , n211286 , n211287 );
buf ( n211289 , n210449 );
buf ( n211290 , n210455 );
xor ( n211291 , n211289 , n211290 );
xor ( n211292 , n203269 , n203273 );
and ( n211293 , n211292 , n30498 );
and ( n211294 , n203269 , n203273 );
or ( n211295 , n211293 , n211294 );
buf ( n211296 , n211295 );
buf ( n211297 , n210444 );
xor ( n211298 , n211296 , n211297 );
buf ( n211299 , n29039 );
buf ( n211300 , n209316 );
xor ( n211301 , n211299 , n211300 );
buf ( n211302 , n211301 );
buf ( n211303 , n211302 );
not ( n211304 , n211303 );
buf ( n211305 , n211304 );
buf ( n211306 , n211305 );
buf ( n211307 , n203282 );
not ( n211308 , n211307 );
buf ( n211309 , n211308 );
buf ( n211310 , n211309 );
and ( n211311 , n211306 , n211310 );
buf ( n211312 , n209348 );
and ( n211313 , n863 , n895 );
buf ( n211314 , n211313 );
buf ( n211315 , n211314 );
nand ( n211316 , n211312 , n211315 );
buf ( n211317 , n211316 );
buf ( n211318 , n211317 );
nor ( n211319 , n211311 , n211318 );
buf ( n211320 , n211319 );
buf ( n211321 , n211320 );
buf ( n211322 , n211305 );
buf ( n211323 , n211309 );
nor ( n211324 , n211322 , n211323 );
buf ( n211325 , n211324 );
buf ( n211326 , n211325 );
nor ( n211327 , n211321 , n211326 );
buf ( n211328 , n211327 );
buf ( n211329 , n211328 );
xor ( n211330 , n203269 , n203273 );
xor ( n211331 , n211330 , n30498 );
buf ( n211332 , n211331 );
and ( n211333 , n211299 , n211300 );
buf ( n211334 , n211333 );
buf ( n211335 , n211334 );
nor ( n211336 , n211332 , n211335 );
buf ( n211337 , n211336 );
buf ( n211338 , n211337 );
or ( n211339 , n211329 , n211338 );
buf ( n211340 , n211331 );
buf ( n211341 , n211334 );
nand ( n211342 , n211340 , n211341 );
buf ( n211343 , n211342 );
buf ( n211344 , n211343 );
nand ( n211345 , n211339 , n211344 );
buf ( n211346 , n211345 );
buf ( n211347 , n211346 );
and ( n211348 , n211298 , n211347 );
and ( n211349 , n211296 , n211297 );
or ( n211350 , n211348 , n211349 );
buf ( n211351 , n211350 );
buf ( n211352 , n211351 );
and ( n211353 , n211291 , n211352 );
and ( n211354 , n211289 , n211290 );
or ( n211355 , n211353 , n211354 );
buf ( n211356 , n211355 );
buf ( n211357 , n211356 );
and ( n211358 , n211288 , n211357 );
and ( n211359 , n211286 , n211287 );
or ( n211360 , n211358 , n211359 );
buf ( n211361 , n211360 );
buf ( n211362 , n211361 );
and ( n211363 , n211282 , n211362 );
and ( n211364 , n211272 , n211281 );
or ( n211365 , n211363 , n211364 );
buf ( n211366 , n211365 );
buf ( n211367 , n211366 );
and ( n211368 , n211271 , n211367 );
and ( n211369 , n211269 , n211270 );
or ( n211370 , n211368 , n211369 );
buf ( n211371 , n211370 );
buf ( n211372 , n211371 );
buf ( n211373 , n211256 );
buf ( n211374 , n211223 );
buf ( n211375 , n211227 );
buf ( n211376 , n210482 );
nor ( n211377 , n211375 , n211376 );
buf ( n211378 , n211377 );
buf ( n211379 , n211378 );
nor ( n211380 , n211374 , n211379 );
buf ( n211381 , n211380 );
buf ( n211382 , n211381 );
buf ( n211383 , n211206 );
and ( n211384 , n211382 , n211383 );
buf ( n211385 , n211384 );
buf ( n211386 , n211385 );
nand ( n211387 , n211372 , n211373 , n211386 );
buf ( n211388 , n211387 );
buf ( n211389 , n211388 );
nand ( n211390 , n211268 , n211389 );
buf ( n211391 , n211390 );
buf ( n211392 , n211391 );
buf ( n211393 , n211179 );
buf ( n211394 , n211137 );
not ( n211395 , n211394 );
buf ( n211396 , n211395 );
buf ( n211397 , n211396 );
nor ( n211398 , n211393 , n211397 );
buf ( n211399 , n211398 );
buf ( n211400 , n211399 );
buf ( n211401 , n211143 );
not ( n211402 , n211401 );
buf ( n211403 , n211402 );
buf ( n211404 , n211403 );
buf ( n211405 , n210510 );
buf ( n211406 , n210504 );
or ( n211407 , n211405 , n211406 );
buf ( n211408 , n211407 );
buf ( n211409 , n211408 );
nand ( n211410 , n211392 , n211400 , n211404 , n211409 );
buf ( n211411 , n211410 );
buf ( n211412 , n211411 );
nand ( n211413 , n211194 , n211412 );
buf ( n211414 , n211413 );
buf ( n211415 , n211414 );
buf ( n211416 , n210543 );
not ( n211417 , n202938 );
buf ( n211418 , n202955 );
not ( n211419 , n211418 );
or ( n211420 , n211417 , n211419 );
or ( n211421 , n211418 , n202938 );
not ( n211422 , n41565 );
not ( n211423 , n211422 );
nand ( n211424 , n211421 , n211423 );
nand ( n211425 , n211420 , n211424 );
buf ( n211426 , n211425 );
or ( n211427 , n211416 , n211426 );
buf ( n211428 , n211427 );
buf ( n211429 , n211428 );
not ( n211430 , n211429 );
xor ( n211431 , n211170 , n211171 );
and ( n211432 , n211431 , n211173 );
and ( n211433 , n211170 , n211171 );
or ( n211434 , n211432 , n211433 );
buf ( n211435 , n211434 );
buf ( n211436 , n211435 );
buf ( n211437 , n202972 );
buf ( n211438 , n27087 );
xor ( n211439 , n211437 , n211438 );
buf ( n211440 , n41609 );
xor ( n211441 , n211439 , n211440 );
buf ( n211442 , n211441 );
buf ( n211443 , n211442 );
nor ( n211444 , n211436 , n211443 );
buf ( n211445 , n211444 );
buf ( n211446 , n211445 );
not ( n211447 , n211446 );
xor ( n211448 , n211418 , n202938 );
not ( n211449 , n35709 );
xor ( n211450 , n211449 , n202982 );
buf ( n211451 , n41700 );
and ( n211452 , n211450 , n211451 );
and ( n211453 , n211449 , n202982 );
or ( n211454 , n211452 , n211453 );
or ( n211455 , n211448 , n211454 , n211423 );
not ( n211456 , n211454 );
nand ( n211457 , n211456 , n211423 , n211448 );
nand ( n211458 , n211455 , n211457 );
not ( n211459 , n211458 );
buf ( n211460 , n211459 );
xor ( n211461 , n211437 , n211438 );
and ( n211462 , n211461 , n211440 );
and ( n211463 , n211437 , n211438 );
or ( n211464 , n211462 , n211463 );
buf ( n211465 , n211464 );
buf ( n211466 , n211465 );
xor ( n211467 , n211449 , n202982 );
xor ( n211468 , n211467 , n211451 );
buf ( n211469 , n211468 );
nor ( n211470 , n211466 , n211469 );
buf ( n211471 , n211470 );
buf ( n211472 , n211471 );
not ( n211473 , n211472 );
buf ( n211474 , n211473 );
buf ( n211475 , n211474 );
nand ( n211476 , n211447 , n211460 , n211475 );
buf ( n211477 , n211476 );
buf ( n211478 , n211477 );
nor ( n211479 , n211430 , n211478 );
buf ( n211480 , n211479 );
buf ( n211481 , n211480 );
and ( n211482 , n211133 , n211415 , n211481 );
buf ( n211483 , n211482 );
buf ( n211484 , n211483 );
buf ( n211485 , n211132 );
buf ( n211486 , n211428 );
not ( n211487 , n211486 );
not ( n211488 , n211471 );
buf ( n211489 , n211435 );
buf ( n211490 , n211442 );
nand ( n211491 , n211489 , n211490 );
buf ( n211492 , n211491 );
not ( n211493 , n211492 );
and ( n211494 , n211488 , n211493 );
buf ( n211495 , n211465 );
buf ( n211496 , n211468 );
and ( n211497 , n211495 , n211496 );
buf ( n211498 , n211497 );
nor ( n211499 , n211494 , n211498 );
buf ( n211500 , n211499 );
buf ( n211501 , n211458 );
or ( n211502 , n211500 , n211501 );
xor ( n211503 , n211423 , n211448 );
buf ( n211504 , n211503 );
buf ( n211505 , n211454 );
nand ( n211506 , n211504 , n211505 );
buf ( n211507 , n211506 );
buf ( n211508 , n211507 );
nand ( n211509 , n211502 , n211508 );
buf ( n211510 , n211509 );
buf ( n211511 , n211510 );
not ( n211512 , n211511 );
or ( n211513 , n211487 , n211512 );
buf ( n211514 , n210543 );
buf ( n211515 , n211425 );
nand ( n211516 , n211514 , n211515 );
buf ( n211517 , n211516 );
buf ( n211518 , n211517 );
nand ( n211519 , n211513 , n211518 );
buf ( n211520 , n211519 );
buf ( n211521 , n211520 );
nand ( n211522 , n211485 , n211521 );
buf ( n211523 , n211522 );
buf ( n211524 , n211117 );
not ( n211525 , n211524 );
buf ( n211526 , n211099 );
buf ( n211527 , n211103 );
buf ( n211528 , n210548 );
nand ( n211529 , n211527 , n211528 );
buf ( n211530 , n211529 );
buf ( n211531 , n211530 );
or ( n211532 , n211526 , n211531 );
buf ( n211533 , n211096 );
buf ( n211534 , n211087 );
nand ( n211535 , n211533 , n211534 );
buf ( n211536 , n211535 );
buf ( n211537 , n211536 );
nand ( n211538 , n211532 , n211537 );
buf ( n211539 , n211538 );
buf ( n211540 , n211539 );
not ( n211541 , n211540 );
or ( n211542 , n211525 , n211541 );
nand ( n211543 , n210554 , n211116 );
buf ( n211544 , n211543 );
nand ( n211545 , n211542 , n211544 );
buf ( n211546 , n211545 );
buf ( n211547 , n211546 );
buf ( n211548 , n211129 );
nand ( n211549 , n211547 , n211548 );
buf ( n211550 , n211549 );
buf ( n211551 , n210559 );
buf ( n211552 , n211125 );
nand ( n211553 , n211551 , n211552 );
buf ( n211554 , n211553 );
nand ( n211555 , n211523 , n211550 , n211554 );
buf ( n211556 , n211555 );
or ( n211557 , n211484 , n211556 );
buf ( n211558 , n210589 );
not ( n211559 , n211558 );
xor ( n211560 , n35539 , n41165 );
not ( n211561 , n36276 );
and ( n211562 , n211560 , n211561 );
and ( n211563 , n35539 , n41165 );
or ( n211564 , n211562 , n211563 );
not ( n211565 , n211564 );
buf ( n211566 , n211565 );
nand ( n211567 , n211559 , n211566 );
buf ( n211568 , n211567 );
buf ( n211569 , n211568 );
xor ( n211570 , n35539 , n41165 );
not ( n211571 , n36276 );
xor ( n211572 , n211570 , n211571 );
buf ( n211573 , n211572 );
buf ( n211574 , n210571 );
or ( n211575 , n211573 , n211574 );
buf ( n211576 , n211575 );
buf ( n211577 , n211576 );
not ( n211578 , n211577 );
buf ( n211579 , n210566 );
buf ( n211580 , n210582 );
nor ( n211581 , n211579 , n211580 );
buf ( n211582 , n211581 );
buf ( n211583 , n211582 );
not ( n211584 , n211583 );
buf ( n211585 , n211584 );
buf ( n211586 , n211585 );
buf ( n211587 , n210577 );
xor ( n211588 , n211119 , n211121 );
and ( n211589 , n211588 , n211123 );
and ( n211590 , n211119 , n211121 );
or ( n211591 , n211589 , n211590 );
buf ( n211592 , n211591 );
buf ( n211593 , n211592 );
or ( n211594 , n211587 , n211593 );
buf ( n211595 , n211594 );
buf ( n211596 , n211595 );
nand ( n211597 , n211586 , n211596 );
buf ( n211598 , n211597 );
buf ( n211599 , n211598 );
nor ( n211600 , n211578 , n211599 );
buf ( n211601 , n211600 );
buf ( n211602 , n211601 );
and ( n211603 , n211569 , n211602 );
buf ( n211604 , n211603 );
buf ( n211605 , n211604 );
nand ( n211606 , n211557 , n211605 );
buf ( n211607 , n211606 );
buf ( n211608 , n211607 );
not ( n211609 , n211608 );
buf ( n211610 , n211576 );
not ( n211611 , n211610 );
buf ( n211612 , n211582 );
buf ( n211613 , n210577 );
buf ( n211614 , n211592 );
nand ( n211615 , n211613 , n211614 );
buf ( n211616 , n211615 );
buf ( n211617 , n211616 );
or ( n211618 , n211612 , n211617 );
buf ( n211619 , n210582 );
buf ( n211620 , n210566 );
nand ( n211621 , n211619 , n211620 );
buf ( n211622 , n211621 );
buf ( n211623 , n211622 );
nand ( n211624 , n211618 , n211623 );
buf ( n211625 , n211624 );
buf ( n211626 , n211625 );
not ( n211627 , n211626 );
or ( n211628 , n211611 , n211627 );
buf ( n211629 , n211572 );
buf ( n211630 , n210571 );
nand ( n211631 , n211629 , n211630 );
buf ( n211632 , n211631 );
buf ( n211633 , n211632 );
nand ( n211634 , n211628 , n211633 );
buf ( n211635 , n211634 );
buf ( n211636 , n211635 );
not ( n211637 , n211636 );
buf ( n211638 , n211568 );
not ( n211639 , n211638 );
or ( n211640 , n211637 , n211639 );
buf ( n211641 , n211565 );
not ( n211642 , n211641 );
buf ( n211643 , n210589 );
nand ( n211644 , n211642 , n211643 );
buf ( n211645 , n211644 );
buf ( n211646 , n211645 );
nand ( n211647 , n211640 , n211646 );
buf ( n211648 , n211647 );
buf ( n211649 , n211648 );
not ( n211650 , n211649 );
buf ( n211651 , n211650 );
buf ( n211652 , n211651 );
not ( n211653 , n211652 );
or ( n211654 , n211609 , n211653 );
buf ( n211655 , n210619 );
not ( n211656 , n211655 );
buf ( n211657 , n210627 );
not ( n211658 , n211657 );
buf ( n211659 , n211658 );
buf ( n211660 , n211659 );
nand ( n211661 , n211656 , n211660 );
buf ( n211662 , n211661 );
buf ( n211663 , n211662 );
buf ( n211664 , n210614 );
buf ( n211665 , n202557 );
buf ( n211666 , n211665 );
buf ( n211667 , n211666 );
buf ( n211668 , n36304 );
buf ( n211669 , n211668 );
xor ( n211670 , n211667 , n211669 );
buf ( n211671 , n208044 );
and ( n211672 , n211670 , n211671 );
and ( n211673 , n211667 , n211669 );
or ( n211674 , n211672 , n211673 );
buf ( n211675 , n211674 );
buf ( n211676 , n211675 );
or ( n211677 , n211664 , n211676 );
buf ( n211678 , n211677 );
buf ( n211679 , n211678 );
nand ( n211680 , n211663 , n211679 );
buf ( n211681 , n211680 );
buf ( n211682 , n211681 );
buf ( n211683 , n210606 );
xor ( n211684 , n211667 , n211669 );
xor ( n211685 , n211684 , n211671 );
buf ( n211686 , n211685 );
buf ( n211687 , n211686 );
nor ( n211688 , n211683 , n211687 );
buf ( n211689 , n211688 );
buf ( n211690 , n211689 );
not ( n211691 , n211690 );
buf ( n211692 , n210601 );
buf ( n211693 , n210594 );
or ( n211694 , n211692 , n211693 );
buf ( n211695 , n211694 );
buf ( n211696 , n211695 );
nand ( n211697 , n211691 , n211696 );
buf ( n211698 , n211697 );
buf ( n211699 , n211698 );
nor ( n211700 , n211682 , n211699 );
buf ( n211701 , n211700 );
buf ( n211702 , n211701 );
nand ( n211703 , n211654 , n211702 );
buf ( n211704 , n211703 );
buf ( n211705 , n211704 );
buf ( n211706 , n211681 );
not ( n211707 , n211706 );
buf ( n211708 , n211707 );
buf ( n211709 , n211708 );
buf ( n211710 , n211689 );
buf ( n211711 , n210594 );
buf ( n211712 , n210601 );
nand ( n211713 , n211711 , n211712 );
buf ( n211714 , n211713 );
buf ( n211715 , n211714 );
or ( n211716 , n211710 , n211715 );
buf ( n211717 , n210606 );
buf ( n211718 , n211686 );
nand ( n211719 , n211717 , n211718 );
buf ( n211720 , n211719 );
buf ( n211721 , n211720 );
nand ( n211722 , n211716 , n211721 );
buf ( n211723 , n211722 );
buf ( n211724 , n211723 );
and ( n211725 , n211709 , n211724 );
buf ( n211726 , n211675 );
buf ( n211727 , n210614 );
and ( n211728 , n211726 , n211727 );
buf ( n211729 , n211728 );
buf ( n211730 , n211729 );
not ( n211731 , n211730 );
buf ( n211732 , n211662 );
not ( n211733 , n211732 );
or ( n211734 , n211731 , n211733 );
buf ( n211735 , n211659 );
not ( n211736 , n211735 );
buf ( n211737 , n210619 );
nand ( n211738 , n211736 , n211737 );
buf ( n211739 , n211738 );
buf ( n211740 , n211739 );
nand ( n211741 , n211734 , n211740 );
buf ( n211742 , n211741 );
buf ( n211743 , n211742 );
nor ( n211744 , n211725 , n211743 );
buf ( n211745 , n211744 );
buf ( n211746 , n211745 );
nand ( n211747 , n211705 , n211746 );
buf ( n211748 , n211747 );
buf ( n211749 , n211748 );
buf ( n211750 , n210651 );
buf ( n211751 , n201310 );
buf ( n211752 , n201305 );
buf ( n211753 , n211752 );
xor ( n211754 , n211751 , n211753 );
buf ( n211755 , n40410 );
and ( n211756 , n211754 , n211755 );
and ( n211757 , n211751 , n211753 );
or ( n211758 , n211756 , n211757 );
buf ( n211759 , n211758 );
buf ( n211760 , n211759 );
nor ( n211761 , n211750 , n211760 );
buf ( n211762 , n211761 );
buf ( n211763 , n211762 );
buf ( n211764 , n210656 );
xor ( n211765 , n200908 , n33637 );
xor ( n211766 , n211765 , n40397 );
buf ( n211767 , n211766 );
nor ( n211768 , n211764 , n211767 );
buf ( n211769 , n211768 );
buf ( n211770 , n211769 );
nor ( n211771 , n211763 , n211770 );
buf ( n211772 , n211771 );
buf ( n211773 , n211772 );
buf ( n211774 , n210662 );
not ( n211775 , n211774 );
xor ( n211776 , n200908 , n33637 );
and ( n211777 , n211776 , n40397 );
and ( n211778 , n200908 , n33637 );
nor ( n211779 , n211777 , n211778 );
buf ( n211780 , n211779 );
nand ( n211781 , n211775 , n211780 );
buf ( n211782 , n211781 );
buf ( n211783 , n211782 );
xor ( n211784 , n210962 , n210963 );
xor ( n211785 , n211784 , n210965 );
buf ( n211786 , n211785 );
buf ( n211787 , n211786 );
buf ( n211788 , n210667 );
or ( n211789 , n211787 , n211788 );
buf ( n211790 , n211789 );
buf ( n211791 , n211790 );
and ( n211792 , n211773 , n211783 , n211791 );
buf ( n211793 , n211792 );
buf ( n211794 , n211793 );
not ( n211795 , n211794 );
buf ( n211796 , n211795 );
buf ( n211797 , n211796 );
buf ( n211798 , n201295 );
buf ( n211799 , n23048 );
xor ( n211800 , n211798 , n211799 );
buf ( n211801 , n207946 );
and ( n211802 , n211800 , n211801 );
and ( n211803 , n211798 , n211799 );
or ( n211804 , n211802 , n211803 );
buf ( n211805 , n211804 );
buf ( n211806 , n211805 );
xor ( n211807 , n211751 , n211753 );
xor ( n211808 , n211807 , n211755 );
buf ( n211809 , n211808 );
buf ( n211810 , n211809 );
or ( n211811 , n211806 , n211810 );
buf ( n211812 , n211811 );
buf ( n211813 , n211812 );
xor ( n211814 , n211798 , n211799 );
xor ( n211815 , n211814 , n211801 );
buf ( n211816 , n211815 );
buf ( n211817 , n211816 );
buf ( n211818 , n210644 );
or ( n211819 , n211817 , n211818 );
buf ( n211820 , n211819 );
buf ( n211821 , n211820 );
and ( n211822 , n211813 , n211821 );
buf ( n211823 , n211822 );
buf ( n211824 , n211823 );
buf ( n211825 , n24888 );
buf ( n211826 , n201288 );
xor ( n211827 , n211825 , n211826 );
buf ( n211828 , n40625 );
xor ( n211829 , n211827 , n211828 );
buf ( n211830 , n211829 );
buf ( n211831 , n211830 );
buf ( n211832 , n210632 );
nor ( n211833 , n211831 , n211832 );
buf ( n211834 , n211833 );
buf ( n211835 , n211834 );
xor ( n211836 , n211825 , n211826 );
and ( n211837 , n211836 , n211828 );
and ( n211838 , n211825 , n211826 );
or ( n211839 , n211837 , n211838 );
buf ( n211840 , n211839 );
buf ( n211841 , n211840 );
buf ( n211842 , n210639 );
nor ( n211843 , n211841 , n211842 );
buf ( n211844 , n211843 );
buf ( n211845 , n211844 );
nor ( n211846 , n211835 , n211845 );
buf ( n211847 , n211846 );
buf ( n211848 , n211847 );
nand ( n211849 , n211824 , n211848 );
buf ( n211850 , n211849 );
buf ( n211851 , n211850 );
nor ( n211852 , n211797 , n211851 );
buf ( n211853 , n211852 );
buf ( n211854 , n211853 );
nand ( n211855 , n211080 , n211749 , n211854 );
buf ( n211856 , n211855 );
buf ( n211857 , n211856 );
buf ( n211858 , n211079 );
buf ( n211859 , n211823 );
not ( n211860 , n211859 );
buf ( n211861 , n211830 );
buf ( n211862 , n210632 );
nand ( n211863 , n211861 , n211862 );
buf ( n211864 , n211863 );
buf ( n211865 , n211864 );
buf ( n211866 , n211844 );
or ( n211867 , n211865 , n211866 );
buf ( n211868 , n211840 );
buf ( n211869 , n210639 );
nand ( n211870 , n211868 , n211869 );
buf ( n211871 , n211870 );
buf ( n211872 , n211871 );
nand ( n211873 , n211867 , n211872 );
buf ( n211874 , n211873 );
buf ( n211875 , n211874 );
not ( n211876 , n211875 );
or ( n211877 , n211860 , n211876 );
buf ( n211878 , n210644 );
buf ( n211879 , n211816 );
and ( n211880 , n211878 , n211879 );
buf ( n211881 , n211880 );
buf ( n211882 , n211881 );
not ( n211883 , n211882 );
buf ( n211884 , n211812 );
not ( n211885 , n211884 );
or ( n211886 , n211883 , n211885 );
buf ( n211887 , n211805 );
buf ( n211888 , n211809 );
nand ( n211889 , n211887 , n211888 );
buf ( n211890 , n211889 );
buf ( n211891 , n211890 );
nand ( n211892 , n211886 , n211891 );
buf ( n211893 , n211892 );
buf ( n211894 , n211893 );
not ( n211895 , n211894 );
buf ( n211896 , n211895 );
buf ( n211897 , n211896 );
nand ( n211898 , n211877 , n211897 );
buf ( n211899 , n211898 );
buf ( n211900 , n211899 );
buf ( n211901 , n211793 );
nand ( n211902 , n211900 , n211901 );
buf ( n211903 , n211902 );
buf ( n211904 , n211903 );
buf ( n211905 , n211782 );
not ( n211906 , n211905 );
buf ( n211907 , n211769 );
buf ( n211908 , n210651 );
buf ( n211909 , n211759 );
nand ( n211910 , n211908 , n211909 );
buf ( n211911 , n211910 );
buf ( n211912 , n211911 );
or ( n211913 , n211907 , n211912 );
buf ( n211914 , n210656 );
buf ( n211915 , n211766 );
nand ( n211916 , n211914 , n211915 );
buf ( n211917 , n211916 );
buf ( n211918 , n211917 );
nand ( n211919 , n211913 , n211918 );
buf ( n211920 , n211919 );
buf ( n211921 , n211920 );
not ( n211922 , n211921 );
or ( n211923 , n211906 , n211922 );
buf ( n211924 , n211779 );
not ( n211925 , n211924 );
buf ( n211926 , n210662 );
nand ( n211927 , n211925 , n211926 );
buf ( n211928 , n211927 );
buf ( n211929 , n211928 );
nand ( n211930 , n211923 , n211929 );
buf ( n211931 , n211930 );
buf ( n211932 , n211931 );
buf ( n211933 , n211790 );
nand ( n211934 , n211932 , n211933 );
buf ( n211935 , n211934 );
buf ( n211936 , n211935 );
buf ( n211937 , n210667 );
buf ( n211938 , n211786 );
nand ( n211939 , n211937 , n211938 );
buf ( n211940 , n211939 );
buf ( n211941 , n211940 );
nand ( n211942 , n211904 , n211936 , n211941 );
buf ( n211943 , n211942 );
buf ( n211944 , n211943 );
nand ( n211945 , n211858 , n211944 );
buf ( n211946 , n211945 );
buf ( n211947 , n211946 );
nand ( n211948 , n211065 , n211857 , n211947 );
buf ( n211949 , n211948 );
buf ( n211950 , n211949 );
not ( n211951 , n211950 );
or ( n211952 , n210893 , n211951 );
buf ( n211953 , n210816 );
not ( n211954 , n211953 );
buf ( n211955 , n210806 );
not ( n211956 , n211955 );
buf ( n211957 , n210724 );
buf ( n211958 , n210827 );
nand ( n211959 , n211957 , n211958 );
buf ( n211960 , n211959 );
buf ( n211961 , n211960 );
buf ( n211962 , n210840 );
or ( n211963 , n211961 , n211962 );
buf ( n211964 , n210833 );
buf ( n211965 , n210839 );
nand ( n211966 , n211964 , n211965 );
buf ( n211967 , n211966 );
buf ( n211968 , n211967 );
nand ( n211969 , n211963 , n211968 );
buf ( n211970 , n211969 );
buf ( n211971 , n211970 );
not ( n211972 , n211971 );
or ( n211973 , n211956 , n211972 );
buf ( n211974 , n210803 );
not ( n211975 , n211974 );
buf ( n211976 , n210797 );
nand ( n211977 , n211975 , n211976 );
buf ( n211978 , n211977 );
buf ( n211979 , n211978 );
nand ( n211980 , n211973 , n211979 );
buf ( n211981 , n211980 );
buf ( n211982 , n211981 );
not ( n211983 , n211982 );
or ( n211984 , n211954 , n211983 );
buf ( n211985 , n210812 );
buf ( n211986 , n210741 );
nand ( n211987 , n211985 , n211986 );
buf ( n211988 , n211987 );
buf ( n211989 , n211988 );
nand ( n211990 , n211984 , n211989 );
buf ( n211991 , n211990 );
buf ( n211992 , n210888 );
not ( n211993 , n211992 );
buf ( n211994 , n211993 );
and ( n211995 , n211991 , n211994 );
buf ( n211996 , n210882 );
not ( n211997 , n211996 );
buf ( n211998 , n211997 );
buf ( n211999 , n211998 );
not ( n212000 , n211999 );
buf ( n212001 , n210869 );
buf ( n212002 , n210746 );
buf ( n212003 , n210856 );
nand ( n212004 , n212002 , n212003 );
buf ( n212005 , n212004 );
buf ( n212006 , n212005 );
or ( n212007 , n212001 , n212006 );
buf ( n212008 , n210685 );
buf ( n212009 , n210866 );
nand ( n212010 , n212008 , n212009 );
buf ( n212011 , n212010 );
buf ( n212012 , n212011 );
nand ( n212013 , n212007 , n212012 );
buf ( n212014 , n212013 );
buf ( n212015 , n212014 );
not ( n212016 , n212015 );
or ( n212017 , n212000 , n212016 );
buf ( n212018 , n210690 );
buf ( n212019 , n210421 );
nand ( n212020 , n212018 , n212019 );
buf ( n212021 , n212020 );
buf ( n212022 , n212021 );
nand ( n212023 , n212017 , n212022 );
buf ( n212024 , n212023 );
buf ( n212025 , n210877 );
not ( n212026 , n212025 );
buf ( n212027 , n212026 );
and ( n212028 , n212024 , n212027 );
buf ( n212029 , n210730 );
buf ( n212030 , n210426 );
and ( n212031 , n212029 , n212030 );
buf ( n212032 , n212031 );
nor ( n212033 , n211995 , n212028 , n212032 );
buf ( n212034 , n212033 );
nand ( n212035 , n211952 , n212034 );
buf ( n212036 , n212035 );
buf ( n212037 , n212036 );
buf ( n212038 , n210410 );
buf ( n212039 , n210735 );
or ( n212040 , n212038 , n212039 );
buf ( n212041 , n212040 );
buf ( n212042 , n212041 );
nand ( n212043 , n212037 , n212042 );
buf ( n212044 , n212043 );
buf ( n212045 , n210399 );
buf ( n212046 , n210415 );
nor ( n212047 , n212045 , n212046 );
buf ( n212048 , n212047 );
not ( n212049 , n212048 );
buf ( n212050 , n210404 );
buf ( n212051 , n210433 );
or ( n212052 , n212050 , n212051 );
buf ( n212053 , n212052 );
buf ( n212054 , n210438 );
buf ( n212055 , n210756 );
or ( n212056 , n212054 , n212055 );
buf ( n212057 , n212056 );
nand ( n212058 , n212049 , n212053 , n212057 );
or ( n212059 , n212044 , n212058 );
buf ( n212060 , n212053 );
not ( n212061 , n212060 );
buf ( n212062 , n210410 );
buf ( n212063 , n210735 );
nand ( n212064 , n212062 , n212063 );
buf ( n212065 , n212064 );
or ( n212066 , n212048 , n212065 );
buf ( n212067 , n210399 );
buf ( n212068 , n210415 );
nand ( n212069 , n212067 , n212068 );
buf ( n212070 , n212069 );
nand ( n212071 , n212066 , n212070 );
buf ( n212072 , n212071 );
not ( n212073 , n212072 );
or ( n212074 , n212061 , n212073 );
buf ( n212075 , n210404 );
buf ( n212076 , n210433 );
nand ( n212077 , n212075 , n212076 );
buf ( n212078 , n212077 );
buf ( n212079 , n212078 );
nand ( n212080 , n212074 , n212079 );
buf ( n212081 , n212080 );
and ( n212082 , n212081 , n212057 );
buf ( n212083 , n210438 );
buf ( n212084 , n210756 );
and ( n212085 , n212083 , n212084 );
buf ( n212086 , n212085 );
nor ( n212087 , n212082 , n212086 );
nand ( n212088 , n212059 , n212087 );
buf ( n212089 , n212088 );
not ( n212090 , n212089 );
or ( n212091 , n210791 , n212090 );
buf ( n212092 , n210758 );
buf ( n212093 , n210750 );
nand ( n212094 , n212092 , n212093 );
buf ( n212095 , n212094 );
buf ( n212096 , n212095 );
not ( n212097 , n212096 );
buf ( n212098 , n210786 );
not ( n212099 , n212098 );
and ( n212100 , n212097 , n212099 );
buf ( n212101 , n210752 );
buf ( n212102 , n210762 );
and ( n212103 , n212101 , n212102 );
buf ( n212104 , n212103 );
buf ( n212105 , n212104 );
nor ( n212106 , n212100 , n212105 );
buf ( n212107 , n212106 );
buf ( n212108 , n212107 );
nand ( n212109 , n212091 , n212108 );
buf ( n212110 , n212109 );
buf ( n212111 , n212110 );
xor ( n212112 , n210775 , n210776 );
xor ( n212113 , n212112 , n212111 );
buf ( n212114 , n212113 );
xor ( n212115 , n210775 , n210776 );
and ( n212116 , n212115 , n212111 );
and ( n212117 , n210775 , n210776 );
or ( n212118 , n212116 , n212117 );
buf ( n212119 , n212118 );
buf ( n212120 , n212086 );
not ( n212121 , n212120 );
buf ( n212122 , n212057 );
nand ( n212123 , n212121 , n212122 );
buf ( n212124 , n212123 );
buf ( n212125 , n212124 );
buf ( n212126 , n212124 );
not ( n212127 , n212126 );
buf ( n212128 , n212127 );
buf ( n212129 , n212128 );
buf ( n212130 , n212053 );
not ( n212131 , n212130 );
or ( n212132 , n212044 , n212048 );
not ( n212133 , n212071 );
nand ( n212134 , n212132 , n212133 );
buf ( n212135 , n212134 );
not ( n212136 , n212135 );
or ( n212137 , n212131 , n212136 );
buf ( n212138 , n212078 );
nand ( n212139 , n212137 , n212138 );
buf ( n212140 , n212139 );
buf ( n212141 , n212140 );
and ( n212142 , n212141 , n212129 );
not ( n212143 , n212141 );
and ( n212144 , n212143 , n212125 );
nor ( n212145 , n212142 , n212144 );
buf ( n212146 , n212145 );
buf ( n212147 , n210939 );
buf ( n212148 , n210914 );
not ( n212149 , n212148 );
buf ( n212150 , n211076 );
not ( n212151 , n212150 );
buf ( n212152 , n211796 );
buf ( n212153 , n211850 );
not ( n212154 , n212153 );
buf ( n212155 , n211748 );
nand ( n212156 , n212154 , n212155 );
buf ( n212157 , n212156 );
buf ( n212158 , n212157 );
or ( n212159 , n212152 , n212158 );
buf ( n212160 , n211943 );
not ( n212161 , n212160 );
buf ( n212162 , n212161 );
buf ( n212163 , n212162 );
nand ( n212164 , n212159 , n212163 );
buf ( n212165 , n212164 );
buf ( n212166 , n212165 );
not ( n212167 , n212166 );
or ( n212168 , n212151 , n212167 );
buf ( n212169 , n211011 );
not ( n212170 , n212169 );
buf ( n212171 , n212170 );
buf ( n212172 , n212171 );
nand ( n212173 , n212168 , n212172 );
buf ( n212174 , n212173 );
buf ( n212175 , n212174 );
not ( n212176 , n212175 );
or ( n212177 , n212149 , n212176 );
buf ( n212178 , n211035 );
not ( n212179 , n212178 );
buf ( n212180 , n212179 );
buf ( n212181 , n212180 );
nand ( n212182 , n212177 , n212181 );
buf ( n212183 , n212182 );
buf ( n212184 , n212183 );
buf ( n212185 , n211043 );
not ( n212186 , n212147 );
not ( n212187 , n212184 );
or ( n212188 , n212186 , n212187 );
nand ( n212189 , n212188 , n212185 );
buf ( n212190 , n212189 );
buf ( n212191 , n210995 );
not ( n212192 , n211073 );
and ( n212193 , n212165 , n211068 );
not ( n212194 , n212193 );
or ( n212195 , n212192 , n212194 );
buf ( n212196 , n210985 );
not ( n212197 , n212196 );
buf ( n212198 , n212197 );
nand ( n212199 , n212195 , n212198 );
buf ( n212200 , n212199 );
buf ( n212201 , n210999 );
not ( n212202 , n212191 );
not ( n212203 , n212200 );
or ( n212204 , n212202 , n212203 );
nand ( n212205 , n212204 , n212201 );
buf ( n212206 , n212205 );
buf ( n212207 , n210859 );
not ( n212208 , n212207 );
buf ( n212209 , n212208 );
buf ( n212210 , n212209 );
buf ( n212211 , n210846 );
not ( n212212 , n212211 );
buf ( n212213 , n212212 );
buf ( n212214 , n212213 );
not ( n212215 , n212214 );
buf ( n212216 , n211949 );
not ( n212217 , n212216 );
or ( n212218 , n212215 , n212217 );
buf ( n212219 , n211991 );
not ( n212220 , n212219 );
buf ( n212221 , n212220 );
buf ( n212222 , n212221 );
nand ( n212223 , n212218 , n212222 );
buf ( n212224 , n212223 );
buf ( n212225 , n212224 );
buf ( n212226 , n212005 );
not ( n212227 , n212210 );
not ( n212228 , n212225 );
or ( n212229 , n212227 , n212228 );
nand ( n212230 , n212229 , n212226 );
buf ( n212231 , n212230 );
buf ( n212232 , n210911 );
not ( n212233 , n212232 );
buf ( n212234 , n212233 );
buf ( n212235 , n212234 );
buf ( n212236 , n212174 );
buf ( n212237 , n211020 );
not ( n212238 , n212237 );
buf ( n212239 , n212238 );
buf ( n212240 , n212239 );
not ( n212241 , n212235 );
not ( n212242 , n212236 );
or ( n212243 , n212241 , n212242 );
nand ( n212244 , n212243 , n212240 );
buf ( n212245 , n212244 );
buf ( n212246 , n210872 );
buf ( n212247 , n212224 );
buf ( n212248 , n212014 );
not ( n212249 , n212248 );
buf ( n212250 , n212249 );
buf ( n212251 , n212250 );
not ( n212252 , n212246 );
not ( n212253 , n212247 );
or ( n212254 , n212252 , n212253 );
nand ( n212255 , n212254 , n212251 );
buf ( n212256 , n212255 );
buf ( n212257 , n210806 );
buf ( n212258 , n210843 );
not ( n212259 , n212258 );
buf ( n212260 , n211949 );
not ( n212261 , n212260 );
or ( n212262 , n212259 , n212261 );
buf ( n212263 , n211970 );
not ( n212264 , n212263 );
buf ( n212265 , n212264 );
buf ( n212266 , n212265 );
nand ( n212267 , n212262 , n212266 );
buf ( n212268 , n212267 );
buf ( n212269 , n212268 );
buf ( n212270 , n211978 );
not ( n212271 , n212257 );
not ( n212272 , n212269 );
or ( n212273 , n212271 , n212272 );
nand ( n212274 , n212273 , n212270 );
buf ( n212275 , n212274 );
buf ( n212276 , n211782 );
buf ( n212277 , n211772 );
not ( n212278 , n212277 );
buf ( n212279 , n211899 );
not ( n212280 , n212279 );
buf ( n212281 , n212157 );
nand ( n212282 , n212280 , n212281 );
buf ( n212283 , n212282 );
buf ( n212284 , n212283 );
not ( n212285 , n212284 );
or ( n212286 , n212278 , n212285 );
buf ( n212287 , n211920 );
not ( n212288 , n212287 );
buf ( n212289 , n212288 );
buf ( n212290 , n212289 );
nand ( n212291 , n212286 , n212290 );
buf ( n212292 , n212291 );
buf ( n212293 , n212292 );
buf ( n212294 , n211928 );
not ( n212295 , n212276 );
not ( n212296 , n212293 );
or ( n212297 , n212295 , n212296 );
nand ( n212298 , n212297 , n212294 );
buf ( n212299 , n212298 );
buf ( n212300 , n210830 );
not ( n212301 , n212300 );
buf ( n212302 , n212301 );
buf ( n212303 , n212302 );
buf ( n212304 , n211949 );
buf ( n212305 , n211960 );
not ( n212306 , n212303 );
not ( n212307 , n212304 );
or ( n212308 , n212306 , n212307 );
nand ( n212309 , n212308 , n212305 );
buf ( n212310 , n212309 );
buf ( n212311 , n211762 );
not ( n212312 , n212311 );
buf ( n212313 , n212312 );
buf ( n212314 , n212313 );
buf ( n212315 , n212283 );
buf ( n212316 , n211911 );
not ( n212317 , n212314 );
not ( n212318 , n212315 );
or ( n212319 , n212317 , n212318 );
nand ( n212320 , n212319 , n212316 );
buf ( n212321 , n212320 );
buf ( n212322 , n211678 );
buf ( n212323 , n211604 );
not ( n212324 , n212323 );
buf ( n212325 , n211132 );
not ( n212326 , n212325 );
buf ( n212327 , n211480 );
not ( n212328 , n212327 );
buf ( n212329 , n211414 );
not ( n212330 , n212329 );
buf ( n212331 , n212330 );
buf ( n212332 , n212331 );
nor ( n212333 , n212328 , n212332 );
buf ( n212334 , n212333 );
buf ( n212335 , n212334 );
not ( n212336 , n212335 );
or ( n212337 , n212326 , n212336 );
not ( n212338 , n211555 );
buf ( n212339 , n212338 );
nand ( n212340 , n212337 , n212339 );
buf ( n212341 , n212340 );
buf ( n212342 , n212341 );
not ( n212343 , n212342 );
or ( n212344 , n212324 , n212343 );
buf ( n212345 , n211651 );
nand ( n212346 , n212344 , n212345 );
buf ( n212347 , n212346 );
buf ( n212348 , n212347 );
buf ( n212349 , n211695 );
nand ( n212350 , n212348 , n212349 );
buf ( n212351 , n212350 );
buf ( n212352 , n212351 );
buf ( n212353 , n211689 );
or ( n212354 , n212352 , n212353 );
buf ( n212355 , n211723 );
not ( n212356 , n212355 );
buf ( n212357 , n212356 );
buf ( n212358 , n212357 );
nand ( n212359 , n212354 , n212358 );
buf ( n212360 , n212359 );
buf ( n212361 , n212360 );
buf ( n212362 , n211729 );
not ( n212363 , n212362 );
buf ( n212364 , n212363 );
buf ( n212365 , n212364 );
not ( n212366 , n212322 );
not ( n212367 , n212361 );
or ( n212368 , n212366 , n212367 );
nand ( n212369 , n212368 , n212365 );
buf ( n212370 , n212369 );
buf ( n212371 , n211847 );
buf ( n212372 , n211748 );
buf ( n212373 , n211874 );
not ( n212374 , n212373 );
buf ( n212375 , n212374 );
buf ( n212376 , n212375 );
not ( n212377 , n212371 );
not ( n212378 , n212372 );
or ( n212379 , n212377 , n212378 );
nand ( n212380 , n212379 , n212376 );
buf ( n212381 , n212380 );
buf ( n212382 , n211834 );
not ( n212383 , n212382 );
buf ( n212384 , n212383 );
buf ( n212385 , n212384 );
buf ( n212386 , n211748 );
buf ( n212387 , n211864 );
not ( n212388 , n212385 );
not ( n212389 , n212386 );
or ( n212390 , n212388 , n212389 );
nand ( n212391 , n212390 , n212387 );
buf ( n212392 , n212391 );
buf ( n212393 , n212384 );
buf ( n212394 , n211864 );
nand ( n212395 , n212393 , n212394 );
buf ( n212396 , n212395 );
buf ( n212397 , n212396 );
buf ( n212398 , n211748 );
buf ( n212399 , n212396 );
buf ( n212400 , n211748 );
not ( n212401 , n212397 );
not ( n212402 , n212398 );
or ( n212403 , n212401 , n212402 );
or ( n212404 , n212399 , n212400 );
nand ( n212405 , n212403 , n212404 );
buf ( n212406 , n212405 );
buf ( n212407 , n211576 );
buf ( n212408 , n211598 );
not ( n212409 , n212408 );
buf ( n212410 , n212409 );
buf ( n212411 , n212410 );
not ( n212412 , n212411 );
buf ( n212413 , n212341 );
not ( n212414 , n212413 );
or ( n212415 , n212412 , n212414 );
buf ( n212416 , n211625 );
not ( n212417 , n212416 );
buf ( n212418 , n212417 );
buf ( n212419 , n212418 );
nand ( n212420 , n212415 , n212419 );
buf ( n212421 , n212420 );
buf ( n212422 , n212421 );
buf ( n212423 , n211632 );
not ( n212424 , n212407 );
not ( n212425 , n212422 );
or ( n212426 , n212424 , n212425 );
nand ( n212427 , n212426 , n212423 );
buf ( n212428 , n212427 );
buf ( n212429 , n211595 );
buf ( n212430 , n212341 );
buf ( n212431 , n211616 );
not ( n212432 , n212429 );
not ( n212433 , n212430 );
or ( n212434 , n212432 , n212433 );
nand ( n212435 , n212434 , n212431 );
buf ( n212436 , n212435 );
buf ( n212437 , n211595 );
buf ( n212438 , n211616 );
nand ( n212439 , n212437 , n212438 );
buf ( n212440 , n212439 );
buf ( n212441 , n212440 );
buf ( n212442 , n212341 );
buf ( n212443 , n212440 );
buf ( n212444 , n212341 );
not ( n212445 , n212441 );
not ( n212446 , n212442 );
or ( n212447 , n212445 , n212446 );
or ( n212448 , n212443 , n212444 );
nand ( n212449 , n212447 , n212448 );
buf ( n212450 , n212449 );
buf ( n212451 , n211474 );
not ( n212452 , n212451 );
buf ( n212453 , n212331 );
buf ( n212454 , n211445 );
nor ( n212455 , n212453 , n212454 );
buf ( n212456 , n212455 );
buf ( n212457 , n212456 );
not ( n212458 , n212457 );
or ( n212459 , n212452 , n212458 );
buf ( n212460 , n211499 );
nand ( n212461 , n212459 , n212460 );
buf ( n212462 , n212461 );
buf ( n212463 , n212462 );
buf ( n212464 , n211459 );
buf ( n212465 , n211507 );
nand ( n212466 , n212464 , n212465 );
buf ( n212467 , n212466 );
buf ( n212468 , n212467 );
buf ( n212469 , n212467 );
buf ( n212470 , n212462 );
not ( n212471 , n212463 );
not ( n212472 , n212468 );
or ( n212473 , n212471 , n212472 );
or ( n212474 , n212469 , n212470 );
nand ( n212475 , n212473 , n212474 );
buf ( n212476 , n212475 );
buf ( n212477 , n211107 );
not ( n212478 , n212477 );
buf ( n212479 , n212478 );
buf ( n212480 , n212479 );
buf ( n212481 , n212334 );
buf ( n212482 , n211520 );
or ( n212483 , n212481 , n212482 );
buf ( n212484 , n212483 );
buf ( n212485 , n212484 );
buf ( n212486 , n211530 );
not ( n212487 , n212480 );
not ( n212488 , n212485 );
or ( n212489 , n212487 , n212488 );
nand ( n212490 , n212489 , n212486 );
buf ( n212491 , n212490 );
buf ( n212492 , n212479 );
buf ( n212493 , n211530 );
nand ( n212494 , n212492 , n212493 );
buf ( n212495 , n212494 );
buf ( n212496 , n212495 );
buf ( n212497 , n212484 );
buf ( n212498 , n212495 );
buf ( n212499 , n212484 );
not ( n212500 , n212496 );
not ( n212501 , n212497 );
or ( n212502 , n212500 , n212501 );
or ( n212503 , n212498 , n212499 );
nand ( n212504 , n212502 , n212503 );
buf ( n212505 , n212504 );
buf ( n212506 , n212456 );
not ( n212507 , n212506 );
buf ( n212508 , n211492 );
nand ( n212509 , n212507 , n212508 );
buf ( n212510 , n212509 );
buf ( n212511 , n212510 );
buf ( n212512 , n211498 );
not ( n212513 , n212512 );
buf ( n212514 , n211474 );
nand ( n212515 , n212513 , n212514 );
buf ( n212516 , n212515 );
buf ( n212517 , n212516 );
buf ( n212518 , n212516 );
buf ( n212519 , n212510 );
not ( n212520 , n212511 );
not ( n212521 , n212517 );
or ( n212522 , n212520 , n212521 );
or ( n212523 , n212518 , n212519 );
nand ( n212524 , n212522 , n212523 );
buf ( n212525 , n212524 );
buf ( n212526 , n211182 );
buf ( n212527 , n211189 );
nand ( n212528 , n212526 , n212527 );
buf ( n212529 , n212528 );
buf ( n212530 , n212529 );
buf ( n212531 , n211391 );
buf ( n212532 , n211408 );
and ( n212533 , n212531 , n212532 );
buf ( n212534 , n212533 );
and ( n212535 , n212534 , n211403 );
nor ( n212536 , n212535 , n211157 );
buf ( n212537 , n212536 );
buf ( n212538 , n211396 );
or ( n212539 , n212537 , n212538 );
buf ( n212540 , n211164 );
nand ( n212541 , n212539 , n212540 );
buf ( n212542 , n212541 );
buf ( n212543 , n212542 );
buf ( n212544 , n212529 );
buf ( n212545 , n212542 );
not ( n212546 , n212530 );
not ( n212547 , n212543 );
or ( n212548 , n212546 , n212547 );
or ( n212549 , n212544 , n212545 );
nand ( n212550 , n212548 , n212549 );
buf ( n212551 , n212550 );
buf ( n212552 , n211492 );
not ( n212553 , n212552 );
buf ( n212554 , n211445 );
nor ( n212555 , n212553 , n212554 );
buf ( n212556 , n212555 );
buf ( n212557 , n212556 );
buf ( n212558 , n212331 );
buf ( n212559 , n212556 );
buf ( n212560 , n212331 );
not ( n212561 , n212557 );
not ( n212562 , n212558 );
or ( n212563 , n212561 , n212562 );
or ( n212564 , n212559 , n212560 );
nand ( n212565 , n212563 , n212564 );
buf ( n212566 , n212565 );
buf ( n212567 , n212536 );
buf ( n212568 , n211137 );
buf ( n212569 , n211164 );
and ( n212570 , n212568 , n212569 );
buf ( n212571 , n212570 );
buf ( n212572 , n212571 );
buf ( n212573 , n212571 );
buf ( n212574 , n212536 );
not ( n212575 , n212567 );
not ( n212576 , n212572 );
or ( n212577 , n212575 , n212576 );
or ( n212578 , n212573 , n212574 );
nand ( n212579 , n212577 , n212578 );
buf ( n212580 , n212579 );
buf ( n212581 , n211403 );
buf ( n212582 , n211154 );
nand ( n212583 , n212581 , n212582 );
buf ( n212584 , n212583 );
buf ( n212585 , n212584 );
buf ( n212586 , n212534 );
not ( n212587 , n212586 );
buf ( n212588 , n211148 );
nand ( n212589 , n212587 , n212588 );
buf ( n212590 , n212589 );
buf ( n212591 , n212590 );
buf ( n212592 , n212584 );
buf ( n212593 , n212590 );
not ( n212594 , n212585 );
not ( n212595 , n212591 );
or ( n212596 , n212594 , n212595 );
or ( n212597 , n212592 , n212593 );
nand ( n212598 , n212596 , n212597 );
buf ( n212599 , n212598 );
buf ( n212600 , n211256 );
buf ( n212601 , n211263 );
nand ( n212602 , n212600 , n212601 );
buf ( n212603 , n212602 );
buf ( n212604 , n212603 );
buf ( n212605 , n211371 );
buf ( n212606 , n211381 );
and ( n212607 , n212605 , n212606 );
buf ( n212608 , n211240 );
nor ( n212609 , n212607 , n212608 );
buf ( n212610 , n212609 );
buf ( n212611 , n212610 );
buf ( n212612 , n211206 );
not ( n212613 , n212612 );
buf ( n212614 , n212613 );
buf ( n212615 , n212614 );
or ( n212616 , n212611 , n212615 );
buf ( n212617 , n211247 );
nand ( n212618 , n212616 , n212617 );
buf ( n212619 , n212618 );
buf ( n212620 , n212619 );
buf ( n212621 , n212603 );
buf ( n212622 , n212619 );
not ( n212623 , n212604 );
not ( n212624 , n212620 );
or ( n212625 , n212623 , n212624 );
or ( n212626 , n212621 , n212622 );
nand ( n212627 , n212625 , n212626 );
buf ( n212628 , n212627 );
buf ( n212629 , n211408 );
buf ( n212630 , n211148 );
nand ( n212631 , n212629 , n212630 );
buf ( n212632 , n212631 );
buf ( n212633 , n212632 );
buf ( n212634 , n211391 );
buf ( n212635 , n212632 );
buf ( n212636 , n211391 );
not ( n212637 , n212633 );
not ( n212638 , n212634 );
or ( n212639 , n212637 , n212638 );
or ( n212640 , n212635 , n212636 );
nand ( n212641 , n212639 , n212640 );
buf ( n212642 , n212641 );
buf ( n212643 , n212610 );
buf ( n212644 , n211206 );
buf ( n212645 , n211247 );
and ( n212646 , n212644 , n212645 );
buf ( n212647 , n212646 );
buf ( n212648 , n212647 );
buf ( n212649 , n212647 );
buf ( n212650 , n212610 );
not ( n212651 , n212643 );
not ( n212652 , n212648 );
or ( n212653 , n212651 , n212652 );
or ( n212654 , n212649 , n212650 );
nand ( n212655 , n212653 , n212654 );
buf ( n212656 , n212655 );
buf ( n212657 , n211223 );
not ( n212658 , n212657 );
buf ( n212659 , n211237 );
nand ( n212660 , n212658 , n212659 );
buf ( n212661 , n212660 );
buf ( n212662 , n212661 );
buf ( n212663 , n211378 );
not ( n212664 , n212663 );
buf ( n212665 , n212664 );
buf ( n212666 , n212665 );
not ( n212667 , n212666 );
buf ( n212668 , n211371 );
not ( n212669 , n212668 );
or ( n212670 , n212667 , n212669 );
buf ( n212671 , n211231 );
nand ( n212672 , n212670 , n212671 );
buf ( n212673 , n212672 );
buf ( n212674 , n212673 );
buf ( n212675 , n212661 );
buf ( n212676 , n212673 );
not ( n212677 , n212662 );
not ( n212678 , n212674 );
or ( n212679 , n212677 , n212678 );
or ( n212680 , n212675 , n212676 );
nand ( n212681 , n212679 , n212680 );
buf ( n212682 , n212681 );
buf ( n212683 , n212665 );
buf ( n212684 , n211231 );
nand ( n212685 , n212683 , n212684 );
buf ( n212686 , n212685 );
buf ( n212687 , n212686 );
buf ( n212688 , n211371 );
buf ( n212689 , n212686 );
buf ( n212690 , n211371 );
not ( n212691 , n212687 );
not ( n212692 , n212688 );
or ( n212693 , n212691 , n212692 );
or ( n212694 , n212689 , n212690 );
nand ( n212695 , n212693 , n212694 );
buf ( n212696 , n212695 );
xor ( n212697 , n211269 , n211270 );
xor ( n212698 , n212697 , n211367 );
buf ( n212699 , n212698 );
xor ( n212700 , n211272 , n211281 );
xor ( n212701 , n212700 , n211362 );
buf ( n212702 , n212701 );
xor ( n212703 , n211286 , n211287 );
xor ( n212704 , n212703 , n211357 );
buf ( n212705 , n212704 );
xor ( n212706 , n211289 , n211290 );
xor ( n212707 , n212706 , n211352 );
buf ( n212708 , n212707 );
xor ( n212709 , n211296 , n211297 );
xor ( n212710 , n212709 , n211347 );
buf ( n212711 , n212710 );
buf ( n212712 , n211343 );
not ( n212713 , n212712 );
buf ( n212714 , n211337 );
nor ( n212715 , n212713 , n212714 );
buf ( n212716 , n212715 );
buf ( n212717 , n212716 );
buf ( n212718 , n211328 );
buf ( n212719 , n211328 );
buf ( n212720 , n212716 );
not ( n212721 , n212717 );
not ( n212722 , n212718 );
or ( n212723 , n212721 , n212722 );
or ( n212724 , n212719 , n212720 );
nand ( n212725 , n212723 , n212724 );
buf ( n212726 , n212725 );
buf ( n212727 , n211317 );
not ( n212728 , n212727 );
buf ( n212729 , n212728 );
buf ( n212730 , n212729 );
buf ( n212731 , n211305 );
buf ( n212732 , n211309 );
and ( n212733 , n212731 , n212732 );
buf ( n212734 , n211325 );
nor ( n212735 , n212733 , n212734 );
buf ( n212736 , n212735 );
buf ( n212737 , n212736 );
not ( n212738 , n212737 );
buf ( n212739 , n212738 );
buf ( n212740 , n212739 );
buf ( n212741 , n212729 );
buf ( n212742 , n212739 );
not ( n212743 , n212730 );
not ( n212744 , n212740 );
or ( n212745 , n212743 , n212744 );
or ( n212746 , n212741 , n212742 );
nand ( n212747 , n212745 , n212746 );
buf ( n212748 , n212747 );
buf ( n212749 , n211539 );
not ( n212750 , n212749 );
buf ( n212751 , n212750 );
buf ( n212752 , n212234 );
buf ( n212753 , n212239 );
nand ( n212754 , n212752 , n212753 );
buf ( n212755 , n212754 );
buf ( n212756 , n210958 );
buf ( n212757 , n211008 );
nand ( n212758 , n212756 , n212757 );
buf ( n212759 , n212758 );
buf ( n212760 , n211068 );
buf ( n212761 , n210972 );
nand ( n212762 , n212760 , n212761 );
buf ( n212763 , n212762 );
buf ( n212764 , n211790 );
buf ( n212765 , n211940 );
nand ( n212766 , n212764 , n212765 );
buf ( n212767 , n212766 );
buf ( n212768 , n211568 );
buf ( n212769 , n211645 );
nand ( n212770 , n212768 , n212769 );
buf ( n212771 , n212770 );
buf ( n212772 , n211099 );
buf ( n212773 , n211536 );
not ( n212774 , n212772 );
nand ( n212775 , n212774 , n212773 );
buf ( n212776 , n212775 );
buf ( n212777 , n212313 );
buf ( n212778 , n211911 );
nand ( n212779 , n212777 , n212778 );
buf ( n212780 , n212779 );
buf ( n212781 , n211820 );
buf ( n212782 , n211881 );
not ( n212783 , n212782 );
buf ( n212784 , n212783 );
buf ( n212785 , n212784 );
nand ( n212786 , n212781 , n212785 );
buf ( n212787 , n212786 );
buf ( n212788 , n211844 );
buf ( n212789 , n211871 );
not ( n212790 , n212788 );
nand ( n212791 , n212790 , n212789 );
buf ( n212792 , n212791 );
buf ( n212793 , n211695 );
buf ( n212794 , n211714 );
nand ( n212795 , n212793 , n212794 );
buf ( n212796 , n212795 );
buf ( n212797 , n211117 );
buf ( n212798 , n211543 );
nand ( n212799 , n212797 , n212798 );
buf ( n212800 , n212799 );
buf ( n212801 , n211782 );
buf ( n212802 , n211928 );
nand ( n212803 , n212801 , n212802 );
buf ( n212804 , n212803 );
buf ( n212805 , n211678 );
buf ( n212806 , n212364 );
nand ( n212807 , n212805 , n212806 );
buf ( n212808 , n212807 );
buf ( n212809 , n210928 );
buf ( n212810 , n211054 );
nand ( n212811 , n212809 , n212810 );
buf ( n212812 , n212811 );
buf ( n212813 , n211025 );
buf ( n212814 , n211032 );
nand ( n212815 , n212813 , n212814 );
buf ( n212816 , n212815 );
buf ( n212817 , n211576 );
buf ( n212818 , n211632 );
nand ( n212819 , n212817 , n212818 );
buf ( n212820 , n212819 );
buf ( n212821 , n211769 );
buf ( n212822 , n211917 );
not ( n212823 , n212821 );
nand ( n212824 , n212823 , n212822 );
buf ( n212825 , n212824 );
buf ( n212826 , n211073 );
buf ( n212827 , n210984 );
nand ( n212828 , n212826 , n212827 );
buf ( n212829 , n212828 );
buf ( n212830 , n211662 );
buf ( n212831 , n211739 );
nand ( n212832 , n212830 , n212831 );
buf ( n212833 , n212832 );
buf ( n212834 , n210939 );
buf ( n212835 , n211043 );
nand ( n212836 , n212834 , n212835 );
buf ( n212837 , n212836 );
buf ( n212838 , n210780 );
buf ( n212839 , n212095 );
nand ( n212840 , n212838 , n212839 );
buf ( n212841 , n212840 );
buf ( n212842 , n212053 );
buf ( n212843 , n212078 );
nand ( n212844 , n212842 , n212843 );
buf ( n212845 , n212844 );
buf ( n212846 , n212041 );
buf ( n212847 , n212065 );
nand ( n212848 , n212846 , n212847 );
buf ( n212849 , n212848 );
buf ( n212850 , n211998 );
buf ( n212851 , n212021 );
nand ( n212852 , n212850 , n212851 );
buf ( n212853 , n212852 );
buf ( n212854 , n210869 );
buf ( n212855 , n212011 );
not ( n212856 , n212854 );
nand ( n212857 , n212856 , n212855 );
buf ( n212858 , n212857 );
buf ( n212859 , n211129 );
buf ( n212860 , n211554 );
nand ( n212861 , n212859 , n212860 );
buf ( n212862 , n212861 );
buf ( n212863 , n212209 );
buf ( n212864 , n212005 );
nand ( n212865 , n212863 , n212864 );
buf ( n212866 , n212865 );
buf ( n212867 , n210816 );
buf ( n212868 , n211988 );
nand ( n212869 , n212867 , n212868 );
buf ( n212870 , n212869 );
buf ( n212871 , n210806 );
buf ( n212872 , n211978 );
nand ( n212873 , n212871 , n212872 );
buf ( n212874 , n212873 );
buf ( n212875 , n210840 );
buf ( n212876 , n211967 );
not ( n212877 , n212875 );
nand ( n212878 , n212877 , n212876 );
buf ( n212879 , n212878 );
buf ( n212880 , n212302 );
buf ( n212881 , n211960 );
nand ( n212882 , n212880 , n212881 );
buf ( n212883 , n212882 );
buf ( n212884 , n211585 );
buf ( n212885 , n211622 );
nand ( n212886 , n212884 , n212885 );
buf ( n212887 , n212886 );
buf ( n212888 , n210770 );
buf ( n212889 , n210774 );
buf ( n212890 , n210770 );
buf ( n212891 , n210774 );
not ( n212892 , n212888 );
not ( n212893 , n212889 );
and ( n212894 , n212892 , n212893 );
and ( n212895 , n212890 , n212891 );
nor ( n212896 , n212894 , n212895 );
buf ( n212897 , n212896 );
buf ( n212898 , n212134 );
buf ( n212899 , n212845 );
xnor ( n212900 , n212898 , n212899 );
buf ( n212901 , n212900 );
buf ( n212902 , n212193 );
buf ( n212903 , n210972 );
not ( n212904 , n212902 );
nand ( n212905 , n212904 , n212903 );
buf ( n212906 , n212905 );
buf ( n212907 , n212360 );
buf ( n212908 , n212808 );
xnor ( n212909 , n212907 , n212908 );
buf ( n212910 , n212909 );
buf ( n212911 , n212174 );
buf ( n212912 , n212755 );
xnor ( n212913 , n212911 , n212912 );
buf ( n212914 , n212913 );
buf ( n212915 , n212206 );
buf ( n212916 , n212759 );
xnor ( n212917 , n212915 , n212916 );
buf ( n212918 , n212917 );
buf ( n212919 , n212299 );
buf ( n212920 , n212767 );
xnor ( n212921 , n212919 , n212920 );
buf ( n212922 , n212921 );
buf ( n212923 , n212428 );
buf ( n212924 , n212771 );
xnor ( n212925 , n212923 , n212924 );
buf ( n212926 , n212925 );
buf ( n212927 , n212491 );
buf ( n212928 , n212776 );
xnor ( n212929 , n212927 , n212928 );
buf ( n212930 , n212929 );
buf ( n212931 , n212283 );
buf ( n212932 , n212780 );
xnor ( n212933 , n212931 , n212932 );
buf ( n212934 , n212933 );
buf ( n212935 , n212381 );
buf ( n212936 , n212787 );
xnor ( n212937 , n212935 , n212936 );
buf ( n212938 , n212937 );
buf ( n212939 , n212392 );
buf ( n212940 , n212792 );
xnor ( n212941 , n212939 , n212940 );
buf ( n212942 , n212941 );
buf ( n212943 , n212347 );
buf ( n212944 , n212796 );
xnor ( n212945 , n212943 , n212944 );
buf ( n212946 , n212945 );
not ( n212947 , n211110 );
not ( n212948 , n212484 );
or ( n212949 , n212947 , n212948 );
nand ( n212950 , n212949 , n212751 );
buf ( n212951 , n212950 );
buf ( n212952 , n212800 );
xnor ( n212953 , n212951 , n212952 );
buf ( n212954 , n212953 );
buf ( n212955 , n212292 );
buf ( n212956 , n212804 );
xnor ( n212957 , n212955 , n212956 );
buf ( n212958 , n212957 );
buf ( n212959 , n212190 );
buf ( n212960 , n212812 );
xnor ( n212961 , n212959 , n212960 );
buf ( n212962 , n212961 );
buf ( n212963 , n212245 );
buf ( n212964 , n212816 );
xnor ( n212965 , n212963 , n212964 );
buf ( n212966 , n212965 );
buf ( n212967 , n212421 );
buf ( n212968 , n212820 );
xnor ( n212969 , n212967 , n212968 );
buf ( n212970 , n212969 );
buf ( n212971 , n212321 );
buf ( n212972 , n212825 );
xnor ( n212973 , n212971 , n212972 );
buf ( n212974 , n212973 );
buf ( n212975 , n212906 );
buf ( n212976 , n212829 );
xnor ( n212977 , n212975 , n212976 );
buf ( n212978 , n212977 );
buf ( n212979 , n212370 );
buf ( n212980 , n212833 );
xnor ( n212981 , n212979 , n212980 );
buf ( n212982 , n212981 );
buf ( n212983 , n212183 );
buf ( n212984 , n212837 );
xnor ( n212985 , n212983 , n212984 );
buf ( n212986 , n212985 );
buf ( n212987 , n212088 );
buf ( n212988 , n212841 );
xnor ( n212989 , n212987 , n212988 );
buf ( n212990 , n212989 );
buf ( n212991 , n212036 );
buf ( n212992 , n212849 );
xnor ( n212993 , n212991 , n212992 );
buf ( n212994 , n212993 );
buf ( n212995 , n212256 );
buf ( n212996 , n212853 );
xnor ( n212997 , n212995 , n212996 );
buf ( n212998 , n212997 );
buf ( n212999 , n212231 );
buf ( n213000 , n212858 );
xnor ( n213001 , n212999 , n213000 );
buf ( n213002 , n213001 );
not ( n213003 , n211117 );
not ( n213004 , n212950 );
or ( n213005 , n213003 , n213004 );
nand ( n213006 , n213005 , n211543 );
buf ( n213007 , n213006 );
buf ( n213008 , n212862 );
xnor ( n213009 , n213007 , n213008 );
buf ( n213010 , n213009 );
buf ( n213011 , n212224 );
buf ( n213012 , n212866 );
xnor ( n213013 , n213011 , n213012 );
buf ( n213014 , n213013 );
buf ( n213015 , n212275 );
buf ( n213016 , n212870 );
xnor ( n213017 , n213015 , n213016 );
buf ( n213018 , n213017 );
buf ( n213019 , n212268 );
buf ( n213020 , n212874 );
xnor ( n213021 , n213019 , n213020 );
buf ( n213022 , n213021 );
buf ( n213023 , n212310 );
buf ( n213024 , n212879 );
xnor ( n213025 , n213023 , n213024 );
buf ( n213026 , n213025 );
buf ( n213027 , n211949 );
buf ( n213028 , n212883 );
xnor ( n213029 , n213027 , n213028 );
buf ( n213030 , n213029 );
buf ( n213031 , n212436 );
buf ( n213032 , n212887 );
xnor ( n213033 , n213031 , n213032 );
buf ( n213034 , n213033 );
not ( n213035 , n37569 );
not ( n213036 , n213035 );
not ( n213037 , n37566 );
not ( n213038 , n213037 );
or ( n213039 , n213036 , n213038 );
nand ( n213040 , n213039 , n37570 );
buf ( n213041 , n213040 );
not ( n213042 , n213041 );
or ( n213043 , n37502 , n37501 );
nand ( n213044 , n213043 , n37503 );
not ( n213045 , n213044 );
not ( n213046 , n213045 );
or ( n213047 , n213042 , n213046 );
not ( n213048 , n213041 );
nand ( n213049 , n213044 , n213048 );
nand ( n213050 , n213047 , n213049 );
buf ( n213051 , n209375 );
and ( n213052 , n213050 , n213051 );
not ( n213053 , n37698 );
and ( n213054 , n37684 , n213053 );
not ( n213055 , n37684 );
and ( n213056 , n213055 , n37698 );
nor ( n213057 , n213054 , n213056 );
not ( n213058 , n213057 );
not ( n213059 , n213058 );
buf ( n213060 , n213040 );
not ( n213061 , n213060 );
not ( n213062 , n30666 );
not ( n213063 , n213062 );
or ( n213064 , n213061 , n213063 );
not ( n213065 , n213040 );
nand ( n213066 , n213065 , n30666 );
nand ( n213067 , n213064 , n213066 );
not ( n213068 , n213067 );
or ( n213069 , n213059 , n213068 );
not ( n213070 , n213040 );
nand ( n213071 , n213070 , n213053 );
not ( n213072 , n213071 );
nand ( n213073 , n213040 , n37698 );
nand ( n213074 , n213073 , n213057 );
nor ( n213075 , n213072 , n213074 );
buf ( n213076 , n213075 );
not ( n213077 , n168522 );
or ( n213078 , n213040 , n213077 );
nand ( n213079 , n213077 , n213040 );
nand ( n213080 , n213078 , n213079 );
nand ( n213081 , n213076 , n213080 );
nand ( n213082 , n213069 , n213081 );
xor ( n213083 , n213052 , n213082 );
not ( n213084 , n209375 );
nand ( n213085 , n213053 , n213084 );
not ( n213086 , n37684 );
not ( n213087 , n213086 );
and ( n213088 , n213085 , n213087 );
and ( n213089 , n37698 , n213051 );
nor ( n213090 , n213088 , n213089 , n213065 );
xnor ( n213091 , n213084 , n213040 );
not ( n213092 , n213091 );
not ( n213093 , n213075 );
or ( n213094 , n213092 , n213093 );
not ( n213095 , n213057 );
nand ( n213096 , n213095 , n213080 );
nand ( n213097 , n213094 , n213096 );
and ( n213098 , n213090 , n213097 );
xor ( n213099 , n213083 , n213098 );
xor ( n213100 , n213052 , n213082 );
and ( n213101 , n213100 , n213098 );
and ( n213102 , n213052 , n213082 );
or ( n213103 , n213101 , n213102 );
not ( n213104 , n213051 );
xnor ( n213105 , n37496 , n37610 );
not ( n213106 , n213105 );
and ( n213107 , n213104 , n213106 );
not ( n213108 , n213104 );
not ( n213109 , n213106 );
and ( n213110 , n213108 , n213109 );
nor ( n213111 , n213107 , n213110 );
not ( n213112 , n213111 );
and ( n213113 , n213105 , n213044 );
not ( n213114 , n213105 );
and ( n213115 , n213114 , n213045 );
nor ( n213116 , n213113 , n213115 );
not ( n213117 , n213041 );
not ( n213118 , n213044 );
or ( n213119 , n213117 , n213118 );
nand ( n213120 , n213045 , n213048 );
nand ( n213121 , n213119 , n213120 );
and ( n213122 , n213116 , n213121 );
not ( n213123 , n213122 );
or ( n213124 , n213112 , n213123 );
not ( n213125 , n213121 );
not ( n213126 , n213077 );
not ( n213127 , n213126 );
not ( n213128 , n213106 );
or ( n213129 , n213127 , n213128 );
buf ( n213130 , n213105 );
nand ( n213131 , n213130 , n213077 );
nand ( n213132 , n213129 , n213131 );
nand ( n213133 , n213125 , n213132 );
nand ( n213134 , n213124 , n213133 );
not ( n213135 , n213045 );
or ( n213136 , n213135 , n213051 );
buf ( n213137 , n213060 );
nand ( n213138 , n213136 , n213137 );
not ( n213139 , n213104 );
nand ( n213140 , n213135 , n213139 );
and ( n213141 , n213109 , n213138 , n213140 );
not ( n213142 , n213057 );
not ( n213143 , n213142 );
not ( n213144 , n30643 );
and ( n213145 , n213144 , n213137 );
not ( n213146 , n213144 );
not ( n213147 , n213060 );
and ( n213148 , n213146 , n213147 );
or ( n213149 , n213145 , n213148 );
not ( n213150 , n213149 );
or ( n213151 , n213143 , n213150 );
buf ( n213152 , n213076 );
nand ( n213153 , n213067 , n213152 );
nand ( n213154 , n213151 , n213153 );
xor ( n213155 , n213141 , n213154 );
xor ( n213156 , n213134 , n213155 );
not ( n213157 , n211314 );
not ( n213158 , n209348 );
and ( n213159 , n213158 , n213087 );
not ( n213160 , n213158 );
and ( n213161 , n213160 , n213086 );
or ( n213162 , n213159 , n213161 );
not ( n213163 , n213162 );
or ( n213164 , n213157 , n213163 );
not ( n213165 , n213087 );
not ( n213166 , n209360 );
not ( n213167 , n213166 );
or ( n213168 , n213165 , n213167 );
nand ( n213169 , n209360 , n213086 );
nand ( n213170 , n213168 , n213169 );
not ( n213171 , n211314 );
nand ( n213172 , n213171 , n37684 );
not ( n213173 , n213172 );
nand ( n213174 , n213170 , n213173 );
nand ( n213175 , n213164 , n213174 );
xor ( n213176 , n213156 , n213175 );
xor ( n213177 , n213134 , n213155 );
and ( n213178 , n213177 , n213175 );
and ( n213179 , n213134 , n213155 );
or ( n213180 , n213178 , n213179 );
not ( n213181 , n213132 );
not ( n213182 , n213122 );
or ( n213183 , n213181 , n213182 );
not ( n213184 , n213106 );
not ( n213185 , n30666 );
or ( n213186 , n213184 , n213185 );
not ( n213187 , n213106 );
not ( n213188 , n30666 );
nand ( n213189 , n213187 , n213188 );
nand ( n213190 , n213186 , n213189 );
nand ( n213191 , n213190 , n213050 );
nand ( n213192 , n213183 , n213191 );
nand ( n213193 , n36149 , n36151 );
nand ( n213194 , n36014 , n37589 );
not ( n213195 , n213194 );
and ( n213196 , n213193 , n213195 );
not ( n213197 , n213193 );
and ( n213198 , n213197 , n213194 );
nor ( n213199 , n213196 , n213198 );
not ( n213200 , n213199 );
and ( n213201 , n213106 , n213200 );
not ( n213202 , n213106 );
and ( n213203 , n213202 , n213199 );
nor ( n213204 , n213201 , n213203 );
not ( n213205 , n213204 );
not ( n213206 , n213205 );
and ( n213207 , n213206 , n213051 );
xor ( n213208 , n213192 , n213207 );
not ( n213209 , n213058 );
not ( n213210 , n213137 );
not ( n213211 , n213166 );
or ( n213212 , n213210 , n213211 );
nand ( n213213 , n209360 , n213147 );
nand ( n213214 , n213212 , n213213 );
not ( n213215 , n213214 );
or ( n213216 , n213209 , n213215 );
buf ( n213217 , n213076 );
nand ( n213218 , n213149 , n213217 );
nand ( n213219 , n213216 , n213218 );
xor ( n213220 , n213208 , n213219 );
xor ( n213221 , n213192 , n213207 );
and ( n213222 , n213221 , n213219 );
and ( n213223 , n213192 , n213207 );
or ( n213224 , n213222 , n213223 );
and ( n213225 , n213141 , n213154 );
xor ( n213226 , n213225 , n213220 );
not ( n213227 , n211314 );
not ( n213228 , n213087 );
not ( n213229 , n209316 );
not ( n213230 , n213229 );
or ( n213231 , n213228 , n213230 );
not ( n213232 , n213229 );
nand ( n213233 , n213232 , n213086 );
nand ( n213234 , n213231 , n213233 );
not ( n213235 , n213234 );
or ( n213236 , n213227 , n213235 );
nand ( n213237 , n213162 , n213173 );
nand ( n213238 , n213236 , n213237 );
xor ( n213239 , n213226 , n213238 );
xor ( n213240 , n213225 , n213220 );
and ( n213241 , n213240 , n213238 );
and ( n213242 , n213225 , n213220 );
or ( n213243 , n213241 , n213242 );
not ( n213244 , n213139 );
not ( n213245 , n37628 );
and ( n213246 , n35963 , n36013 );
nand ( n213247 , n213246 , n37676 , n37502 );
not ( n213248 , n36148 );
not ( n213249 , n37675 );
or ( n213250 , n213248 , n213249 );
nand ( n213251 , n213250 , n35961 );
nand ( n213252 , n213247 , n213251 , n36151 );
not ( n213253 , n213252 );
not ( n213254 , n213253 );
or ( n213255 , n213245 , n213254 );
nand ( n213256 , n37627 , n213252 );
nand ( n213257 , n213255 , n213256 );
not ( n213258 , n213257 );
not ( n213259 , n213258 );
or ( n213260 , n213244 , n213259 );
buf ( n213261 , n213257 );
nand ( n213262 , n213261 , n213104 );
nand ( n213263 , n213260 , n213262 );
not ( n213264 , n213263 );
not ( n213265 , n213204 );
not ( n213266 , n213257 );
not ( n213267 , n213200 );
or ( n213268 , n213266 , n213267 );
or ( n213269 , n213257 , n213200 );
nand ( n213270 , n213268 , n213269 );
nand ( n213271 , n213265 , n213270 );
not ( n213272 , n213271 );
not ( n213273 , n213272 );
or ( n213274 , n213264 , n213273 );
not ( n213275 , n213126 );
not ( n213276 , n213258 );
or ( n213277 , n213275 , n213276 );
not ( n213278 , n213258 );
nand ( n213279 , n213278 , n213077 );
nand ( n213280 , n213277 , n213279 );
nand ( n213281 , n213206 , n213280 );
nand ( n213282 , n213274 , n213281 );
not ( n213283 , n213190 );
not ( n213284 , n213122 );
or ( n213285 , n213283 , n213284 );
not ( n213286 , n30643 );
not ( n213287 , n213106 );
or ( n213288 , n213286 , n213287 );
nand ( n213289 , n213144 , n213130 );
nand ( n213290 , n213288 , n213289 );
nand ( n213291 , n213290 , n213050 );
nand ( n213292 , n213285 , n213291 );
not ( n213293 , n213261 );
buf ( n213294 , n213199 );
nor ( n213295 , n213294 , n213139 );
or ( n213296 , n213295 , n213106 );
nand ( n213297 , n213294 , n213051 );
nand ( n213298 , n213296 , n213297 );
nor ( n213299 , n213293 , n213298 );
xor ( n213300 , n213292 , n213299 );
xor ( n213301 , n213282 , n213300 );
not ( n213302 , n213214 );
not ( n213303 , n213217 );
or ( n213304 , n213302 , n213303 );
not ( n213305 , n213147 );
not ( n213306 , n209348 );
and ( n213307 , n213305 , n213306 );
buf ( n213308 , n209348 );
and ( n213309 , n213308 , n213147 );
nor ( n213310 , n213307 , n213309 );
or ( n213311 , n213310 , n213057 );
nand ( n213312 , n213304 , n213311 );
xor ( n213313 , n213301 , n213312 );
xor ( n213314 , n213282 , n213300 );
and ( n213315 , n213314 , n213312 );
and ( n213316 , n213282 , n213300 );
or ( n213317 , n213315 , n213316 );
not ( n213318 , n211314 );
not ( n213319 , n213086 );
not ( n213320 , n30498 );
or ( n213321 , n213319 , n213320 );
not ( n213322 , n30498 );
nand ( n213323 , n213322 , n213087 );
nand ( n213324 , n213321 , n213323 );
not ( n213325 , n213324 );
or ( n213326 , n213318 , n213325 );
nand ( n213327 , n213234 , n213173 );
nand ( n213328 , n213326 , n213327 );
xor ( n213329 , n213224 , n213328 );
xor ( n213330 , n213329 , n213313 );
xor ( n213331 , n213224 , n213328 );
and ( n213332 , n213331 , n213313 );
and ( n213333 , n213224 , n213328 );
or ( n213334 , n213332 , n213333 );
not ( n213335 , n213050 );
and ( n213336 , n209359 , n213106 );
not ( n213337 , n209359 );
and ( n213338 , n213337 , n213130 );
or ( n213339 , n213336 , n213338 );
not ( n213340 , n213339 );
or ( n213341 , n213335 , n213340 );
nand ( n213342 , n213122 , n213290 );
nand ( n213343 , n213341 , n213342 );
not ( n213344 , n213280 );
not ( n213345 , n213272 );
or ( n213346 , n213344 , n213345 );
not ( n213347 , n213188 );
and ( n213348 , n213258 , n213347 );
not ( n213349 , n213258 );
and ( n213350 , n213349 , n213188 );
or ( n213351 , n213348 , n213350 );
nand ( n213352 , n213351 , n213206 );
nand ( n213353 , n213346 , n213352 );
xor ( n213354 , n213343 , n213353 );
xor ( n213355 , n37029 , n37674 );
xnor ( n213356 , n213278 , n213355 );
nor ( n213357 , n213356 , n213104 );
xor ( n213358 , n213354 , n213357 );
xor ( n213359 , n213343 , n213353 );
and ( n213360 , n213359 , n213357 );
and ( n213361 , n213343 , n213353 );
or ( n213362 , n213360 , n213361 );
and ( n213363 , n213292 , n213299 );
not ( n213364 , n213142 );
and ( n213365 , n213229 , n213137 );
not ( n213366 , n213229 );
and ( n213367 , n213366 , n213147 );
or ( n213368 , n213365 , n213367 );
not ( n213369 , n213368 );
or ( n213370 , n213364 , n213369 );
not ( n213371 , n213310 );
nand ( n213372 , n213371 , n213217 );
nand ( n213373 , n213370 , n213372 );
xor ( n213374 , n213363 , n213373 );
xor ( n213375 , n213374 , n213317 );
xor ( n213376 , n213363 , n213373 );
and ( n213377 , n213376 , n213317 );
and ( n213378 , n213363 , n213373 );
or ( n213379 , n213377 , n213378 );
not ( n213380 , n211314 );
buf ( n213381 , n213086 );
not ( n213382 , n213381 );
not ( n213383 , n213382 );
not ( n213384 , n30412 );
not ( n213385 , n213384 );
or ( n213386 , n213383 , n213385 );
nand ( n213387 , n30412 , n213381 );
nand ( n213388 , n213386 , n213387 );
not ( n213389 , n213388 );
or ( n213390 , n213380 , n213389 );
nand ( n213391 , n213324 , n213173 );
nand ( n213392 , n213390 , n213391 );
xor ( n213393 , n213358 , n213392 );
xor ( n213394 , n213393 , n213375 );
xor ( n213395 , n213358 , n213392 );
and ( n213396 , n213395 , n213375 );
and ( n213397 , n213358 , n213392 );
or ( n213398 , n213396 , n213397 );
buf ( n213399 , n37096 );
not ( n213400 , n213399 );
buf ( n213401 , n213355 );
nand ( n213402 , n213401 , n213139 );
not ( n213403 , n213261 );
and ( n213404 , n213402 , n213403 );
nor ( n213405 , n213401 , n213139 );
nor ( n213406 , n213404 , n213405 );
nor ( n213407 , n213400 , n213406 );
not ( n213408 , n213050 );
and ( n213409 , n209347 , n213106 );
not ( n213410 , n209347 );
and ( n213411 , n213410 , n213109 );
or ( n213412 , n213409 , n213411 );
not ( n213413 , n213412 );
or ( n213414 , n213408 , n213413 );
nand ( n213415 , n213122 , n213339 );
nand ( n213416 , n213414 , n213415 );
not ( n213417 , n213351 );
not ( n213418 , n213272 );
or ( n213419 , n213417 , n213418 );
not ( n213420 , n213403 );
buf ( n213421 , n30643 );
not ( n213422 , n213421 );
or ( n213423 , n213420 , n213422 );
not ( n213424 , n213421 );
nand ( n213425 , n213261 , n213424 );
nand ( n213426 , n213423 , n213425 );
nand ( n213427 , n213426 , n213206 );
nand ( n213428 , n213419 , n213427 );
xor ( n213429 , n213416 , n213428 );
xor ( n213430 , n213407 , n213429 );
xor ( n213431 , n213430 , n213362 );
xor ( n213432 , n213407 , n213429 );
and ( n213433 , n213432 , n213362 );
and ( n213434 , n213407 , n213429 );
or ( n213435 , n213433 , n213434 );
not ( n213436 , n213142 );
not ( n213437 , n213147 );
not ( n213438 , n30498 );
or ( n213439 , n213437 , n213438 );
nand ( n213440 , n213322 , n213137 );
nand ( n213441 , n213439 , n213440 );
not ( n213442 , n213441 );
or ( n213443 , n213436 , n213442 );
nand ( n213444 , n213368 , n213217 );
nand ( n213445 , n213443 , n213444 );
and ( n213446 , n213051 , n213399 );
not ( n213447 , n213051 );
not ( n213448 , n213399 );
and ( n213449 , n213447 , n213448 );
nor ( n213450 , n213446 , n213449 );
not ( n213451 , n213450 );
or ( n213452 , n213401 , n37096 );
nand ( n213453 , n213401 , n37096 );
and ( n213454 , n213452 , n213453 , n213356 );
not ( n213455 , n213454 );
or ( n213456 , n213451 , n213455 );
not ( n213457 , n213126 );
not ( n213458 , n37096 );
not ( n213459 , n213458 );
or ( n213460 , n213457 , n213459 );
nand ( n213461 , n213399 , n213077 );
nand ( n213462 , n213460 , n213461 );
not ( n213463 , n213356 );
nand ( n213464 , n213462 , n213463 );
nand ( n213465 , n213456 , n213464 );
xor ( n213466 , n213445 , n213465 );
xor ( n213467 , n213466 , n213431 );
xor ( n213468 , n213445 , n213465 );
and ( n213469 , n213468 , n213431 );
and ( n213470 , n213445 , n213465 );
or ( n213471 , n213469 , n213470 );
not ( n213472 , n211314 );
not ( n213473 , n30610 );
and ( n213474 , n213381 , n213473 );
not ( n213475 , n213381 );
and ( n213476 , n213475 , n41981 );
nor ( n213477 , n213474 , n213476 );
not ( n213478 , n213477 );
or ( n213479 , n213472 , n213478 );
nand ( n213480 , n213388 , n213173 );
nand ( n213481 , n213479 , n213480 );
xor ( n213482 , n213481 , n213379 );
xor ( n213483 , n213482 , n213467 );
xor ( n213484 , n213481 , n213379 );
and ( n213485 , n213484 , n213467 );
and ( n213486 , n213481 , n213379 );
or ( n213487 , n213485 , n213486 );
not ( n213488 , n213426 );
not ( n213489 , n213272 );
or ( n213490 , n213488 , n213489 );
not ( n213491 , n209360 );
not ( n213492 , n213403 );
or ( n213493 , n213491 , n213492 );
nand ( n213494 , n213278 , n213166 );
nand ( n213495 , n213493 , n213494 );
nand ( n213496 , n213495 , n213206 );
nand ( n213497 , n213490 , n213496 );
buf ( n213498 , n213050 );
not ( n213499 , n213498 );
and ( n213500 , n209316 , n213106 );
not ( n213501 , n209316 );
and ( n213502 , n213501 , n213109 );
or ( n213503 , n213500 , n213502 );
not ( n213504 , n213503 );
or ( n213505 , n213499 , n213504 );
nand ( n213506 , n213412 , n213122 );
nand ( n213507 , n213505 , n213506 );
xor ( n213508 , n213497 , n213507 );
not ( n213509 , n37084 );
not ( n213510 , n213509 );
not ( n213511 , n213399 );
and ( n213512 , n213510 , n213511 );
not ( n213513 , n213458 );
and ( n213514 , n213509 , n213513 );
nor ( n213515 , n213512 , n213514 );
nor ( n213516 , n213515 , n213104 );
xor ( n213517 , n213508 , n213516 );
xor ( n213518 , n213497 , n213507 );
and ( n213519 , n213518 , n213516 );
and ( n213520 , n213497 , n213507 );
or ( n213521 , n213519 , n213520 );
and ( n213522 , n213416 , n213428 );
not ( n213523 , n213462 );
not ( n213524 , n213454 );
or ( n213525 , n213523 , n213524 );
not ( n213526 , n213347 );
not ( n213527 , n213448 );
or ( n213528 , n213526 , n213527 );
nand ( n213529 , n213399 , n213188 );
nand ( n213530 , n213528 , n213529 );
nand ( n213531 , n213530 , n213463 );
nand ( n213532 , n213525 , n213531 );
xor ( n213533 , n213522 , n213532 );
not ( n213534 , n213142 );
not ( n213535 , n213060 );
not ( n213536 , n213384 );
or ( n213537 , n213535 , n213536 );
nand ( n213538 , n30412 , n213147 );
nand ( n213539 , n213537 , n213538 );
not ( n213540 , n213539 );
or ( n213541 , n213534 , n213540 );
nand ( n213542 , n213441 , n213217 );
nand ( n213543 , n213541 , n213542 );
xor ( n213544 , n213533 , n213543 );
xor ( n213545 , n213522 , n213532 );
and ( n213546 , n213545 , n213543 );
and ( n213547 , n213522 , n213532 );
or ( n213548 , n213546 , n213547 );
not ( n213549 , n211314 );
and ( n213550 , n41978 , n213381 );
not ( n213551 , n41978 );
and ( n213552 , n213551 , n213382 );
or ( n213553 , n213550 , n213552 );
not ( n213554 , n213553 );
or ( n213555 , n213549 , n213554 );
nand ( n213556 , n213173 , n213477 );
nand ( n213557 , n213555 , n213556 );
xor ( n213558 , n213517 , n213557 );
xor ( n213559 , n213558 , n213435 );
xor ( n213560 , n213517 , n213557 );
and ( n213561 , n213560 , n213435 );
and ( n213562 , n213517 , n213557 );
or ( n213563 , n213561 , n213562 );
xor ( n213564 , n213544 , n213471 );
xor ( n213565 , n213564 , n213559 );
xor ( n213566 , n213544 , n213471 );
and ( n213567 , n213566 , n213559 );
and ( n213568 , n213544 , n213471 );
or ( n213569 , n213567 , n213568 );
not ( n213570 , n213498 );
and ( n213571 , n30498 , n213106 );
not ( n213572 , n30498 );
and ( n213573 , n213572 , n213109 );
or ( n213574 , n213571 , n213573 );
not ( n213575 , n213574 );
or ( n213576 , n213570 , n213575 );
buf ( n213577 , n213122 );
nand ( n213578 , n213503 , n213577 );
nand ( n213579 , n213576 , n213578 );
not ( n213580 , n213530 );
not ( n213581 , n213454 );
or ( n213582 , n213580 , n213581 );
not ( n213583 , n213424 );
not ( n213584 , n213583 );
not ( n213585 , n213458 );
or ( n213586 , n213584 , n213585 );
nand ( n213587 , n213399 , n213424 );
nand ( n213588 , n213586 , n213587 );
nand ( n213589 , n213463 , n213588 );
nand ( n213590 , n213582 , n213589 );
xor ( n213591 , n213579 , n213590 );
not ( n213592 , n213495 );
not ( n213593 , n213272 );
or ( n213594 , n213592 , n213593 );
not ( n213595 , n213261 );
not ( n213596 , n213158 );
or ( n213597 , n213595 , n213596 );
nand ( n213598 , n213308 , n213403 );
nand ( n213599 , n213597 , n213598 );
nand ( n213600 , n213206 , n213599 );
nand ( n213601 , n213594 , n213600 );
nand ( n213602 , n213509 , n213104 );
nand ( n213603 , n213399 , n213602 );
not ( n213604 , n36262 );
nor ( n213605 , n213604 , n37606 );
and ( n213606 , n37426 , n213605 );
not ( n213607 , n37426 );
and ( n213608 , n213607 , n37608 );
nor ( n213609 , n213606 , n213608 );
not ( n213610 , n213609 );
not ( n213611 , n213610 );
nand ( n213612 , n37084 , n213051 );
and ( n213613 , n213603 , n213611 , n213612 );
xor ( n213614 , n213601 , n213613 );
xor ( n213615 , n213591 , n213614 );
xor ( n213616 , n213579 , n213590 );
and ( n213617 , n213616 , n213614 );
and ( n213618 , n213579 , n213590 );
or ( n213619 , n213617 , n213618 );
and ( n213620 , n213051 , n213611 );
not ( n213621 , n213051 );
buf ( n213622 , n213610 );
and ( n213623 , n213621 , n213622 );
nor ( n213624 , n213620 , n213623 );
not ( n213625 , n213624 );
not ( n213626 , n37084 );
not ( n213627 , n213610 );
or ( n213628 , n213626 , n213627 );
nand ( n213629 , n213609 , n213509 );
nand ( n213630 , n213628 , n213629 );
and ( n213631 , n213515 , n213630 );
not ( n213632 , n213631 );
or ( n213633 , n213625 , n213632 );
not ( n213634 , n213126 );
not ( n213635 , n213611 );
not ( n213636 , n213635 );
or ( n213637 , n213634 , n213636 );
nand ( n213638 , n213611 , n213077 );
nand ( n213639 , n213637 , n213638 );
and ( n213640 , n213509 , n213399 );
not ( n213641 , n213509 );
and ( n213642 , n213641 , n213448 );
nor ( n213643 , n213640 , n213642 );
not ( n213644 , n213643 );
nand ( n213645 , n213639 , n213644 );
nand ( n213646 , n213633 , n213645 );
xor ( n213647 , n213646 , n213521 );
not ( n213648 , n213142 );
not ( n213649 , n213060 );
not ( n213650 , n213473 );
or ( n213651 , n213649 , n213650 );
nand ( n213652 , n41981 , n213147 );
nand ( n213653 , n213651 , n213652 );
not ( n213654 , n213653 );
or ( n213655 , n213648 , n213654 );
nand ( n213656 , n213539 , n213217 );
nand ( n213657 , n213655 , n213656 );
xor ( n213658 , n213647 , n213657 );
xor ( n213659 , n213646 , n213521 );
and ( n213660 , n213659 , n213657 );
and ( n213661 , n213646 , n213521 );
or ( n213662 , n213660 , n213661 );
not ( n213663 , n213173 );
not ( n213664 , n213553 );
or ( n213665 , n213663 , n213664 );
or ( n213666 , n30384 , n213381 );
nand ( n213667 , n30384 , n213381 );
nand ( n213668 , n213666 , n213667 );
nand ( n213669 , n211314 , n213668 );
nand ( n213670 , n213665 , n213669 );
xor ( n213671 , n213670 , n213615 );
xor ( n213672 , n213671 , n213548 );
xor ( n213673 , n213670 , n213615 );
and ( n213674 , n213673 , n213548 );
and ( n213675 , n213670 , n213615 );
or ( n213676 , n213674 , n213675 );
xor ( n213677 , n213658 , n213563 );
xor ( n213678 , n213677 , n213672 );
xor ( n213679 , n213658 , n213563 );
and ( n213680 , n213679 , n213672 );
and ( n213681 , n213658 , n213563 );
or ( n213682 , n213680 , n213681 );
not ( n213683 , n213206 );
and ( n213684 , n213261 , n213229 );
not ( n213685 , n213261 );
and ( n213686 , n213685 , n213232 );
or ( n213687 , n213684 , n213686 );
not ( n213688 , n213687 );
or ( n213689 , n213683 , n213688 );
nand ( n213690 , n213272 , n213599 );
nand ( n213691 , n213689 , n213690 );
not ( n213692 , n213588 );
not ( n213693 , n213454 );
or ( n213694 , n213692 , n213693 );
not ( n213695 , n209360 );
not ( n213696 , n213458 );
or ( n213697 , n213695 , n213696 );
buf ( n213698 , n213166 );
nand ( n213699 , n213513 , n213698 );
nand ( n213700 , n213697 , n213699 );
nand ( n213701 , n213700 , n213463 );
nand ( n213702 , n213694 , n213701 );
xor ( n213703 , n213691 , n213702 );
and ( n213704 , n213601 , n213613 );
xor ( n213705 , n213703 , n213704 );
xor ( n213706 , n213691 , n213702 );
and ( n213707 , n213706 , n213704 );
and ( n213708 , n213691 , n213702 );
or ( n213709 , n213707 , n213708 );
not ( n213710 , n213639 );
nand ( n213711 , n213399 , n37084 );
not ( n213712 , n213711 );
not ( n213713 , n213399 );
nand ( n213714 , n213713 , n213509 );
not ( n213715 , n213714 );
or ( n213716 , n213712 , n213715 );
nand ( n213717 , n213716 , n213630 );
not ( n213718 , n213717 );
not ( n213719 , n213718 );
or ( n213720 , n213710 , n213719 );
not ( n213721 , n213347 );
buf ( n213722 , n213609 );
not ( n213723 , n213722 );
not ( n213724 , n213723 );
or ( n213725 , n213721 , n213724 );
not ( n213726 , n213622 );
nand ( n213727 , n213726 , n213188 );
nand ( n213728 , n213725 , n213727 );
nand ( n213729 , n213728 , n213644 );
nand ( n213730 , n213720 , n213729 );
not ( n213731 , n213498 );
buf ( n213732 , n213106 );
and ( n213733 , n30412 , n213732 );
not ( n213734 , n30412 );
not ( n213735 , n213732 );
and ( n213736 , n213734 , n213735 );
or ( n213737 , n213733 , n213736 );
not ( n213738 , n213737 );
or ( n213739 , n213731 , n213738 );
nand ( n213740 , n213574 , n213577 );
nand ( n213741 , n213739 , n213740 );
xor ( n213742 , n213730 , n213741 );
nor ( n213743 , n37026 , n36220 );
and ( n213744 , n213743 , n37614 );
not ( n213745 , n213743 );
and ( n213746 , n213745 , n37615 );
nor ( n213747 , n213744 , n213746 );
xnor ( n213748 , n213611 , n213747 );
buf ( n213749 , n213748 );
buf ( n213750 , n213051 );
not ( n213751 , n213750 );
nor ( n213752 , n213749 , n213751 );
xor ( n213753 , n213742 , n213752 );
xor ( n213754 , n213730 , n213741 );
and ( n213755 , n213754 , n213752 );
and ( n213756 , n213730 , n213741 );
or ( n213757 , n213755 , n213756 );
buf ( n213758 , n213076 );
not ( n213759 , n213758 );
not ( n213760 , n213653 );
or ( n213761 , n213759 , n213760 );
not ( n213762 , n213060 );
not ( n213763 , n41978 );
not ( n213764 , n213763 );
or ( n213765 , n213762 , n213764 );
nand ( n213766 , n41979 , n213147 );
nand ( n213767 , n213765 , n213766 );
nand ( n213768 , n213142 , n213767 );
nand ( n213769 , n213761 , n213768 );
xor ( n213770 , n213769 , n213619 );
xor ( n213771 , n213770 , n213705 );
xor ( n213772 , n213769 , n213619 );
and ( n213773 , n213772 , n213705 );
and ( n213774 , n213769 , n213619 );
or ( n213775 , n213773 , n213774 );
xor ( n213776 , n213662 , n213753 );
not ( n213777 , n211314 );
and ( n213778 , n30292 , n213381 );
not ( n213779 , n30292 );
and ( n213780 , n213779 , n213382 );
or ( n213781 , n213778 , n213780 );
not ( n213782 , n213781 );
or ( n213783 , n213777 , n213782 );
buf ( n213784 , n213173 );
nand ( n213785 , n213668 , n213784 );
nand ( n213786 , n213783 , n213785 );
xor ( n213787 , n213776 , n213786 );
xor ( n213788 , n213662 , n213753 );
and ( n213789 , n213788 , n213786 );
and ( n213790 , n213662 , n213753 );
or ( n213791 , n213789 , n213790 );
xor ( n213792 , n213676 , n213771 );
xor ( n213793 , n213792 , n213787 );
xor ( n213794 , n213676 , n213771 );
and ( n213795 , n213794 , n213787 );
and ( n213796 , n213676 , n213771 );
or ( n213797 , n213795 , n213796 );
not ( n213798 , n213728 );
not ( n213799 , n213718 );
or ( n213800 , n213798 , n213799 );
not ( n213801 , n213583 );
not ( n213802 , n213635 );
or ( n213803 , n213801 , n213802 );
nand ( n213804 , n213611 , n213424 );
nand ( n213805 , n213803 , n213804 );
nand ( n213806 , n213805 , n213644 );
nand ( n213807 , n213800 , n213806 );
buf ( n213808 , n213747 );
not ( n213809 , n213808 );
nand ( n213810 , n213809 , n213104 );
not ( n213811 , n213810 );
not ( n213812 , n213051 );
not ( n213813 , n213808 );
or ( n213814 , n213812 , n213813 );
buf ( n213815 , n213610 );
nand ( n213816 , n213814 , n213815 );
not ( n213817 , n213816 );
or ( n213818 , n213811 , n213817 );
not ( n213819 , n37039 );
buf ( n213820 , n213819 );
not ( n213821 , n213820 );
nand ( n213822 , n213818 , n213821 );
not ( n213823 , n213822 );
xor ( n213824 , n213807 , n213823 );
not ( n213825 , n213498 );
not ( n213826 , n213732 );
not ( n213827 , n41981 );
or ( n213828 , n213826 , n213827 );
nand ( n213829 , n213473 , n213735 );
nand ( n213830 , n213828 , n213829 );
not ( n213831 , n213830 );
or ( n213832 , n213825 , n213831 );
nand ( n213833 , n213737 , n213577 );
nand ( n213834 , n213832 , n213833 );
xor ( n213835 , n213824 , n213834 );
xor ( n213836 , n213807 , n213823 );
and ( n213837 , n213836 , n213834 );
and ( n213838 , n213807 , n213823 );
or ( n213839 , n213837 , n213838 );
not ( n213840 , n213206 );
not ( n213841 , n213261 );
not ( n213842 , n213322 );
or ( n213843 , n213841 , n213842 );
nand ( n213844 , n30498 , n213403 );
nand ( n213845 , n213843 , n213844 );
not ( n213846 , n213845 );
or ( n213847 , n213840 , n213846 );
nand ( n213848 , n213687 , n213272 );
nand ( n213849 , n213847 , n213848 );
not ( n213850 , n213700 );
not ( n213851 , n213454 );
or ( n213852 , n213850 , n213851 );
not ( n213853 , n213458 );
not ( n213854 , n213308 );
or ( n213855 , n213853 , n213854 );
not ( n213856 , n213308 );
nand ( n213857 , n213399 , n213856 );
nand ( n213858 , n213855 , n213857 );
nand ( n213859 , n213463 , n213858 );
nand ( n213860 , n213852 , n213859 );
xor ( n213861 , n213849 , n213860 );
xor ( n213862 , n213861 , n213709 );
not ( n213863 , n213142 );
buf ( n213864 , n213060 );
not ( n213865 , n213864 );
not ( n213866 , n30384 );
not ( n213867 , n213866 );
or ( n213868 , n213865 , n213867 );
buf ( n213869 , n213147 );
nand ( n213870 , n30384 , n213869 );
nand ( n213871 , n213868 , n213870 );
not ( n213872 , n213871 );
or ( n213873 , n213863 , n213872 );
buf ( n213874 , n213758 );
nand ( n213875 , n213874 , n213767 );
nand ( n213876 , n213873 , n213875 );
xor ( n213877 , n213862 , n213876 );
xor ( n213878 , n213861 , n213709 );
and ( n213879 , n213878 , n213876 );
and ( n213880 , n213861 , n213709 );
or ( n213881 , n213879 , n213880 );
not ( n213882 , n213750 );
not ( n213883 , n37039 );
not ( n213884 , n213883 );
or ( n213885 , n213882 , n213884 );
not ( n213886 , n213883 );
nand ( n213887 , n213886 , n213751 );
nand ( n213888 , n213885 , n213887 );
not ( n213889 , n213888 );
nand ( n213890 , n213883 , n213809 );
not ( n213891 , n213819 );
nand ( n213892 , n213891 , n213808 );
nand ( n213893 , n213890 , n213748 , n213892 );
not ( n213894 , n213893 );
not ( n213895 , n213894 );
or ( n213896 , n213889 , n213895 );
not ( n213897 , n213126 );
not ( n213898 , n213820 );
or ( n213899 , n213897 , n213898 );
nand ( n213900 , n213886 , n213077 );
nand ( n213901 , n213899 , n213900 );
not ( n213902 , n213749 );
nand ( n213903 , n213901 , n213902 );
nand ( n213904 , n213896 , n213903 );
xor ( n213905 , n213904 , n213757 );
xor ( n213906 , n213905 , n213835 );
xor ( n213907 , n213904 , n213757 );
and ( n213908 , n213907 , n213835 );
and ( n213909 , n213904 , n213757 );
or ( n213910 , n213908 , n213909 );
not ( n213911 , n211314 );
not ( n213912 , n213911 );
not ( n213913 , n213912 );
not ( n213914 , n213382 );
not ( n213915 , n209248 );
or ( n213916 , n213914 , n213915 );
not ( n213917 , n41966 );
not ( n213918 , n213917 );
nand ( n213919 , n213918 , n213381 );
nand ( n213920 , n213916 , n213919 );
not ( n213921 , n213920 );
or ( n213922 , n213913 , n213921 );
nand ( n213923 , n213781 , n213784 );
nand ( n213924 , n213922 , n213923 );
xor ( n213925 , n213924 , n213877 );
xor ( n213926 , n213925 , n213775 );
xor ( n213927 , n213924 , n213877 );
and ( n213928 , n213927 , n213775 );
and ( n213929 , n213924 , n213877 );
or ( n213930 , n213928 , n213929 );
xor ( n213931 , n213906 , n213791 );
xor ( n213932 , n213931 , n213926 );
xor ( n213933 , n213906 , n213791 );
and ( n213934 , n213933 , n213926 );
and ( n213935 , n213906 , n213791 );
or ( n213936 , n213934 , n213935 );
not ( n213937 , n213858 );
not ( n213938 , n213454 );
or ( n213939 , n213937 , n213938 );
not ( n213940 , n213232 );
not ( n213941 , n213448 );
or ( n213942 , n213940 , n213941 );
nand ( n213943 , n213513 , n213229 );
nand ( n213944 , n213942 , n213943 );
nand ( n213945 , n213944 , n213463 );
nand ( n213946 , n213939 , n213945 );
not ( n213947 , n213805 );
not ( n213948 , n213631 );
or ( n213949 , n213947 , n213948 );
not ( n213950 , n209360 );
buf ( n213951 , n213610 );
not ( n213952 , n213951 );
or ( n213953 , n213950 , n213952 );
nand ( n213954 , n213611 , n213698 );
nand ( n213955 , n213953 , n213954 );
nand ( n213956 , n213955 , n213644 );
nand ( n213957 , n213949 , n213956 );
xor ( n213958 , n213946 , n213957 );
not ( n213959 , n213206 );
buf ( n213960 , n213261 );
not ( n213961 , n213960 );
not ( n213962 , n213384 );
or ( n213963 , n213961 , n213962 );
not ( n213964 , n213261 );
nand ( n213965 , n30412 , n213964 );
nand ( n213966 , n213963 , n213965 );
not ( n213967 , n213966 );
or ( n213968 , n213959 , n213967 );
nand ( n213969 , n213845 , n213272 );
nand ( n213970 , n213968 , n213969 );
xor ( n213971 , n213958 , n213970 );
xor ( n213972 , n213946 , n213957 );
and ( n213973 , n213972 , n213970 );
and ( n213974 , n213946 , n213957 );
or ( n213975 , n213973 , n213974 );
not ( n213976 , n37039 );
and ( n213977 , n37072 , n213976 );
not ( n213978 , n37072 );
and ( n213979 , n213978 , n213891 );
nor ( n213980 , n213977 , n213979 );
nor ( n213981 , n213980 , n213104 );
and ( n213982 , n213860 , n213849 );
xor ( n213983 , n213981 , n213982 );
not ( n213984 , n213577 );
not ( n213985 , n213830 );
or ( n213986 , n213984 , n213985 );
not ( n213987 , n213735 );
not ( n213988 , n213763 );
or ( n213989 , n213987 , n213988 );
nand ( n213990 , n41978 , n213732 );
nand ( n213991 , n213989 , n213990 );
nand ( n213992 , n213991 , n213498 );
nand ( n213993 , n213986 , n213992 );
xor ( n213994 , n213983 , n213993 );
xor ( n213995 , n213981 , n213982 );
and ( n213996 , n213995 , n213993 );
and ( n213997 , n213981 , n213982 );
or ( n213998 , n213996 , n213997 );
not ( n213999 , n213901 );
and ( n214000 , n213890 , n213892 , n213748 );
not ( n214001 , n214000 );
or ( n214002 , n213999 , n214001 );
not ( n214003 , n213347 );
not ( n214004 , n213976 );
or ( n214005 , n214003 , n214004 );
nand ( n214006 , n213886 , n213188 );
nand ( n214007 , n214005 , n214006 );
nand ( n214008 , n214007 , n213902 );
nand ( n214009 , n214002 , n214008 );
xor ( n214010 , n214009 , n213971 );
not ( n214011 , n213142 );
and ( n214012 , n30292 , n213869 );
not ( n214013 , n30292 );
and ( n214014 , n214013 , n213864 );
or ( n214015 , n214012 , n214014 );
not ( n214016 , n214015 );
or ( n214017 , n214011 , n214016 );
nand ( n214018 , n213871 , n213758 );
nand ( n214019 , n214017 , n214018 );
xor ( n214020 , n214010 , n214019 );
xor ( n214021 , n214009 , n213971 );
and ( n214022 , n214021 , n214019 );
and ( n214023 , n214009 , n213971 );
or ( n214024 , n214022 , n214023 );
not ( n214025 , n213784 );
not ( n214026 , n213920 );
or ( n214027 , n214025 , n214026 );
not ( n214028 , n213382 );
not ( n214029 , n41894 );
not ( n214030 , n214029 );
or ( n214031 , n214028 , n214030 );
nand ( n214032 , n41894 , n213381 );
nand ( n214033 , n214031 , n214032 );
nand ( n214034 , n214033 , n213912 );
nand ( n214035 , n214027 , n214034 );
xor ( n214036 , n213839 , n214035 );
xor ( n214037 , n214036 , n213994 );
xor ( n214038 , n213839 , n214035 );
and ( n214039 , n214038 , n213994 );
and ( n214040 , n213839 , n214035 );
or ( n214041 , n214039 , n214040 );
xor ( n214042 , n213881 , n214020 );
xor ( n214043 , n214042 , n213910 );
xor ( n214044 , n213881 , n214020 );
and ( n214045 , n214044 , n213910 );
and ( n214046 , n213881 , n214020 );
or ( n214047 , n214045 , n214046 );
xor ( n214048 , n213930 , n214037 );
xor ( n214049 , n214048 , n214043 );
xor ( n214050 , n213930 , n214037 );
and ( n214051 , n214050 , n214043 );
and ( n214052 , n213930 , n214037 );
or ( n214053 , n214051 , n214052 );
or ( n214054 , n37026 , n36220 );
and ( n214055 , n214054 , n37700 );
not ( n214056 , n37065 );
not ( n214057 , n36238 );
or ( n214058 , n214056 , n214057 );
nand ( n214059 , n214058 , n37066 );
nor ( n214060 , n214055 , n214059 );
nand ( n214061 , n36226 , n36242 );
nor ( n214062 , n214060 , n214061 );
not ( n214063 , n214062 );
nand ( n214064 , n214054 , n37700 );
not ( n214065 , n214059 );
nand ( n214066 , n214064 , n214065 , n214061 );
nand ( n214067 , n214063 , n214066 );
not ( n214068 , n214067 );
not ( n214069 , n37072 );
nand ( n214070 , n214069 , n213104 );
not ( n214071 , n213051 );
not ( n214072 , n37072 );
or ( n214073 , n214071 , n214072 );
nand ( n214074 , n214073 , n213976 );
nand ( n214075 , n214070 , n214074 );
and ( n214076 , n214068 , n214075 );
not ( n214077 , n213206 );
not ( n214078 , n213960 );
not ( n214079 , n213473 );
or ( n214080 , n214078 , n214079 );
nand ( n214081 , n41981 , n213964 );
nand ( n214082 , n214080 , n214081 );
not ( n214083 , n214082 );
or ( n214084 , n214077 , n214083 );
not ( n214085 , n213272 );
not ( n214086 , n214085 );
nand ( n214087 , n213966 , n214086 );
nand ( n214088 , n214084 , n214087 );
xor ( n214089 , n214076 , n214088 );
not ( n214090 , n213944 );
not ( n214091 , n213454 );
or ( n214092 , n214090 , n214091 );
not ( n214093 , n209264 );
not ( n214094 , n213448 );
or ( n214095 , n214093 , n214094 );
nand ( n214096 , n213399 , n213322 );
nand ( n214097 , n214095 , n214096 );
nand ( n214098 , n214097 , n213463 );
nand ( n214099 , n214092 , n214098 );
not ( n214100 , n213955 );
not ( n214101 , n213631 );
or ( n214102 , n214100 , n214101 );
not ( n214103 , n213308 );
not ( n214104 , n213951 );
or ( n214105 , n214103 , n214104 );
nand ( n214106 , n213722 , n213856 );
nand ( n214107 , n214105 , n214106 );
nand ( n214108 , n214107 , n213644 );
nand ( n214109 , n214102 , n214108 );
xor ( n214110 , n214099 , n214109 );
xor ( n214111 , n214089 , n214110 );
xor ( n214112 , n214076 , n214088 );
and ( n214113 , n214112 , n214110 );
and ( n214114 , n214076 , n214088 );
or ( n214115 , n214113 , n214114 );
not ( n214116 , n213498 );
not ( n214117 , n213735 );
not ( n214118 , n213866 );
or ( n214119 , n214117 , n214118 );
nand ( n214120 , n30384 , n213732 );
nand ( n214121 , n214119 , n214120 );
not ( n214122 , n214121 );
or ( n214123 , n214116 , n214122 );
nand ( n214124 , n213991 , n213577 );
nand ( n214125 , n214123 , n214124 );
not ( n214126 , n214007 );
not ( n214127 , n214000 );
or ( n214128 , n214126 , n214127 );
not ( n214129 , n213583 );
not ( n214130 , n213976 );
not ( n214131 , n214130 );
not ( n214132 , n214131 );
or ( n214133 , n214129 , n214132 );
not ( n214134 , n213583 );
nand ( n214135 , n213886 , n214134 );
nand ( n214136 , n214133 , n214135 );
nand ( n214137 , n214136 , n213902 );
nand ( n214138 , n214128 , n214137 );
xor ( n214139 , n214125 , n214138 );
and ( n214140 , n213051 , n214067 );
not ( n214141 , n213051 );
not ( n214142 , n214062 );
nand ( n214143 , n214142 , n214066 );
not ( n214144 , n214143 );
buf ( n214145 , n214144 );
and ( n214146 , n214141 , n214145 );
or ( n214147 , n214140 , n214146 );
not ( n214148 , n214147 );
not ( n214149 , n214143 );
not ( n214150 , n37072 );
or ( n214151 , n214149 , n214150 );
nand ( n214152 , n214144 , n214069 );
nand ( n214153 , n214151 , n214152 );
buf ( n214154 , n213980 );
nand ( n214155 , n214153 , n214154 );
not ( n214156 , n214155 );
not ( n214157 , n214156 );
or ( n214158 , n214148 , n214157 );
not ( n214159 , n213126 );
not ( n214160 , n214143 );
or ( n214161 , n214159 , n214160 );
nand ( n214162 , n214068 , n213077 );
nand ( n214163 , n214161 , n214162 );
not ( n214164 , n214154 );
nand ( n214165 , n214163 , n214164 );
nand ( n214166 , n214158 , n214165 );
xor ( n214167 , n214139 , n214166 );
xor ( n214168 , n214125 , n214138 );
and ( n214169 , n214168 , n214166 );
and ( n214170 , n214125 , n214138 );
or ( n214171 , n214169 , n214170 );
xor ( n214172 , n213975 , n213998 );
xor ( n214173 , n214172 , n214111 );
xor ( n214174 , n213975 , n213998 );
and ( n214175 , n214174 , n214111 );
and ( n214176 , n213975 , n213998 );
or ( n214177 , n214175 , n214176 );
not ( n214178 , n213142 );
not ( n214179 , n213864 );
not ( n214180 , n213917 );
or ( n214181 , n214179 , n214180 );
nand ( n214182 , n41966 , n213869 );
nand ( n214183 , n214181 , n214182 );
not ( n214184 , n214183 );
or ( n214185 , n214178 , n214184 );
nand ( n214186 , n214015 , n213758 );
nand ( n214187 , n214185 , n214186 );
not ( n214188 , n213912 );
not ( n214189 , n213382 );
not ( n214190 , n209110 );
not ( n214191 , n214190 );
or ( n214192 , n214189 , n214191 );
nand ( n214193 , n209110 , n213381 );
nand ( n214194 , n214192 , n214193 );
not ( n214195 , n214194 );
or ( n214196 , n214188 , n214195 );
nand ( n214197 , n214033 , n213784 );
nand ( n214198 , n214196 , n214197 );
xor ( n214199 , n214187 , n214198 );
xor ( n214200 , n214199 , n214167 );
xor ( n214201 , n214187 , n214198 );
and ( n214202 , n214201 , n214167 );
and ( n214203 , n214187 , n214198 );
or ( n214204 , n214202 , n214203 );
xor ( n214205 , n214024 , n214173 );
xor ( n214206 , n214205 , n214041 );
xor ( n214207 , n214024 , n214173 );
and ( n214208 , n214207 , n214041 );
and ( n214209 , n214024 , n214173 );
or ( n214210 , n214208 , n214209 );
xor ( n214211 , n214047 , n214200 );
xor ( n214212 , n214211 , n214206 );
xor ( n214213 , n214047 , n214200 );
and ( n214214 , n214213 , n214206 );
and ( n214215 , n214047 , n214200 );
or ( n214216 , n214214 , n214215 );
not ( n214217 , n214107 );
not ( n214218 , n213631 );
or ( n214219 , n214217 , n214218 );
not ( n214220 , n213232 );
not ( n214221 , n213723 );
or ( n214222 , n214220 , n214221 );
nand ( n214223 , n213722 , n213229 );
nand ( n214224 , n214222 , n214223 );
nand ( n214225 , n214224 , n213644 );
nand ( n214226 , n214219 , n214225 );
not ( n214227 , n213463 );
not ( n214228 , n213399 );
not ( n214229 , n213384 );
or ( n214230 , n214228 , n214229 );
nand ( n214231 , n30412 , n213448 );
nand ( n214232 , n214230 , n214231 );
not ( n214233 , n214232 );
or ( n214234 , n214227 , n214233 );
buf ( n214235 , n213454 );
nand ( n214236 , n214235 , n214097 );
nand ( n214237 , n214234 , n214236 );
xor ( n214238 , n214226 , n214237 );
not ( n214239 , n213206 );
not ( n214240 , n213960 );
not ( n214241 , n213763 );
or ( n214242 , n214240 , n214241 );
nand ( n214243 , n41978 , n213964 );
nand ( n214244 , n214242 , n214243 );
not ( n214245 , n214244 );
or ( n214246 , n214239 , n214245 );
nand ( n214247 , n214082 , n214086 );
nand ( n214248 , n214246 , n214247 );
xor ( n214249 , n214238 , n214248 );
xor ( n214250 , n214226 , n214237 );
and ( n214251 , n214250 , n214248 );
and ( n214252 , n214226 , n214237 );
or ( n214253 , n214251 , n214252 );
and ( n214254 , n214099 , n214109 );
not ( n214255 , n214136 );
not ( n214256 , n214000 );
or ( n214257 , n214255 , n214256 );
not ( n214258 , n209360 );
not ( n214259 , n213820 );
or ( n214260 , n214258 , n214259 );
nand ( n214261 , n214130 , n213166 );
nand ( n214262 , n214260 , n214261 );
nand ( n214263 , n214262 , n213902 );
nand ( n214264 , n214257 , n214263 );
xor ( n214265 , n214254 , n214264 );
not ( n214266 , n213347 );
not ( n214267 , n214143 );
or ( n214268 , n214266 , n214267 );
nand ( n214269 , n214068 , n213188 );
nand ( n214270 , n214268 , n214269 );
not ( n214271 , n214270 );
not ( n214272 , n214164 );
or ( n214273 , n214271 , n214272 );
nand ( n214274 , n214156 , n214163 );
nand ( n214275 , n214273 , n214274 );
xor ( n214276 , n214265 , n214275 );
xor ( n214277 , n214254 , n214264 );
and ( n214278 , n214277 , n214275 );
and ( n214279 , n214254 , n214264 );
or ( n214280 , n214278 , n214279 );
not ( n214281 , n37046 );
and ( n214282 , n214067 , n214281 );
not ( n214283 , n214067 );
and ( n214284 , n214283 , n37046 );
nor ( n214285 , n214282 , n214284 );
and ( n214286 , n214285 , n213750 );
not ( n214287 , n213498 );
and ( n214288 , n30292 , n213732 );
not ( n214289 , n30292 );
and ( n214290 , n214289 , n213735 );
or ( n214291 , n214288 , n214290 );
not ( n214292 , n214291 );
or ( n214293 , n214287 , n214292 );
nand ( n214294 , n214121 , n213577 );
nand ( n214295 , n214293 , n214294 );
xor ( n214296 , n214286 , n214295 );
xor ( n214297 , n214296 , n214115 );
xor ( n214298 , n214286 , n214295 );
and ( n214299 , n214298 , n214115 );
and ( n214300 , n214286 , n214295 );
or ( n214301 , n214299 , n214300 );
not ( n214302 , n213142 );
not ( n214303 , n213864 );
not ( n214304 , n41894 );
not ( n214305 , n214304 );
or ( n214306 , n214303 , n214305 );
nand ( n214307 , n41894 , n213869 );
nand ( n214308 , n214306 , n214307 );
not ( n214309 , n214308 );
or ( n214310 , n214302 , n214309 );
nand ( n214311 , n214183 , n213758 );
nand ( n214312 , n214310 , n214311 );
xor ( n214313 , n214249 , n214312 );
xor ( n214314 , n214313 , n214171 );
xor ( n214315 , n214249 , n214312 );
and ( n214316 , n214315 , n214171 );
and ( n214317 , n214249 , n214312 );
or ( n214318 , n214316 , n214317 );
buf ( n214319 , n211314 );
not ( n214320 , n214319 );
xor ( n214321 , n213382 , n30997 );
not ( n214322 , n214321 );
or ( n214323 , n214320 , n214322 );
nand ( n214324 , n214194 , n213784 );
nand ( n214325 , n214323 , n214324 );
xor ( n214326 , n214276 , n214325 );
xor ( n214327 , n214326 , n214177 );
xor ( n214328 , n214276 , n214325 );
and ( n214329 , n214328 , n214177 );
and ( n214330 , n214276 , n214325 );
or ( n214331 , n214329 , n214330 );
xor ( n214332 , n214297 , n214204 );
xor ( n214333 , n214332 , n214314 );
xor ( n214334 , n214297 , n214204 );
and ( n214335 , n214334 , n214314 );
and ( n214336 , n214297 , n214204 );
or ( n214337 , n214335 , n214336 );
xor ( n214338 , n214210 , n214327 );
xor ( n214339 , n214338 , n214333 );
xor ( n214340 , n214210 , n214327 );
and ( n214341 , n214340 , n214333 );
and ( n214342 , n214210 , n214327 );
or ( n214343 , n214341 , n214342 );
not ( n214344 , n213206 );
not ( n214345 , n213960 );
not ( n214346 , n213866 );
or ( n214347 , n214345 , n214346 );
nand ( n214348 , n30384 , n213964 );
nand ( n214349 , n214347 , n214348 );
not ( n214350 , n214349 );
or ( n214351 , n214344 , n214350 );
nand ( n214352 , n214244 , n214086 );
nand ( n214353 , n214351 , n214352 );
not ( n214354 , n214262 );
not ( n214355 , n213894 );
or ( n214356 , n214354 , n214355 );
buf ( n214357 , n213308 );
xnor ( n214358 , n214357 , n213820 );
nand ( n214359 , n214358 , n213902 );
nand ( n214360 , n214356 , n214359 );
xor ( n214361 , n214353 , n214360 );
not ( n214362 , n214270 );
not ( n214363 , n214156 );
or ( n214364 , n214362 , n214363 );
not ( n214365 , n213583 );
not ( n214366 , n214067 );
or ( n214367 , n214365 , n214366 );
nand ( n214368 , n214145 , n214134 );
nand ( n214369 , n214367 , n214368 );
not ( n214370 , n214154 );
nand ( n214371 , n214369 , n214370 );
nand ( n214372 , n214364 , n214371 );
xor ( n214373 , n214361 , n214372 );
xor ( n214374 , n214353 , n214360 );
and ( n214375 , n214374 , n214372 );
and ( n214376 , n214353 , n214360 );
or ( n214377 , n214375 , n214376 );
not ( n214378 , n213463 );
not ( n214379 , n213513 );
not ( n214380 , n213473 );
or ( n214381 , n214379 , n214380 );
nand ( n214382 , n41981 , n213458 );
nand ( n214383 , n214381 , n214382 );
not ( n214384 , n214383 );
or ( n214385 , n214378 , n214384 );
nand ( n214386 , n214232 , n214235 );
nand ( n214387 , n214385 , n214386 );
not ( n214388 , n214224 );
not ( n214389 , n213718 );
or ( n214390 , n214388 , n214389 );
not ( n214391 , n209264 );
not ( n214392 , n213622 );
or ( n214393 , n214391 , n214392 );
nand ( n214394 , n213726 , n213322 );
nand ( n214395 , n214393 , n214394 );
nand ( n214396 , n214395 , n213644 );
nand ( n214397 , n214390 , n214396 );
xor ( n214398 , n214387 , n214397 );
nand ( n214399 , n214281 , n213751 );
not ( n214400 , n214399 );
not ( n214401 , n213051 );
not ( n214402 , n37046 );
or ( n214403 , n214401 , n214402 );
buf ( n214404 , n214143 );
nand ( n214405 , n214403 , n214404 );
not ( n214406 , n214405 );
or ( n214407 , n214400 , n214406 );
not ( n214408 , n37040 );
not ( n214409 , n36268 );
or ( n214410 , n214408 , n214409 );
nand ( n214411 , n214410 , n35696 );
and ( n214412 , n214411 , n37594 );
not ( n214413 , n214411 );
and ( n214414 , n214413 , n37593 );
nor ( n214415 , n214412 , n214414 );
buf ( n214416 , n214415 );
not ( n214417 , n214416 );
not ( n214418 , n214417 );
nand ( n214419 , n214407 , n214418 );
not ( n214420 , n214419 );
xor ( n214421 , n214398 , n214420 );
xor ( n214422 , n214421 , n214253 );
xor ( n214423 , n214398 , n214420 );
and ( n214424 , n214423 , n214253 );
and ( n214425 , n214398 , n214420 );
or ( n214426 , n214424 , n214425 );
not ( n214427 , n213498 );
not ( n214428 , n213735 );
not ( n214429 , n213917 );
or ( n214430 , n214428 , n214429 );
nand ( n214431 , n41972 , n213732 );
nand ( n214432 , n214430 , n214431 );
not ( n214433 , n214432 );
or ( n214434 , n214427 , n214433 );
nand ( n214435 , n214291 , n213577 );
nand ( n214436 , n214434 , n214435 );
not ( n214437 , n213750 );
not ( n214438 , n214417 );
or ( n214439 , n214437 , n214438 );
nand ( n214440 , n214418 , n213751 );
nand ( n214441 , n214439 , n214440 );
not ( n214442 , n214441 );
and ( n214443 , n214416 , n37046 );
not ( n214444 , n214416 );
and ( n214445 , n214444 , n214281 );
nor ( n214446 , n214443 , n214445 );
not ( n214447 , n214285 );
nand ( n214448 , n214446 , n214447 );
not ( n214449 , n214448 );
not ( n214450 , n214449 );
or ( n214451 , n214442 , n214450 );
not ( n214452 , n213126 );
not ( n214453 , n214417 );
or ( n214454 , n214452 , n214453 );
nand ( n214455 , n214418 , n213077 );
nand ( n214456 , n214454 , n214455 );
not ( n214457 , n214447 );
buf ( n214458 , n214457 );
nand ( n214459 , n214456 , n214458 );
nand ( n214460 , n214451 , n214459 );
xor ( n214461 , n214436 , n214460 );
not ( n214462 , n213142 );
not ( n214463 , n213864 );
not ( n214464 , n41834 );
not ( n214465 , n214464 );
or ( n214466 , n214463 , n214465 );
not ( n214467 , n209110 );
not ( n214468 , n214467 );
nand ( n214469 , n214468 , n213869 );
nand ( n214470 , n214466 , n214469 );
not ( n214471 , n214470 );
or ( n214472 , n214462 , n214471 );
nand ( n214473 , n214308 , n213758 );
nand ( n214474 , n214472 , n214473 );
xor ( n214475 , n214461 , n214474 );
xor ( n214476 , n214436 , n214460 );
and ( n214477 , n214476 , n214474 );
and ( n214478 , n214436 , n214460 );
or ( n214479 , n214477 , n214478 );
xor ( n214480 , n214280 , n214373 );
xor ( n214481 , n214480 , n214422 );
xor ( n214482 , n214280 , n214373 );
and ( n214483 , n214482 , n214422 );
and ( n214484 , n214280 , n214373 );
or ( n214485 , n214483 , n214484 );
not ( n214486 , n213912 );
not ( n214487 , n213382 );
not ( n214488 , n41725 );
not ( n214489 , n214488 );
or ( n214490 , n214487 , n214489 );
nand ( n214491 , n41725 , n213381 );
nand ( n214492 , n214490 , n214491 );
not ( n214493 , n214492 );
or ( n214494 , n214486 , n214493 );
nand ( n214495 , n214321 , n213784 );
nand ( n214496 , n214494 , n214495 );
xor ( n214497 , n214301 , n214496 );
xor ( n214498 , n214497 , n214318 );
xor ( n214499 , n214301 , n214496 );
and ( n214500 , n214499 , n214318 );
and ( n214501 , n214301 , n214496 );
or ( n214502 , n214500 , n214501 );
xor ( n214503 , n214481 , n214475 );
xor ( n214504 , n214503 , n214331 );
xor ( n214505 , n214481 , n214475 );
and ( n214506 , n214505 , n214331 );
and ( n214507 , n214481 , n214475 );
or ( n214508 , n214506 , n214507 );
xor ( n214509 , n214337 , n214498 );
xor ( n214510 , n214509 , n214504 );
xor ( n214511 , n214337 , n214498 );
and ( n214512 , n214511 , n214504 );
and ( n214513 , n214337 , n214498 );
or ( n214514 , n214512 , n214513 );
not ( n214515 , n213644 );
and ( n214516 , n30412 , n213951 );
not ( n214517 , n30412 );
and ( n214518 , n214517 , n213722 );
or ( n214519 , n214516 , n214518 );
not ( n214520 , n214519 );
or ( n214521 , n214515 , n214520 );
nand ( n214522 , n214395 , n213718 );
nand ( n214523 , n214521 , n214522 );
not ( n214524 , n214235 );
not ( n214525 , n214383 );
or ( n214526 , n214524 , n214525 );
and ( n214527 , n41978 , n213458 );
not ( n214528 , n41978 );
and ( n214529 , n214528 , n213513 );
or ( n214530 , n214527 , n214529 );
nand ( n214531 , n214530 , n213463 );
nand ( n214532 , n214526 , n214531 );
xor ( n214533 , n214523 , n214532 );
not ( n214534 , n214358 );
not ( n214535 , n214000 );
or ( n214536 , n214534 , n214535 );
buf ( n214537 , n213232 );
and ( n214538 , n214537 , n213820 );
not ( n214539 , n214537 );
and ( n214540 , n214539 , n213886 );
or ( n214541 , n214538 , n214540 );
nand ( n214542 , n214541 , n213902 );
nand ( n214543 , n214536 , n214542 );
xor ( n214544 , n214533 , n214543 );
xor ( n214545 , n214523 , n214532 );
and ( n214546 , n214545 , n214543 );
and ( n214547 , n214523 , n214532 );
or ( n214548 , n214546 , n214547 );
not ( n214549 , n214369 );
nand ( n214550 , n214153 , n214154 );
not ( n214551 , n214550 );
not ( n214552 , n214551 );
or ( n214553 , n214549 , n214552 );
not ( n214554 , n209360 );
not ( n214555 , n214404 );
or ( n214556 , n214554 , n214555 );
nand ( n214557 , n214145 , n213166 );
nand ( n214558 , n214556 , n214557 );
nand ( n214559 , n214558 , n214370 );
nand ( n214560 , n214553 , n214559 );
and ( n214561 , n214387 , n214397 );
xor ( n214562 , n214560 , n214561 );
not ( n214563 , n213206 );
not ( n214564 , n214563 );
not ( n214565 , n214564 );
not ( n214566 , n213960 );
not ( n214567 , n30292 );
not ( n214568 , n214567 );
or ( n214569 , n214566 , n214568 );
not ( n214570 , n213960 );
nand ( n214571 , n30292 , n214570 );
nand ( n214572 , n214569 , n214571 );
not ( n214573 , n214572 );
or ( n214574 , n214565 , n214573 );
nand ( n214575 , n214349 , n214086 );
nand ( n214576 , n214574 , n214575 );
xor ( n214577 , n214562 , n214576 );
xor ( n214578 , n214560 , n214561 );
and ( n214579 , n214578 , n214576 );
and ( n214580 , n214560 , n214561 );
or ( n214581 , n214579 , n214580 );
not ( n214582 , n214416 );
not ( n214583 , n36971 );
not ( n214584 , n214583 );
or ( n214585 , n214582 , n214584 );
not ( n214586 , n214416 );
nand ( n214587 , n36971 , n214586 );
nand ( n214588 , n214585 , n214587 );
and ( n214589 , n214588 , n213750 );
xor ( n214590 , n214544 , n214589 );
not ( n214591 , n213577 );
not ( n214592 , n214432 );
or ( n214593 , n214591 , n214592 );
not ( n214594 , n213735 );
not ( n214595 , n214029 );
or ( n214596 , n214594 , n214595 );
not ( n214597 , n41894 );
not ( n214598 , n214597 );
nand ( n214599 , n214598 , n213732 );
nand ( n214600 , n214596 , n214599 );
nand ( n214601 , n214600 , n213498 );
nand ( n214602 , n214593 , n214601 );
xor ( n214603 , n214590 , n214602 );
xor ( n214604 , n214544 , n214589 );
and ( n214605 , n214604 , n214602 );
and ( n214606 , n214544 , n214589 );
or ( n214607 , n214605 , n214606 );
not ( n214608 , n214456 );
buf ( n214609 , n214448 );
not ( n214610 , n214609 );
not ( n214611 , n214610 );
or ( n214612 , n214608 , n214611 );
not ( n214613 , n213347 );
not ( n214614 , n214417 );
or ( n214615 , n214613 , n214614 );
not ( n214616 , n213347 );
nand ( n214617 , n214418 , n214616 );
nand ( n214618 , n214615 , n214617 );
nand ( n214619 , n214618 , n214458 );
nand ( n214620 , n214612 , n214619 );
xor ( n214621 , n214620 , n214377 );
xor ( n214622 , n214621 , n214426 );
xor ( n214623 , n214620 , n214377 );
and ( n214624 , n214623 , n214426 );
and ( n214625 , n214620 , n214377 );
or ( n214626 , n214624 , n214625 );
not ( n214627 , n213142 );
not ( n214628 , n30997 );
and ( n214629 , n213869 , n214628 );
not ( n214630 , n213869 );
and ( n214631 , n214630 , n30997 );
nor ( n214632 , n214629 , n214631 );
not ( n214633 , n214632 );
or ( n214634 , n214627 , n214633 );
nand ( n214635 , n213758 , n214470 );
nand ( n214636 , n214634 , n214635 );
xor ( n214637 , n214577 , n214636 );
not ( n214638 , n213784 );
not ( n214639 , n214492 );
or ( n214640 , n214638 , n214639 );
not ( n214641 , n213382 );
not ( n214642 , n41716 );
not ( n214643 , n214642 );
or ( n214644 , n214641 , n214643 );
nand ( n214645 , n41716 , n213381 );
nand ( n214646 , n214644 , n214645 );
nand ( n214647 , n214646 , n213912 );
nand ( n214648 , n214640 , n214647 );
xor ( n214649 , n214637 , n214648 );
xor ( n214650 , n214577 , n214636 );
and ( n214651 , n214650 , n214648 );
and ( n214652 , n214577 , n214636 );
or ( n214653 , n214651 , n214652 );
xor ( n214654 , n214479 , n214603 );
xor ( n214655 , n214654 , n214622 );
xor ( n214656 , n214479 , n214603 );
and ( n214657 , n214656 , n214622 );
and ( n214658 , n214479 , n214603 );
or ( n214659 , n214657 , n214658 );
xor ( n214660 , n214485 , n214649 );
xor ( n214661 , n214660 , n214502 );
xor ( n214662 , n214485 , n214649 );
and ( n214663 , n214662 , n214502 );
and ( n214664 , n214485 , n214649 );
or ( n214665 , n214663 , n214664 );
xor ( n214666 , n214655 , n214508 );
xor ( n214667 , n214666 , n214661 );
xor ( n214668 , n214655 , n214508 );
and ( n214669 , n214668 , n214661 );
and ( n214670 , n214655 , n214508 );
or ( n214671 , n214669 , n214670 );
not ( n214672 , n214541 );
not ( n214673 , n213894 );
or ( n214674 , n214672 , n214673 );
not ( n214675 , n209264 );
not ( n214676 , n213820 );
or ( n214677 , n214675 , n214676 );
not ( n214678 , n209264 );
nand ( n214679 , n213886 , n214678 );
nand ( n214680 , n214677 , n214679 );
nand ( n214681 , n214680 , n213902 );
nand ( n214682 , n214674 , n214681 );
not ( n214683 , n214558 );
not ( n214684 , n214551 );
or ( n214685 , n214683 , n214684 );
and ( n214686 , n214357 , n214404 );
not ( n214687 , n214357 );
not ( n214688 , n214404 );
and ( n214689 , n214687 , n214688 );
or ( n214690 , n214686 , n214689 );
nand ( n214691 , n214690 , n214164 );
nand ( n214692 , n214685 , n214691 );
xor ( n214693 , n214682 , n214692 );
buf ( n214694 , n213644 );
not ( n214695 , n214694 );
not ( n214696 , n213722 );
not ( n214697 , n213473 );
or ( n214698 , n214696 , n214697 );
not ( n214699 , n41981 );
not ( n214700 , n214699 );
buf ( n214701 , n213635 );
nand ( n214702 , n214700 , n214701 );
nand ( n214703 , n214698 , n214702 );
not ( n214704 , n214703 );
or ( n214705 , n214695 , n214704 );
nand ( n214706 , n214519 , n213718 );
nand ( n214707 , n214705 , n214706 );
not ( n214708 , n213463 );
not ( n214709 , n213399 );
not ( n214710 , n213866 );
or ( n214711 , n214709 , n214710 );
not ( n214712 , n213399 );
nand ( n214713 , n30384 , n214712 );
nand ( n214714 , n214711 , n214713 );
not ( n214715 , n214714 );
or ( n214716 , n214708 , n214715 );
buf ( n214717 , n214235 );
nand ( n214718 , n214530 , n214717 );
nand ( n214719 , n214716 , n214718 );
xor ( n214720 , n214707 , n214719 );
xor ( n214721 , n214693 , n214720 );
xor ( n214722 , n214682 , n214692 );
and ( n214723 , n214722 , n214720 );
and ( n214724 , n214682 , n214692 );
or ( n214725 , n214723 , n214724 );
not ( n214726 , n214564 );
not ( n214727 , n213960 );
not ( n214728 , n209248 );
or ( n214729 , n214727 , n214728 );
nand ( n214730 , n213918 , n214570 );
nand ( n214731 , n214729 , n214730 );
not ( n214732 , n214731 );
or ( n214733 , n214726 , n214732 );
nand ( n214734 , n214572 , n214086 );
nand ( n214735 , n214733 , n214734 );
not ( n214736 , n214583 );
nand ( n214737 , n214736 , n213750 );
not ( n214738 , n214737 );
not ( n214739 , n214417 );
or ( n214740 , n214738 , n214739 );
nand ( n214741 , n214583 , n213751 );
nand ( n214742 , n214740 , n214741 );
and ( n214743 , n37055 , n37621 );
not ( n214744 , n37055 );
and ( n214745 , n214744 , n37622 );
nor ( n214746 , n214743 , n214745 );
buf ( n214747 , n214746 );
and ( n214748 , n214742 , n214747 );
xor ( n214749 , n214735 , n214748 );
xor ( n214750 , n214749 , n214548 );
xor ( n214751 , n214735 , n214748 );
and ( n214752 , n214751 , n214548 );
and ( n214753 , n214735 , n214748 );
or ( n214754 , n214752 , n214753 );
not ( n214755 , n214618 );
not ( n214756 , n214610 );
or ( n214757 , n214755 , n214756 );
not ( n214758 , n213583 );
buf ( n214759 , n214416 );
not ( n214760 , n214759 );
not ( n214761 , n214760 );
or ( n214762 , n214758 , n214761 );
nand ( n214763 , n214759 , n214134 );
nand ( n214764 , n214762 , n214763 );
nand ( n214765 , n214764 , n214458 );
nand ( n214766 , n214757 , n214765 );
not ( n214767 , n213498 );
not ( n214768 , n213735 );
not ( n214769 , n214464 );
or ( n214770 , n214768 , n214769 );
or ( n214771 , n214467 , n213735 );
nand ( n214772 , n214770 , n214771 );
not ( n214773 , n214772 );
or ( n214774 , n214767 , n214773 );
nand ( n214775 , n214600 , n213577 );
nand ( n214776 , n214774 , n214775 );
xor ( n214777 , n214766 , n214776 );
xor ( n214778 , n214777 , n214721 );
xor ( n214779 , n214766 , n214776 );
and ( n214780 , n214779 , n214721 );
and ( n214781 , n214766 , n214776 );
or ( n214782 , n214780 , n214781 );
not ( n214783 , n214747 );
and ( n214784 , n213751 , n214783 );
not ( n214785 , n213751 );
buf ( n214786 , n214747 );
and ( n214787 , n214785 , n214786 );
nor ( n214788 , n214784 , n214787 );
not ( n214789 , n214788 );
and ( n214790 , n214416 , n214583 );
not ( n214791 , n214416 );
and ( n214792 , n214791 , n214736 );
nor ( n214793 , n214790 , n214792 );
not ( n214794 , n214746 );
or ( n214795 , n214736 , n214794 );
nand ( n214796 , n214794 , n36971 );
nand ( n214797 , n214795 , n214796 );
nand ( n214798 , n214793 , n214797 );
not ( n214799 , n214798 );
not ( n214800 , n214799 );
or ( n214801 , n214789 , n214800 );
not ( n214802 , n213126 );
not ( n214803 , n214747 );
not ( n214804 , n214803 );
or ( n214805 , n214802 , n214804 );
nand ( n214806 , n214786 , n213077 );
nand ( n214807 , n214805 , n214806 );
buf ( n214808 , n214588 );
nand ( n214809 , n214807 , n214808 );
nand ( n214810 , n214801 , n214809 );
xor ( n214811 , n214810 , n214581 );
xor ( n214812 , n214811 , n214607 );
xor ( n214813 , n214810 , n214581 );
and ( n214814 , n214813 , n214607 );
and ( n214815 , n214810 , n214581 );
or ( n214816 , n214814 , n214815 );
not ( n214817 , n213058 );
not ( n214818 , n213147 );
not ( n214819 , n214818 );
not ( n214820 , n31991 );
buf ( n214821 , n214820 );
not ( n214822 , n214821 );
or ( n214823 , n214819 , n214822 );
not ( n214824 , n214818 );
nand ( n214825 , n41725 , n214824 );
nand ( n214826 , n214823 , n214825 );
not ( n214827 , n214826 );
or ( n214828 , n214817 , n214827 );
nand ( n214829 , n214632 , n213758 );
nand ( n214830 , n214828 , n214829 );
xor ( n214831 , n214750 , n214830 );
not ( n214832 , n213912 );
not ( n214833 , n213382 );
not ( n214834 , n30962 );
not ( n214835 , n214834 );
or ( n214836 , n214833 , n214835 );
buf ( n214837 , n30962 );
nand ( n214838 , n214837 , n213381 );
nand ( n214839 , n214836 , n214838 );
not ( n214840 , n214839 );
or ( n214841 , n214832 , n214840 );
nand ( n214842 , n213784 , n214646 );
nand ( n214843 , n214841 , n214842 );
xor ( n214844 , n214831 , n214843 );
xor ( n214845 , n214750 , n214830 );
and ( n214846 , n214845 , n214843 );
and ( n214847 , n214750 , n214830 );
or ( n214848 , n214846 , n214847 );
xor ( n214849 , n214626 , n214778 );
xor ( n214850 , n214849 , n214812 );
xor ( n214851 , n214626 , n214778 );
and ( n214852 , n214851 , n214812 );
and ( n214853 , n214626 , n214778 );
or ( n214854 , n214852 , n214853 );
xor ( n214855 , n214653 , n214659 );
xor ( n214856 , n214855 , n214844 );
xor ( n214857 , n214653 , n214659 );
and ( n214858 , n214857 , n214844 );
and ( n214859 , n214653 , n214659 );
or ( n214860 , n214858 , n214859 );
xor ( n214861 , n214850 , n214665 );
xor ( n214862 , n214861 , n214856 );
xor ( n214863 , n214850 , n214665 );
and ( n214864 , n214863 , n214856 );
and ( n214865 , n214850 , n214665 );
or ( n214866 , n214864 , n214865 );
not ( n214867 , n213718 );
not ( n214868 , n214703 );
or ( n214869 , n214867 , n214868 );
not ( n214870 , n214701 );
not ( n214871 , n214870 );
not ( n214872 , n213763 );
or ( n214873 , n214871 , n214872 );
nand ( n214874 , n214701 , n41979 );
nand ( n214875 , n214873 , n214874 );
nand ( n214876 , n214875 , n214694 );
nand ( n214877 , n214869 , n214876 );
not ( n214878 , n214680 );
not ( n214879 , n213894 );
or ( n214880 , n214878 , n214879 );
buf ( n214881 , n30412 );
not ( n214882 , n214881 );
not ( n214883 , n213820 );
or ( n214884 , n214882 , n214883 );
not ( n214885 , n214881 );
nand ( n214886 , n213821 , n214885 );
nand ( n214887 , n214884 , n214886 );
not ( n214888 , n213749 );
nand ( n214889 , n214887 , n214888 );
nand ( n214890 , n214880 , n214889 );
xor ( n214891 , n214877 , n214890 );
not ( n214892 , n214690 );
not ( n214893 , n214550 );
not ( n214894 , n214893 );
or ( n214895 , n214892 , n214894 );
not ( n214896 , n214537 );
not ( n214897 , n214404 );
or ( n214898 , n214896 , n214897 );
not ( n214899 , n214537 );
nand ( n214900 , n214688 , n214899 );
nand ( n214901 , n214898 , n214900 );
nand ( n214902 , n214901 , n214164 );
nand ( n214903 , n214895 , n214902 );
xor ( n214904 , n214891 , n214903 );
xor ( n214905 , n214877 , n214890 );
and ( n214906 , n214905 , n214903 );
and ( n214907 , n214877 , n214890 );
or ( n214908 , n214906 , n214907 );
and ( n214909 , n214719 , n214707 );
not ( n214910 , n213463 );
not ( n214911 , n213399 );
not ( n214912 , n214567 );
or ( n214913 , n214911 , n214912 );
nand ( n214914 , n30292 , n214712 );
nand ( n214915 , n214913 , n214914 );
not ( n214916 , n214915 );
or ( n214917 , n214910 , n214916 );
nand ( n214918 , n214714 , n214717 );
nand ( n214919 , n214917 , n214918 );
xor ( n214920 , n214909 , n214919 );
not ( n214921 , n214086 );
not ( n214922 , n214731 );
or ( n214923 , n214921 , n214922 );
not ( n214924 , n213960 );
not ( n214925 , n214597 );
or ( n214926 , n214924 , n214925 );
buf ( n214927 , n41894 );
nand ( n214928 , n214927 , n214570 );
nand ( n214929 , n214926 , n214928 );
nand ( n214930 , n214564 , n214929 );
nand ( n214931 , n214923 , n214930 );
xor ( n214932 , n214920 , n214931 );
xor ( n214933 , n214909 , n214919 );
and ( n214934 , n214933 , n214931 );
and ( n214935 , n214909 , n214919 );
or ( n214936 , n214934 , n214935 );
not ( n214937 , n214746 );
and ( n214938 , n37060 , n37604 );
not ( n214939 , n37060 );
not ( n214940 , n37604 );
and ( n214941 , n214939 , n214940 );
or ( n214942 , n214938 , n214941 );
not ( n214943 , n214942 );
or ( n214944 , n214937 , n214943 );
and ( n214945 , n37060 , n37604 );
not ( n214946 , n37060 );
and ( n214947 , n214946 , n214940 );
nor ( n214948 , n214945 , n214947 );
nand ( n214949 , n214948 , n214794 );
nand ( n214950 , n214944 , n214949 );
buf ( n214951 , n214950 );
nor ( n214952 , n214951 , n213751 );
not ( n214953 , n214764 );
not ( n214954 , n214610 );
or ( n214955 , n214953 , n214954 );
buf ( n214956 , n209360 );
not ( n214957 , n214956 );
not ( n214958 , n214417 );
or ( n214959 , n214957 , n214958 );
not ( n214960 , n214956 );
nand ( n214961 , n214759 , n214960 );
nand ( n214962 , n214959 , n214961 );
nand ( n214963 , n214962 , n214458 );
nand ( n214964 , n214955 , n214963 );
xor ( n214965 , n214952 , n214964 );
xor ( n214966 , n214965 , n214904 );
xor ( n214967 , n214952 , n214964 );
and ( n214968 , n214967 , n214904 );
and ( n214969 , n214952 , n214964 );
or ( n214970 , n214968 , n214969 );
not ( n214971 , n214807 );
not ( n214972 , n214799 );
or ( n214973 , n214971 , n214972 );
not ( n214974 , n213347 );
not ( n214975 , n214783 );
or ( n214976 , n214974 , n214975 );
nand ( n214977 , n214786 , n214616 );
nand ( n214978 , n214976 , n214977 );
nand ( n214979 , n214978 , n214808 );
nand ( n214980 , n214973 , n214979 );
xor ( n214981 , n214980 , n214725 );
xor ( n214982 , n214981 , n214932 );
xor ( n214983 , n214980 , n214725 );
and ( n214984 , n214983 , n214932 );
and ( n214985 , n214980 , n214725 );
or ( n214986 , n214984 , n214985 );
not ( n214987 , n213498 );
not ( n214988 , n213735 );
not ( n214989 , n30997 );
not ( n214990 , n214989 );
or ( n214991 , n214988 , n214990 );
nand ( n214992 , n30997 , n213732 );
nand ( n214993 , n214991 , n214992 );
not ( n214994 , n214993 );
or ( n214995 , n214987 , n214994 );
nand ( n214996 , n214772 , n213577 );
nand ( n214997 , n214995 , n214996 );
xor ( n214998 , n214997 , n214754 );
not ( n214999 , n213758 );
not ( n215000 , n214826 );
or ( n215001 , n214999 , n215000 );
not ( n215002 , n214818 );
not ( n215003 , n214642 );
or ( n215004 , n215002 , n215003 );
nand ( n215005 , n41716 , n213147 );
nand ( n215006 , n215004 , n215005 );
nand ( n215007 , n215006 , n213058 );
nand ( n215008 , n215001 , n215007 );
xor ( n215009 , n214998 , n215008 );
xor ( n215010 , n214997 , n214754 );
and ( n215011 , n215010 , n215008 );
and ( n215012 , n214997 , n214754 );
or ( n215013 , n215011 , n215012 );
not ( n215014 , n213784 );
not ( n215015 , n214839 );
or ( n215016 , n215014 , n215015 );
not ( n215017 , n213382 );
not ( n215018 , n208725 );
not ( n215019 , n215018 );
or ( n215020 , n215017 , n215019 );
nand ( n215021 , n208725 , n213381 );
nand ( n215022 , n215020 , n215021 );
nand ( n215023 , n215022 , n211314 );
nand ( n215024 , n215016 , n215023 );
xor ( n215025 , n215024 , n214782 );
xor ( n215026 , n215025 , n214966 );
xor ( n215027 , n215024 , n214782 );
and ( n215028 , n215027 , n214966 );
and ( n215029 , n215024 , n214782 );
or ( n215030 , n215028 , n215029 );
xor ( n215031 , n214816 , n214982 );
xor ( n215032 , n215031 , n215009 );
xor ( n215033 , n214816 , n214982 );
and ( n215034 , n215033 , n215009 );
and ( n215035 , n214816 , n214982 );
or ( n215036 , n215034 , n215035 );
xor ( n215037 , n214848 , n215026 );
xor ( n215038 , n215037 , n214854 );
xor ( n215039 , n214848 , n215026 );
and ( n215040 , n215039 , n214854 );
and ( n215041 , n214848 , n215026 );
or ( n215042 , n215040 , n215041 );
xor ( n215043 , n215032 , n214860 );
xor ( n215044 , n215043 , n215038 );
xor ( n215045 , n215032 , n214860 );
and ( n215046 , n215045 , n215038 );
and ( n215047 , n215032 , n214860 );
or ( n215048 , n215046 , n215047 );
not ( n215049 , n214164 );
buf ( n215050 , n209264 );
not ( n215051 , n215050 );
not ( n215052 , n214404 );
or ( n215053 , n215051 , n215052 );
buf ( n215054 , n214068 );
nand ( n215055 , n215054 , n214678 );
nand ( n215056 , n215053 , n215055 );
not ( n215057 , n215056 );
or ( n215058 , n215049 , n215057 );
nand ( n215059 , n214901 , n214893 );
nand ( n215060 , n215058 , n215059 );
not ( n215061 , n214694 );
not ( n215062 , n214870 );
not ( n215063 , n213866 );
or ( n215064 , n215062 , n215063 );
nand ( n215065 , n30384 , n214701 );
nand ( n215066 , n215064 , n215065 );
not ( n215067 , n215066 );
or ( n215068 , n215061 , n215067 );
nand ( n215069 , n214875 , n213718 );
nand ( n215070 , n215068 , n215069 );
not ( n215071 , n215070 );
not ( n215072 , n214887 );
not ( n215073 , n213894 );
or ( n215074 , n215072 , n215073 );
not ( n215075 , n213473 );
not ( n215076 , n215075 );
not ( n215077 , n213820 );
or ( n215078 , n215076 , n215077 );
not ( n215079 , n213820 );
nand ( n215080 , n215079 , n214699 );
nand ( n215081 , n215078 , n215080 );
nand ( n215082 , n215081 , n214888 );
nand ( n215083 , n215074 , n215082 );
not ( n215084 , n215083 );
not ( n215085 , n215084 );
or ( n215086 , n215071 , n215085 );
or ( n215087 , n215084 , n215070 );
nand ( n215088 , n215086 , n215087 );
xor ( n215089 , n215060 , n215088 );
nand ( n215090 , n214942 , n213750 );
nand ( n215091 , n215090 , n214783 );
not ( n215092 , n213750 );
nand ( n215093 , n215092 , n214948 );
and ( n215094 , n215091 , n215093 );
buf ( n215095 , n35611 );
nand ( n215096 , n35738 , n215095 );
not ( n215097 , n215096 );
not ( n215098 , n215097 );
not ( n215099 , n37017 );
not ( n215100 , n215099 );
or ( n215101 , n215098 , n215100 );
nand ( n215102 , n37017 , n215096 );
nand ( n215103 , n215101 , n215102 );
buf ( n215104 , n215103 );
not ( n215105 , n215104 );
nor ( n215106 , n215094 , n215105 );
xor ( n215107 , n215089 , n215106 );
xor ( n215108 , n215060 , n215088 );
and ( n215109 , n215108 , n215106 );
and ( n215110 , n215060 , n215088 );
or ( n215111 , n215109 , n215110 );
not ( n215112 , n213463 );
not ( n215113 , n214712 );
not ( n215114 , n215113 );
not ( n215115 , n209248 );
or ( n215116 , n215114 , n215115 );
not ( n215117 , n213917 );
buf ( n215118 , n214712 );
nand ( n215119 , n215117 , n215118 );
nand ( n215120 , n215116 , n215119 );
not ( n215121 , n215120 );
or ( n215122 , n215112 , n215121 );
nand ( n215123 , n214915 , n214717 );
nand ( n215124 , n215122 , n215123 );
not ( n215125 , n214962 );
not ( n215126 , n214610 );
or ( n215127 , n215125 , n215126 );
not ( n215128 , n214357 );
not ( n215129 , n214417 );
or ( n215130 , n215128 , n215129 );
not ( n215131 , n214357 );
nand ( n215132 , n214418 , n215131 );
nand ( n215133 , n215130 , n215132 );
nand ( n215134 , n215133 , n214458 );
nand ( n215135 , n215127 , n215134 );
xor ( n215136 , n215124 , n215135 );
not ( n215137 , n214563 );
not ( n215138 , n215137 );
not ( n215139 , n213960 );
not ( n215140 , n214464 );
or ( n215141 , n215139 , n215140 );
nand ( n215142 , n214570 , n214468 );
nand ( n215143 , n215141 , n215142 );
not ( n215144 , n215143 );
or ( n215145 , n215138 , n215144 );
nand ( n215146 , n214929 , n214086 );
nand ( n215147 , n215145 , n215146 );
xor ( n215148 , n215136 , n215147 );
xor ( n215149 , n215124 , n215135 );
and ( n215150 , n215149 , n215147 );
and ( n215151 , n215124 , n215135 );
or ( n215152 , n215150 , n215151 );
not ( n215153 , n214978 );
not ( n215154 , n214799 );
or ( n215155 , n215153 , n215154 );
not ( n215156 , n213583 );
not ( n215157 , n214783 );
or ( n215158 , n215156 , n215157 );
nand ( n215159 , n214786 , n214134 );
nand ( n215160 , n215158 , n215159 );
nand ( n215161 , n215160 , n214808 );
nand ( n215162 , n215155 , n215161 );
xor ( n215163 , n214908 , n215162 );
not ( n215164 , n215104 );
not ( n215165 , n215164 );
and ( n215166 , n213750 , n215165 );
not ( n215167 , n213750 );
and ( n215168 , n215167 , n215164 );
nor ( n215169 , n215166 , n215168 );
not ( n215170 , n215169 );
not ( n215171 , n215097 );
not ( n215172 , n215099 );
or ( n215173 , n215171 , n215172 );
nand ( n215174 , n215173 , n215102 );
nand ( n215175 , n214948 , n215174 );
not ( n215176 , n215175 );
not ( n215177 , n215174 );
nand ( n215178 , n215177 , n214942 );
not ( n215179 , n215178 );
or ( n215180 , n215176 , n215179 );
nand ( n215181 , n215180 , n214950 );
not ( n215182 , n215181 );
buf ( n215183 , n215182 );
not ( n215184 , n215183 );
or ( n215185 , n215170 , n215184 );
not ( n215186 , n213126 );
not ( n215187 , n215164 );
or ( n215188 , n215186 , n215187 );
nand ( n215189 , n215104 , n213077 );
nand ( n215190 , n215188 , n215189 );
not ( n215191 , n214951 );
nand ( n215192 , n215190 , n215191 );
nand ( n215193 , n215185 , n215192 );
xor ( n215194 , n215163 , n215193 );
xor ( n215195 , n214908 , n215162 );
and ( n215196 , n215195 , n215193 );
and ( n215197 , n214908 , n215162 );
or ( n215198 , n215196 , n215197 );
xor ( n215199 , n215107 , n214936 );
not ( n215200 , n213758 );
not ( n215201 , n215006 );
or ( n215202 , n215200 , n215201 );
not ( n215203 , n213864 );
not ( n215204 , n214834 );
or ( n215205 , n215203 , n215204 );
nand ( n215206 , n30962 , n213869 );
nand ( n215207 , n215205 , n215206 );
nand ( n215208 , n215207 , n213058 );
nand ( n215209 , n215202 , n215208 );
xor ( n215210 , n215199 , n215209 );
xor ( n215211 , n215107 , n214936 );
and ( n215212 , n215211 , n215209 );
and ( n215213 , n215107 , n214936 );
or ( n215214 , n215212 , n215213 );
not ( n215215 , n211314 );
and ( n215216 , n41608 , n213381 );
not ( n215217 , n41608 );
and ( n215218 , n215217 , n213382 );
or ( n215219 , n215216 , n215218 );
not ( n215220 , n215219 );
or ( n215221 , n215215 , n215220 );
nand ( n215222 , n215022 , n213784 );
nand ( n215223 , n215221 , n215222 );
not ( n215224 , n213498 );
not ( n215225 , n213735 );
not ( n215226 , n214488 );
or ( n215227 , n215225 , n215226 );
not ( n215228 , n214820 );
nand ( n215229 , n215228 , n213732 );
nand ( n215230 , n215227 , n215229 );
not ( n215231 , n215230 );
or ( n215232 , n215224 , n215231 );
nand ( n215233 , n214993 , n213577 );
nand ( n215234 , n215232 , n215233 );
xor ( n215235 , n215223 , n215234 );
xor ( n215236 , n215235 , n214970 );
xor ( n215237 , n215223 , n215234 );
and ( n215238 , n215237 , n214970 );
and ( n215239 , n215223 , n215234 );
or ( n215240 , n215238 , n215239 );
xor ( n215241 , n215148 , n214986 );
xor ( n215242 , n215241 , n215194 );
xor ( n215243 , n215148 , n214986 );
and ( n215244 , n215243 , n215194 );
and ( n215245 , n215148 , n214986 );
or ( n215246 , n215244 , n215245 );
xor ( n215247 , n215013 , n215210 );
xor ( n215248 , n215247 , n215030 );
xor ( n215249 , n215013 , n215210 );
and ( n215250 , n215249 , n215030 );
and ( n215251 , n215013 , n215210 );
or ( n215252 , n215250 , n215251 );
xor ( n215253 , n215236 , n215242 );
xor ( n215254 , n215253 , n215036 );
xor ( n215255 , n215236 , n215242 );
and ( n215256 , n215255 , n215036 );
and ( n215257 , n215236 , n215242 );
or ( n215258 , n215256 , n215257 );
xor ( n215259 , n215248 , n215042 );
xor ( n215260 , n215259 , n215254 );
xor ( n215261 , n215248 , n215042 );
and ( n215262 , n215261 , n215254 );
and ( n215263 , n215248 , n215042 );
or ( n215264 , n215262 , n215263 );
not ( n215265 , n215081 );
not ( n215266 , n213894 );
or ( n215267 , n215265 , n215266 );
not ( n215268 , n213763 );
not ( n215269 , n215268 );
not ( n215270 , n213820 );
or ( n215271 , n215269 , n215270 );
not ( n215272 , n213820 );
nand ( n215273 , n215272 , n213763 );
nand ( n215274 , n215271 , n215273 );
nand ( n215275 , n215274 , n214888 );
nand ( n215276 , n215267 , n215275 );
not ( n215277 , n215056 );
not ( n215278 , n214893 );
or ( n215279 , n215277 , n215278 );
not ( n215280 , n214881 );
not ( n215281 , n214067 );
or ( n215282 , n215280 , n215281 );
nand ( n215283 , n214885 , n214144 );
nand ( n215284 , n215282 , n215283 );
nand ( n215285 , n215284 , n214164 );
nand ( n215286 , n215279 , n215285 );
xor ( n215287 , n215276 , n215286 );
not ( n215288 , n214694 );
buf ( n215289 , n213815 );
not ( n215290 , n215289 );
not ( n215291 , n215290 );
not ( n215292 , n30292 );
not ( n215293 , n215292 );
or ( n215294 , n215291 , n215293 );
nand ( n215295 , n30292 , n215289 );
nand ( n215296 , n215294 , n215295 );
not ( n215297 , n215296 );
or ( n215298 , n215288 , n215297 );
nand ( n215299 , n215066 , n213718 );
nand ( n215300 , n215298 , n215299 );
xor ( n215301 , n215287 , n215300 );
xor ( n215302 , n215276 , n215286 );
and ( n215303 , n215302 , n215300 );
and ( n215304 , n215276 , n215286 );
or ( n215305 , n215303 , n215304 );
not ( n215306 , n215070 );
nor ( n215307 , n215306 , n215084 );
not ( n215308 , n215103 );
not ( n215309 , n215308 );
not ( n215310 , n36659 );
not ( n215311 , n35759 );
nor ( n215312 , n215311 , n36652 );
not ( n215313 , n215312 );
or ( n215314 , n215310 , n215313 );
nand ( n215315 , n215314 , n37682 );
nand ( n215316 , n36980 , n35625 );
and ( n215317 , n215315 , n215316 );
not ( n215318 , n215315 );
not ( n215319 , n215316 );
and ( n215320 , n215318 , n215319 );
nor ( n215321 , n215317 , n215320 );
not ( n215322 , n215321 );
or ( n215323 , n215309 , n215322 );
not ( n215324 , n215321 );
nand ( n215325 , n215103 , n215324 );
nand ( n215326 , n215323 , n215325 );
not ( n215327 , n215326 );
and ( n215328 , n215327 , n213750 );
xor ( n215329 , n215307 , n215328 );
not ( n215330 , n214717 );
not ( n215331 , n215120 );
or ( n215332 , n215330 , n215331 );
not ( n215333 , n215118 );
not ( n215334 , n215333 );
not ( n215335 , n214029 );
or ( n215336 , n215334 , n215335 );
not ( n215337 , n214304 );
nand ( n215338 , n215337 , n215118 );
nand ( n215339 , n215336 , n215338 );
nand ( n215340 , n215339 , n213463 );
nand ( n215341 , n215332 , n215340 );
xor ( n215342 , n215329 , n215341 );
xor ( n215343 , n215307 , n215328 );
and ( n215344 , n215343 , n215341 );
and ( n215345 , n215307 , n215328 );
or ( n215346 , n215344 , n215345 );
not ( n215347 , n215133 );
not ( n215348 , n214610 );
or ( n215349 , n215347 , n215348 );
not ( n215350 , n214537 );
not ( n215351 , n214586 );
or ( n215352 , n215350 , n215351 );
nand ( n215353 , n214418 , n214899 );
nand ( n215354 , n215352 , n215353 );
nand ( n215355 , n215354 , n214458 );
nand ( n215356 , n215349 , n215355 );
not ( n215357 , n215160 );
not ( n215358 , n214799 );
or ( n215359 , n215357 , n215358 );
not ( n215360 , n214956 );
not ( n215361 , n214803 );
or ( n215362 , n215360 , n215361 );
nand ( n215363 , n214786 , n214960 );
nand ( n215364 , n215362 , n215363 );
nand ( n215365 , n215364 , n214808 );
nand ( n215366 , n215359 , n215365 );
xor ( n215367 , n215356 , n215366 );
xor ( n215368 , n215367 , n215301 );
xor ( n215369 , n215356 , n215366 );
and ( n215370 , n215369 , n215301 );
and ( n215371 , n215356 , n215366 );
or ( n215372 , n215370 , n215371 );
not ( n215373 , n215190 );
not ( n215374 , n215183 );
or ( n215375 , n215373 , n215374 );
not ( n215376 , n213347 );
not ( n215377 , n215164 );
or ( n215378 , n215376 , n215377 );
nand ( n215379 , n215104 , n214616 );
nand ( n215380 , n215378 , n215379 );
nand ( n215381 , n215380 , n215191 );
nand ( n215382 , n215375 , n215381 );
buf ( n215383 , n213206 );
not ( n215384 , n215383 );
not ( n215385 , n213960 );
not ( n215386 , n214628 );
or ( n215387 , n215385 , n215386 );
not ( n215388 , n213960 );
nand ( n215389 , n30997 , n215388 );
nand ( n215390 , n215387 , n215389 );
not ( n215391 , n215390 );
or ( n215392 , n215384 , n215391 );
nand ( n215393 , n215143 , n214086 );
nand ( n215394 , n215392 , n215393 );
xor ( n215395 , n215382 , n215394 );
xor ( n215396 , n215395 , n215111 );
xor ( n215397 , n215382 , n215394 );
and ( n215398 , n215397 , n215111 );
and ( n215399 , n215382 , n215394 );
or ( n215400 , n215398 , n215399 );
not ( n215401 , n213758 );
not ( n215402 , n215207 );
or ( n215403 , n215401 , n215402 );
not ( n215404 , n213864 );
not ( n215405 , n215018 );
or ( n215406 , n215404 , n215405 );
nand ( n215407 , n208725 , n213869 );
nand ( n215408 , n215406 , n215407 );
nand ( n215409 , n215408 , n213142 );
nand ( n215410 , n215403 , n215409 );
xor ( n215411 , n215410 , n215342 );
xor ( n215412 , n215411 , n215152 );
xor ( n215413 , n215410 , n215342 );
and ( n215414 , n215413 , n215152 );
and ( n215415 , n215410 , n215342 );
or ( n215416 , n215414 , n215415 );
not ( n215417 , n213577 );
not ( n215418 , n215230 );
or ( n215419 , n215417 , n215418 );
and ( n215420 , n41716 , n213732 );
not ( n215421 , n41716 );
and ( n215422 , n215421 , n213735 );
or ( n215423 , n215420 , n215422 );
nand ( n215424 , n215423 , n213498 );
nand ( n215425 , n215419 , n215424 );
not ( n215426 , n211314 );
not ( n215427 , n213382 );
not ( n215428 , n211451 );
not ( n215429 , n215428 );
or ( n215430 , n215427 , n215429 );
nand ( n215431 , n41701 , n213381 );
nand ( n215432 , n215430 , n215431 );
not ( n215433 , n215432 );
or ( n215434 , n215426 , n215433 );
nand ( n215435 , n215219 , n213784 );
nand ( n215436 , n215434 , n215435 );
xor ( n215437 , n215425 , n215436 );
xor ( n215438 , n215437 , n215198 );
xor ( n215439 , n215425 , n215436 );
and ( n215440 , n215439 , n215198 );
and ( n215441 , n215425 , n215436 );
or ( n215442 , n215440 , n215441 );
xor ( n215443 , n215368 , n215240 );
xor ( n215444 , n215443 , n215396 );
xor ( n215445 , n215368 , n215240 );
and ( n215446 , n215445 , n215396 );
and ( n215447 , n215368 , n215240 );
or ( n215448 , n215446 , n215447 );
xor ( n215449 , n215214 , n215438 );
xor ( n215450 , n215449 , n215412 );
xor ( n215451 , n215214 , n215438 );
and ( n215452 , n215451 , n215412 );
and ( n215453 , n215214 , n215438 );
or ( n215454 , n215452 , n215453 );
xor ( n215455 , n215246 , n215444 );
xor ( n215456 , n215455 , n215252 );
xor ( n215457 , n215246 , n215444 );
and ( n215458 , n215457 , n215252 );
and ( n215459 , n215246 , n215444 );
or ( n215460 , n215458 , n215459 );
xor ( n215461 , n215450 , n215258 );
xor ( n215462 , n215461 , n215456 );
xor ( n215463 , n215450 , n215258 );
and ( n215464 , n215463 , n215456 );
and ( n215465 , n215450 , n215258 );
or ( n215466 , n215464 , n215465 );
not ( n215467 , n214694 );
not ( n215468 , n213918 );
not ( n215469 , n215289 );
or ( n215470 , n215468 , n215469 );
nand ( n215471 , n215290 , n209248 );
nand ( n215472 , n215470 , n215471 );
not ( n215473 , n215472 );
or ( n215474 , n215467 , n215473 );
nand ( n215475 , n215296 , n213718 );
nand ( n215476 , n215474 , n215475 );
not ( n215477 , n215274 );
not ( n215478 , n213894 );
or ( n215479 , n215477 , n215478 );
not ( n215480 , n214130 );
not ( n215481 , n30384 );
not ( n215482 , n215481 );
or ( n215483 , n215480 , n215482 );
nand ( n215484 , n30384 , n213883 );
nand ( n215485 , n215483 , n215484 );
nand ( n215486 , n215485 , n213902 );
nand ( n215487 , n215479 , n215486 );
not ( n215488 , n215284 );
not ( n215489 , n214551 );
or ( n215490 , n215488 , n215489 );
and ( n215491 , n214145 , n213473 );
not ( n215492 , n214145 );
and ( n215493 , n215492 , n215075 );
or ( n215494 , n215491 , n215493 );
nand ( n215495 , n215494 , n214370 );
nand ( n215496 , n215490 , n215495 );
xor ( n215497 , n215487 , n215496 );
xor ( n215498 , n215476 , n215497 );
not ( n215499 , n213750 );
not ( n215500 , n215321 );
not ( n215501 , n215500 );
or ( n215502 , n215499 , n215501 );
nand ( n215503 , n215502 , n215105 );
buf ( n215504 , n215321 );
nand ( n215505 , n215504 , n213751 );
and ( n215506 , n215503 , n215505 );
not ( n215507 , n37616 );
not ( n215508 , n37018 );
or ( n215509 , n215507 , n215508 );
nand ( n215510 , n215509 , n36985 );
buf ( n215511 , n215510 );
not ( n215512 , n215511 );
nor ( n215513 , n215506 , n215512 );
xor ( n215514 , n215498 , n215513 );
xor ( n215515 , n215476 , n215497 );
and ( n215516 , n215515 , n215513 );
and ( n215517 , n215476 , n215497 );
or ( n215518 , n215516 , n215517 );
not ( n215519 , n215354 );
not ( n215520 , n214449 );
or ( n215521 , n215519 , n215520 );
not ( n215522 , n215050 );
not ( n215523 , n214417 );
or ( n215524 , n215522 , n215523 );
nand ( n215525 , n214759 , n214678 );
nand ( n215526 , n215524 , n215525 );
nand ( n215527 , n215526 , n214457 );
nand ( n215528 , n215521 , n215527 );
not ( n215529 , n213463 );
not ( n215530 , n215113 );
not ( n215531 , n214190 );
or ( n215532 , n215530 , n215531 );
not ( n215533 , n214467 );
nand ( n215534 , n215533 , n214712 );
nand ( n215535 , n215532 , n215534 );
not ( n215536 , n215535 );
or ( n215537 , n215529 , n215536 );
nand ( n215538 , n215339 , n214717 );
nand ( n215539 , n215537 , n215538 );
xor ( n215540 , n215528 , n215539 );
not ( n215541 , n215380 );
not ( n215542 , n215182 );
or ( n215543 , n215541 , n215542 );
not ( n215544 , n213583 );
not ( n215545 , n215104 );
not ( n215546 , n215545 );
or ( n215547 , n215544 , n215546 );
nand ( n215548 , n215104 , n214134 );
nand ( n215549 , n215547 , n215548 );
not ( n215550 , n214951 );
nand ( n215551 , n215549 , n215550 );
nand ( n215552 , n215543 , n215551 );
xor ( n215553 , n215540 , n215552 );
xor ( n215554 , n215528 , n215539 );
and ( n215555 , n215554 , n215552 );
and ( n215556 , n215528 , n215539 );
or ( n215557 , n215555 , n215556 );
not ( n215558 , n215364 );
not ( n215559 , n214799 );
or ( n215560 , n215558 , n215559 );
not ( n215561 , n214357 );
not ( n215562 , n214803 );
or ( n215563 , n215561 , n215562 );
nand ( n215564 , n214786 , n215131 );
nand ( n215565 , n215563 , n215564 );
nand ( n215566 , n215565 , n214588 );
nand ( n215567 , n215560 , n215566 );
not ( n215568 , n213750 );
not ( n215569 , n215511 );
not ( n215570 , n215569 );
or ( n215571 , n215568 , n215570 );
not ( n215572 , n215569 );
nand ( n215573 , n215572 , n213751 );
nand ( n215574 , n215571 , n215573 );
not ( n215575 , n215574 );
xor ( n215576 , n215510 , n215500 );
nand ( n215577 , n215576 , n215326 );
not ( n215578 , n215577 );
not ( n215579 , n215578 );
or ( n215580 , n215575 , n215579 );
not ( n215581 , n213126 );
not ( n215582 , n215512 );
or ( n215583 , n215581 , n215582 );
nand ( n215584 , n215511 , n213077 );
nand ( n215585 , n215583 , n215584 );
not ( n215586 , n215327 );
not ( n215587 , n215586 );
nand ( n215588 , n215585 , n215587 );
nand ( n215589 , n215580 , n215588 );
xor ( n215590 , n215567 , n215589 );
xor ( n215591 , n215590 , n215305 );
xor ( n215592 , n215567 , n215589 );
and ( n215593 , n215592 , n215305 );
and ( n215594 , n215567 , n215589 );
or ( n215595 , n215593 , n215594 );
not ( n215596 , n215137 );
not ( n215597 , n213960 );
not ( n215598 , n214488 );
or ( n215599 , n215597 , n215598 );
not ( n215600 , n213960 );
nand ( n215601 , n215228 , n215600 );
nand ( n215602 , n215599 , n215601 );
not ( n215603 , n215602 );
or ( n215604 , n215596 , n215603 );
not ( n215605 , n214085 );
nand ( n215606 , n215390 , n215605 );
nand ( n215607 , n215604 , n215606 );
xor ( n215608 , n215346 , n215607 );
not ( n215609 , n213784 );
not ( n215610 , n215432 );
or ( n215611 , n215609 , n215610 );
not ( n215612 , n213382 );
not ( n215613 , n41564 );
not ( n215614 , n215613 );
or ( n215615 , n215612 , n215614 );
not ( n215616 , n41563 );
nand ( n215617 , n215616 , n213381 );
nand ( n215618 , n215615 , n215617 );
nand ( n215619 , n215618 , n211314 );
nand ( n215620 , n215611 , n215619 );
xor ( n215621 , n215608 , n215620 );
xor ( n215622 , n215346 , n215607 );
and ( n215623 , n215622 , n215620 );
and ( n215624 , n215346 , n215607 );
or ( n215625 , n215623 , n215624 );
not ( n215626 , n213142 );
not ( n215627 , n213864 );
not ( n215628 , n41608 );
not ( n215629 , n215628 );
or ( n215630 , n215627 , n215629 );
nand ( n215631 , n41608 , n213869 );
nand ( n215632 , n215630 , n215631 );
not ( n215633 , n215632 );
or ( n215634 , n215626 , n215633 );
nand ( n215635 , n215408 , n213758 );
nand ( n215636 , n215634 , n215635 );
xor ( n215637 , n215636 , n215514 );
not ( n215638 , n213498 );
not ( n215639 , n213735 );
not ( n215640 , n214834 );
or ( n215641 , n215639 , n215640 );
not ( n215642 , n214834 );
nand ( n215643 , n215642 , n213732 );
nand ( n215644 , n215641 , n215643 );
not ( n215645 , n215644 );
or ( n215646 , n215638 , n215645 );
nand ( n215647 , n215423 , n213577 );
nand ( n215648 , n215646 , n215647 );
xor ( n215649 , n215637 , n215648 );
xor ( n215650 , n215636 , n215514 );
and ( n215651 , n215650 , n215648 );
and ( n215652 , n215636 , n215514 );
or ( n215653 , n215651 , n215652 );
xor ( n215654 , n215372 , n215553 );
xor ( n215655 , n215654 , n215591 );
xor ( n215656 , n215372 , n215553 );
and ( n215657 , n215656 , n215591 );
and ( n215658 , n215372 , n215553 );
or ( n215659 , n215657 , n215658 );
xor ( n215660 , n215400 , n215416 );
xor ( n215661 , n215660 , n215649 );
xor ( n215662 , n215400 , n215416 );
and ( n215663 , n215662 , n215649 );
and ( n215664 , n215400 , n215416 );
or ( n215665 , n215663 , n215664 );
xor ( n215666 , n215442 , n215621 );
xor ( n215667 , n215666 , n215655 );
xor ( n215668 , n215442 , n215621 );
and ( n215669 , n215668 , n215655 );
and ( n215670 , n215442 , n215621 );
or ( n215671 , n215669 , n215670 );
xor ( n215672 , n215448 , n215661 );
xor ( n215673 , n215672 , n215454 );
xor ( n215674 , n215448 , n215661 );
and ( n215675 , n215674 , n215454 );
and ( n215676 , n215448 , n215661 );
or ( n215677 , n215675 , n215676 );
xor ( n215678 , n215667 , n215460 );
xor ( n215679 , n215678 , n215673 );
xor ( n215680 , n215667 , n215460 );
and ( n215681 , n215680 , n215673 );
and ( n215682 , n215667 , n215460 );
or ( n215683 , n215681 , n215682 );
not ( n215684 , n215494 );
not ( n215685 , n214551 );
or ( n215686 , n215684 , n215685 );
not ( n215687 , n215268 );
not ( n215688 , n214067 );
or ( n215689 , n215687 , n215688 );
nand ( n215690 , n214144 , n213763 );
nand ( n215691 , n215689 , n215690 );
nand ( n215692 , n214370 , n215691 );
nand ( n215693 , n215686 , n215692 );
not ( n215694 , n214888 );
not ( n215695 , n215272 );
not ( n215696 , n30292 );
not ( n215697 , n215696 );
or ( n215698 , n215695 , n215697 );
nand ( n215699 , n30292 , n214131 );
nand ( n215700 , n215698 , n215699 );
not ( n215701 , n215700 );
or ( n215702 , n215694 , n215701 );
nand ( n215703 , n215485 , n213894 );
nand ( n215704 , n215702 , n215703 );
xor ( n215705 , n215693 , n215704 );
not ( n215706 , n213718 );
not ( n215707 , n215472 );
or ( n215708 , n215706 , n215707 );
not ( n215709 , n215290 );
not ( n215710 , n214029 );
or ( n215711 , n215709 , n215710 );
nand ( n215712 , n41894 , n215289 );
nand ( n215713 , n215711 , n215712 );
nand ( n215714 , n215713 , n214694 );
nand ( n215715 , n215708 , n215714 );
xor ( n215716 , n215705 , n215715 );
xor ( n215717 , n215693 , n215704 );
and ( n215718 , n215717 , n215715 );
and ( n215719 , n215693 , n215704 );
or ( n215720 , n215718 , n215719 );
and ( n215721 , n215487 , n215496 );
not ( n215722 , n215526 );
not ( n215723 , n214610 );
or ( n215724 , n215722 , n215723 );
not ( n215725 , n214881 );
not ( n215726 , n214417 );
or ( n215727 , n215725 , n215726 );
nand ( n215728 , n214759 , n214885 );
nand ( n215729 , n215727 , n215728 );
nand ( n215730 , n215729 , n214458 );
nand ( n215731 , n215724 , n215730 );
xor ( n215732 , n215721 , n215731 );
not ( n215733 , n215565 );
not ( n215734 , n214799 );
or ( n215735 , n215733 , n215734 );
not ( n215736 , n214537 );
not ( n215737 , n214783 );
or ( n215738 , n215736 , n215737 );
nand ( n215739 , n214747 , n214899 );
nand ( n215740 , n215738 , n215739 );
nand ( n215741 , n214808 , n215740 );
nand ( n215742 , n215735 , n215741 );
xor ( n215743 , n215732 , n215742 );
xor ( n215744 , n215721 , n215731 );
and ( n215745 , n215744 , n215742 );
and ( n215746 , n215721 , n215731 );
or ( n215747 , n215745 , n215746 );
xor ( n215748 , n215557 , n215595 );
xor ( n215749 , n215748 , n215743 );
xor ( n215750 , n215749 , n215659 );
not ( n215751 , n215549 );
not ( n215752 , n215182 );
or ( n215753 , n215751 , n215752 );
not ( n215754 , n214956 );
not ( n215755 , n215545 );
or ( n215756 , n215754 , n215755 );
nand ( n215757 , n215104 , n214960 );
nand ( n215758 , n215756 , n215757 );
nand ( n215759 , n215758 , n215550 );
nand ( n215760 , n215753 , n215759 );
buf ( n215761 , n215326 );
not ( n215762 , n215761 );
not ( n215763 , n215762 );
not ( n215764 , n214616 );
not ( n215765 , n215510 );
not ( n215766 , n215765 );
not ( n215767 , n215766 );
or ( n215768 , n215764 , n215767 );
nand ( n215769 , n215569 , n213347 );
nand ( n215770 , n215768 , n215769 );
not ( n215771 , n215770 );
or ( n215772 , n215763 , n215771 );
not ( n215773 , n215577 );
nand ( n215774 , n215773 , n215585 );
nand ( n215775 , n215772 , n215774 );
xor ( n215776 , n215760 , n215775 );
and ( n215777 , n37490 , n36272 );
not ( n215778 , n215777 );
not ( n215779 , n36999 );
or ( n215780 , n215778 , n215779 );
or ( n215781 , n215777 , n36999 );
nand ( n215782 , n215780 , n215781 );
not ( n215783 , n215782 );
and ( n215784 , n215783 , n215511 );
not ( n215785 , n215783 );
and ( n215786 , n215785 , n215765 );
nor ( n215787 , n215784 , n215786 );
not ( n215788 , n215787 );
buf ( n215789 , n215788 );
nor ( n215790 , n215789 , n213751 );
xor ( n215791 , n215776 , n215790 );
not ( n215792 , n213382 );
not ( n215793 , n208717 );
not ( n215794 , n215793 );
or ( n215795 , n215792 , n215794 );
buf ( n215796 , n208717 );
nand ( n215797 , n215796 , n213381 );
nand ( n215798 , n215795 , n215797 );
not ( n215799 , n215798 );
not ( n215800 , n211314 );
or ( n215801 , n215799 , n215800 );
nand ( n215802 , n215618 , n213784 );
nand ( n215803 , n215801 , n215802 );
xor ( n215804 , n215791 , n215803 );
not ( n215805 , n213463 );
not ( n215806 , n30997 );
xor ( n215807 , n214712 , n215806 );
not ( n215808 , n215807 );
or ( n215809 , n215805 , n215808 );
nand ( n215810 , n215535 , n214717 );
nand ( n215811 , n215809 , n215810 );
xor ( n215812 , n215716 , n215811 );
xor ( n215813 , n215812 , n215518 );
xor ( n215814 , n215804 , n215813 );
xor ( n215815 , n215750 , n215814 );
xor ( n215816 , n215815 , n215677 );
xor ( n215817 , n215653 , n215625 );
not ( n215818 , n213142 );
not ( n215819 , n213864 );
not ( n215820 , n41700 );
not ( n215821 , n215820 );
or ( n215822 , n215819 , n215821 );
nand ( n215823 , n211451 , n213869 );
nand ( n215824 , n215822 , n215823 );
not ( n215825 , n215824 );
or ( n215826 , n215818 , n215825 );
nand ( n215827 , n215632 , n213758 );
nand ( n215828 , n215826 , n215827 );
not ( n215829 , n214086 );
not ( n215830 , n215602 );
or ( n215831 , n215829 , n215830 );
not ( n215832 , n213960 );
not ( n215833 , n41716 );
not ( n215834 , n215833 );
or ( n215835 , n215832 , n215834 );
nand ( n215836 , n41716 , n215600 );
nand ( n215837 , n215835 , n215836 );
nand ( n215838 , n215837 , n215137 );
nand ( n215839 , n215831 , n215838 );
xor ( n215840 , n215828 , n215839 );
not ( n215841 , n213577 );
not ( n215842 , n215644 );
or ( n215843 , n215841 , n215842 );
not ( n215844 , n213735 );
not ( n215845 , n208725 );
not ( n215846 , n215845 );
or ( n215847 , n215844 , n215846 );
nand ( n215848 , n208725 , n213732 );
nand ( n215849 , n215847 , n215848 );
nand ( n215850 , n215849 , n213498 );
nand ( n215851 , n215843 , n215850 );
xor ( n215852 , n215840 , n215851 );
xor ( n215853 , n215817 , n215852 );
xor ( n215854 , n215853 , n215665 );
xor ( n215855 , n215854 , n215671 );
xor ( n215856 , n215816 , n215855 );
xor ( n215857 , n215815 , n215677 );
and ( n215858 , n215857 , n215855 );
and ( n215859 , n215815 , n215677 );
or ( n215860 , n215858 , n215859 );
xor ( n215861 , n215760 , n215775 );
and ( n215862 , n215861 , n215790 );
and ( n215863 , n215760 , n215775 );
or ( n215864 , n215862 , n215863 );
xor ( n215865 , n215716 , n215811 );
and ( n215866 , n215865 , n215518 );
and ( n215867 , n215716 , n215811 );
or ( n215868 , n215866 , n215867 );
xor ( n215869 , n215828 , n215839 );
and ( n215870 , n215869 , n215851 );
and ( n215871 , n215828 , n215839 );
or ( n215872 , n215870 , n215871 );
xor ( n215873 , n215557 , n215595 );
and ( n215874 , n215873 , n215743 );
and ( n215875 , n215557 , n215595 );
or ( n215876 , n215874 , n215875 );
xor ( n215877 , n215791 , n215803 );
and ( n215878 , n215877 , n215813 );
and ( n215879 , n215791 , n215803 );
or ( n215880 , n215878 , n215879 );
xor ( n215881 , n215653 , n215625 );
and ( n215882 , n215881 , n215852 );
and ( n215883 , n215653 , n215625 );
or ( n215884 , n215882 , n215883 );
xor ( n215885 , n215749 , n215659 );
and ( n215886 , n215885 , n215814 );
and ( n215887 , n215749 , n215659 );
or ( n215888 , n215886 , n215887 );
xor ( n215889 , n215853 , n215665 );
and ( n215890 , n215889 , n215671 );
and ( n215891 , n215853 , n215665 );
or ( n215892 , n215890 , n215891 );
not ( n215893 , n215729 );
not ( n215894 , n214610 );
or ( n215895 , n215893 , n215894 );
not ( n215896 , n215075 );
not ( n215897 , n214417 );
or ( n215898 , n215896 , n215897 );
not ( n215899 , n215075 );
nand ( n215900 , n214418 , n215899 );
nand ( n215901 , n215898 , n215900 );
nand ( n215902 , n215901 , n214458 );
nand ( n215903 , n215895 , n215902 );
not ( n215904 , n214694 );
not ( n215905 , n215290 );
not ( n215906 , n214190 );
or ( n215907 , n215905 , n215906 );
nand ( n215908 , n215289 , n214468 );
nand ( n215909 , n215907 , n215908 );
not ( n215910 , n215909 );
or ( n215911 , n215904 , n215910 );
nand ( n215912 , n215713 , n213718 );
nand ( n215913 , n215911 , n215912 );
xor ( n215914 , n215903 , n215913 );
not ( n215915 , n215740 );
not ( n215916 , n214799 );
or ( n215917 , n215915 , n215916 );
not ( n215918 , n215050 );
not ( n215919 , n214803 );
or ( n215920 , n215918 , n215919 );
not ( n215921 , n214783 );
nand ( n215922 , n215921 , n214678 );
nand ( n215923 , n215920 , n215922 );
nand ( n215924 , n215923 , n214808 );
nand ( n215925 , n215917 , n215924 );
xor ( n215926 , n215914 , n215925 );
xor ( n215927 , n215903 , n215913 );
and ( n215928 , n215927 , n215925 );
and ( n215929 , n215903 , n215913 );
or ( n215930 , n215928 , n215929 );
not ( n215931 , n215758 );
not ( n215932 , n215182 );
or ( n215933 , n215931 , n215932 );
not ( n215934 , n214357 );
not ( n215935 , n215164 );
or ( n215936 , n215934 , n215935 );
nand ( n215937 , n215104 , n215131 );
nand ( n215938 , n215936 , n215937 );
nand ( n215939 , n215938 , n215550 );
nand ( n215940 , n215933 , n215939 );
not ( n215941 , n215770 );
not ( n215942 , n215578 );
or ( n215943 , n215941 , n215942 );
not ( n215944 , n213583 );
not ( n215945 , n215512 );
or ( n215946 , n215944 , n215945 );
nand ( n215947 , n215511 , n214134 );
nand ( n215948 , n215946 , n215947 );
nand ( n215949 , n215948 , n215762 );
nand ( n215950 , n215943 , n215949 );
xor ( n215951 , n215940 , n215950 );
not ( n215952 , n214164 );
not ( n215953 , n215481 );
not ( n215954 , n215953 );
buf ( n215955 , n214688 );
not ( n215956 , n215955 );
not ( n215957 , n215956 );
or ( n215958 , n215954 , n215957 );
nand ( n215959 , n215955 , n215481 );
nand ( n215960 , n215958 , n215959 );
not ( n215961 , n215960 );
or ( n215962 , n215952 , n215961 );
not ( n215963 , n214550 );
nand ( n215964 , n215963 , n215691 );
nand ( n215965 , n215962 , n215964 );
not ( n215966 , n213749 );
not ( n215967 , n215966 );
not ( n215968 , n215272 );
not ( n215969 , n209248 );
or ( n215970 , n215968 , n215969 );
not ( n215971 , n215272 );
nand ( n215972 , n41972 , n215971 );
nand ( n215973 , n215970 , n215972 );
not ( n215974 , n215973 );
or ( n215975 , n215967 , n215974 );
nand ( n215976 , n215700 , n213894 );
nand ( n215977 , n215975 , n215976 );
xor ( n215978 , n215965 , n215977 );
xor ( n215979 , n215951 , n215978 );
xor ( n215980 , n215940 , n215950 );
and ( n215981 , n215980 , n215978 );
and ( n215982 , n215940 , n215950 );
or ( n215983 , n215981 , n215982 );
xor ( n215984 , n215926 , n215868 );
xor ( n215985 , n215984 , n215979 );
xor ( n215986 , n215985 , n215880 );
not ( n215987 , n211314 );
not ( n215988 , n213382 );
not ( n215989 , n41396 );
not ( n215990 , n215989 );
or ( n215991 , n215988 , n215990 );
nand ( n215992 , n41397 , n213381 );
nand ( n215993 , n215991 , n215992 );
not ( n215994 , n215993 );
or ( n215995 , n215987 , n215994 );
nand ( n215996 , n215798 , n213784 );
nand ( n215997 , n215995 , n215996 );
xor ( n215998 , n215997 , n215872 );
not ( n215999 , n213751 );
and ( n216000 , n215783 , n215999 );
nor ( n216001 , n216000 , n215766 );
nor ( n216002 , n215783 , n213750 );
or ( n216003 , n216001 , n216002 );
not ( n216004 , n37673 );
buf ( n216005 , n36272 );
nand ( n216006 , n37491 , n37022 , n216005 );
not ( n216007 , n216006 );
or ( n216008 , n216004 , n216007 );
not ( n216009 , n216005 );
nor ( n216010 , n216009 , n37673 );
nand ( n216011 , n37491 , n37022 , n216010 );
nand ( n216012 , n216008 , n216011 );
not ( n216013 , n216012 );
buf ( n216014 , n216013 );
not ( n216015 , n216014 );
nand ( n216016 , n216003 , n216015 );
not ( n216017 , n216016 );
xor ( n216018 , n216017 , n215720 );
not ( n216019 , n215383 );
not ( n216020 , n213960 );
not ( n216021 , n214834 );
or ( n216022 , n216020 , n216021 );
nand ( n216023 , n30962 , n215388 );
nand ( n216024 , n216022 , n216023 );
not ( n216025 , n216024 );
or ( n216026 , n216019 , n216025 );
nand ( n216027 , n215837 , n214086 );
nand ( n216028 , n216026 , n216027 );
xor ( n216029 , n216018 , n216028 );
xor ( n216030 , n215998 , n216029 );
xor ( n216031 , n215986 , n216030 );
xor ( n216032 , n216031 , n215892 );
not ( n216033 , n213463 );
not ( n216034 , n215333 );
not ( n216035 , n214820 );
or ( n216036 , n216034 , n216035 );
not ( n216037 , n215113 );
nand ( n216038 , n41725 , n216037 );
nand ( n216039 , n216036 , n216038 );
not ( n216040 , n216039 );
or ( n216041 , n216033 , n216040 );
nand ( n216042 , n215807 , n214717 );
nand ( n216043 , n216041 , n216042 );
not ( n216044 , n213498 );
not ( n216045 , n213735 );
not ( n216046 , n41608 );
not ( n216047 , n216046 );
or ( n216048 , n216045 , n216047 );
not ( n216049 , n215628 );
nand ( n216050 , n216049 , n213732 );
nand ( n216051 , n216048 , n216050 );
not ( n216052 , n216051 );
or ( n216053 , n216044 , n216052 );
nand ( n216054 , n215849 , n213577 );
nand ( n216055 , n216053 , n216054 );
xor ( n216056 , n216043 , n216055 );
not ( n216057 , n215783 );
buf ( n216058 , n216012 );
not ( n216059 , n216058 );
not ( n216060 , n216059 );
or ( n216061 , n216057 , n216060 );
nand ( n216062 , n216058 , n215782 );
nand ( n216063 , n216061 , n216062 );
nand ( n216064 , n216063 , n215788 );
not ( n216065 , n216064 );
not ( n216066 , n216065 );
not ( n216067 , n216058 );
not ( n216068 , n216067 );
and ( n216069 , n216068 , n213751 );
not ( n216070 , n216068 );
and ( n216071 , n216070 , n213750 );
nor ( n216072 , n216069 , n216071 );
or ( n216073 , n216066 , n216072 );
not ( n216074 , n216067 );
not ( n216075 , n216074 );
buf ( n216076 , n213077 );
not ( n216077 , n216076 );
and ( n216078 , n216075 , n216077 );
and ( n216079 , n216015 , n213077 );
nor ( n216080 , n216078 , n216079 );
or ( n216081 , n216080 , n215789 );
nand ( n216082 , n216073 , n216081 );
xor ( n216083 , n216056 , n216082 );
xor ( n216084 , n216083 , n215876 );
not ( n216085 , n213142 );
not ( n216086 , n213864 );
not ( n216087 , n41563 );
or ( n216088 , n216086 , n216087 );
not ( n216089 , n41563 );
nand ( n216090 , n216089 , n213869 );
nand ( n216091 , n216088 , n216090 );
not ( n216092 , n216091 );
or ( n216093 , n216085 , n216092 );
nand ( n216094 , n215824 , n213758 );
nand ( n216095 , n216093 , n216094 );
xor ( n216096 , n216095 , n215747 );
xor ( n216097 , n216096 , n215864 );
xor ( n216098 , n216084 , n216097 );
xor ( n216099 , n215884 , n216098 );
xor ( n216100 , n216099 , n215888 );
xor ( n216101 , n216032 , n216100 );
xor ( n216102 , n216031 , n215892 );
and ( n216103 , n216102 , n216100 );
and ( n216104 , n216031 , n215892 );
or ( n216105 , n216103 , n216104 );
xor ( n216106 , n216017 , n215720 );
and ( n216107 , n216106 , n216028 );
and ( n216108 , n216017 , n215720 );
or ( n216109 , n216107 , n216108 );
xor ( n216110 , n216043 , n216055 );
and ( n216111 , n216110 , n216082 );
and ( n216112 , n216043 , n216055 );
or ( n216113 , n216111 , n216112 );
xor ( n216114 , n216095 , n215747 );
and ( n216115 , n216114 , n215864 );
and ( n216116 , n216095 , n215747 );
or ( n216117 , n216115 , n216116 );
xor ( n216118 , n215926 , n215868 );
and ( n216119 , n216118 , n215979 );
and ( n216120 , n215926 , n215868 );
or ( n216121 , n216119 , n216120 );
xor ( n216122 , n215997 , n215872 );
and ( n216123 , n216122 , n216029 );
and ( n216124 , n215997 , n215872 );
or ( n216125 , n216123 , n216124 );
xor ( n216126 , n216083 , n215876 );
and ( n216127 , n216126 , n216097 );
and ( n216128 , n216083 , n215876 );
or ( n216129 , n216127 , n216128 );
xor ( n216130 , n215985 , n215880 );
and ( n216131 , n216130 , n216030 );
and ( n216132 , n215985 , n215880 );
or ( n216133 , n216131 , n216132 );
xor ( n216134 , n215884 , n216098 );
and ( n216135 , n216134 , n215888 );
and ( n216136 , n215884 , n216098 );
or ( n216137 , n216135 , n216136 );
not ( n216138 , n214164 );
not ( n216139 , n30292 );
and ( n216140 , n215054 , n216139 );
not ( n216141 , n215054 );
not ( n216142 , n216139 );
and ( n216143 , n216141 , n216142 );
or ( n216144 , n216140 , n216143 );
not ( n216145 , n216144 );
or ( n216146 , n216138 , n216145 );
nand ( n216147 , n214893 , n215960 );
nand ( n216148 , n216146 , n216147 );
not ( n216149 , n213894 );
not ( n216150 , n215973 );
or ( n216151 , n216149 , n216150 );
not ( n216152 , n214304 );
not ( n216153 , n216152 );
not ( n216154 , n214131 );
and ( n216155 , n216153 , n216154 );
and ( n216156 , n214927 , n215971 );
nor ( n216157 , n216155 , n216156 );
not ( n216158 , n216157 );
nand ( n216159 , n216158 , n215966 );
nand ( n216160 , n216151 , n216159 );
xor ( n216161 , n216148 , n216160 );
not ( n216162 , n215901 );
not ( n216163 , n214610 );
or ( n216164 , n216162 , n216163 );
not ( n216165 , n215268 );
buf ( n216166 , n214418 );
not ( n216167 , n216166 );
not ( n216168 , n216167 );
or ( n216169 , n216165 , n216168 );
not ( n216170 , n215268 );
nand ( n216171 , n216166 , n216170 );
nand ( n216172 , n216169 , n216171 );
nand ( n216173 , n216172 , n214458 );
nand ( n216174 , n216164 , n216173 );
xor ( n216175 , n216161 , n216174 );
xor ( n216176 , n216148 , n216160 );
and ( n216177 , n216176 , n216174 );
and ( n216178 , n216148 , n216160 );
or ( n216179 , n216177 , n216178 );
not ( n216180 , n37706 );
not ( n216181 , n216180 );
not ( n216182 , n37019 );
buf ( n216183 , n35598 );
nand ( n216184 , n216182 , n36658 , n216183 );
not ( n216185 , n36647 );
nand ( n216186 , n216185 , n216183 );
not ( n216187 , n36993 );
nand ( n216188 , n216184 , n216186 , n216187 );
not ( n216189 , n216188 );
or ( n216190 , n216181 , n216189 );
nand ( n216191 , n216184 , n216186 , n216187 , n37706 );
nand ( n216192 , n216190 , n216191 );
not ( n216193 , n216192 );
and ( n216194 , n216193 , n216013 );
not ( n216195 , n216193 );
not ( n216196 , n216012 );
not ( n216197 , n216196 );
and ( n216198 , n216195 , n216197 );
nor ( n216199 , n216194 , n216198 );
buf ( n216200 , n216199 );
not ( n216201 , n216200 );
and ( n216202 , n216201 , n213750 );
not ( n216203 , n215923 );
buf ( n216204 , n214799 );
not ( n216205 , n216204 );
or ( n216206 , n216203 , n216205 );
buf ( n216207 , n214885 );
not ( n216208 , n216207 );
and ( n216209 , n216208 , n214786 );
not ( n216210 , n216208 );
and ( n216211 , n216210 , n214783 );
nor ( n216212 , n216209 , n216211 );
nand ( n216213 , n214808 , n216212 );
nand ( n216214 , n216206 , n216213 );
xor ( n216215 , n216202 , n216214 );
not ( n216216 , n215938 );
not ( n216217 , n215183 );
or ( n216218 , n216216 , n216217 );
nand ( n216219 , n215104 , n214899 );
nand ( n216220 , n214537 , n215105 );
nand ( n216221 , n216219 , n216220 );
nand ( n216222 , n215550 , n216221 );
nand ( n216223 , n216218 , n216222 );
xor ( n216224 , n216215 , n216223 );
xor ( n216225 , n216202 , n216214 );
and ( n216226 , n216225 , n216223 );
and ( n216227 , n216202 , n216214 );
or ( n216228 , n216226 , n216227 );
not ( n216229 , n214086 );
not ( n216230 , n216024 );
or ( n216231 , n216229 , n216230 );
not ( n216232 , n213960 );
not ( n216233 , n208726 );
or ( n216234 , n216232 , n216233 );
nand ( n216235 , n208725 , n215388 );
nand ( n216236 , n216234 , n216235 );
nand ( n216237 , n216236 , n215137 );
nand ( n216238 , n216231 , n216237 );
buf ( n216239 , n213463 );
not ( n216240 , n216239 );
not ( n216241 , n215333 );
not ( n216242 , n215833 );
or ( n216243 , n216241 , n216242 );
nand ( n216244 , n41716 , n216037 );
nand ( n216245 , n216243 , n216244 );
not ( n216246 , n216245 );
or ( n216247 , n216240 , n216246 );
nand ( n216248 , n216039 , n214717 );
nand ( n216249 , n216247 , n216248 );
xor ( n216250 , n216238 , n216249 );
xor ( n216251 , n216250 , n216175 );
xor ( n216252 , n216251 , n216121 );
xor ( n216253 , n216252 , n216125 );
xor ( n216254 , n216129 , n216253 );
xor ( n216255 , n216254 , n216133 );
xor ( n216256 , n216129 , n216253 );
and ( n216257 , n216256 , n216133 );
and ( n216258 , n216129 , n216253 );
or ( n216259 , n216257 , n216258 );
not ( n216260 , n213058 );
not ( n216261 , n208717 );
buf ( n216262 , n213060 );
and ( n216263 , n216261 , n216262 );
not ( n216264 , n216261 );
buf ( n216265 , n213147 );
and ( n216266 , n216264 , n216265 );
or ( n216267 , n216263 , n216266 );
not ( n216268 , n216267 );
or ( n216269 , n216260 , n216268 );
nand ( n216270 , n216091 , n213874 );
nand ( n216271 , n216269 , n216270 );
xor ( n216272 , n215983 , n216271 );
not ( n216273 , n215948 );
not ( n216274 , n215773 );
or ( n216275 , n216273 , n216274 );
not ( n216276 , n214956 );
not ( n216277 , n215766 );
not ( n216278 , n216277 );
or ( n216279 , n216276 , n216278 );
not ( n216280 , n215511 );
not ( n216281 , n216280 );
nand ( n216282 , n216281 , n214960 );
nand ( n216283 , n216279 , n216282 );
nand ( n216284 , n216283 , n215762 );
nand ( n216285 , n216275 , n216284 );
and ( n216286 , n215965 , n215977 );
xor ( n216287 , n216285 , n216286 );
not ( n216288 , n214694 );
not ( n216289 , n215290 );
not ( n216290 , n30997 );
not ( n216291 , n216290 );
or ( n216292 , n216289 , n216291 );
buf ( n216293 , n30997 );
nand ( n216294 , n216293 , n215289 );
nand ( n216295 , n216292 , n216294 );
not ( n216296 , n216295 );
or ( n216297 , n216288 , n216296 );
not ( n216298 , n213718 );
not ( n216299 , n216298 );
nand ( n216300 , n215909 , n216299 );
nand ( n216301 , n216297 , n216300 );
xor ( n216302 , n216287 , n216301 );
xor ( n216303 , n216272 , n216302 );
not ( n216304 , n213912 );
not ( n216305 , n213382 );
not ( n216306 , n208594 );
not ( n216307 , n216306 );
not ( n216308 , n216307 );
or ( n216309 , n216305 , n216308 );
not ( n216310 , n41316 );
buf ( n216311 , n216310 );
nand ( n216312 , n216311 , n213381 );
nand ( n216313 , n216309 , n216312 );
not ( n216314 , n216313 );
or ( n216315 , n216304 , n216314 );
nand ( n216316 , n215993 , n213784 );
nand ( n216317 , n216315 , n216316 );
xor ( n216318 , n216224 , n216317 );
xor ( n216319 , n216318 , n216109 );
xor ( n216320 , n216303 , n216319 );
xor ( n216321 , n216113 , n216117 );
not ( n216322 , n216080 );
not ( n216323 , n216322 );
not ( n216324 , n216064 );
not ( n216325 , n216324 );
or ( n216326 , n216323 , n216325 );
not ( n216327 , n216059 );
and ( n216328 , n213347 , n216327 );
not ( n216329 , n213347 );
and ( n216330 , n216329 , n216014 );
nor ( n216331 , n216328 , n216330 );
not ( n216332 , n215789 );
nand ( n216333 , n216331 , n216332 );
nand ( n216334 , n216326 , n216333 );
buf ( n216335 , n213121 );
not ( n216336 , n216335 );
not ( n216337 , n216336 );
not ( n216338 , n213735 );
not ( n216339 , n211451 );
not ( n216340 , n216339 );
or ( n216341 , n216338 , n216340 );
nand ( n216342 , n211451 , n213732 );
nand ( n216343 , n216341 , n216342 );
not ( n216344 , n216343 );
or ( n216345 , n216337 , n216344 );
nand ( n216346 , n216051 , n213577 );
nand ( n216347 , n216345 , n216346 );
xor ( n216348 , n216334 , n216347 );
xor ( n216349 , n216348 , n215930 );
xor ( n216350 , n216321 , n216349 );
xor ( n216351 , n216320 , n216350 );
xor ( n216352 , n216351 , n216137 );
xor ( n216353 , n216352 , n216255 );
xor ( n216354 , n216351 , n216137 );
and ( n216355 , n216354 , n216255 );
and ( n216356 , n216351 , n216137 );
or ( n216357 , n216355 , n216356 );
xor ( n216358 , n216285 , n216286 );
and ( n216359 , n216358 , n216301 );
and ( n216360 , n216285 , n216286 );
or ( n216361 , n216359 , n216360 );
xor ( n216362 , n216238 , n216249 );
and ( n216363 , n216362 , n216175 );
and ( n216364 , n216238 , n216249 );
or ( n216365 , n216363 , n216364 );
xor ( n216366 , n216334 , n216347 );
and ( n216367 , n216366 , n215930 );
and ( n216368 , n216334 , n216347 );
or ( n216369 , n216367 , n216368 );
xor ( n216370 , n215983 , n216271 );
and ( n216371 , n216370 , n216302 );
and ( n216372 , n215983 , n216271 );
or ( n216373 , n216371 , n216372 );
xor ( n216374 , n216224 , n216317 );
and ( n216375 , n216374 , n216109 );
and ( n216376 , n216224 , n216317 );
or ( n216377 , n216375 , n216376 );
xor ( n216378 , n216113 , n216117 );
and ( n216379 , n216378 , n216349 );
and ( n216380 , n216113 , n216117 );
or ( n216381 , n216379 , n216380 );
xor ( n216382 , n216251 , n216121 );
and ( n216383 , n216382 , n216125 );
and ( n216384 , n216251 , n216121 );
or ( n216385 , n216383 , n216384 );
xor ( n216386 , n216303 , n216319 );
and ( n216387 , n216386 , n216350 );
and ( n216388 , n216303 , n216319 );
or ( n216389 , n216387 , n216388 );
not ( n216390 , n216172 );
not ( n216391 , n214610 );
or ( n216392 , n216390 , n216391 );
not ( n216393 , n215953 );
not ( n216394 , n214417 );
or ( n216395 , n216393 , n216394 );
nand ( n216396 , n214416 , n215481 );
nand ( n216397 , n216395 , n216396 );
nand ( n216398 , n216397 , n214458 );
nand ( n216399 , n216392 , n216398 );
nand ( n216400 , n216193 , n213750 );
not ( n216401 , n216400 );
buf ( n216402 , n216196 );
not ( n216403 , n216402 );
not ( n216404 , n216403 );
not ( n216405 , n216404 );
or ( n216406 , n216401 , n216405 );
not ( n216407 , n216193 );
nand ( n216408 , n216407 , n213751 );
nand ( n216409 , n216406 , n216408 );
buf ( n216410 , n36289 );
nand ( n216411 , n216410 , n36292 );
not ( n216412 , n216411 );
not ( n216413 , n216412 );
not ( n216414 , n36997 );
not ( n216415 , n216414 );
or ( n216416 , n216413 , n216415 );
nand ( n216417 , n36997 , n216411 );
nand ( n216418 , n216416 , n216417 );
buf ( n216419 , n216418 );
not ( n216420 , n216419 );
not ( n216421 , n216420 );
buf ( n216422 , n216421 );
and ( n216423 , n216409 , n216422 );
xor ( n216424 , n216399 , n216423 );
not ( n216425 , n216212 );
not ( n216426 , n214798 );
not ( n216427 , n216426 );
or ( n216428 , n216425 , n216427 );
and ( n216429 , n214803 , n215075 );
not ( n216430 , n214803 );
and ( n216431 , n216430 , n215899 );
or ( n216432 , n216429 , n216431 );
nand ( n216433 , n214808 , n216432 );
nand ( n216434 , n216428 , n216433 );
xor ( n216435 , n216424 , n216434 );
xor ( n216436 , n216399 , n216423 );
and ( n216437 , n216436 , n216434 );
and ( n216438 , n216399 , n216423 );
or ( n216439 , n216437 , n216438 );
not ( n216440 , n216221 );
not ( n216441 , n215182 );
or ( n216442 , n216440 , n216441 );
not ( n216443 , n215050 );
not ( n216444 , n215545 );
or ( n216445 , n216443 , n216444 );
nand ( n216446 , n215104 , n214678 );
nand ( n216447 , n216445 , n216446 );
nand ( n216448 , n216447 , n215191 );
nand ( n216449 , n216442 , n216448 );
not ( n216450 , n216283 );
not ( n216451 , n215773 );
or ( n216452 , n216450 , n216451 );
not ( n216453 , n214357 );
not ( n216454 , n215512 );
or ( n216455 , n216453 , n216454 );
nand ( n216456 , n215511 , n215131 );
nand ( n216457 , n216455 , n216456 );
buf ( n216458 , n215327 );
nand ( n216459 , n216457 , n216458 );
nand ( n216460 , n216452 , n216459 );
xor ( n216461 , n216449 , n216460 );
not ( n216462 , n214164 );
not ( n216463 , n213917 );
not ( n216464 , n214145 );
and ( n216465 , n216463 , n216464 );
and ( n216466 , n209248 , n215054 );
nor ( n216467 , n216465 , n216466 );
not ( n216468 , n216467 );
not ( n216469 , n216468 );
or ( n216470 , n216462 , n216469 );
nand ( n216471 , n216144 , n214893 );
nand ( n216472 , n216470 , n216471 );
not ( n216473 , n216472 );
not ( n216474 , n216473 );
not ( n216475 , n215272 );
not ( n216476 , n214190 );
or ( n216477 , n216475 , n216476 );
nand ( n216478 , n214468 , n214131 );
nand ( n216479 , n216477 , n216478 );
and ( n216480 , n216479 , n215966 );
not ( n216481 , n213894 );
nor ( n216482 , n216481 , n216157 );
nor ( n216483 , n216480 , n216482 );
not ( n216484 , n216483 );
not ( n216485 , n216484 );
or ( n216486 , n216474 , n216485 );
or ( n216487 , n216473 , n216484 );
nand ( n216488 , n216486 , n216487 );
xor ( n216489 , n216461 , n216488 );
xor ( n216490 , n216449 , n216460 );
and ( n216491 , n216490 , n216488 );
and ( n216492 , n216449 , n216460 );
or ( n216493 , n216491 , n216492 );
xor ( n216494 , n216373 , n216377 );
xor ( n216495 , n216361 , n216489 );
not ( n216496 , n213874 );
not ( n216497 , n216267 );
or ( n216498 , n216496 , n216497 );
not ( n216499 , n216262 );
not ( n216500 , n41396 );
not ( n216501 , n216500 );
or ( n216502 , n216499 , n216501 );
nand ( n216503 , n41396 , n216265 );
nand ( n216504 , n216502 , n216503 );
nand ( n216505 , n216504 , n213058 );
nand ( n216506 , n216498 , n216505 );
xor ( n216507 , n216495 , n216506 );
xor ( n216508 , n216494 , n216507 );
xor ( n216509 , n216385 , n216508 );
xor ( n216510 , n216509 , n216389 );
xor ( n216511 , n216385 , n216508 );
and ( n216512 , n216511 , n216389 );
and ( n216513 , n216385 , n216508 );
or ( n216514 , n216512 , n216513 );
not ( n216515 , n213784 );
not ( n216516 , n216313 );
or ( n216517 , n216515 , n216516 );
not ( n216518 , n213382 );
not ( n216519 , n41249 );
not ( n216520 , n216519 );
not ( n216521 , n216520 );
or ( n216522 , n216518 , n216521 );
nand ( n216523 , n216519 , n213381 );
nand ( n216524 , n216522 , n216523 );
nand ( n216525 , n216524 , n213912 );
nand ( n216526 , n216517 , n216525 );
xor ( n216527 , n216365 , n216526 );
not ( n216528 , n216239 );
not ( n216529 , n215333 );
not ( n216530 , n30962 );
not ( n216531 , n216530 );
or ( n216532 , n216529 , n216531 );
nand ( n216533 , n30962 , n216037 );
nand ( n216534 , n216532 , n216533 );
not ( n216535 , n216534 );
or ( n216536 , n216528 , n216535 );
nand ( n216537 , n216245 , n214717 );
nand ( n216538 , n216536 , n216537 );
not ( n216539 , n213498 );
not ( n216540 , n213735 );
not ( n216541 , n208839 );
buf ( n216542 , n216541 );
not ( n216543 , n216542 );
not ( n216544 , n216543 );
or ( n216545 , n216540 , n216544 );
nand ( n216546 , n215616 , n213732 );
nand ( n216547 , n216545 , n216546 );
not ( n216548 , n216547 );
or ( n216549 , n216539 , n216548 );
nand ( n216550 , n216343 , n213577 );
nand ( n216551 , n216549 , n216550 );
xor ( n216552 , n216538 , n216551 );
not ( n216553 , n214694 );
not ( n216554 , n215290 );
not ( n216555 , n215228 );
not ( n216556 , n216555 );
or ( n216557 , n216554 , n216556 );
nand ( n216558 , n215228 , n215289 );
nand ( n216559 , n216557 , n216558 );
not ( n216560 , n216559 );
or ( n216561 , n216553 , n216560 );
not ( n216562 , n216298 );
nand ( n216563 , n216295 , n216562 );
nand ( n216564 , n216561 , n216563 );
xor ( n216565 , n216552 , n216564 );
xor ( n216566 , n216527 , n216565 );
xor ( n216567 , n216381 , n216566 );
not ( n216568 , n216418 );
buf ( n216569 , n216568 );
and ( n216570 , n213751 , n216569 );
not ( n216571 , n213751 );
buf ( n216572 , n216419 );
and ( n216573 , n216571 , n216572 );
nor ( n216574 , n216570 , n216573 );
not ( n216575 , n216574 );
not ( n216576 , n216412 );
not ( n216577 , n216414 );
or ( n216578 , n216576 , n216577 );
nand ( n216579 , n216578 , n216417 );
and ( n216580 , n216193 , n216579 );
not ( n216581 , n216193 );
and ( n216582 , n216581 , n216568 );
nor ( n216583 , n216580 , n216582 );
nand ( n216584 , n216199 , n216583 );
buf ( n216585 , n216584 );
not ( n216586 , n216585 );
not ( n216587 , n216586 );
or ( n216588 , n216575 , n216587 );
and ( n216589 , n213126 , n216569 );
not ( n216590 , n213126 );
buf ( n216591 , n216579 );
not ( n216592 , n216591 );
buf ( n216593 , n216592 );
not ( n216594 , n216593 );
and ( n216595 , n216590 , n216594 );
nor ( n216596 , n216589 , n216595 );
not ( n216597 , n216596 );
not ( n216598 , n216200 );
nand ( n216599 , n216597 , n216598 );
nand ( n216600 , n216588 , n216599 );
xor ( n216601 , n216600 , n216179 );
not ( n216602 , n213206 );
not ( n216603 , n216046 );
not ( n216604 , n216603 );
not ( n216605 , n215388 );
and ( n216606 , n216604 , n216605 );
not ( n216607 , n41608 );
not ( n216608 , n216607 );
and ( n216609 , n216608 , n215600 );
nor ( n216610 , n216606 , n216609 );
not ( n216611 , n216610 );
not ( n216612 , n216611 );
or ( n216613 , n216602 , n216612 );
nand ( n216614 , n216236 , n215605 );
nand ( n216615 , n216613 , n216614 );
xor ( n216616 , n216601 , n216615 );
xor ( n216617 , n216369 , n216616 );
not ( n216618 , n216331 );
not ( n216619 , n216066 );
not ( n216620 , n216619 );
or ( n216621 , n216618 , n216620 );
not ( n216622 , n213583 );
not ( n216623 , n216067 );
not ( n216624 , n216623 );
not ( n216625 , n216624 );
or ( n216626 , n216622 , n216625 );
not ( n216627 , n216014 );
nand ( n216628 , n216627 , n214134 );
nand ( n216629 , n216626 , n216628 );
not ( n216630 , n215788 );
nand ( n216631 , n216629 , n216630 );
nand ( n216632 , n216621 , n216631 );
xor ( n216633 , n216632 , n216228 );
xor ( n216634 , n216633 , n216435 );
xor ( n216635 , n216617 , n216634 );
xor ( n216636 , n216567 , n216635 );
xor ( n216637 , n216636 , n216259 );
xor ( n216638 , n216637 , n216510 );
xor ( n216639 , n216636 , n216259 );
and ( n216640 , n216639 , n216510 );
and ( n216641 , n216636 , n216259 );
or ( n216642 , n216640 , n216641 );
xor ( n216643 , n216600 , n216179 );
and ( n216644 , n216643 , n216615 );
and ( n216645 , n216600 , n216179 );
or ( n216646 , n216644 , n216645 );
xor ( n216647 , n216538 , n216551 );
and ( n216648 , n216647 , n216564 );
and ( n216649 , n216538 , n216551 );
or ( n216650 , n216648 , n216649 );
xor ( n216651 , n216632 , n216228 );
and ( n216652 , n216651 , n216435 );
and ( n216653 , n216632 , n216228 );
or ( n216654 , n216652 , n216653 );
xor ( n216655 , n216361 , n216489 );
and ( n216656 , n216655 , n216506 );
and ( n216657 , n216361 , n216489 );
or ( n216658 , n216656 , n216657 );
xor ( n216659 , n216365 , n216526 );
and ( n216660 , n216659 , n216565 );
and ( n216661 , n216365 , n216526 );
or ( n216662 , n216660 , n216661 );
xor ( n216663 , n216369 , n216616 );
and ( n216664 , n216663 , n216634 );
and ( n216665 , n216369 , n216616 );
or ( n216666 , n216664 , n216665 );
xor ( n216667 , n216373 , n216377 );
and ( n216668 , n216667 , n216507 );
and ( n216669 , n216373 , n216377 );
or ( n216670 , n216668 , n216669 );
xor ( n216671 , n216381 , n216566 );
and ( n216672 , n216671 , n216635 );
and ( n216673 , n216381 , n216566 );
or ( n216674 , n216672 , n216673 );
not ( n216675 , n214370 );
and ( n216676 , n41894 , n214404 );
not ( n216677 , n41894 );
and ( n216678 , n216677 , n214688 );
or ( n216679 , n216676 , n216678 );
not ( n216680 , n216679 );
or ( n216681 , n216675 , n216680 );
not ( n216682 , n214551 );
or ( n216683 , n216467 , n216682 );
nand ( n216684 , n216681 , n216683 );
not ( n216685 , n216397 );
not ( n216686 , n214449 );
or ( n216687 , n216685 , n216686 );
and ( n216688 , n30292 , n214586 );
not ( n216689 , n30292 );
and ( n216690 , n216689 , n214759 );
or ( n216691 , n216688 , n216690 );
nand ( n216692 , n216691 , n214457 );
nand ( n216693 , n216687 , n216692 );
xor ( n216694 , n216684 , n216693 );
not ( n216695 , n213750 );
and ( n216696 , n216418 , n36670 );
not ( n216697 , n216418 );
not ( n216698 , n36670 );
and ( n216699 , n216697 , n216698 );
nor ( n216700 , n216696 , n216699 );
not ( n216701 , n216700 );
nor ( n216702 , n216695 , n216701 );
xor ( n216703 , n216694 , n216702 );
xor ( n216704 , n216684 , n216693 );
and ( n216705 , n216704 , n216702 );
and ( n216706 , n216684 , n216693 );
or ( n216707 , n216705 , n216706 );
not ( n216708 , n216432 );
not ( n216709 , n214799 );
or ( n216710 , n216708 , n216709 );
not ( n216711 , n215268 );
not ( n216712 , n214783 );
or ( n216713 , n216711 , n216712 );
nand ( n216714 , n214786 , n216170 );
nand ( n216715 , n216713 , n216714 );
nand ( n216716 , n214808 , n216715 );
nand ( n216717 , n216710 , n216716 );
not ( n216718 , n216447 );
not ( n216719 , n215183 );
or ( n216720 , n216718 , n216719 );
not ( n216721 , n216208 );
not ( n216722 , n215164 );
or ( n216723 , n216721 , n216722 );
nand ( n216724 , n215104 , n216207 );
nand ( n216725 , n216723 , n216724 );
nand ( n216726 , n216725 , n215191 );
nand ( n216727 , n216720 , n216726 );
xor ( n216728 , n216717 , n216727 );
not ( n216729 , n216457 );
not ( n216730 , n215773 );
not ( n216731 , n216730 );
not ( n216732 , n216731 );
or ( n216733 , n216729 , n216732 );
not ( n216734 , n214537 );
not ( n216735 , n215765 );
or ( n216736 , n216734 , n216735 );
nand ( n216737 , n215766 , n214899 );
nand ( n216738 , n216736 , n216737 );
nand ( n216739 , n216738 , n215762 );
nand ( n216740 , n216733 , n216739 );
xor ( n216741 , n216728 , n216740 );
xor ( n216742 , n216717 , n216727 );
and ( n216743 , n216742 , n216740 );
and ( n216744 , n216717 , n216727 );
or ( n216745 , n216743 , n216744 );
not ( n216746 , n215966 );
and ( n216747 , n30997 , n214131 );
not ( n216748 , n30997 );
and ( n216749 , n216748 , n215272 );
or ( n216750 , n216747 , n216749 );
not ( n216751 , n216750 );
or ( n216752 , n216746 , n216751 );
nand ( n216753 , n216479 , n213894 );
nand ( n216754 , n216752 , n216753 );
not ( n216755 , n216472 );
nor ( n216756 , n216755 , n216483 );
xor ( n216757 , n216754 , n216756 );
or ( n216758 , n216585 , n216596 );
not ( n216759 , n213347 );
not ( n216760 , n216420 );
or ( n216761 , n216759 , n216760 );
not ( n216762 , n216569 );
nand ( n216763 , n216762 , n214616 );
nand ( n216764 , n216761 , n216763 );
not ( n216765 , n216764 );
or ( n216766 , n216765 , n216200 );
nand ( n216767 , n216758 , n216766 );
xor ( n216768 , n216757 , n216767 );
xor ( n216769 , n216650 , n216768 );
not ( n216770 , n214717 );
not ( n216771 , n216534 );
or ( n216772 , n216770 , n216771 );
not ( n216773 , n215113 );
not ( n216774 , n215845 );
or ( n216775 , n216773 , n216774 );
nand ( n216776 , n208725 , n216037 );
nand ( n216777 , n216775 , n216776 );
nand ( n216778 , n216777 , n216239 );
nand ( n216779 , n216772 , n216778 );
not ( n216780 , n214564 );
not ( n216781 , n213960 );
not ( n216782 , n41700 );
not ( n216783 , n216782 );
or ( n216784 , n216781 , n216783 );
nand ( n216785 , n41700 , n214570 );
nand ( n216786 , n216784 , n216785 );
not ( n216787 , n216786 );
or ( n216788 , n216780 , n216787 );
or ( n216789 , n216610 , n214085 );
nand ( n216790 , n216788 , n216789 );
xor ( n216791 , n216779 , n216790 );
not ( n216792 , n216629 );
not ( n216793 , n216324 );
or ( n216794 , n216792 , n216793 );
not ( n216795 , n216630 );
not ( n216796 , n216795 );
not ( n216797 , n214960 );
not ( n216798 , n216068 );
or ( n216799 , n216797 , n216798 );
nand ( n216800 , n216014 , n214956 );
nand ( n216801 , n216799 , n216800 );
nand ( n216802 , n216796 , n216801 );
nand ( n216803 , n216794 , n216802 );
xor ( n216804 , n216791 , n216803 );
xor ( n216805 , n216769 , n216804 );
xor ( n216806 , n216805 , n216666 );
not ( n216807 , n216299 );
not ( n216808 , n216559 );
or ( n216809 , n216807 , n216808 );
not ( n216810 , n215289 );
not ( n216811 , n216810 );
not ( n216812 , n215833 );
or ( n216813 , n216811 , n216812 );
nand ( n216814 , n41716 , n215289 );
nand ( n216815 , n216813 , n216814 );
nand ( n216816 , n216815 , n214694 );
nand ( n216817 , n216809 , n216816 );
xor ( n216818 , n216817 , n216703 );
xor ( n216819 , n216818 , n216439 );
xor ( n216820 , n216654 , n216819 );
not ( n216821 , n213498 );
not ( n216822 , n213735 );
not ( n216823 , n216261 );
or ( n216824 , n216822 , n216823 );
nand ( n216825 , n215796 , n213732 );
nand ( n216826 , n216824 , n216825 );
not ( n216827 , n216826 );
or ( n216828 , n216821 , n216827 );
nand ( n216829 , n216547 , n213577 );
nand ( n216830 , n216828 , n216829 );
xor ( n216831 , n216493 , n216830 );
xor ( n216832 , n216831 , n216741 );
xor ( n216833 , n216820 , n216832 );
xor ( n216834 , n216806 , n216833 );
xor ( n216835 , n216805 , n216666 );
and ( n216836 , n216835 , n216833 );
and ( n216837 , n216805 , n216666 );
or ( n216838 , n216836 , n216837 );
xor ( n216839 , n216670 , n216674 );
xor ( n216840 , n216658 , n216662 );
not ( n216841 , n213058 );
not ( n216842 , n216262 );
not ( n216843 , n216307 );
or ( n216844 , n216842 , n216843 );
nand ( n216845 , n216311 , n216265 );
nand ( n216846 , n216844 , n216845 );
not ( n216847 , n216846 );
or ( n216848 , n216841 , n216847 );
nand ( n216849 , n216504 , n213874 );
nand ( n216850 , n216848 , n216849 );
not ( n216851 , n213784 );
not ( n216852 , n216524 );
or ( n216853 , n216851 , n216852 );
not ( n216854 , n213382 );
not ( n216855 , n208164 );
not ( n216856 , n216855 );
or ( n216857 , n216854 , n216856 );
not ( n216858 , n40886 );
not ( n216859 , n216858 );
nand ( n216860 , n216859 , n213381 );
nand ( n216861 , n216857 , n216860 );
nand ( n216862 , n216861 , n213912 );
nand ( n216863 , n216853 , n216862 );
xor ( n216864 , n216850 , n216863 );
xor ( n216865 , n216864 , n216646 );
xor ( n216866 , n216840 , n216865 );
xor ( n216867 , n216839 , n216866 );
xor ( n216868 , n216670 , n216674 );
and ( n216869 , n216868 , n216866 );
and ( n216870 , n216670 , n216674 );
or ( n216871 , n216869 , n216870 );
xor ( n216872 , n216834 , n216514 );
xor ( n216873 , n216872 , n216867 );
xor ( n216874 , n216834 , n216514 );
and ( n216875 , n216874 , n216867 );
and ( n216876 , n216834 , n216514 );
or ( n216877 , n216875 , n216876 );
xor ( n216878 , n216754 , n216756 );
and ( n216879 , n216878 , n216767 );
and ( n216880 , n216754 , n216756 );
or ( n216881 , n216879 , n216880 );
xor ( n216882 , n216779 , n216790 );
and ( n216883 , n216882 , n216803 );
and ( n216884 , n216779 , n216790 );
or ( n216885 , n216883 , n216884 );
xor ( n216886 , n216817 , n216703 );
and ( n216887 , n216886 , n216439 );
and ( n216888 , n216817 , n216703 );
or ( n216889 , n216887 , n216888 );
xor ( n216890 , n216493 , n216830 );
and ( n216891 , n216890 , n216741 );
and ( n216892 , n216493 , n216830 );
or ( n216893 , n216891 , n216892 );
xor ( n216894 , n216850 , n216863 );
and ( n216895 , n216894 , n216646 );
and ( n216896 , n216850 , n216863 );
or ( n216897 , n216895 , n216896 );
xor ( n216898 , n216650 , n216768 );
and ( n216899 , n216898 , n216804 );
and ( n216900 , n216650 , n216768 );
or ( n216901 , n216899 , n216900 );
xor ( n216902 , n216654 , n216819 );
and ( n216903 , n216902 , n216832 );
and ( n216904 , n216654 , n216819 );
or ( n216905 , n216903 , n216904 );
xor ( n216906 , n216658 , n216662 );
and ( n216907 , n216906 , n216865 );
and ( n216908 , n216658 , n216662 );
or ( n216909 , n216907 , n216908 );
not ( n216910 , n216698 );
nand ( n216911 , n216910 , n213750 );
not ( n216912 , n216911 );
not ( n216913 , n216569 );
or ( n216914 , n216912 , n216913 );
nand ( n216915 , n216698 , n213751 );
nand ( n216916 , n216914 , n216915 );
not ( n216917 , n37500 );
nand ( n216918 , n216917 , n37492 , n37004 );
buf ( n216919 , n36305 );
buf ( n216920 , n35282 );
nand ( n216921 , n216919 , n216920 );
not ( n216922 , n216921 );
and ( n216923 , n216918 , n216922 );
not ( n216924 , n216918 );
and ( n216925 , n216924 , n216921 );
nor ( n216926 , n216923 , n216925 );
buf ( n216927 , n216926 );
buf ( n216928 , n216927 );
buf ( n216929 , n216928 );
and ( n216930 , n216916 , n216929 );
not ( n216931 , n216715 );
not ( n216932 , n216204 );
or ( n216933 , n216931 , n216932 );
buf ( n216934 , n215953 );
not ( n216935 , n216934 );
not ( n216936 , n214783 );
or ( n216937 , n216935 , n216936 );
buf ( n216938 , n214803 );
not ( n216939 , n216938 );
not ( n216940 , n216934 );
nand ( n216941 , n216939 , n216940 );
nand ( n216942 , n216937 , n216941 );
nand ( n216943 , n214808 , n216942 );
nand ( n216944 , n216933 , n216943 );
xor ( n216945 , n216930 , n216944 );
not ( n216946 , n216725 );
not ( n216947 , n215183 );
or ( n216948 , n216946 , n216947 );
not ( n216949 , n215075 );
not ( n216950 , n215105 );
or ( n216951 , n216949 , n216950 );
nand ( n216952 , n215104 , n215899 );
nand ( n216953 , n216951 , n216952 );
nand ( n216954 , n215550 , n216953 );
nand ( n216955 , n216948 , n216954 );
xor ( n216956 , n216945 , n216955 );
xor ( n216957 , n216930 , n216944 );
and ( n216958 , n216957 , n216955 );
and ( n216959 , n216930 , n216944 );
or ( n216960 , n216958 , n216959 );
not ( n216961 , n216738 );
not ( n216962 , n215773 );
or ( n216963 , n216961 , n216962 );
not ( n216964 , n214678 );
not ( n216965 , n216964 );
not ( n216966 , n215569 );
or ( n216967 , n216965 , n216966 );
not ( n216968 , n215765 );
nand ( n216969 , n216968 , n214678 );
nand ( n216970 , n216967 , n216969 );
nand ( n216971 , n215327 , n216970 );
nand ( n216972 , n216963 , n216971 );
not ( n216973 , n216764 );
not ( n216974 , n216586 );
or ( n216975 , n216973 , n216974 );
not ( n216976 , n213583 );
not ( n216977 , n216420 );
or ( n216978 , n216976 , n216977 );
nand ( n216979 , n216591 , n214134 );
nand ( n216980 , n216978 , n216979 );
nand ( n216981 , n216980 , n216201 );
nand ( n216982 , n216975 , n216981 );
xor ( n216983 , n216972 , n216982 );
not ( n216984 , n214164 );
buf ( n216985 , n215054 );
not ( n216986 , n216985 );
not ( n216987 , n214464 );
or ( n216988 , n216986 , n216987 );
not ( n216989 , n215955 );
nand ( n216990 , n214468 , n216989 );
nand ( n216991 , n216988 , n216990 );
not ( n216992 , n216991 );
or ( n216993 , n216984 , n216992 );
nand ( n216994 , n216679 , n215963 );
nand ( n216995 , n216993 , n216994 );
not ( n216996 , n216691 );
not ( n216997 , n214449 );
or ( n216998 , n216996 , n216997 );
not ( n216999 , n215117 );
not ( n217000 , n214417 );
or ( n217001 , n216999 , n217000 );
not ( n217002 , n214760 );
nand ( n217003 , n217002 , n213917 );
nand ( n217004 , n217001 , n217003 );
nand ( n217005 , n217004 , n214458 );
nand ( n217006 , n216998 , n217005 );
xor ( n217007 , n216995 , n217006 );
xor ( n217008 , n216983 , n217007 );
xor ( n217009 , n216972 , n216982 );
and ( n217010 , n217009 , n217007 );
and ( n217011 , n216972 , n216982 );
or ( n217012 , n217010 , n217011 );
not ( n217013 , n215966 );
not ( n217014 , n214820 );
not ( n217015 , n214130 );
or ( n217016 , n217014 , n217015 );
not ( n217017 , n215971 );
not ( n217018 , n217017 );
nand ( n217019 , n217018 , n215228 );
nand ( n217020 , n217016 , n217019 );
not ( n217021 , n217020 );
or ( n217022 , n217013 , n217021 );
buf ( n217023 , n213894 );
nand ( n217024 , n216750 , n217023 );
nand ( n217025 , n217022 , n217024 );
not ( n217026 , n214694 );
not ( n217027 , n216810 );
not ( n217028 , n216530 );
or ( n217029 , n217027 , n217028 );
nand ( n217030 , n30962 , n215289 );
nand ( n217031 , n217029 , n217030 );
not ( n217032 , n217031 );
or ( n217033 , n217026 , n217032 );
nand ( n217034 , n216815 , n213718 );
nand ( n217035 , n217033 , n217034 );
xor ( n217036 , n217025 , n217035 );
not ( n217037 , n216801 );
not ( n217038 , n216324 );
or ( n217039 , n217037 , n217038 );
not ( n217040 , n215131 );
not ( n217041 , n216068 );
or ( n217042 , n217040 , n217041 );
not ( n217043 , n216403 );
not ( n217044 , n215131 );
nand ( n217045 , n217043 , n217044 );
nand ( n217046 , n217042 , n217045 );
not ( n217047 , n215788 );
nand ( n217048 , n217046 , n217047 );
nand ( n217049 , n217039 , n217048 );
xor ( n217050 , n217036 , n217049 );
not ( n217051 , n215137 );
not ( n217052 , n213960 );
not ( n217053 , n41563 );
or ( n217054 , n217052 , n217053 );
nand ( n217055 , n216541 , n214570 );
nand ( n217056 , n217054 , n217055 );
not ( n217057 , n217056 );
or ( n217058 , n217051 , n217057 );
nand ( n217059 , n216786 , n214086 );
nand ( n217060 , n217058 , n217059 );
xor ( n217061 , n217060 , n216707 );
not ( n217062 , n214717 );
not ( n217063 , n216777 );
or ( n217064 , n217062 , n217063 );
not ( n217065 , n215333 );
not ( n217066 , n41608 );
not ( n217067 , n217066 );
or ( n217068 , n217065 , n217067 );
nand ( n217069 , n216608 , n216037 );
nand ( n217070 , n217068 , n217069 );
nand ( n217071 , n217070 , n216239 );
nand ( n217072 , n217064 , n217071 );
xor ( n217073 , n217061 , n217072 );
xor ( n217074 , n217050 , n217073 );
xor ( n217075 , n217074 , n216889 );
not ( n217076 , n216928 );
and ( n217077 , n213751 , n217076 );
not ( n217078 , n213751 );
not ( n217079 , n216927 );
not ( n217080 , n217079 );
and ( n217081 , n217078 , n217080 );
nor ( n217082 , n217077 , n217081 );
not ( n217083 , n217082 );
not ( n217084 , n216927 );
nand ( n217085 , n217084 , n216698 );
nand ( n217086 , n216927 , n216910 );
nand ( n217087 , n217085 , n217086 , n216701 );
buf ( n217088 , n217087 );
not ( n217089 , n217088 );
not ( n217090 , n217089 );
or ( n217091 , n217083 , n217090 );
not ( n217092 , n213126 );
buf ( n217093 , n217084 );
not ( n217094 , n217093 );
or ( n217095 , n217092 , n217094 );
nand ( n217096 , n216928 , n216076 );
nand ( n217097 , n217095 , n217096 );
buf ( n217098 , n216701 );
not ( n217099 , n217098 );
nand ( n217100 , n217097 , n217099 );
nand ( n217101 , n217091 , n217100 );
xor ( n217102 , n217101 , n216745 );
xor ( n217103 , n217102 , n216881 );
xor ( n217104 , n217103 , n216893 );
xor ( n217105 , n217104 , n216897 );
xor ( n217106 , n217075 , n217105 );
xor ( n217107 , n217106 , n216905 );
xor ( n217108 , n217075 , n217105 );
and ( n217109 , n217108 , n216905 );
and ( n217110 , n217075 , n217105 );
or ( n217111 , n217109 , n217110 );
not ( n217112 , n213912 );
not ( n217113 , n213382 );
not ( n217114 , n208258 );
not ( n217115 , n217114 );
buf ( n217116 , n217115 );
not ( n217117 , n217116 );
or ( n217118 , n217113 , n217117 );
not ( n217119 , n217114 );
not ( n217120 , n217119 );
nand ( n217121 , n217120 , n213381 );
nand ( n217122 , n217118 , n217121 );
not ( n217123 , n217122 );
or ( n217124 , n217112 , n217123 );
nand ( n217125 , n216861 , n213784 );
nand ( n217126 , n217124 , n217125 );
xor ( n217127 , n217126 , n216885 );
not ( n217128 , n216336 );
not ( n217129 , n213735 );
not ( n217130 , n41397 );
not ( n217131 , n217130 );
or ( n217132 , n217129 , n217131 );
not ( n217133 , n215989 );
nand ( n217134 , n217133 , n213732 );
nand ( n217135 , n217132 , n217134 );
not ( n217136 , n217135 );
or ( n217137 , n217128 , n217136 );
nand ( n217138 , n216826 , n213577 );
nand ( n217139 , n217137 , n217138 );
xor ( n217140 , n217127 , n217139 );
xor ( n217141 , n217140 , n216901 );
buf ( n217142 , n213058 );
not ( n217143 , n217142 );
not ( n217144 , n216262 );
not ( n217145 , n41249 );
or ( n217146 , n217144 , n217145 );
buf ( n217147 , n41249 );
not ( n217148 , n217147 );
nand ( n217149 , n217148 , n216265 );
nand ( n217150 , n217146 , n217149 );
not ( n217151 , n217150 );
or ( n217152 , n217143 , n217151 );
nand ( n217153 , n216846 , n213874 );
nand ( n217154 , n217152 , n217153 );
xor ( n217155 , n216956 , n217154 );
xor ( n217156 , n217155 , n217008 );
xor ( n217157 , n217141 , n217156 );
xor ( n217158 , n216909 , n217157 );
xor ( n217159 , n217158 , n216838 );
xor ( n217160 , n216909 , n217157 );
and ( n217161 , n217160 , n216838 );
and ( n217162 , n216909 , n217157 );
or ( n217163 , n217161 , n217162 );
xor ( n217164 , n217107 , n216871 );
xor ( n217165 , n217164 , n217159 );
xor ( n217166 , n217107 , n216871 );
and ( n217167 , n217166 , n217159 );
and ( n217168 , n217107 , n216871 );
or ( n217169 , n217167 , n217168 );
xor ( n217170 , n217060 , n216707 );
and ( n217171 , n217170 , n217072 );
and ( n217172 , n217060 , n216707 );
or ( n217173 , n217171 , n217172 );
xor ( n217174 , n217025 , n217035 );
and ( n217175 , n217174 , n217049 );
and ( n217176 , n217025 , n217035 );
or ( n217177 , n217175 , n217176 );
xor ( n217178 , n217101 , n216745 );
and ( n217179 , n217178 , n216881 );
and ( n217180 , n217101 , n216745 );
or ( n217181 , n217179 , n217180 );
xor ( n217182 , n216956 , n217154 );
and ( n217183 , n217182 , n217008 );
and ( n217184 , n216956 , n217154 );
or ( n217185 , n217183 , n217184 );
xor ( n217186 , n217126 , n216885 );
and ( n217187 , n217186 , n217139 );
and ( n217188 , n217126 , n216885 );
or ( n217189 , n217187 , n217188 );
xor ( n217190 , n217050 , n217073 );
and ( n217191 , n217190 , n216889 );
and ( n217192 , n217050 , n217073 );
or ( n217193 , n217191 , n217192 );
xor ( n217194 , n217103 , n216893 );
and ( n217195 , n217194 , n216897 );
and ( n217196 , n217103 , n216893 );
or ( n217197 , n217195 , n217196 );
xor ( n217198 , n217140 , n216901 );
and ( n217199 , n217198 , n217156 );
and ( n217200 , n217140 , n216901 );
or ( n217201 , n217199 , n217200 );
not ( n217202 , n217004 );
not ( n217203 , n214610 );
or ( n217204 , n217202 , n217203 );
and ( n217205 , n41894 , n214418 );
not ( n217206 , n41894 );
and ( n217207 , n217206 , n214417 );
nor ( n217208 , n217205 , n217207 );
nand ( n217209 , n214458 , n217208 );
nand ( n217210 , n217204 , n217209 );
not ( n217211 , n216942 );
not ( n217212 , n216426 );
or ( n217213 , n217211 , n217212 );
not ( n217214 , n30292 );
not ( n217215 , n214783 );
or ( n217216 , n217214 , n217215 );
nand ( n217217 , n214786 , n216139 );
nand ( n217218 , n217216 , n217217 );
nand ( n217219 , n214808 , n217218 );
nand ( n217220 , n217213 , n217219 );
xor ( n217221 , n217210 , n217220 );
and ( n217222 , n37686 , n37600 );
not ( n217223 , n37686 );
and ( n217224 , n217223 , n37599 );
nor ( n217225 , n217222 , n217224 );
and ( n217226 , n217225 , n217084 );
not ( n217227 , n217225 );
and ( n217228 , n217227 , n216927 );
nor ( n217229 , n217226 , n217228 );
not ( n217230 , n217229 );
and ( n217231 , n217230 , n213750 );
xor ( n217232 , n217221 , n217231 );
xor ( n217233 , n217210 , n217220 );
and ( n217234 , n217233 , n217231 );
and ( n217235 , n217210 , n217220 );
or ( n217236 , n217234 , n217235 );
not ( n217237 , n216953 );
not ( n217238 , n215183 );
or ( n217239 , n217237 , n217238 );
not ( n217240 , n215268 );
not ( n217241 , n215105 );
or ( n217242 , n217240 , n217241 );
nand ( n217243 , n215165 , n216170 );
nand ( n217244 , n217242 , n217243 );
nand ( n217245 , n217244 , n215191 );
nand ( n217246 , n217239 , n217245 );
not ( n217247 , n216970 );
not ( n217248 , n215773 );
or ( n217249 , n217247 , n217248 );
and ( n217250 , n216208 , n216968 );
not ( n217251 , n216208 );
and ( n217252 , n217251 , n215512 );
nor ( n217253 , n217250 , n217252 );
nand ( n217254 , n216458 , n217253 );
nand ( n217255 , n217249 , n217254 );
xor ( n217256 , n217246 , n217255 );
and ( n217257 , n216995 , n217006 );
xor ( n217258 , n217256 , n217257 );
xor ( n217259 , n217246 , n217255 );
and ( n217260 , n217259 , n217257 );
and ( n217261 , n217246 , n217255 );
or ( n217262 , n217260 , n217261 );
not ( n217263 , n216336 );
not ( n217264 , n213735 );
not ( n217265 , n216307 );
or ( n217266 , n217264 , n217265 );
nand ( n217267 , n216311 , n213732 );
nand ( n217268 , n217266 , n217267 );
not ( n217269 , n217268 );
or ( n217270 , n217263 , n217269 );
nand ( n217271 , n217135 , n213577 );
nand ( n217272 , n217270 , n217271 );
xor ( n217273 , n217173 , n217272 );
not ( n217274 , n214164 );
not ( n217275 , n215955 );
not ( n217276 , n216290 );
or ( n217277 , n217275 , n217276 );
not ( n217278 , n30997 );
not ( n217279 , n217278 );
not ( n217280 , n216985 );
nand ( n217281 , n217279 , n217280 );
nand ( n217282 , n217277 , n217281 );
not ( n217283 , n217282 );
or ( n217284 , n217274 , n217283 );
nand ( n217285 , n216991 , n215963 );
nand ( n217286 , n217284 , n217285 );
not ( n217287 , n216980 );
not ( n217288 , n216584 );
buf ( n217289 , n217288 );
not ( n217290 , n217289 );
or ( n217291 , n217287 , n217290 );
not ( n217292 , n214956 );
not ( n217293 , n216420 );
or ( n217294 , n217292 , n217293 );
nand ( n217295 , n216419 , n214960 );
nand ( n217296 , n217294 , n217295 );
nand ( n217297 , n216598 , n217296 );
nand ( n217298 , n217291 , n217297 );
xor ( n217299 , n217286 , n217298 );
not ( n217300 , n214717 );
not ( n217301 , n217070 );
or ( n217302 , n217300 , n217301 );
not ( n217303 , n215333 );
not ( n217304 , n215820 );
or ( n217305 , n217303 , n217304 );
nand ( n217306 , n41701 , n216037 );
nand ( n217307 , n217305 , n217306 );
nand ( n217308 , n217307 , n216239 );
nand ( n217309 , n217302 , n217308 );
xor ( n217310 , n217299 , n217309 );
xor ( n217311 , n217273 , n217310 );
not ( n217312 , n217142 );
not ( n217313 , n216262 );
not ( n217314 , n216859 );
not ( n217315 , n217314 );
or ( n217316 , n217313 , n217315 );
not ( n217317 , n208164 );
not ( n217318 , n217317 );
nand ( n217319 , n217318 , n216265 );
nand ( n217320 , n217316 , n217319 );
not ( n217321 , n217320 );
or ( n217322 , n217312 , n217321 );
nand ( n217323 , n217150 , n213874 );
nand ( n217324 , n217322 , n217323 );
xor ( n217325 , n217177 , n217324 );
not ( n217326 , n213784 );
not ( n217327 , n217122 );
or ( n217328 , n217326 , n217327 );
not ( n217329 , n213381 );
not ( n217330 , n41069 );
not ( n217331 , n217330 );
not ( n217332 , n217331 );
or ( n217333 , n217329 , n217332 );
nand ( n217334 , n217330 , n213382 );
nand ( n217335 , n217333 , n217334 );
nand ( n217336 , n217335 , n213912 );
nand ( n217337 , n217328 , n217336 );
xor ( n217338 , n217325 , n217337 );
xor ( n217339 , n217311 , n217338 );
xor ( n217340 , n217339 , n217193 );
xor ( n217341 , n217311 , n217338 );
and ( n217342 , n217341 , n217193 );
and ( n217343 , n217311 , n217338 );
or ( n217344 , n217342 , n217343 );
not ( n217345 , n214694 );
not ( n217346 , n216810 );
not ( n217347 , n208726 );
or ( n217348 , n217346 , n217347 );
nand ( n217349 , n208725 , n215289 );
nand ( n217350 , n217348 , n217349 );
not ( n217351 , n217350 );
or ( n217352 , n217345 , n217351 );
nand ( n217353 , n217031 , n213718 );
nand ( n217354 , n217352 , n217353 );
not ( n217355 , n217046 );
not ( n217356 , n216065 );
or ( n217357 , n217355 , n217356 );
not ( n217358 , n214537 );
not ( n217359 , n216624 );
or ( n217360 , n217358 , n217359 );
nand ( n217361 , n216015 , n214899 );
nand ( n217362 , n217360 , n217361 );
nand ( n217363 , n216332 , n217362 );
nand ( n217364 , n217357 , n217363 );
xor ( n217365 , n217354 , n217364 );
not ( n217366 , n217020 );
not ( n217367 , n217023 );
or ( n217368 , n217366 , n217367 );
not ( n217369 , n217017 );
not ( n217370 , n214642 );
or ( n217371 , n217369 , n217370 );
nand ( n217372 , n41716 , n215971 );
nand ( n217373 , n217371 , n217372 );
not ( n217374 , n217373 );
or ( n217375 , n217374 , n213749 );
nand ( n217376 , n217368 , n217375 );
xor ( n217377 , n217365 , n217376 );
xor ( n217378 , n217377 , n217181 );
not ( n217379 , n217097 );
not ( n217380 , n217088 );
not ( n217381 , n217380 );
or ( n217382 , n217379 , n217381 );
not ( n217383 , n213347 );
not ( n217384 , n217093 );
or ( n217385 , n217383 , n217384 );
nand ( n217386 , n216929 , n214616 );
nand ( n217387 , n217385 , n217386 );
buf ( n217388 , n217099 );
nand ( n217389 , n217387 , n217388 );
nand ( n217390 , n217382 , n217389 );
xor ( n217391 , n217390 , n216960 );
not ( n217392 , n213206 );
not ( n217393 , n213960 );
not ( n217394 , n215796 );
not ( n217395 , n217394 );
or ( n217396 , n217393 , n217395 );
not ( n217397 , n213261 );
nand ( n217398 , n215796 , n217397 );
nand ( n217399 , n217396 , n217398 );
not ( n217400 , n217399 );
or ( n217401 , n217392 , n217400 );
nand ( n217402 , n217056 , n215605 );
nand ( n217403 , n217401 , n217402 );
xor ( n217404 , n217391 , n217403 );
xor ( n217405 , n217378 , n217404 );
xor ( n217406 , n217197 , n217405 );
xor ( n217407 , n217406 , n217201 );
xor ( n217408 , n217197 , n217405 );
and ( n217409 , n217408 , n217201 );
and ( n217410 , n217197 , n217405 );
or ( n217411 , n217409 , n217410 );
xor ( n217412 , n217012 , n217258 );
xor ( n217413 , n217412 , n217232 );
xor ( n217414 , n217413 , n217189 );
xor ( n217415 , n217414 , n217185 );
xor ( n217416 , n217415 , n217340 );
xor ( n217417 , n217416 , n217111 );
xor ( n217418 , n217415 , n217340 );
and ( n217419 , n217418 , n217111 );
and ( n217420 , n217415 , n217340 );
or ( n217421 , n217419 , n217420 );
xor ( n217422 , n217407 , n217417 );
xor ( n217423 , n217422 , n217163 );
xor ( n217424 , n217407 , n217417 );
and ( n217425 , n217424 , n217163 );
and ( n217426 , n217407 , n217417 );
or ( n217427 , n217425 , n217426 );
xor ( n217428 , n217286 , n217298 );
and ( n217429 , n217428 , n217309 );
and ( n217430 , n217286 , n217298 );
or ( n217431 , n217429 , n217430 );
xor ( n217432 , n217354 , n217364 );
and ( n217433 , n217432 , n217376 );
and ( n217434 , n217354 , n217364 );
or ( n217435 , n217433 , n217434 );
xor ( n217436 , n217390 , n216960 );
and ( n217437 , n217436 , n217403 );
and ( n217438 , n217390 , n216960 );
or ( n217439 , n217437 , n217438 );
xor ( n217440 , n217012 , n217258 );
and ( n217441 , n217440 , n217232 );
and ( n217442 , n217012 , n217258 );
or ( n217443 , n217441 , n217442 );
xor ( n217444 , n217177 , n217324 );
and ( n217445 , n217444 , n217337 );
and ( n217446 , n217177 , n217324 );
or ( n217447 , n217445 , n217446 );
xor ( n217448 , n217173 , n217272 );
and ( n217449 , n217448 , n217310 );
and ( n217450 , n217173 , n217272 );
or ( n217451 , n217449 , n217450 );
xor ( n217452 , n217377 , n217181 );
and ( n217453 , n217452 , n217404 );
and ( n217454 , n217377 , n217181 );
or ( n217455 , n217453 , n217454 );
xor ( n217456 , n217413 , n217189 );
and ( n217457 , n217456 , n217185 );
and ( n217458 , n217413 , n217189 );
or ( n217459 , n217457 , n217458 );
not ( n217460 , n213750 );
not ( n217461 , n217225 );
or ( n217462 , n217460 , n217461 );
nand ( n217463 , n217462 , n217084 );
not ( n217464 , n217225 );
nand ( n217465 , n217464 , n213751 );
and ( n217466 , n217463 , n217465 );
not ( n217467 , n37613 );
not ( n217468 , n36729 );
or ( n217469 , n217467 , n217468 );
nand ( n217470 , n36728 , n37612 );
nand ( n217471 , n217469 , n217470 );
buf ( n217472 , n217471 );
not ( n217473 , n217472 );
nor ( n217474 , n217466 , n217473 );
not ( n217475 , n217244 );
not ( n217476 , n215183 );
or ( n217477 , n217475 , n217476 );
not ( n217478 , n216934 );
and ( n217479 , n215104 , n217478 );
not ( n217480 , n215104 );
and ( n217481 , n217480 , n216934 );
or ( n217482 , n217479 , n217481 );
nand ( n217483 , n217482 , n215191 );
nand ( n217484 , n217477 , n217483 );
xor ( n217485 , n217474 , n217484 );
buf ( n217486 , n215773 );
not ( n217487 , n217486 );
not ( n217488 , n217253 );
or ( n217489 , n217487 , n217488 );
not ( n217490 , n215075 );
not ( n217491 , n216277 );
or ( n217492 , n217490 , n217491 );
not ( n217493 , n215075 );
nand ( n217494 , n217493 , n216281 );
nand ( n217495 , n217492 , n217494 );
not ( n217496 , n217495 );
or ( n217497 , n217496 , n215586 );
nand ( n217498 , n217489 , n217497 );
xor ( n217499 , n217485 , n217498 );
xor ( n217500 , n217474 , n217484 );
and ( n217501 , n217500 , n217498 );
and ( n217502 , n217474 , n217484 );
or ( n217503 , n217501 , n217502 );
not ( n217504 , n217296 );
buf ( n217505 , n217289 );
not ( n217506 , n217505 );
or ( n217507 , n217504 , n217506 );
not ( n217508 , n217044 );
not ( n217509 , n216593 );
or ( n217510 , n217508 , n217509 );
not ( n217511 , n216569 );
nand ( n217512 , n217511 , n215131 );
nand ( n217513 , n217510 , n217512 );
nand ( n217514 , n216598 , n217513 );
nand ( n217515 , n217507 , n217514 );
not ( n217516 , n217208 );
not ( n217517 , n214449 );
or ( n217518 , n217516 , n217517 );
not ( n217519 , n214759 );
not ( n217520 , n214467 );
or ( n217521 , n217519 , n217520 );
nand ( n217522 , n41834 , n214417 );
nand ( n217523 , n217521 , n217522 );
nand ( n217524 , n217523 , n214457 );
nand ( n217525 , n217518 , n217524 );
not ( n217526 , n217525 );
not ( n217527 , n217526 );
not ( n217528 , n217527 );
and ( n217529 , n214799 , n217218 );
not ( n217530 , n215117 );
not ( n217531 , n214803 );
or ( n217532 , n217530 , n217531 );
nand ( n217533 , n213917 , n214786 );
nand ( n217534 , n217532 , n217533 );
and ( n217535 , n217534 , n214588 );
nor ( n217536 , n217529 , n217535 );
not ( n217537 , n217536 );
or ( n217538 , n217528 , n217537 );
or ( n217539 , n217527 , n217536 );
nand ( n217540 , n217538 , n217539 );
xor ( n217541 , n217515 , n217540 );
not ( n217542 , n216989 );
not ( n217543 , n217542 );
not ( n217544 , n214488 );
or ( n217545 , n217543 , n217544 );
nand ( n217546 , n215228 , n216989 );
nand ( n217547 , n217545 , n217546 );
not ( n217548 , n217547 );
not ( n217549 , n214164 );
or ( n217550 , n217548 , n217549 );
not ( n217551 , n215963 );
not ( n217552 , n217551 );
nand ( n217553 , n217282 , n217552 );
nand ( n217554 , n217550 , n217553 );
xor ( n217555 , n217541 , n217554 );
xor ( n217556 , n217515 , n217540 );
and ( n217557 , n217556 , n217554 );
and ( n217558 , n217515 , n217540 );
or ( n217559 , n217557 , n217558 );
not ( n217560 , n217142 );
not ( n217561 , n216262 );
not ( n217562 , n217119 );
or ( n217563 , n217561 , n217562 );
not ( n217564 , n217116 );
nand ( n217565 , n217564 , n214824 );
nand ( n217566 , n217563 , n217565 );
not ( n217567 , n217566 );
or ( n217568 , n217560 , n217567 );
nand ( n217569 , n217320 , n213874 );
nand ( n217570 , n217568 , n217569 );
buf ( n217571 , n213206 );
not ( n217572 , n217571 );
not ( n217573 , n217397 );
not ( n217574 , n217573 );
not ( n217575 , n215989 );
or ( n217576 , n217574 , n217575 );
not ( n217577 , n213960 );
nand ( n217578 , n217577 , n217133 );
nand ( n217579 , n217576 , n217578 );
not ( n217580 , n217579 );
or ( n217581 , n217572 , n217580 );
nand ( n217582 , n217399 , n215605 );
nand ( n217583 , n217581 , n217582 );
xor ( n217584 , n217570 , n217583 );
xor ( n217585 , n217584 , n217431 );
xor ( n217586 , n217585 , n217455 );
not ( n217587 , n215966 );
not ( n217588 , n217017 );
not ( n217589 , n214834 );
or ( n217590 , n217588 , n217589 );
nand ( n217591 , n30962 , n215971 );
nand ( n217592 , n217590 , n217591 );
not ( n217593 , n217592 );
or ( n217594 , n217587 , n217593 );
nand ( n217595 , n217373 , n217023 );
nand ( n217596 , n217594 , n217595 );
not ( n217597 , n217387 );
not ( n217598 , n217380 );
or ( n217599 , n217597 , n217598 );
not ( n217600 , n217098 );
not ( n217601 , n213583 );
not ( n217602 , n216928 );
not ( n217603 , n217602 );
or ( n217604 , n217601 , n217603 );
not ( n217605 , n217084 );
nand ( n217606 , n217605 , n214134 );
nand ( n217607 , n217604 , n217606 );
nand ( n217608 , n217600 , n217607 );
nand ( n217609 , n217599 , n217608 );
xor ( n217610 , n217596 , n217609 );
not ( n217611 , n217472 );
and ( n217612 , n213751 , n217611 );
not ( n217613 , n213751 );
buf ( n217614 , n217472 );
not ( n217615 , n217614 );
not ( n217616 , n217615 );
and ( n217617 , n217613 , n217616 );
nor ( n217618 , n217612 , n217617 );
not ( n217619 , n217618 );
not ( n217620 , n217464 );
not ( n217621 , n216927 );
and ( n217622 , n217620 , n217621 );
and ( n217623 , n217464 , n216927 );
nor ( n217624 , n217622 , n217623 );
and ( n217625 , n217472 , n217225 );
not ( n217626 , n217472 );
and ( n217627 , n217626 , n217464 );
nor ( n217628 , n217625 , n217627 );
nand ( n217629 , n217624 , n217628 );
buf ( n217630 , n217629 );
not ( n217631 , n217630 );
not ( n217632 , n217631 );
or ( n217633 , n217619 , n217632 );
not ( n217634 , n217473 );
and ( n217635 , n216076 , n217634 );
not ( n217636 , n216076 );
not ( n217637 , n217614 );
and ( n217638 , n217636 , n217637 );
or ( n217639 , n217635 , n217638 );
buf ( n217640 , n217229 );
not ( n217641 , n217640 );
nand ( n217642 , n217639 , n217641 );
nand ( n217643 , n217633 , n217642 );
xor ( n217644 , n217610 , n217643 );
not ( n217645 , n216239 );
not ( n217646 , n215113 );
not ( n217647 , n41563 );
or ( n217648 , n217646 , n217647 );
nand ( n217649 , n216089 , n215118 );
nand ( n217650 , n217648 , n217649 );
not ( n217651 , n217650 );
or ( n217652 , n217645 , n217651 );
nand ( n217653 , n217307 , n214717 );
nand ( n217654 , n217652 , n217653 );
not ( n217655 , n216562 );
not ( n217656 , n217350 );
or ( n217657 , n217655 , n217656 );
not ( n217658 , n215290 );
not ( n217659 , n215628 );
or ( n217660 , n217658 , n217659 );
nand ( n217661 , n41608 , n215289 );
nand ( n217662 , n217660 , n217661 );
nand ( n217663 , n217662 , n214694 );
nand ( n217664 , n217657 , n217663 );
xor ( n217665 , n217654 , n217664 );
not ( n217666 , n217362 );
not ( n217667 , n216619 );
or ( n217668 , n217666 , n217667 );
not ( n217669 , n216964 );
not ( n217670 , n216014 );
or ( n217671 , n217669 , n217670 );
nand ( n217672 , n216068 , n214678 );
nand ( n217673 , n217671 , n217672 );
nand ( n217674 , n217673 , n216630 );
nand ( n217675 , n217668 , n217674 );
xor ( n217676 , n217665 , n217675 );
xor ( n217677 , n217644 , n217676 );
xor ( n217678 , n217677 , n217555 );
xor ( n217679 , n217586 , n217678 );
xor ( n217680 , n217585 , n217455 );
and ( n217681 , n217680 , n217678 );
and ( n217682 , n217585 , n217455 );
or ( n217683 , n217681 , n217682 );
xor ( n217684 , n217439 , n217443 );
xor ( n217685 , n217236 , n217262 );
xor ( n217686 , n217685 , n217499 );
xor ( n217687 , n217684 , n217686 );
xor ( n217688 , n217459 , n217687 );
xor ( n217689 , n217688 , n217344 );
xor ( n217690 , n217459 , n217687 );
and ( n217691 , n217690 , n217344 );
and ( n217692 , n217459 , n217687 );
or ( n217693 , n217691 , n217692 );
xor ( n217694 , n217451 , n217447 );
not ( n217695 , n216336 );
not ( n217696 , n213735 );
not ( n217697 , n41250 );
not ( n217698 , n217697 );
or ( n217699 , n217696 , n217698 );
not ( n217700 , n217147 );
nand ( n217701 , n217700 , n213732 );
nand ( n217702 , n217699 , n217701 );
not ( n217703 , n217702 );
or ( n217704 , n217695 , n217703 );
nand ( n217705 , n217268 , n213577 );
nand ( n217706 , n217704 , n217705 );
xor ( n217707 , n217435 , n217706 );
not ( n217708 , n213912 );
not ( n217709 , n213382 );
not ( n217710 , n41165 );
not ( n217711 , n217710 );
or ( n217712 , n217709 , n217711 );
not ( n217713 , n41164 );
not ( n217714 , n217713 );
not ( n217715 , n213382 );
nand ( n217716 , n217714 , n217715 );
nand ( n217717 , n217712 , n217716 );
not ( n217718 , n217717 );
or ( n217719 , n217708 , n217718 );
nand ( n217720 , n217335 , n213784 );
nand ( n217721 , n217719 , n217720 );
xor ( n217722 , n217707 , n217721 );
xor ( n217723 , n217694 , n217722 );
xor ( n217724 , n217723 , n217679 );
xor ( n217725 , n217724 , n217689 );
xor ( n217726 , n217723 , n217679 );
and ( n217727 , n217726 , n217689 );
and ( n217728 , n217723 , n217679 );
or ( n217729 , n217727 , n217728 );
xor ( n217730 , n217411 , n217421 );
xor ( n217731 , n217730 , n217725 );
xor ( n217732 , n217411 , n217421 );
and ( n217733 , n217732 , n217725 );
and ( n217734 , n217411 , n217421 );
or ( n217735 , n217733 , n217734 );
xor ( n217736 , n217654 , n217664 );
and ( n217737 , n217736 , n217675 );
and ( n217738 , n217654 , n217664 );
or ( n217739 , n217737 , n217738 );
xor ( n217740 , n217596 , n217609 );
and ( n217741 , n217740 , n217643 );
and ( n217742 , n217596 , n217609 );
or ( n217743 , n217741 , n217742 );
xor ( n217744 , n217236 , n217262 );
and ( n217745 , n217744 , n217499 );
and ( n217746 , n217236 , n217262 );
or ( n217747 , n217745 , n217746 );
xor ( n217748 , n217570 , n217583 );
and ( n217749 , n217748 , n217431 );
and ( n217750 , n217570 , n217583 );
or ( n217751 , n217749 , n217750 );
xor ( n217752 , n217435 , n217706 );
and ( n217753 , n217752 , n217721 );
and ( n217754 , n217435 , n217706 );
or ( n217755 , n217753 , n217754 );
xor ( n217756 , n217644 , n217676 );
and ( n217757 , n217756 , n217555 );
and ( n217758 , n217644 , n217676 );
or ( n217759 , n217757 , n217758 );
xor ( n217760 , n217439 , n217443 );
and ( n217761 , n217760 , n217686 );
and ( n217762 , n217439 , n217443 );
or ( n217763 , n217761 , n217762 );
xor ( n217764 , n217451 , n217447 );
and ( n217765 , n217764 , n217722 );
and ( n217766 , n217451 , n217447 );
or ( n217767 , n217765 , n217766 );
not ( n217768 , n217534 );
not ( n217769 , n214799 );
or ( n217770 , n217768 , n217769 );
not ( n217771 , n214598 );
not ( n217772 , n214783 );
or ( n217773 , n217771 , n217772 );
nand ( n217774 , n214786 , n214304 );
nand ( n217775 , n217773 , n217774 );
nand ( n217776 , n214588 , n217775 );
nand ( n217777 , n217770 , n217776 );
not ( n217778 , n217482 );
not ( n217779 , n215183 );
or ( n217780 , n217778 , n217779 );
not ( n217781 , n216142 );
not ( n217782 , n215545 );
or ( n217783 , n217781 , n217782 );
nand ( n217784 , n215104 , n215292 );
nand ( n217785 , n217783 , n217784 );
nand ( n217786 , n217785 , n215191 );
nand ( n217787 , n217780 , n217786 );
xor ( n217788 , n217777 , n217787 );
not ( n217789 , n217495 );
not ( n217790 , n216731 );
or ( n217791 , n217789 , n217790 );
not ( n217792 , n215268 );
not ( n217793 , n216280 );
or ( n217794 , n217792 , n217793 );
nand ( n217795 , n216968 , n216170 );
nand ( n217796 , n217794 , n217795 );
nand ( n217797 , n217796 , n215762 );
nand ( n217798 , n217791 , n217797 );
xor ( n217799 , n217788 , n217798 );
xor ( n217800 , n217777 , n217787 );
and ( n217801 , n217800 , n217798 );
and ( n217802 , n217777 , n217787 );
or ( n217803 , n217801 , n217802 );
not ( n217804 , n214458 );
not ( n217805 , n216166 );
not ( n217806 , n214989 );
or ( n217807 , n217805 , n217806 );
not ( n217808 , n216166 );
nand ( n217809 , n217808 , n30997 );
nand ( n217810 , n217807 , n217809 );
not ( n217811 , n217810 );
or ( n217812 , n217804 , n217811 );
nand ( n217813 , n214610 , n217523 );
nand ( n217814 , n217812 , n217813 );
not ( n217815 , n217513 );
not ( n217816 , n217289 );
or ( n217817 , n217815 , n217816 );
not ( n217818 , n214537 );
not ( n217819 , n216592 );
or ( n217820 , n217818 , n217819 );
nand ( n217821 , n216419 , n214899 );
nand ( n217822 , n217820 , n217821 );
not ( n217823 , n216199 );
buf ( n217824 , n217823 );
nand ( n217825 , n217822 , n217824 );
nand ( n217826 , n217817 , n217825 );
xor ( n217827 , n217814 , n217826 );
not ( n217828 , n214164 );
not ( n217829 , n215955 );
not ( n217830 , n215833 );
or ( n217831 , n217829 , n217830 );
nand ( n217832 , n41716 , n217280 );
nand ( n217833 , n217831 , n217832 );
not ( n217834 , n217833 );
or ( n217835 , n217828 , n217834 );
nand ( n217836 , n217547 , n215963 );
nand ( n217837 , n217835 , n217836 );
xor ( n217838 , n217827 , n217837 );
xor ( n217839 , n217814 , n217826 );
and ( n217840 , n217839 , n217837 );
and ( n217841 , n217814 , n217826 );
or ( n217842 , n217840 , n217841 );
xor ( n217843 , n217799 , n217838 );
xor ( n217844 , n217843 , n217739 );
xor ( n217845 , n217844 , n217755 );
xor ( n217846 , n217845 , n217759 );
xor ( n217847 , n217844 , n217755 );
and ( n217848 , n217847 , n217759 );
and ( n217849 , n217844 , n217755 );
or ( n217850 , n217848 , n217849 );
not ( n217851 , n213577 );
not ( n217852 , n217702 );
or ( n217853 , n217851 , n217852 );
and ( n217854 , n213735 , n208164 );
not ( n217855 , n213735 );
not ( n217856 , n208164 );
and ( n217857 , n217855 , n217856 );
nor ( n217858 , n217854 , n217857 );
nand ( n217859 , n217858 , n216336 );
nand ( n217860 , n217853 , n217859 );
xor ( n217861 , n217860 , n217743 );
not ( n217862 , n217673 );
nand ( n217863 , n216063 , n215788 );
not ( n217864 , n217863 );
not ( n217865 , n217864 );
or ( n217866 , n217862 , n217865 );
not ( n217867 , n216208 );
not ( n217868 , n216014 );
or ( n217869 , n217867 , n217868 );
nand ( n217870 , n216403 , n216207 );
nand ( n217871 , n217869 , n217870 );
nand ( n217872 , n216630 , n217871 );
nand ( n217873 , n217866 , n217872 );
not ( n217874 , n217607 );
not ( n217875 , n217087 );
not ( n217876 , n217875 );
not ( n217877 , n217876 );
not ( n217878 , n217877 );
or ( n217879 , n217874 , n217878 );
not ( n217880 , n214956 );
not ( n217881 , n217084 );
or ( n217882 , n217880 , n217881 );
nand ( n217883 , n216928 , n214960 );
nand ( n217884 , n217882 , n217883 );
not ( n217885 , n217098 );
nand ( n217886 , n217884 , n217885 );
nand ( n217887 , n217879 , n217886 );
xor ( n217888 , n217873 , n217887 );
not ( n217889 , n217639 );
not ( n217890 , n217630 );
not ( n217891 , n217890 );
or ( n217892 , n217889 , n217891 );
not ( n217893 , n213347 );
not ( n217894 , n217473 );
or ( n217895 , n217893 , n217894 );
nand ( n217896 , n217614 , n214616 );
nand ( n217897 , n217895 , n217896 );
nand ( n217898 , n217897 , n217641 );
nand ( n217899 , n217892 , n217898 );
xor ( n217900 , n217888 , n217899 );
xor ( n217901 , n217861 , n217900 );
nor ( n217902 , n217536 , n217526 );
not ( n217903 , n214694 );
not ( n217904 , n215290 );
not ( n217905 , n216782 );
or ( n217906 , n217904 , n217905 );
nand ( n217907 , n213815 , n41700 );
nand ( n217908 , n217906 , n217907 );
not ( n217909 , n217908 );
or ( n217910 , n217903 , n217909 );
nand ( n217911 , n217662 , n213718 );
nand ( n217912 , n217910 , n217911 );
xor ( n217913 , n217902 , n217912 );
not ( n217914 , n217023 );
not ( n217915 , n217592 );
or ( n217916 , n217914 , n217915 );
and ( n217917 , n208725 , n215971 );
not ( n217918 , n208725 );
and ( n217919 , n217918 , n217017 );
or ( n217920 , n217917 , n217919 );
nand ( n217921 , n217920 , n215966 );
nand ( n217922 , n217916 , n217921 );
xor ( n217923 , n217913 , n217922 );
not ( n217924 , n37630 );
not ( n217925 , n217924 );
not ( n217926 , n36320 );
not ( n217927 , n217926 );
or ( n217928 , n217925 , n217927 );
nand ( n217929 , n36320 , n37630 );
nand ( n217930 , n217928 , n217929 );
not ( n217931 , n217930 );
and ( n217932 , n217472 , n217931 );
not ( n217933 , n217472 );
and ( n217934 , n217933 , n217930 );
nor ( n217935 , n217932 , n217934 );
buf ( n217936 , n217935 );
nor ( n217937 , n217936 , n213751 );
xor ( n217938 , n217937 , n217503 );
not ( n217939 , n216239 );
not ( n217940 , n215113 );
not ( n217941 , n208717 );
not ( n217942 , n217941 );
or ( n217943 , n217940 , n217942 );
buf ( n217944 , n216037 );
nand ( n217945 , n208717 , n217944 );
nand ( n217946 , n217943 , n217945 );
not ( n217947 , n217946 );
or ( n217948 , n217939 , n217947 );
nand ( n217949 , n217650 , n214717 );
nand ( n217950 , n217948 , n217949 );
xor ( n217951 , n217938 , n217950 );
xor ( n217952 , n217923 , n217951 );
xor ( n217953 , n217952 , n217747 );
xor ( n217954 , n217901 , n217953 );
xor ( n217955 , n217954 , n217763 );
xor ( n217956 , n217901 , n217953 );
and ( n217957 , n217956 , n217763 );
and ( n217958 , n217901 , n217953 );
or ( n217959 , n217957 , n217958 );
not ( n217960 , n213912 );
not ( n217961 , n213381 );
not ( n217962 , n40724 );
or ( n217963 , n217961 , n217962 );
not ( n217964 , n40724 );
nand ( n217965 , n217964 , n213382 );
nand ( n217966 , n217963 , n217965 );
not ( n217967 , n217966 );
or ( n217968 , n217960 , n217967 );
buf ( n217969 , n213784 );
nand ( n217970 , n217717 , n217969 );
nand ( n217971 , n217968 , n217970 );
xor ( n217972 , n217971 , n217751 );
not ( n217973 , n213874 );
not ( n217974 , n217566 );
or ( n217975 , n217973 , n217974 );
not ( n217976 , n214818 );
not ( n217977 , n41069 );
not ( n217978 , n217977 );
or ( n217979 , n217976 , n217978 );
or ( n217980 , n217977 , n214818 );
nand ( n217981 , n217979 , n217980 );
nand ( n217982 , n217981 , n213058 );
nand ( n217983 , n217975 , n217982 );
not ( n217984 , n213206 );
not ( n217985 , n213960 );
not ( n217986 , n41318 );
or ( n217987 , n217985 , n217986 );
nand ( n217988 , n216311 , n217397 );
nand ( n217989 , n217987 , n217988 );
not ( n217990 , n217989 );
or ( n217991 , n217984 , n217990 );
nand ( n217992 , n217579 , n215605 );
nand ( n217993 , n217991 , n217992 );
xor ( n217994 , n217983 , n217993 );
xor ( n217995 , n217994 , n217559 );
xor ( n217996 , n217972 , n217995 );
xor ( n217997 , n217767 , n217996 );
xor ( n217998 , n217997 , n217846 );
xor ( n217999 , n217767 , n217996 );
and ( n218000 , n217999 , n217846 );
and ( n218001 , n217767 , n217996 );
or ( n218002 , n218000 , n218001 );
xor ( n218003 , n217683 , n217693 );
xor ( n218004 , n218003 , n217955 );
xor ( n218005 , n217683 , n217693 );
and ( n218006 , n218005 , n217955 );
and ( n218007 , n217683 , n217693 );
or ( n218008 , n218006 , n218007 );
xor ( n218009 , n217998 , n217729 );
xor ( n218010 , n218009 , n218004 );
xor ( n218011 , n217998 , n217729 );
and ( n218012 , n218011 , n218004 );
and ( n218013 , n217998 , n217729 );
or ( n218014 , n218012 , n218013 );
xor ( n218015 , n217902 , n217912 );
and ( n218016 , n218015 , n217922 );
and ( n218017 , n217902 , n217912 );
or ( n218018 , n218016 , n218017 );
xor ( n218019 , n217873 , n217887 );
and ( n218020 , n218019 , n217899 );
and ( n218021 , n217873 , n217887 );
or ( n218022 , n218020 , n218021 );
xor ( n218023 , n217937 , n217503 );
and ( n218024 , n218023 , n217950 );
and ( n218025 , n217937 , n217503 );
or ( n218026 , n218024 , n218025 );
xor ( n218027 , n217799 , n217838 );
and ( n218028 , n218027 , n217739 );
and ( n218029 , n217799 , n217838 );
or ( n218030 , n218028 , n218029 );
xor ( n218031 , n217983 , n217993 );
and ( n218032 , n218031 , n217559 );
and ( n218033 , n217983 , n217993 );
or ( n218034 , n218032 , n218033 );
xor ( n218035 , n217860 , n217743 );
and ( n218036 , n218035 , n217900 );
and ( n218037 , n217860 , n217743 );
or ( n218038 , n218036 , n218037 );
xor ( n218039 , n217923 , n217951 );
and ( n218040 , n218039 , n217747 );
and ( n218041 , n217923 , n217951 );
or ( n218042 , n218040 , n218041 );
xor ( n218043 , n217971 , n217751 );
and ( n218044 , n218043 , n217995 );
and ( n218045 , n217971 , n217751 );
or ( n218046 , n218044 , n218045 );
not ( n218047 , n217796 );
nand ( n218048 , n215326 , n215576 );
not ( n218049 , n218048 );
not ( n218050 , n218049 );
or ( n218051 , n218047 , n218050 );
not ( n218052 , n215953 );
not ( n218053 , n216280 );
or ( n218054 , n218052 , n218053 );
nand ( n218055 , n215511 , n215481 );
nand ( n218056 , n218054 , n218055 );
nand ( n218057 , n218056 , n215587 );
nand ( n218058 , n218051 , n218057 );
not ( n218059 , n217822 );
not ( n218060 , n217288 );
or ( n218061 , n218059 , n218060 );
not ( n218062 , n216964 );
not ( n218063 , n216592 );
or ( n218064 , n218062 , n218063 );
not ( n218065 , n215050 );
nand ( n218066 , n218065 , n216591 );
nand ( n218067 , n218064 , n218066 );
nand ( n218068 , n218067 , n217823 );
nand ( n218069 , n218061 , n218068 );
xor ( n218070 , n218058 , n218069 );
not ( n218071 , n216166 );
not ( n218072 , n214820 );
or ( n218073 , n218071 , n218072 );
nand ( n218074 , n41725 , n217808 );
nand ( n218075 , n218073 , n218074 );
not ( n218076 , n218075 );
buf ( n218077 , n214285 );
not ( n218078 , n218077 );
or ( n218079 , n218076 , n218078 );
nand ( n218080 , n217810 , n214610 );
nand ( n218081 , n218079 , n218080 );
xor ( n218082 , n218070 , n218081 );
xor ( n218083 , n218058 , n218069 );
and ( n218084 , n218083 , n218081 );
and ( n218085 , n218058 , n218069 );
or ( n218086 , n218084 , n218085 );
not ( n218087 , n217785 );
not ( n218088 , n215182 );
or ( n218089 , n218087 , n218088 );
not ( n218090 , n213918 );
not ( n218091 , n215545 );
or ( n218092 , n218090 , n218091 );
nand ( n218093 , n215104 , n209248 );
nand ( n218094 , n218092 , n218093 );
nand ( n218095 , n218094 , n215191 );
nand ( n218096 , n218089 , n218095 );
not ( n218097 , n217775 );
not ( n218098 , n214799 );
or ( n218099 , n218097 , n218098 );
not ( n218100 , n214786 );
not ( n218101 , n214467 );
or ( n218102 , n218100 , n218101 );
nand ( n218103 , n41834 , n214783 );
nand ( n218104 , n218102 , n218103 );
nand ( n218105 , n218104 , n214588 );
nand ( n218106 , n218099 , n218105 );
xor ( n218107 , n218096 , n218106 );
not ( n218108 , n214694 );
not ( n218109 , n215289 );
not ( n218110 , n41564 );
or ( n218111 , n218109 , n218110 );
nand ( n218112 , n41563 , n216810 );
nand ( n218113 , n218111 , n218112 );
not ( n218114 , n218113 );
or ( n218115 , n218108 , n218114 );
nand ( n218116 , n213718 , n217908 );
nand ( n218117 , n218115 , n218116 );
xor ( n218118 , n218107 , n218117 );
not ( n218119 , n217833 );
or ( n218120 , n218119 , n217551 );
and ( n218121 , n214834 , n217542 );
not ( n218122 , n214834 );
and ( n218123 , n218122 , n215956 );
or ( n218124 , n218121 , n218123 );
not ( n218125 , n218124 );
or ( n218126 , n218125 , n217549 );
nand ( n218127 , n218120 , n218126 );
xor ( n218128 , n218118 , n218127 );
xor ( n218129 , n218107 , n218117 );
and ( n218130 , n218129 , n218127 );
and ( n218131 , n218107 , n218117 );
or ( n218132 , n218130 , n218131 );
not ( n218133 , n213498 );
not ( n218134 , n213735 );
not ( n218135 , n217115 );
or ( n218136 , n218134 , n218135 );
not ( n218137 , n217119 );
nand ( n218138 , n218137 , n213732 );
nand ( n218139 , n218136 , n218138 );
not ( n218140 , n218139 );
or ( n218141 , n218133 , n218140 );
nand ( n218142 , n217858 , n213577 );
nand ( n218143 , n218141 , n218142 );
xor ( n218144 , n218018 , n218143 );
xor ( n218145 , n218144 , n218082 );
not ( n218146 , n217981 );
not ( n218147 , n213874 );
or ( n218148 , n218146 , n218147 );
xor ( n218149 , n217710 , n214818 );
not ( n218150 , n217142 );
or ( n218151 , n218149 , n218150 );
nand ( n218152 , n218148 , n218151 );
xor ( n218153 , n218022 , n218152 );
not ( n218154 , n217023 );
not ( n218155 , n217920 );
or ( n218156 , n218154 , n218155 );
not ( n218157 , n215272 );
not ( n218158 , n215628 );
or ( n218159 , n218157 , n218158 );
not ( n218160 , n215272 );
nand ( n218161 , n218160 , n41608 );
nand ( n218162 , n218159 , n218161 );
nand ( n218163 , n218162 , n215966 );
nand ( n218164 , n218156 , n218163 );
not ( n218165 , n217871 );
not ( n218166 , n217864 );
or ( n218167 , n218165 , n218166 );
not ( n218168 , n215075 );
not ( n218169 , n216014 );
or ( n218170 , n218168 , n218169 );
nand ( n218171 , n216068 , n215899 );
nand ( n218172 , n218170 , n218171 );
nand ( n218173 , n218172 , n216630 );
nand ( n218174 , n218167 , n218173 );
xor ( n218175 , n218164 , n218174 );
not ( n218176 , n217884 );
not ( n218177 , n217877 );
or ( n218178 , n218176 , n218177 );
not ( n218179 , n217044 );
not ( n218180 , n217079 );
or ( n218181 , n218179 , n218180 );
nand ( n218182 , n217080 , n215131 );
nand ( n218183 , n218181 , n218182 );
nand ( n218184 , n218183 , n217885 );
nand ( n218185 , n218178 , n218184 );
xor ( n218186 , n218175 , n218185 );
xor ( n218187 , n218153 , n218186 );
xor ( n218188 , n218145 , n218187 );
xor ( n218189 , n218188 , n218042 );
xor ( n218190 , n218145 , n218187 );
and ( n218191 , n218190 , n218042 );
and ( n218192 , n218145 , n218187 );
or ( n218193 , n218191 , n218192 );
buf ( n218194 , n33682 );
buf ( n218195 , n218194 );
nand ( n218196 , n218195 , n36398 );
not ( n218197 , n218196 );
not ( n218198 , n218197 );
not ( n218199 , n36589 );
not ( n218200 , n218199 );
or ( n218201 , n218198 , n218200 );
nand ( n218202 , n36589 , n218196 );
nand ( n218203 , n218201 , n218202 );
not ( n218204 , n218203 );
not ( n218205 , n218204 );
and ( n218206 , n215999 , n218205 );
not ( n218207 , n215999 );
not ( n218208 , n218204 );
not ( n218209 , n218208 );
and ( n218210 , n218207 , n218209 );
nor ( n218211 , n218206 , n218210 );
not ( n218212 , n218211 );
nand ( n218213 , n217931 , n218204 );
not ( n218214 , n218197 );
not ( n218215 , n218199 );
or ( n218216 , n218214 , n218215 );
nand ( n218217 , n218216 , n218202 );
nand ( n218218 , n218217 , n217930 );
nand ( n218219 , n218213 , n218218 , n217935 );
buf ( n218220 , n218219 );
not ( n218221 , n218220 );
not ( n218222 , n218221 );
or ( n218223 , n218212 , n218222 );
not ( n218224 , n216076 );
not ( n218225 , n218224 );
not ( n218226 , n218203 );
not ( n218227 , n218226 );
or ( n218228 , n218225 , n218227 );
nand ( n218229 , n218208 , n216076 );
nand ( n218230 , n218228 , n218229 );
not ( n218231 , n217936 );
buf ( n218232 , n218231 );
nand ( n218233 , n218230 , n218232 );
nand ( n218234 , n218223 , n218233 );
xor ( n218235 , n218128 , n218234 );
xor ( n218236 , n218235 , n218026 );
xor ( n218237 , n218236 , n217850 );
not ( n218238 , n217897 );
not ( n218239 , n217629 );
not ( n218240 , n218239 );
or ( n218241 , n218238 , n218240 );
not ( n218242 , n213583 );
not ( n218243 , n217611 );
or ( n218244 , n218242 , n218243 );
nand ( n218245 , n217614 , n214134 );
nand ( n218246 , n218244 , n218245 );
nand ( n218247 , n218246 , n217230 );
nand ( n218248 , n218241 , n218247 );
not ( n218249 , n217930 );
not ( n218250 , n213750 );
and ( n218251 , n218249 , n218250 );
nand ( n218252 , n217930 , n213750 );
not ( n218253 , n217614 );
and ( n218254 , n218252 , n218253 );
nor ( n218255 , n218251 , n218254 );
buf ( n218256 , n218204 );
nor ( n218257 , n218255 , n218256 );
xor ( n218258 , n218248 , n218257 );
xor ( n218259 , n218258 , n217803 );
xor ( n218260 , n218259 , n218034 );
xor ( n218261 , n218260 , n218030 );
xor ( n218262 , n218237 , n218261 );
xor ( n218263 , n218236 , n217850 );
and ( n218264 , n218263 , n218261 );
and ( n218265 , n218236 , n217850 );
or ( n218266 , n218264 , n218265 );
not ( n218267 , n214319 );
not ( n218268 , n40710 );
and ( n218269 , n213382 , n218268 );
not ( n218270 , n213382 );
and ( n218271 , n218270 , n40710 );
or ( n218272 , n218269 , n218271 );
not ( n218273 , n218272 );
or ( n218274 , n218267 , n218273 );
nand ( n218275 , n217966 , n217969 );
nand ( n218276 , n218274 , n218275 );
not ( n218277 , n215605 );
not ( n218278 , n217989 );
or ( n218279 , n218277 , n218278 );
not ( n218280 , n213960 );
not ( n218281 , n41249 );
or ( n218282 , n218280 , n218281 );
not ( n218283 , n41249 );
nand ( n218284 , n218283 , n217397 );
nand ( n218285 , n218282 , n218284 );
nand ( n218286 , n218285 , n213206 );
nand ( n218287 , n218279 , n218286 );
not ( n218288 , n216239 );
not ( n218289 , n215113 );
not ( n218290 , n41396 );
not ( n218291 , n218290 );
or ( n218292 , n218289 , n218291 );
nand ( n218293 , n41396 , n217944 );
nand ( n218294 , n218292 , n218293 );
not ( n218295 , n218294 );
or ( n218296 , n218288 , n218295 );
nand ( n218297 , n217946 , n214717 );
nand ( n218298 , n218296 , n218297 );
xor ( n218299 , n218287 , n218298 );
xor ( n218300 , n218299 , n217842 );
xor ( n218301 , n218276 , n218300 );
xor ( n218302 , n218301 , n218038 );
xor ( n218303 , n218046 , n218302 );
xor ( n218304 , n218303 , n218189 );
xor ( n218305 , n218046 , n218302 );
and ( n218306 , n218305 , n218189 );
and ( n218307 , n218046 , n218302 );
or ( n218308 , n218306 , n218307 );
xor ( n218309 , n217959 , n218002 );
xor ( n218310 , n218309 , n218262 );
xor ( n218311 , n217959 , n218002 );
and ( n218312 , n218311 , n218262 );
and ( n218313 , n217959 , n218002 );
or ( n218314 , n218312 , n218313 );
xor ( n218315 , n218304 , n218008 );
xor ( n218316 , n218315 , n218310 );
xor ( n218317 , n218304 , n218008 );
and ( n218318 , n218317 , n218310 );
and ( n218319 , n218304 , n218008 );
or ( n218320 , n218318 , n218319 );
xor ( n218321 , n218164 , n218174 );
and ( n218322 , n218321 , n218185 );
and ( n218323 , n218164 , n218174 );
or ( n218324 , n218322 , n218323 );
xor ( n218325 , n218248 , n218257 );
and ( n218326 , n218325 , n217803 );
and ( n218327 , n218248 , n218257 );
or ( n218328 , n218326 , n218327 );
xor ( n218329 , n218287 , n218298 );
and ( n218330 , n218329 , n217842 );
and ( n218331 , n218287 , n218298 );
or ( n218332 , n218330 , n218331 );
xor ( n218333 , n218018 , n218143 );
and ( n218334 , n218333 , n218082 );
and ( n218335 , n218018 , n218143 );
or ( n218336 , n218334 , n218335 );
xor ( n218337 , n218022 , n218152 );
and ( n218338 , n218337 , n218186 );
and ( n218339 , n218022 , n218152 );
or ( n218340 , n218338 , n218339 );
xor ( n218341 , n218128 , n218234 );
and ( n218342 , n218341 , n218026 );
and ( n218343 , n218128 , n218234 );
or ( n218344 , n218342 , n218343 );
xor ( n218345 , n218259 , n218034 );
and ( n218346 , n218345 , n218030 );
and ( n218347 , n218259 , n218034 );
or ( n218348 , n218346 , n218347 );
xor ( n218349 , n218276 , n218300 );
and ( n218350 , n218349 , n218038 );
and ( n218351 , n218276 , n218300 );
or ( n218352 , n218350 , n218351 );
not ( n218353 , n218094 );
not ( n218354 , n215182 );
or ( n218355 , n218353 , n218354 );
not ( n218356 , n214927 );
not ( n218357 , n215105 );
or ( n218358 , n218356 , n218357 );
nand ( n218359 , n215104 , n214304 );
nand ( n218360 , n218358 , n218359 );
nand ( n218361 , n218360 , n215191 );
nand ( n218362 , n218355 , n218361 );
not ( n218363 , n218056 );
or ( n218364 , n218048 , n218363 );
not ( n218365 , n216142 );
not ( n218366 , n215765 );
or ( n218367 , n218365 , n218366 );
nand ( n218368 , n215511 , n215292 );
nand ( n218369 , n218367 , n218368 );
not ( n218370 , n218369 );
or ( n218371 , n218370 , n215586 );
nand ( n218372 , n218364 , n218371 );
xor ( n218373 , n218362 , n218372 );
not ( n218374 , n214808 );
not ( n218375 , n214786 );
not ( n218376 , n214628 );
or ( n218377 , n218375 , n218376 );
not ( n218378 , n214786 );
nand ( n218379 , n218378 , n30997 );
nand ( n218380 , n218377 , n218379 );
not ( n218381 , n218380 );
or ( n218382 , n218374 , n218381 );
nand ( n218383 , n214799 , n218104 );
nand ( n218384 , n218382 , n218383 );
xor ( n218385 , n218373 , n218384 );
xor ( n218386 , n218362 , n218372 );
and ( n218387 , n218386 , n218384 );
and ( n218388 , n218362 , n218372 );
or ( n218389 , n218387 , n218388 );
not ( n218390 , n218067 );
not ( n218391 , n217288 );
or ( n218392 , n218390 , n218391 );
not ( n218393 , n216208 );
not ( n218394 , n216569 );
or ( n218395 , n218393 , n218394 );
nand ( n218396 , n216207 , n216419 );
nand ( n218397 , n218395 , n218396 );
nand ( n218398 , n218397 , n217823 );
nand ( n218399 , n218392 , n218398 );
not ( n218400 , n214458 );
and ( n218401 , n41716 , n216167 );
not ( n218402 , n41716 );
and ( n218403 , n218402 , n216166 );
or ( n218404 , n218401 , n218403 );
not ( n218405 , n218404 );
or ( n218406 , n218400 , n218405 );
nand ( n218407 , n218075 , n214610 );
nand ( n218408 , n218406 , n218407 );
xor ( n218409 , n218399 , n218408 );
and ( n218410 , n218096 , n218106 );
xor ( n218411 , n218409 , n218410 );
xor ( n218412 , n218399 , n218408 );
and ( n218413 , n218412 , n218410 );
and ( n218414 , n218399 , n218408 );
or ( n218415 , n218413 , n218414 );
not ( n218416 , n213577 );
not ( n218417 , n218139 );
or ( n218418 , n218416 , n218417 );
not ( n218419 , n213735 );
not ( n218420 , n41069 );
not ( n218421 , n218420 );
or ( n218422 , n218419 , n218421 );
nand ( n218423 , n41069 , n213732 );
nand ( n218424 , n218422 , n218423 );
nand ( n218425 , n218424 , n213498 );
nand ( n218426 , n218418 , n218425 );
xor ( n218427 , n218324 , n218426 );
xor ( n218428 , n218427 , n218328 );
not ( n218429 , n214694 );
not ( n218430 , n215290 );
not ( n218431 , n217941 );
or ( n218432 , n218430 , n218431 );
not ( n218433 , n215793 );
nand ( n218434 , n218433 , n215289 );
nand ( n218435 , n218432 , n218434 );
not ( n218436 , n218435 );
or ( n218437 , n218429 , n218436 );
nand ( n218438 , n218113 , n216562 );
nand ( n218439 , n218437 , n218438 );
not ( n218440 , n37601 );
not ( n218441 , n36374 );
or ( n218442 , n218440 , n218441 );
nand ( n218443 , n218442 , n37586 );
nand ( n218444 , n36395 , n36402 );
not ( n218445 , n218444 );
and ( n218446 , n218443 , n218445 );
not ( n218447 , n218443 );
and ( n218448 , n218447 , n218444 );
nor ( n218449 , n218446 , n218448 );
and ( n218450 , n218217 , n218449 );
not ( n218451 , n218217 );
not ( n218452 , n218449 );
and ( n218453 , n218451 , n218452 );
nor ( n218454 , n218450 , n218453 );
buf ( n218455 , n218454 );
not ( n218456 , n218455 );
nor ( n218457 , n218456 , n213751 );
xor ( n218458 , n218439 , n218457 );
not ( n218459 , n217571 );
not ( n218460 , n213960 );
not ( n218461 , n216855 );
or ( n218462 , n218460 , n218461 );
nand ( n218463 , n216859 , n217397 );
nand ( n218464 , n218462 , n218463 );
not ( n218465 , n218464 );
or ( n218466 , n218459 , n218465 );
not ( n218467 , n214085 );
nand ( n218468 , n218285 , n218467 );
nand ( n218469 , n218466 , n218468 );
xor ( n218470 , n218458 , n218469 );
xor ( n218471 , n218428 , n218470 );
not ( n218472 , n218294 );
not ( n218473 , n214717 );
or ( n218474 , n218472 , n218473 );
not ( n218475 , n215113 );
not ( n218476 , n208594 );
or ( n218477 , n218475 , n218476 );
nand ( n218478 , n216310 , n216037 );
nand ( n218479 , n218477 , n218478 );
nand ( n218480 , n218479 , n216239 );
nand ( n218481 , n218474 , n218480 );
xor ( n218482 , n218481 , n218086 );
xor ( n218483 , n218482 , n218132 );
xor ( n218484 , n218471 , n218483 );
xor ( n218485 , n218428 , n218470 );
and ( n218486 , n218485 , n218483 );
and ( n218487 , n218428 , n218470 );
or ( n218488 , n218486 , n218487 );
not ( n218489 , n215966 );
not ( n218490 , n214130 );
not ( n218491 , n215820 );
or ( n218492 , n218490 , n218491 );
nand ( n218493 , n41700 , n215971 );
nand ( n218494 , n218492 , n218493 );
not ( n218495 , n218494 );
or ( n218496 , n218489 , n218495 );
nand ( n218497 , n218162 , n213894 );
nand ( n218498 , n218496 , n218497 );
not ( n218499 , n215963 );
not ( n218500 , n218124 );
or ( n218501 , n218499 , n218500 );
not ( n218502 , n216985 );
not ( n218503 , n208725 );
not ( n218504 , n218503 );
or ( n218505 , n218502 , n218504 );
nand ( n218506 , n215956 , n208725 );
nand ( n218507 , n218505 , n218506 );
nand ( n218508 , n218507 , n214164 );
nand ( n218509 , n218501 , n218508 );
xor ( n218510 , n218498 , n218509 );
not ( n218511 , n218172 );
not ( n218512 , n216065 );
or ( n218513 , n218511 , n218512 );
not ( n218514 , n216170 );
not ( n218515 , n218514 );
not ( n218516 , n216014 );
or ( n218517 , n218515 , n218516 );
nand ( n218518 , n216327 , n216170 );
nand ( n218519 , n218517 , n218518 );
nand ( n218520 , n217047 , n218519 );
nand ( n218521 , n218513 , n218520 );
xor ( n218522 , n218510 , n218521 );
xor ( n218523 , n218522 , n218411 );
not ( n218524 , n218230 );
not ( n218525 , n218220 );
not ( n218526 , n218525 );
or ( n218527 , n218524 , n218526 );
not ( n218528 , n213347 );
not ( n218529 , n218226 );
or ( n218530 , n218528 , n218529 );
nand ( n218531 , n218208 , n214616 );
nand ( n218532 , n218530 , n218531 );
not ( n218533 , n217936 );
nand ( n218534 , n218532 , n218533 );
nand ( n218535 , n218527 , n218534 );
xor ( n218536 , n218523 , n218535 );
xor ( n218537 , n218536 , n218344 );
xor ( n218538 , n218537 , n218348 );
xor ( n218539 , n218536 , n218344 );
and ( n218540 , n218539 , n218348 );
and ( n218541 , n218536 , n218344 );
or ( n218542 , n218540 , n218541 );
not ( n218543 , n218183 );
not ( n218544 , n217088 );
not ( n218545 , n218544 );
or ( n218546 , n218543 , n218545 );
not ( n218547 , n214537 );
not ( n218548 , n217602 );
or ( n218549 , n218547 , n218548 );
nand ( n218550 , n217080 , n214899 );
nand ( n218551 , n218549 , n218550 );
nand ( n218552 , n218551 , n217885 );
nand ( n218553 , n218546 , n218552 );
not ( n218554 , n218246 );
not ( n218555 , n217890 );
or ( n218556 , n218554 , n218555 );
not ( n218557 , n214956 );
not ( n218558 , n217611 );
or ( n218559 , n218557 , n218558 );
not ( n218560 , n217611 );
nand ( n218561 , n218560 , n214960 );
nand ( n218562 , n218559 , n218561 );
nand ( n218563 , n218562 , n217230 );
nand ( n218564 , n218556 , n218563 );
xor ( n218565 , n218553 , n218564 );
xor ( n218566 , n218565 , n218385 );
xor ( n218567 , n218566 , n218336 );
xor ( n218568 , n218567 , n218332 );
xor ( n218569 , n218568 , n218352 );
xor ( n218570 , n218569 , n218484 );
xor ( n218571 , n218568 , n218352 );
and ( n218572 , n218571 , n218484 );
and ( n218573 , n218568 , n218352 );
or ( n218574 , n218572 , n218573 );
not ( n218575 , n217142 );
not ( n218576 , n214824 );
not ( n218577 , n40724 );
or ( n218578 , n218576 , n218577 );
nand ( n218579 , n217964 , n216262 );
nand ( n218580 , n218578 , n218579 );
not ( n218581 , n218580 );
or ( n218582 , n218575 , n218581 );
not ( n218583 , n218149 );
nand ( n218584 , n218583 , n213874 );
nand ( n218585 , n218582 , n218584 );
xor ( n218586 , n218585 , n218340 );
not ( n218587 , n218272 );
not ( n218588 , n217969 );
or ( n218589 , n218587 , n218588 );
not ( n218590 , n208042 );
xor ( n218591 , n218590 , n213382 );
not ( n218592 , n218591 );
or ( n218593 , n218592 , n213171 );
nand ( n218594 , n218589 , n218593 );
xor ( n218595 , n218586 , n218594 );
xor ( n218596 , n218193 , n218595 );
xor ( n218597 , n218596 , n218538 );
xor ( n218598 , n218193 , n218595 );
and ( n218599 , n218598 , n218538 );
and ( n218600 , n218193 , n218595 );
or ( n218601 , n218599 , n218600 );
xor ( n218602 , n218266 , n218570 );
xor ( n218603 , n218602 , n218308 );
xor ( n218604 , n218266 , n218570 );
and ( n218605 , n218604 , n218308 );
and ( n218606 , n218266 , n218570 );
or ( n218607 , n218605 , n218606 );
xor ( n218608 , n218597 , n218314 );
xor ( n218609 , n218608 , n218603 );
xor ( n218610 , n218597 , n218314 );
and ( n218611 , n218610 , n218603 );
and ( n218612 , n218597 , n218314 );
or ( n218613 , n218611 , n218612 );
xor ( n218614 , n218498 , n218509 );
and ( n218615 , n218614 , n218521 );
and ( n218616 , n218498 , n218509 );
or ( n218617 , n218615 , n218616 );
xor ( n218618 , n218553 , n218564 );
and ( n218619 , n218618 , n218385 );
and ( n218620 , n218553 , n218564 );
or ( n218621 , n218619 , n218620 );
xor ( n218622 , n218439 , n218457 );
and ( n218623 , n218622 , n218469 );
and ( n218624 , n218439 , n218457 );
or ( n218625 , n218623 , n218624 );
xor ( n218626 , n218481 , n218086 );
and ( n218627 , n218626 , n218132 );
and ( n218628 , n218481 , n218086 );
or ( n218629 , n218627 , n218628 );
xor ( n218630 , n218324 , n218426 );
and ( n218631 , n218630 , n218328 );
and ( n218632 , n218324 , n218426 );
or ( n218633 , n218631 , n218632 );
xor ( n218634 , n218522 , n218411 );
and ( n218635 , n218634 , n218535 );
and ( n218636 , n218522 , n218411 );
or ( n218637 , n218635 , n218636 );
xor ( n218638 , n218566 , n218336 );
and ( n218639 , n218638 , n218332 );
and ( n218640 , n218566 , n218336 );
or ( n218641 , n218639 , n218640 );
xor ( n218642 , n218585 , n218340 );
and ( n218643 , n218642 , n218594 );
and ( n218644 , n218585 , n218340 );
or ( n218645 , n218643 , n218644 );
not ( n218646 , n218397 );
not ( n218647 , n216585 );
not ( n218648 , n218647 );
or ( n218649 , n218646 , n218648 );
not ( n218650 , n215075 );
not ( n218651 , n216593 );
or ( n218652 , n218650 , n218651 );
nand ( n218653 , n216572 , n215899 );
nand ( n218654 , n218652 , n218653 );
nand ( n218655 , n218654 , n217824 );
nand ( n218656 , n218649 , n218655 );
not ( n218657 , n215966 );
not ( n218658 , n217017 );
not ( n218659 , n41563 );
or ( n218660 , n218658 , n218659 );
buf ( n218661 , n215971 );
nand ( n218662 , n41564 , n218661 );
nand ( n218663 , n218660 , n218662 );
not ( n218664 , n218663 );
or ( n218665 , n218657 , n218664 );
nand ( n218666 , n218494 , n217023 );
nand ( n218667 , n218665 , n218666 );
xor ( n218668 , n218656 , n218667 );
not ( n218669 , n218077 );
not ( n218670 , n214837 );
and ( n218671 , n216166 , n218670 );
not ( n218672 , n216166 );
and ( n218673 , n218672 , n214837 );
or ( n218674 , n218671 , n218673 );
not ( n218675 , n218674 );
or ( n218676 , n218669 , n218675 );
buf ( n218677 , n214609 );
not ( n218678 , n218677 );
nand ( n218679 , n218404 , n218678 );
nand ( n218680 , n218676 , n218679 );
xor ( n218681 , n218668 , n218680 );
xor ( n218682 , n218656 , n218667 );
and ( n218683 , n218682 , n218680 );
and ( n218684 , n218656 , n218667 );
or ( n218685 , n218683 , n218684 );
not ( n218686 , n218369 );
not ( n218687 , n218049 );
or ( n218688 , n218686 , n218687 );
not ( n218689 , n215117 );
not ( n218690 , n215569 );
or ( n218691 , n218689 , n218690 );
nand ( n218692 , n216968 , n213917 );
nand ( n218693 , n218691 , n218692 );
nand ( n218694 , n218693 , n215327 );
nand ( n218695 , n218688 , n218694 );
not ( n218696 , n215191 );
not ( n218697 , n215104 );
not ( n218698 , n214467 );
or ( n218699 , n218697 , n218698 );
nand ( n218700 , n215545 , n214468 );
nand ( n218701 , n218699 , n218700 );
not ( n218702 , n218701 );
or ( n218703 , n218696 , n218702 );
nand ( n218704 , n218360 , n215182 );
nand ( n218705 , n218703 , n218704 );
xor ( n218706 , n218695 , n218705 );
not ( n218707 , n214164 );
and ( n218708 , n41608 , n215956 );
not ( n218709 , n41608 );
and ( n218710 , n218709 , n216985 );
or ( n218711 , n218708 , n218710 );
not ( n218712 , n218711 );
or ( n218713 , n218707 , n218712 );
nand ( n218714 , n218507 , n215963 );
nand ( n218715 , n218713 , n218714 );
xor ( n218716 , n218706 , n218715 );
not ( n218717 , n214808 );
not ( n218718 , n214747 );
not ( n218719 , n214488 );
or ( n218720 , n218718 , n218719 );
nand ( n218721 , n41725 , n216938 );
nand ( n218722 , n218720 , n218721 );
not ( n218723 , n218722 );
or ( n218724 , n218717 , n218723 );
nand ( n218725 , n218380 , n216426 );
nand ( n218726 , n218724 , n218725 );
xor ( n218727 , n218716 , n218726 );
xor ( n218728 , n218706 , n218715 );
and ( n218729 , n218728 , n218726 );
and ( n218730 , n218706 , n218715 );
or ( n218731 , n218729 , n218730 );
not ( n218732 , n218519 );
not ( n218733 , n216065 );
or ( n218734 , n218732 , n218733 );
not ( n218735 , n216934 );
not ( n218736 , n216074 );
not ( n218737 , n218736 );
or ( n218738 , n218735 , n218737 );
nand ( n218739 , n216403 , n217478 );
nand ( n218740 , n218738 , n218739 );
nand ( n218741 , n216332 , n218740 );
nand ( n218742 , n218734 , n218741 );
not ( n218743 , n218551 );
not ( n218744 , n217380 );
or ( n218745 , n218743 , n218744 );
not ( n218746 , n216964 );
not ( n218747 , n217076 );
or ( n218748 , n218746 , n218747 );
nand ( n218749 , n216929 , n214678 );
nand ( n218750 , n218748 , n218749 );
nand ( n218751 , n218750 , n217099 );
nand ( n218752 , n218745 , n218751 );
xor ( n218753 , n218742 , n218752 );
not ( n218754 , n218562 );
not ( n218755 , n217890 );
or ( n218756 , n218754 , n218755 );
not ( n218757 , n217044 );
not ( n218758 , n217611 );
or ( n218759 , n218757 , n218758 );
nand ( n218760 , n217634 , n215131 );
nand ( n218761 , n218759 , n218760 );
not ( n218762 , n217229 );
nand ( n218763 , n218761 , n218762 );
nand ( n218764 , n218756 , n218763 );
xor ( n218765 , n218753 , n218764 );
xor ( n218766 , n218765 , n218727 );
not ( n218767 , n218532 );
not ( n218768 , n218221 );
or ( n218769 , n218767 , n218768 );
not ( n218770 , n213583 );
buf ( n218771 , n218217 );
not ( n218772 , n218771 );
not ( n218773 , n218772 );
or ( n218774 , n218770 , n218773 );
not ( n218775 , n218226 );
nand ( n218776 , n218775 , n214134 );
nand ( n218777 , n218774 , n218776 );
nand ( n218778 , n218777 , n218232 );
nand ( n218779 , n218769 , n218778 );
xor ( n218780 , n218766 , n218779 );
xor ( n218781 , n218637 , n218780 );
not ( n218782 , n214694 );
not ( n218783 , n216810 );
not ( n218784 , n217130 );
or ( n218785 , n218783 , n218784 );
not ( n218786 , n216500 );
nand ( n218787 , n218786 , n215289 );
nand ( n218788 , n218785 , n218787 );
not ( n218789 , n218788 );
or ( n218790 , n218782 , n218789 );
nand ( n218791 , n216299 , n218435 );
nand ( n218792 , n218790 , n218791 );
xor ( n218793 , n218792 , n218681 );
not ( n218794 , n216336 );
not ( n218795 , n213735 );
not ( n218796 , n217710 );
or ( n218797 , n218795 , n218796 );
nand ( n218798 , n41165 , n213732 );
nand ( n218799 , n218797 , n218798 );
not ( n218800 , n218799 );
or ( n218801 , n218794 , n218800 );
nand ( n218802 , n218424 , n213577 );
nand ( n218803 , n218801 , n218802 );
xor ( n218804 , n218793 , n218803 );
xor ( n218805 , n218781 , n218804 );
xor ( n218806 , n218637 , n218780 );
and ( n218807 , n218806 , n218804 );
and ( n218808 , n218637 , n218780 );
or ( n218809 , n218807 , n218808 );
not ( n218810 , n37623 );
not ( n218811 , n36641 );
or ( n218812 , n218810 , n218811 );
nand ( n218813 , n218812 , n36408 );
not ( n218814 , n218813 );
not ( n218815 , n218814 );
and ( n218816 , n215999 , n218815 );
not ( n218817 , n215999 );
buf ( n218818 , n218814 );
and ( n218819 , n218817 , n218818 );
nor ( n218820 , n218816 , n218819 );
not ( n218821 , n218820 );
not ( n218822 , n218217 );
not ( n218823 , n218452 );
or ( n218824 , n218822 , n218823 );
nand ( n218825 , n218204 , n218449 );
nand ( n218826 , n218824 , n218825 );
not ( n218827 , n218449 );
not ( n218828 , n218813 );
or ( n218829 , n218827 , n218828 );
not ( n218830 , n218813 );
nand ( n218831 , n218830 , n218452 );
nand ( n218832 , n218829 , n218831 );
nor ( n218833 , n218826 , n218832 );
not ( n218834 , n218833 );
not ( n218835 , n218834 );
not ( n218836 , n218835 );
or ( n218837 , n218821 , n218836 );
not ( n218838 , n218224 );
not ( n218839 , n218814 );
or ( n218840 , n218838 , n218839 );
nand ( n218841 , n218815 , n216076 );
nand ( n218842 , n218840 , n218841 );
buf ( n218843 , n218455 );
nand ( n218844 , n218842 , n218843 );
nand ( n218845 , n218837 , n218844 );
xor ( n218846 , n218845 , n218621 );
xor ( n218847 , n218846 , n218625 );
xor ( n218848 , n218641 , n218847 );
xor ( n218849 , n218848 , n218645 );
xor ( n218850 , n218641 , n218847 );
and ( n218851 , n218850 , n218645 );
and ( n218852 , n218641 , n218847 );
or ( n218853 , n218851 , n218852 );
not ( n218854 , n216239 );
not ( n218855 , n217944 );
not ( n218856 , n218855 );
not ( n218857 , n216520 );
or ( n218858 , n218856 , n218857 );
nand ( n218859 , n216519 , n217944 );
nand ( n218860 , n218858 , n218859 );
not ( n218861 , n218860 );
or ( n218862 , n218854 , n218861 );
nand ( n218863 , n218479 , n214717 );
nand ( n218864 , n218862 , n218863 );
xor ( n218865 , n218389 , n218864 );
not ( n218866 , n218208 );
nand ( n218867 , n218449 , n215999 );
nand ( n218868 , n218866 , n218867 );
nand ( n218869 , n218452 , n213751 );
and ( n218870 , n218868 , n218869 );
not ( n218871 , n37623 );
not ( n218872 , n36641 );
or ( n218873 , n218871 , n218872 );
nand ( n218874 , n218873 , n36408 );
not ( n218875 , n218874 );
buf ( n218876 , n218875 );
nor ( n218877 , n218870 , n218876 );
xor ( n218878 , n218865 , n218877 );
xor ( n218879 , n218629 , n218878 );
not ( n218880 , n217142 );
not ( n218881 , n214818 );
buf ( n218882 , n207986 );
not ( n218883 , n218882 );
buf ( n218884 , n218883 );
not ( n218885 , n218884 );
or ( n218886 , n218881 , n218885 );
not ( n218887 , n216262 );
nand ( n218888 , n40710 , n218887 );
nand ( n218889 , n218886 , n218888 );
not ( n218890 , n218889 );
or ( n218891 , n218880 , n218890 );
nand ( n218892 , n218580 , n213874 );
nand ( n218893 , n218891 , n218892 );
xor ( n218894 , n218879 , n218893 );
xor ( n218895 , n218488 , n218894 );
xor ( n218896 , n218415 , n218617 );
not ( n218897 , n217571 );
not ( n218898 , n213960 );
not ( n218899 , n217119 );
or ( n218900 , n218898 , n218899 );
nand ( n218901 , n218137 , n215600 );
nand ( n218902 , n218900 , n218901 );
not ( n218903 , n218902 );
or ( n218904 , n218897 , n218903 );
nand ( n218905 , n218464 , n215605 );
nand ( n218906 , n218904 , n218905 );
xor ( n218907 , n218896 , n218906 );
xor ( n218908 , n218907 , n218633 );
not ( n218909 , n214319 );
not ( n218910 , n213382 );
buf ( n218911 , n208078 );
not ( n218912 , n218911 );
not ( n218913 , n218912 );
or ( n218914 , n218910 , n218913 );
nand ( n218915 , n218911 , n217715 );
nand ( n218916 , n218914 , n218915 );
not ( n218917 , n218916 );
or ( n218918 , n218909 , n218917 );
nand ( n218919 , n218591 , n217969 );
nand ( n218920 , n218918 , n218919 );
xor ( n218921 , n218908 , n218920 );
xor ( n218922 , n218895 , n218921 );
xor ( n218923 , n218488 , n218894 );
and ( n218924 , n218923 , n218921 );
and ( n218925 , n218488 , n218894 );
or ( n218926 , n218924 , n218925 );
xor ( n218927 , n218805 , n218542 );
xor ( n218928 , n218927 , n218849 );
xor ( n218929 , n218805 , n218542 );
and ( n218930 , n218929 , n218849 );
and ( n218931 , n218805 , n218542 );
or ( n218932 , n218930 , n218931 );
xor ( n218933 , n218574 , n218922 );
xor ( n218934 , n218933 , n218601 );
xor ( n218935 , n218574 , n218922 );
and ( n218936 , n218935 , n218601 );
and ( n218937 , n218574 , n218922 );
or ( n218938 , n218936 , n218937 );
xor ( n218939 , n218928 , n218607 );
xor ( n218940 , n218939 , n218934 );
xor ( n218941 , n218928 , n218607 );
and ( n218942 , n218941 , n218934 );
and ( n218943 , n218928 , n218607 );
or ( n218944 , n218942 , n218943 );
xor ( n218945 , n218742 , n218752 );
and ( n218946 , n218945 , n218764 );
and ( n218947 , n218742 , n218752 );
or ( n218948 , n218946 , n218947 );
xor ( n218949 , n218389 , n218864 );
and ( n218950 , n218949 , n218877 );
and ( n218951 , n218389 , n218864 );
or ( n218952 , n218950 , n218951 );
xor ( n218953 , n218415 , n218617 );
and ( n218954 , n218953 , n218906 );
and ( n218955 , n218415 , n218617 );
or ( n218956 , n218954 , n218955 );
xor ( n218957 , n218792 , n218681 );
and ( n218958 , n218957 , n218803 );
and ( n218959 , n218792 , n218681 );
or ( n218960 , n218958 , n218959 );
xor ( n218961 , n218765 , n218727 );
and ( n218962 , n218961 , n218779 );
and ( n218963 , n218765 , n218727 );
or ( n218964 , n218962 , n218963 );
xor ( n218965 , n218845 , n218621 );
and ( n218966 , n218965 , n218625 );
and ( n218967 , n218845 , n218621 );
or ( n218968 , n218966 , n218967 );
xor ( n218969 , n218629 , n218878 );
and ( n218970 , n218969 , n218893 );
and ( n218971 , n218629 , n218878 );
or ( n218972 , n218970 , n218971 );
xor ( n218973 , n218907 , n218633 );
and ( n218974 , n218973 , n218920 );
and ( n218975 , n218907 , n218633 );
or ( n218976 , n218974 , n218975 );
not ( n218977 , n215578 );
not ( n218978 , n218693 );
or ( n218979 , n218977 , n218978 );
buf ( n218980 , n214597 );
not ( n218981 , n218980 );
not ( n218982 , n218981 );
not ( n218983 , n215512 );
or ( n218984 , n218982 , n218983 );
nand ( n218985 , n216968 , n218980 );
nand ( n218986 , n218984 , n218985 );
nand ( n218987 , n218986 , n216458 );
nand ( n218988 , n218979 , n218987 );
not ( n218989 , n215550 );
buf ( n218990 , n215104 );
not ( n218991 , n218990 );
not ( n218992 , n216290 );
or ( n218993 , n218991 , n218992 );
not ( n218994 , n218990 );
nand ( n218995 , n30997 , n218994 );
nand ( n218996 , n218993 , n218995 );
not ( n218997 , n218996 );
or ( n218998 , n218989 , n218997 );
nand ( n218999 , n215183 , n218701 );
nand ( n219000 , n218998 , n218999 );
xor ( n219001 , n218988 , n219000 );
not ( n219002 , n218654 );
not ( n219003 , n217505 );
or ( n219004 , n219002 , n219003 );
not ( n219005 , n218514 );
not ( n219006 , n216593 );
or ( n219007 , n219005 , n219006 );
nand ( n219008 , n216421 , n216170 );
nand ( n219009 , n219007 , n219008 );
nand ( n219010 , n219009 , n216201 );
nand ( n219011 , n219004 , n219010 );
xor ( n219012 , n219001 , n219011 );
xor ( n219013 , n218988 , n219000 );
and ( n219014 , n219013 , n219011 );
and ( n219015 , n218988 , n219000 );
or ( n219016 , n219014 , n219015 );
not ( n219017 , n214164 );
not ( n219018 , n217542 );
not ( n219019 , n215820 );
or ( n219020 , n219018 , n219019 );
nand ( n219021 , n211451 , n216989 );
nand ( n219022 , n219020 , n219021 );
not ( n219023 , n219022 );
or ( n219024 , n219017 , n219023 );
nand ( n219025 , n218711 , n215963 );
nand ( n219026 , n219024 , n219025 );
not ( n219027 , n218678 );
not ( n219028 , n218674 );
or ( n219029 , n219027 , n219028 );
not ( n219030 , n216166 );
not ( n219031 , n208726 );
or ( n219032 , n219030 , n219031 );
buf ( n219033 , n214416 );
not ( n219034 , n219033 );
nand ( n219035 , n219034 , n208725 );
nand ( n219036 , n219032 , n219035 );
nand ( n219037 , n219036 , n214458 );
nand ( n219038 , n219029 , n219037 );
xor ( n219039 , n219026 , n219038 );
and ( n219040 , n218695 , n218705 );
xor ( n219041 , n219039 , n219040 );
xor ( n219042 , n219026 , n219038 );
and ( n219043 , n219042 , n219040 );
and ( n219044 , n219026 , n219038 );
or ( n219045 , n219043 , n219044 );
not ( n219046 , n214717 );
not ( n219047 , n218860 );
or ( n219048 , n219046 , n219047 );
not ( n219049 , n218855 );
not ( n219050 , n216858 );
not ( n219051 , n219050 );
not ( n219052 , n219051 );
or ( n219053 , n219049 , n219052 );
nand ( n219054 , n208164 , n217944 );
nand ( n219055 , n219053 , n219054 );
nand ( n219056 , n219055 , n216239 );
nand ( n219057 , n219048 , n219056 );
buf ( n219058 , n34087 );
not ( n219059 , n219058 );
buf ( n219060 , n33647 );
nor ( n219061 , n219059 , n219060 );
and ( n219062 , n37571 , n219061 );
not ( n219063 , n219062 );
buf ( n219064 , n36319 );
nand ( n219065 , n219064 , n37583 );
not ( n219066 , n219065 );
or ( n219067 , n219063 , n219066 );
not ( n219068 , n219065 );
not ( n219069 , n37571 );
or ( n219070 , n219068 , n219069 );
not ( n219071 , n219061 );
nand ( n219072 , n219070 , n219071 );
nand ( n219073 , n219067 , n219072 );
xnor ( n219074 , n218813 , n219073 );
not ( n219075 , n219074 );
buf ( n219076 , n219075 );
not ( n219077 , n219076 );
nor ( n219078 , n219077 , n213751 );
xor ( n219079 , n219057 , n219078 );
xor ( n219080 , n219079 , n218685 );
xor ( n219081 , n218960 , n219080 );
xor ( n219082 , n219081 , n218964 );
xor ( n219083 , n218960 , n219080 );
and ( n219084 , n219083 , n218964 );
and ( n219085 , n218960 , n219080 );
or ( n219086 , n219084 , n219085 );
xor ( n219087 , n219041 , n218948 );
not ( n219088 , n214808 );
not ( n219089 , n214747 );
not ( n219090 , n214642 );
or ( n219091 , n219089 , n219090 );
not ( n219092 , n214786 );
nand ( n219093 , n41716 , n219092 );
nand ( n219094 , n219091 , n219093 );
not ( n219095 , n219094 );
or ( n219096 , n219088 , n219095 );
nand ( n219097 , n218722 , n214799 );
nand ( n219098 , n219096 , n219097 );
not ( n219099 , n218740 );
not ( n219100 , n216065 );
or ( n219101 , n219099 , n219100 );
not ( n219102 , n216139 );
not ( n219103 , n219102 );
not ( n219104 , n216014 );
or ( n219105 , n219103 , n219104 );
nand ( n219106 , n216623 , n216139 );
nand ( n219107 , n219105 , n219106 );
nand ( n219108 , n219107 , n217047 );
nand ( n219109 , n219101 , n219108 );
xor ( n219110 , n219098 , n219109 );
not ( n219111 , n218750 );
not ( n219112 , n217089 );
or ( n219113 , n219111 , n219112 );
not ( n219114 , n216208 );
not ( n219115 , n217602 );
or ( n219116 , n219114 , n219115 );
nand ( n219117 , n216929 , n216207 );
nand ( n219118 , n219116 , n219117 );
not ( n219119 , n217098 );
nand ( n219120 , n219118 , n219119 );
nand ( n219121 , n219113 , n219120 );
xor ( n219122 , n219110 , n219121 );
xor ( n219123 , n219087 , n219122 );
xor ( n219124 , n219123 , n218968 );
not ( n219125 , n218842 );
not ( n219126 , n218835 );
or ( n219127 , n219125 , n219126 );
not ( n219128 , n218876 );
and ( n219129 , n213347 , n219128 );
not ( n219130 , n213347 );
and ( n219131 , n219130 , n218876 );
nor ( n219132 , n219129 , n219131 );
nand ( n219133 , n219132 , n218843 );
nand ( n219134 , n219127 , n219133 );
not ( n219135 , n218777 );
not ( n219136 , n218221 );
or ( n219137 , n219135 , n219136 );
not ( n219138 , n214956 );
not ( n219139 , n218209 );
or ( n219140 , n219138 , n219139 );
not ( n219141 , n218226 );
nand ( n219142 , n219141 , n214960 );
nand ( n219143 , n219140 , n219142 );
nand ( n219144 , n219143 , n218231 );
nand ( n219145 , n219137 , n219144 );
xor ( n219146 , n219134 , n219145 );
not ( n219147 , n216336 );
not ( n219148 , n213732 );
not ( n219149 , n208002 );
or ( n219150 , n219148 , n219149 );
not ( n219151 , n40724 );
nand ( n219152 , n219151 , n213735 );
nand ( n219153 , n219150 , n219152 );
not ( n219154 , n219153 );
or ( n219155 , n219147 , n219154 );
nand ( n219156 , n218799 , n213577 );
nand ( n219157 , n219155 , n219156 );
xor ( n219158 , n219146 , n219157 );
xor ( n219159 , n219124 , n219158 );
xor ( n219160 , n219123 , n218968 );
and ( n219161 , n219160 , n219158 );
and ( n219162 , n219123 , n218968 );
or ( n219163 , n219161 , n219162 );
xor ( n219164 , n218952 , n218956 );
not ( n219165 , n218761 );
not ( n219166 , n217631 );
or ( n219167 , n219165 , n219166 );
not ( n219168 , n214537 );
not ( n219169 , n217637 );
or ( n219170 , n219168 , n219169 );
nand ( n219171 , n217634 , n214899 );
nand ( n219172 , n219170 , n219171 );
nand ( n219173 , n219172 , n217641 );
nand ( n219174 , n219167 , n219173 );
buf ( n219175 , n215966 );
not ( n219176 , n219175 );
not ( n219177 , n217017 );
not ( n219178 , n217941 );
or ( n219179 , n219177 , n219178 );
nand ( n219180 , n215796 , n215971 );
nand ( n219181 , n219179 , n219180 );
not ( n219182 , n219181 );
or ( n219183 , n219176 , n219182 );
nand ( n219184 , n218663 , n217023 );
nand ( n219185 , n219183 , n219184 );
xor ( n219186 , n219174 , n219185 );
xor ( n219187 , n219186 , n219012 );
xor ( n219188 , n219164 , n219187 );
xor ( n219189 , n218972 , n219188 );
xor ( n219190 , n219189 , n218976 );
xor ( n219191 , n218972 , n219188 );
and ( n219192 , n219191 , n218976 );
and ( n219193 , n218972 , n219188 );
or ( n219194 , n219192 , n219193 );
not ( n219195 , n214086 );
not ( n219196 , n218902 );
or ( n219197 , n219195 , n219196 );
not ( n219198 , n213960 );
not ( n219199 , n41070 );
or ( n219200 , n219198 , n219199 );
buf ( n219201 , n41069 );
nand ( n219202 , n219201 , n215600 );
nand ( n219203 , n219200 , n219202 );
nand ( n219204 , n219203 , n217571 );
nand ( n219205 , n219197 , n219204 );
xor ( n219206 , n218731 , n219205 );
not ( n219207 , n214694 );
not ( n219208 , n216810 );
not ( n219209 , n216307 );
or ( n219210 , n219208 , n219209 );
nand ( n219211 , n216311 , n215289 );
nand ( n219212 , n219210 , n219211 );
not ( n219213 , n219212 );
or ( n219214 , n219207 , n219213 );
nand ( n219215 , n218788 , n216299 );
nand ( n219216 , n219214 , n219215 );
xor ( n219217 , n219206 , n219216 );
not ( n219218 , n217969 );
not ( n219219 , n218916 );
or ( n219220 , n219218 , n219219 );
not ( n219221 , n213382 );
buf ( n219222 , n40559 );
not ( n219223 , n219222 );
not ( n219224 , n219223 );
or ( n219225 , n219221 , n219224 );
buf ( n219226 , n40558 );
nand ( n219227 , n219226 , n213381 );
nand ( n219228 , n219225 , n219227 );
nand ( n219229 , n219228 , n211314 );
nand ( n219230 , n219220 , n219229 );
xor ( n219231 , n219217 , n219230 );
not ( n219232 , n217142 );
not ( n219233 , n214818 );
not ( n219234 , n218590 );
buf ( n219235 , n219234 );
not ( n219236 , n219235 );
or ( n219237 , n219233 , n219236 );
not ( n219238 , n40764 );
not ( n219239 , n219238 );
nand ( n219240 , n219239 , n214824 );
nand ( n219241 , n219237 , n219240 );
not ( n219242 , n219241 );
or ( n219243 , n219232 , n219242 );
nand ( n219244 , n218889 , n213874 );
nand ( n219245 , n219243 , n219244 );
xor ( n219246 , n219231 , n219245 );
xor ( n219247 , n219082 , n219246 );
xor ( n219248 , n219247 , n218809 );
xor ( n219249 , n219082 , n219246 );
and ( n219250 , n219249 , n218809 );
and ( n219251 , n219082 , n219246 );
or ( n219252 , n219250 , n219251 );
xor ( n219253 , n218853 , n219159 );
xor ( n219254 , n219253 , n218926 );
xor ( n219255 , n218853 , n219159 );
and ( n219256 , n219255 , n218926 );
and ( n219257 , n218853 , n219159 );
or ( n219258 , n219256 , n219257 );
xor ( n219259 , n219190 , n219248 );
xor ( n219260 , n219259 , n218932 );
xor ( n219261 , n219190 , n219248 );
and ( n219262 , n219261 , n218932 );
and ( n219263 , n219190 , n219248 );
or ( n219264 , n219262 , n219263 );
xor ( n219265 , n219254 , n218938 );
xor ( n219266 , n219265 , n219260 );
xor ( n219267 , n219254 , n218938 );
and ( n219268 , n219267 , n219260 );
and ( n219269 , n219254 , n218938 );
or ( n219270 , n219268 , n219269 );
xor ( n219271 , n219098 , n219109 );
and ( n219272 , n219271 , n219121 );
and ( n219273 , n219098 , n219109 );
or ( n219274 , n219272 , n219273 );
xor ( n219275 , n219174 , n219185 );
and ( n219276 , n219275 , n219012 );
and ( n219277 , n219174 , n219185 );
or ( n219278 , n219276 , n219277 );
xor ( n219279 , n219057 , n219078 );
and ( n219280 , n219279 , n218685 );
and ( n219281 , n219057 , n219078 );
or ( n219282 , n219280 , n219281 );
xor ( n219283 , n218731 , n219205 );
and ( n219284 , n219283 , n219216 );
and ( n219285 , n218731 , n219205 );
or ( n219286 , n219284 , n219285 );
xor ( n219287 , n219041 , n218948 );
and ( n219288 , n219287 , n219122 );
and ( n219289 , n219041 , n218948 );
or ( n219290 , n219288 , n219289 );
xor ( n219291 , n219134 , n219145 );
and ( n219292 , n219291 , n219157 );
and ( n219293 , n219134 , n219145 );
or ( n219294 , n219292 , n219293 );
xor ( n219295 , n218952 , n218956 );
and ( n219296 , n219295 , n219187 );
and ( n219297 , n218952 , n218956 );
or ( n219298 , n219296 , n219297 );
xor ( n219299 , n219217 , n219230 );
and ( n219300 , n219299 , n219245 );
and ( n219301 , n219217 , n219230 );
or ( n219302 , n219300 , n219301 );
not ( n219303 , n218077 );
not ( n219304 , n216166 );
not ( n219305 , n216608 );
not ( n219306 , n219305 );
or ( n219307 , n219304 , n219306 );
nand ( n219308 , n216603 , n219034 );
nand ( n219309 , n219307 , n219308 );
not ( n219310 , n219309 );
or ( n219311 , n219303 , n219310 );
nand ( n219312 , n219036 , n214449 );
nand ( n219313 , n219311 , n219312 );
buf ( n219314 , n214808 );
not ( n219315 , n219314 );
xor ( n219316 , n216938 , n216530 );
not ( n219317 , n219316 );
or ( n219318 , n219315 , n219317 );
nand ( n219319 , n216426 , n219094 );
nand ( n219320 , n219318 , n219319 );
xor ( n219321 , n219313 , n219320 );
not ( n219322 , n215550 );
not ( n219323 , n215165 );
not ( n219324 , n214820 );
or ( n219325 , n219323 , n219324 );
not ( n219326 , n215165 );
nand ( n219327 , n41725 , n219326 );
nand ( n219328 , n219325 , n219327 );
not ( n219329 , n219328 );
or ( n219330 , n219322 , n219329 );
not ( n219331 , n215182 );
not ( n219332 , n219331 );
nand ( n219333 , n218996 , n219332 );
nand ( n219334 , n219330 , n219333 );
xor ( n219335 , n219321 , n219334 );
xor ( n219336 , n219313 , n219320 );
and ( n219337 , n219336 , n219334 );
and ( n219338 , n219313 , n219320 );
or ( n219339 , n219337 , n219338 );
not ( n219340 , n219107 );
not ( n219341 , n216324 );
or ( n219342 , n219340 , n219341 );
buf ( n219343 , n215117 );
not ( n219344 , n219343 );
not ( n219345 , n218736 );
or ( n219346 , n219344 , n219345 );
not ( n219347 , n216014 );
not ( n219348 , n219343 );
nand ( n219349 , n219347 , n219348 );
nand ( n219350 , n219346 , n219349 );
nand ( n219351 , n217047 , n219350 );
nand ( n219352 , n219342 , n219351 );
not ( n219353 , n217549 );
not ( n219354 , n219353 );
not ( n219355 , n217542 );
not ( n219356 , n216543 );
or ( n219357 , n219355 , n219356 );
not ( n219358 , n215955 );
nand ( n219359 , n41564 , n219358 );
nand ( n219360 , n219357 , n219359 );
not ( n219361 , n219360 );
or ( n219362 , n219354 , n219361 );
nand ( n219363 , n219022 , n215963 );
nand ( n219364 , n219362 , n219363 );
xor ( n219365 , n219352 , n219364 );
not ( n219366 , n219118 );
buf ( n219367 , n217875 );
buf ( n219368 , n219367 );
not ( n219369 , n219368 );
or ( n219370 , n219366 , n219369 );
not ( n219371 , n215075 );
not ( n219372 , n217602 );
or ( n219373 , n219371 , n219372 );
nand ( n219374 , n217080 , n215899 );
nand ( n219375 , n219373 , n219374 );
nand ( n219376 , n219375 , n217388 );
nand ( n219377 , n219370 , n219376 );
xor ( n219378 , n219365 , n219377 );
xor ( n219379 , n219352 , n219364 );
and ( n219380 , n219379 , n219377 );
and ( n219381 , n219352 , n219364 );
or ( n219382 , n219380 , n219381 );
xor ( n219383 , n219335 , n219378 );
not ( n219384 , n215137 );
not ( n219385 , n217573 );
not ( n219386 , n41165 );
not ( n219387 , n219386 );
or ( n219388 , n219385 , n219387 );
buf ( n219389 , n217714 );
not ( n219390 , n213960 );
nand ( n219391 , n219389 , n219390 );
nand ( n219392 , n219388 , n219391 );
not ( n219393 , n219392 );
or ( n219394 , n219384 , n219393 );
nand ( n219395 , n219203 , n218467 );
nand ( n219396 , n219394 , n219395 );
xor ( n219397 , n219383 , n219396 );
xor ( n219398 , n219290 , n219397 );
xor ( n219399 , n219398 , n219294 );
xor ( n219400 , n219290 , n219397 );
and ( n219401 , n219400 , n219294 );
and ( n219402 , n219290 , n219397 );
or ( n219403 , n219401 , n219402 );
not ( n219404 , n213750 );
and ( n219405 , n37583 , n219058 );
not ( n219406 , n219405 );
not ( n219407 , n219064 );
or ( n219408 , n219406 , n219407 );
and ( n219409 , n37548 , n219058 );
nor ( n219410 , n219409 , n219060 );
nand ( n219411 , n219408 , n219410 );
and ( n219412 , n219411 , n37591 );
not ( n219413 , n219411 );
and ( n219414 , n219413 , n37592 );
nor ( n219415 , n219412 , n219414 );
buf ( n219416 , n219415 );
not ( n219417 , n219416 );
not ( n219418 , n219417 );
not ( n219419 , n219418 );
buf ( n219420 , n219419 );
not ( n219421 , n219420 );
or ( n219422 , n219404 , n219421 );
buf ( n219423 , n219417 );
not ( n219424 , n219423 );
nand ( n219425 , n219424 , n213751 );
nand ( n219426 , n219422 , n219425 );
not ( n219427 , n219426 );
and ( n219428 , n219073 , n219416 );
not ( n219429 , n219073 );
not ( n219430 , n219415 );
and ( n219431 , n219429 , n219430 );
nor ( n219432 , n219428 , n219431 );
nand ( n219433 , n219432 , n219074 );
buf ( n219434 , n219433 );
not ( n219435 , n219434 );
not ( n219436 , n219435 );
or ( n219437 , n219427 , n219436 );
not ( n219438 , n218224 );
buf ( n219439 , n219430 );
buf ( n219440 , n219439 );
not ( n219441 , n219440 );
or ( n219442 , n219438 , n219441 );
not ( n219443 , n219440 );
nand ( n219444 , n219443 , n216076 );
nand ( n219445 , n219442 , n219444 );
nand ( n219446 , n219445 , n219076 );
nand ( n219447 , n219437 , n219446 );
not ( n219448 , n219132 );
not ( n219449 , n218834 );
not ( n219450 , n219449 );
or ( n219451 , n219448 , n219450 );
not ( n219452 , n213583 );
not ( n219453 , n218818 );
or ( n219454 , n219452 , n219453 );
nand ( n219455 , n218815 , n214134 );
nand ( n219456 , n219454 , n219455 );
nand ( n219457 , n219456 , n218843 );
nand ( n219458 , n219451 , n219457 );
xor ( n219459 , n219447 , n219458 );
not ( n219460 , n219143 );
buf ( n219461 , n218525 );
not ( n219462 , n219461 );
or ( n219463 , n219460 , n219462 );
and ( n219464 , n214357 , n218771 );
not ( n219465 , n214357 );
and ( n219466 , n219465 , n218772 );
nor ( n219467 , n219464 , n219466 );
nand ( n219468 , n219467 , n218533 );
nand ( n219469 , n219463 , n219468 );
xor ( n219470 , n219459 , n219469 );
xor ( n219471 , n219470 , n219298 );
not ( n219472 , n219172 );
not ( n219473 , n217631 );
or ( n219474 , n219472 , n219473 );
not ( n219475 , n214678 );
not ( n219476 , n219475 );
not ( n219477 , n217637 );
or ( n219478 , n219476 , n219477 );
nand ( n219479 , n217614 , n214678 );
nand ( n219480 , n219478 , n219479 );
nand ( n219481 , n219480 , n217230 );
nand ( n219482 , n219474 , n219481 );
not ( n219483 , n218986 );
not ( n219484 , n215773 );
or ( n219485 , n219483 , n219484 );
not ( n219486 , n214190 );
and ( n219487 , n216280 , n219486 );
not ( n219488 , n216280 );
and ( n219489 , n219488 , n214467 );
or ( n219490 , n219487 , n219489 );
nand ( n219491 , n219490 , n215762 );
nand ( n219492 , n219485 , n219491 );
not ( n219493 , n219009 );
not ( n219494 , n216586 );
or ( n219495 , n219493 , n219494 );
not ( n219496 , n216934 );
not ( n219497 , n216569 );
or ( n219498 , n219496 , n219497 );
nand ( n219499 , n216594 , n217478 );
nand ( n219500 , n219498 , n219499 );
not ( n219501 , n216200 );
nand ( n219502 , n219500 , n219501 );
nand ( n219503 , n219495 , n219502 );
xor ( n219504 , n219492 , n219503 );
xor ( n219505 , n219482 , n219504 );
xor ( n219506 , n219505 , n219016 );
xor ( n219507 , n219506 , n219278 );
xor ( n219508 , n219507 , n219282 );
xor ( n219509 , n219471 , n219508 );
xor ( n219510 , n219470 , n219298 );
and ( n219511 , n219510 , n219508 );
and ( n219512 , n219470 , n219298 );
or ( n219513 , n219511 , n219512 );
not ( n219514 , n217969 );
not ( n219515 , n219228 );
or ( n219516 , n219514 , n219515 );
not ( n219517 , n213382 );
not ( n219518 , n40625 );
not ( n219519 , n219518 );
or ( n219520 , n219517 , n219519 );
not ( n219521 , n40623 );
not ( n219522 , n219521 );
nand ( n219523 , n219522 , n213381 );
nand ( n219524 , n219520 , n219523 );
nand ( n219525 , n219524 , n213912 );
nand ( n219526 , n219516 , n219525 );
not ( n219527 , n213874 );
not ( n219528 , n219241 );
or ( n219529 , n219527 , n219528 );
and ( n219530 , n216262 , n218912 );
not ( n219531 , n216262 );
not ( n219532 , n208078 );
not ( n219533 , n219532 );
and ( n219534 , n219531 , n219533 );
or ( n219535 , n219530 , n219534 );
nand ( n219536 , n219535 , n217142 );
nand ( n219537 , n219529 , n219536 );
xor ( n219538 , n219526 , n219537 );
not ( n219539 , n216239 );
not ( n219540 , n218855 );
not ( n219541 , n217119 );
or ( n219542 , n219540 , n219541 );
nand ( n219543 , n217564 , n216037 );
nand ( n219544 , n219542 , n219543 );
not ( n219545 , n219544 );
or ( n219546 , n219539 , n219545 );
nand ( n219547 , n219055 , n214717 );
nand ( n219548 , n219546 , n219547 );
and ( n219549 , n219073 , n213750 );
nor ( n219550 , n219549 , n218815 );
not ( n219551 , n213751 );
nor ( n219552 , n219551 , n219073 );
or ( n219553 , n219550 , n219552 );
nand ( n219554 , n219553 , n219424 );
not ( n219555 , n219554 );
xor ( n219556 , n219548 , n219555 );
xor ( n219557 , n219556 , n219045 );
xor ( n219558 , n219538 , n219557 );
xor ( n219559 , n219302 , n219558 );
xor ( n219560 , n219559 , n219086 );
xor ( n219561 , n219302 , n219558 );
and ( n219562 , n219561 , n219086 );
and ( n219563 , n219302 , n219558 );
or ( n219564 , n219562 , n219563 );
not ( n219565 , n216299 );
not ( n219566 , n219212 );
or ( n219567 , n219565 , n219566 );
not ( n219568 , n216810 );
not ( n219569 , n217147 );
or ( n219570 , n219568 , n219569 );
nand ( n219571 , n218283 , n215289 );
nand ( n219572 , n219570 , n219571 );
nand ( n219573 , n219572 , n214694 );
nand ( n219574 , n219567 , n219573 );
xor ( n219575 , n219274 , n219574 );
not ( n219576 , n219175 );
not ( n219577 , n218661 );
not ( n219578 , n219577 );
not ( n219579 , n215989 );
or ( n219580 , n219578 , n219579 );
not ( n219581 , n41396 );
not ( n219582 , n219581 );
not ( n219583 , n217017 );
nand ( n219584 , n219582 , n219583 );
nand ( n219585 , n219580 , n219584 );
not ( n219586 , n219585 );
or ( n219587 , n219576 , n219586 );
nand ( n219588 , n219181 , n217023 );
nand ( n219589 , n219587 , n219588 );
xor ( n219590 , n219575 , n219589 );
xor ( n219591 , n219286 , n219590 );
not ( n219592 , n216336 );
not ( n219593 , n213735 );
buf ( n219594 , n218882 );
not ( n219595 , n219594 );
buf ( n219596 , n219595 );
not ( n219597 , n219596 );
or ( n219598 , n219593 , n219597 );
buf ( n219599 , n40710 );
nand ( n219600 , n219599 , n213732 );
nand ( n219601 , n219598 , n219600 );
not ( n219602 , n219601 );
or ( n219603 , n219592 , n219602 );
nand ( n219604 , n219153 , n213577 );
nand ( n219605 , n219603 , n219604 );
xor ( n219606 , n219591 , n219605 );
xor ( n219607 , n219606 , n219399 );
xor ( n219608 , n219607 , n219163 );
xor ( n219609 , n219606 , n219399 );
and ( n219610 , n219609 , n219163 );
and ( n219611 , n219606 , n219399 );
or ( n219612 , n219610 , n219611 );
xor ( n219613 , n219194 , n219509 );
xor ( n219614 , n219613 , n219252 );
xor ( n219615 , n219194 , n219509 );
and ( n219616 , n219615 , n219252 );
and ( n219617 , n219194 , n219509 );
or ( n219618 , n219616 , n219617 );
xor ( n219619 , n219560 , n219608 );
xor ( n219620 , n219619 , n219258 );
xor ( n219621 , n219560 , n219608 );
and ( n219622 , n219621 , n219258 );
and ( n219623 , n219560 , n219608 );
or ( n219624 , n219622 , n219623 );
xor ( n219625 , n219614 , n219264 );
xor ( n219626 , n219625 , n219620 );
xor ( n219627 , n219614 , n219264 );
and ( n219628 , n219627 , n219620 );
and ( n219629 , n219614 , n219264 );
or ( n219630 , n219628 , n219629 );
xor ( n219631 , n219482 , n219504 );
and ( n219632 , n219631 , n219016 );
and ( n219633 , n219482 , n219504 );
or ( n219634 , n219632 , n219633 );
xor ( n219635 , n219548 , n219555 );
and ( n219636 , n219635 , n219045 );
and ( n219637 , n219548 , n219555 );
or ( n219638 , n219636 , n219637 );
xor ( n219639 , n219274 , n219574 );
and ( n219640 , n219639 , n219589 );
and ( n219641 , n219274 , n219574 );
or ( n219642 , n219640 , n219641 );
xor ( n219643 , n219335 , n219378 );
and ( n219644 , n219643 , n219396 );
and ( n219645 , n219335 , n219378 );
or ( n219646 , n219644 , n219645 );
xor ( n219647 , n219447 , n219458 );
and ( n219648 , n219647 , n219469 );
and ( n219649 , n219447 , n219458 );
or ( n219650 , n219648 , n219649 );
xor ( n219651 , n219506 , n219278 );
and ( n219652 , n219651 , n219282 );
and ( n219653 , n219506 , n219278 );
or ( n219654 , n219652 , n219653 );
xor ( n219655 , n219286 , n219590 );
and ( n219656 , n219655 , n219605 );
and ( n219657 , n219286 , n219590 );
or ( n219658 , n219656 , n219657 );
xor ( n219659 , n219526 , n219537 );
and ( n219660 , n219659 , n219557 );
and ( n219661 , n219526 , n219537 );
or ( n219662 , n219660 , n219661 );
not ( n219663 , n215587 );
not ( n219664 , n215766 );
not ( n219665 , n216290 );
or ( n219666 , n219664 , n219665 );
nand ( n219667 , n216293 , n216280 );
nand ( n219668 , n219666 , n219667 );
not ( n219669 , n219668 );
or ( n219670 , n219663 , n219669 );
nand ( n219671 , n216731 , n219490 );
nand ( n219672 , n219670 , n219671 );
not ( n219673 , n219500 );
not ( n219674 , n217289 );
or ( n219675 , n219673 , n219674 );
not ( n219676 , n219102 );
not ( n219677 , n216420 );
or ( n219678 , n219676 , n219677 );
nand ( n219679 , n216421 , n216139 );
nand ( n219680 , n219678 , n219679 );
nand ( n219681 , n219680 , n216598 );
nand ( n219682 , n219675 , n219681 );
xor ( n219683 , n219672 , n219682 );
not ( n219684 , n216426 );
not ( n219685 , n219316 );
or ( n219686 , n219684 , n219685 );
buf ( n219687 , n214786 );
not ( n219688 , n219687 );
not ( n219689 , n218503 );
not ( n219690 , n219689 );
not ( n219691 , n219690 );
or ( n219692 , n219688 , n219691 );
nand ( n219693 , n208725 , n216938 );
nand ( n219694 , n219692 , n219693 );
nand ( n219695 , n219694 , n219314 );
nand ( n219696 , n219686 , n219695 );
xor ( n219697 , n219683 , n219696 );
xor ( n219698 , n219672 , n219682 );
and ( n219699 , n219698 , n219696 );
and ( n219700 , n219672 , n219682 );
or ( n219701 , n219699 , n219700 );
not ( n219702 , n215183 );
not ( n219703 , n219328 );
or ( n219704 , n219702 , n219703 );
and ( n219705 , n41716 , n215545 );
not ( n219706 , n41716 );
and ( n219707 , n219706 , n215104 );
or ( n219708 , n219705 , n219707 );
nand ( n219709 , n215550 , n219708 );
nand ( n219710 , n219704 , n219709 );
not ( n219711 , n219350 );
not ( n219712 , n216324 );
or ( n219713 , n219711 , n219712 );
not ( n219714 , n218981 );
not ( n219715 , n216402 );
or ( n219716 , n219714 , n219715 );
nand ( n219717 , n216015 , n218980 );
nand ( n219718 , n219716 , n219717 );
nand ( n219719 , n217047 , n219718 );
nand ( n219720 , n219713 , n219719 );
xor ( n219721 , n219710 , n219720 );
not ( n219722 , n214458 );
not ( n219723 , n216166 );
not ( n219724 , n41700 );
not ( n219725 , n219724 );
or ( n219726 , n219723 , n219725 );
nand ( n219727 , n41701 , n219034 );
nand ( n219728 , n219726 , n219727 );
not ( n219729 , n219728 );
or ( n219730 , n219722 , n219729 );
buf ( n219731 , n218678 );
nand ( n219732 , n219309 , n219731 );
nand ( n219733 , n219730 , n219732 );
xor ( n219734 , n219721 , n219733 );
xor ( n219735 , n219710 , n219720 );
and ( n219736 , n219735 , n219733 );
and ( n219737 , n219710 , n219720 );
or ( n219738 , n219736 , n219737 );
not ( n219739 , n217969 );
not ( n219740 , n219524 );
or ( n219741 , n219739 , n219740 );
not ( n219742 , n207938 );
and ( n219743 , n213382 , n219742 );
not ( n219744 , n213382 );
and ( n219745 , n219744 , n207936 );
or ( n219746 , n219743 , n219745 );
nand ( n219747 , n219746 , n211314 );
nand ( n219748 , n219741 , n219747 );
not ( n219749 , n213577 );
not ( n219750 , n219601 );
or ( n219751 , n219749 , n219750 );
not ( n219752 , n213735 );
not ( n219753 , n40766 );
or ( n219754 , n219752 , n219753 );
nand ( n219755 , n219239 , n213732 );
nand ( n219756 , n219754 , n219755 );
nand ( n219757 , n219756 , n216336 );
nand ( n219758 , n219751 , n219757 );
xor ( n219759 , n219748 , n219758 );
not ( n219760 , n37585 );
not ( n219761 , n36319 );
or ( n219762 , n219760 , n219761 );
and ( n219763 , n37545 , n37548 );
nor ( n219764 , n219763 , n37551 );
nand ( n219765 , n219762 , n219764 );
nand ( n219766 , n37544 , n34074 );
not ( n219767 , n219766 );
and ( n219768 , n219765 , n219767 );
not ( n219769 , n219765 );
and ( n219770 , n219769 , n219766 );
nor ( n219771 , n219768 , n219770 );
not ( n219772 , n219771 );
not ( n219773 , n219430 );
or ( n219774 , n219772 , n219773 );
not ( n219775 , n219771 );
nand ( n219776 , n219416 , n219775 );
nand ( n219777 , n219774 , n219776 );
buf ( n219778 , n219777 );
buf ( n219779 , n219778 );
not ( n219780 , n219779 );
nor ( n219781 , n219780 , n213751 );
xor ( n219782 , n219781 , n219339 );
xor ( n219783 , n219782 , n219382 );
xor ( n219784 , n219759 , n219783 );
xor ( n219785 , n219748 , n219758 );
and ( n219786 , n219785 , n219783 );
and ( n219787 , n219748 , n219758 );
or ( n219788 , n219786 , n219787 );
xor ( n219789 , n219650 , n219654 );
not ( n219790 , n219445 );
buf ( n219791 , n219434 );
not ( n219792 , n219791 );
not ( n219793 , n219792 );
or ( n219794 , n219790 , n219793 );
not ( n219795 , n213347 );
not ( n219796 , n219419 );
not ( n219797 , n219796 );
not ( n219798 , n219797 );
or ( n219799 , n219795 , n219798 );
not ( n219800 , n219420 );
nand ( n219801 , n219800 , n214616 );
nand ( n219802 , n219799 , n219801 );
nand ( n219803 , n219802 , n219076 );
nand ( n219804 , n219794 , n219803 );
xor ( n219805 , n219804 , n219634 );
xor ( n219806 , n219805 , n219638 );
xor ( n219807 , n219789 , n219806 );
xor ( n219808 , n219650 , n219654 );
and ( n219809 , n219808 , n219806 );
and ( n219810 , n219650 , n219654 );
or ( n219811 , n219809 , n219810 );
not ( n219812 , n219375 );
not ( n219813 , n218544 );
or ( n219814 , n219812 , n219813 );
not ( n219815 , n218514 );
not ( n219816 , n217602 );
or ( n219817 , n219815 , n219816 );
nand ( n219818 , n216928 , n216170 );
nand ( n219819 , n219817 , n219818 );
nand ( n219820 , n219819 , n217099 );
nand ( n219821 , n219814 , n219820 );
not ( n219822 , n219480 );
not ( n219823 , n217890 );
or ( n219824 , n219822 , n219823 );
not ( n219825 , n216208 );
not ( n219826 , n217473 );
or ( n219827 , n219825 , n219826 );
nand ( n219828 , n217614 , n216207 );
nand ( n219829 , n219827 , n219828 );
nand ( n219830 , n219829 , n218762 );
nand ( n219831 , n219824 , n219830 );
xor ( n219832 , n219821 , n219831 );
and ( n219833 , n219492 , n219503 );
xor ( n219834 , n219832 , n219833 );
not ( n219835 , n219467 );
not ( n219836 , n218220 );
not ( n219837 , n219836 );
or ( n219838 , n219835 , n219837 );
not ( n219839 , n214537 );
not ( n219840 , n218209 );
or ( n219841 , n219839 , n219840 );
nand ( n219842 , n218208 , n214899 );
nand ( n219843 , n219841 , n219842 );
nand ( n219844 , n219843 , n218533 );
nand ( n219845 , n219838 , n219844 );
xor ( n219846 , n219834 , n219845 );
not ( n219847 , n219456 );
not ( n219848 , n219449 );
or ( n219849 , n219847 , n219848 );
not ( n219850 , n214956 );
not ( n219851 , n218814 );
or ( n219852 , n219850 , n219851 );
nand ( n219853 , n219128 , n214960 );
nand ( n219854 , n219852 , n219853 );
nand ( n219855 , n218843 , n219854 );
nand ( n219856 , n219849 , n219855 );
xor ( n219857 , n219846 , n219856 );
not ( n219858 , n215137 );
not ( n219859 , n213960 );
not ( n219860 , n219151 );
or ( n219861 , n219859 , n219860 );
nand ( n219862 , n40724 , n215388 );
nand ( n219863 , n219861 , n219862 );
not ( n219864 , n219863 );
or ( n219865 , n219858 , n219864 );
nand ( n219866 , n219392 , n218467 );
nand ( n219867 , n219865 , n219866 );
xor ( n219868 , n219642 , n219867 );
xor ( n219869 , n219868 , n219646 );
xor ( n219870 , n219857 , n219869 );
xor ( n219871 , n219870 , n219662 );
xor ( n219872 , n219857 , n219869 );
and ( n219873 , n219872 , n219662 );
and ( n219874 , n219857 , n219869 );
or ( n219875 , n219873 , n219874 );
not ( n219876 , n213874 );
not ( n219877 , n219535 );
or ( n219878 , n219876 , n219877 );
not ( n219879 , n214818 );
not ( n219880 , n219226 );
not ( n219881 , n219880 );
or ( n219882 , n219879 , n219881 );
nand ( n219883 , n40559 , n218887 );
nand ( n219884 , n219882 , n219883 );
nand ( n219885 , n219884 , n217142 );
nand ( n219886 , n219878 , n219885 );
not ( n219887 , n216299 );
not ( n219888 , n219572 );
or ( n219889 , n219887 , n219888 );
not ( n219890 , n216810 );
not ( n219891 , n216855 );
or ( n219892 , n219890 , n219891 );
nand ( n219893 , n216859 , n215289 );
nand ( n219894 , n219892 , n219893 );
nand ( n219895 , n219894 , n214694 );
nand ( n219896 , n219889 , n219895 );
not ( n219897 , n219175 );
not ( n219898 , n217017 );
not ( n219899 , n216311 );
not ( n219900 , n219899 );
or ( n219901 , n219898 , n219900 );
not ( n219902 , n216307 );
nand ( n219903 , n219902 , n218661 );
nand ( n219904 , n219901 , n219903 );
not ( n219905 , n219904 );
or ( n219906 , n219897 , n219905 );
nand ( n219907 , n219585 , n217023 );
nand ( n219908 , n219906 , n219907 );
xor ( n219909 , n219896 , n219908 );
xor ( n219910 , n219909 , n219734 );
xor ( n219911 , n219886 , n219910 );
not ( n219912 , n219353 );
not ( n219913 , n217542 );
not ( n219914 , n216261 );
or ( n219915 , n219913 , n219914 );
nand ( n219916 , n208717 , n219358 );
nand ( n219917 , n219915 , n219916 );
not ( n219918 , n219917 );
or ( n219919 , n219912 , n219918 );
nand ( n219920 , n219360 , n217552 );
nand ( n219921 , n219919 , n219920 );
not ( n219922 , n214717 );
not ( n219923 , n219544 );
or ( n219924 , n219922 , n219923 );
not ( n219925 , n218855 );
not ( n219926 , n41070 );
or ( n219927 , n219925 , n219926 );
nand ( n219928 , n41069 , n216037 );
nand ( n219929 , n219927 , n219928 );
nand ( n219930 , n219929 , n216239 );
nand ( n219931 , n219924 , n219930 );
xor ( n219932 , n219921 , n219931 );
xor ( n219933 , n219932 , n219697 );
xor ( n219934 , n219911 , n219933 );
xor ( n219935 , n219658 , n219934 );
xor ( n219936 , n219935 , n219784 );
xor ( n219937 , n219658 , n219934 );
and ( n219938 , n219937 , n219784 );
and ( n219939 , n219658 , n219934 );
or ( n219940 , n219938 , n219939 );
xor ( n219941 , n219403 , n219807 );
xor ( n219942 , n219941 , n219513 );
xor ( n219943 , n219403 , n219807 );
and ( n219944 , n219943 , n219513 );
and ( n219945 , n219403 , n219807 );
or ( n219946 , n219944 , n219945 );
xor ( n219947 , n219871 , n219564 );
xor ( n219948 , n219947 , n219936 );
xor ( n219949 , n219871 , n219564 );
and ( n219950 , n219949 , n219936 );
and ( n219951 , n219871 , n219564 );
or ( n219952 , n219950 , n219951 );
xor ( n219953 , n219612 , n219618 );
xor ( n219954 , n219953 , n219942 );
xor ( n219955 , n219612 , n219618 );
and ( n219956 , n219955 , n219942 );
and ( n219957 , n219612 , n219618 );
or ( n219958 , n219956 , n219957 );
xor ( n219959 , n219948 , n219624 );
xor ( n219960 , n219959 , n219954 );
xor ( n219961 , n219948 , n219624 );
and ( n219962 , n219961 , n219954 );
and ( n219963 , n219948 , n219624 );
or ( n219964 , n219962 , n219963 );
xor ( n219965 , n219821 , n219831 );
and ( n219966 , n219965 , n219833 );
and ( n219967 , n219821 , n219831 );
or ( n219968 , n219966 , n219967 );
xor ( n219969 , n219921 , n219931 );
and ( n219970 , n219969 , n219697 );
and ( n219971 , n219921 , n219931 );
or ( n219972 , n219970 , n219971 );
xor ( n219973 , n219781 , n219339 );
and ( n219974 , n219973 , n219382 );
and ( n219975 , n219781 , n219339 );
or ( n219976 , n219974 , n219975 );
xor ( n219977 , n219896 , n219908 );
and ( n219978 , n219977 , n219734 );
and ( n219979 , n219896 , n219908 );
or ( n219980 , n219978 , n219979 );
xor ( n219981 , n219834 , n219845 );
and ( n219982 , n219981 , n219856 );
and ( n219983 , n219834 , n219845 );
or ( n219984 , n219982 , n219983 );
xor ( n219985 , n219804 , n219634 );
and ( n219986 , n219985 , n219638 );
and ( n219987 , n219804 , n219634 );
or ( n219988 , n219986 , n219987 );
xor ( n219989 , n219642 , n219867 );
and ( n219990 , n219989 , n219646 );
and ( n219991 , n219642 , n219867 );
or ( n219992 , n219990 , n219991 );
xor ( n219993 , n219886 , n219910 );
and ( n219994 , n219993 , n219933 );
and ( n219995 , n219886 , n219910 );
or ( n219996 , n219994 , n219995 );
not ( n219997 , n215183 );
not ( n219998 , n219708 );
or ( n219999 , n219997 , n219998 );
or ( n220000 , n30962 , n215105 );
nand ( n220001 , n30962 , n215545 );
nand ( n220002 , n220000 , n220001 );
nand ( n220003 , n220002 , n215191 );
nand ( n220004 , n219999 , n220003 );
not ( n220005 , n214449 );
not ( n220006 , n219728 );
or ( n220007 , n220005 , n220006 );
not ( n220008 , n219033 );
not ( n220009 , n41563 );
or ( n220010 , n220008 , n220009 );
nand ( n220011 , n216089 , n216167 );
nand ( n220012 , n220010 , n220011 );
nand ( n220013 , n220012 , n214458 );
nand ( n220014 , n220007 , n220013 );
xor ( n220015 , n220004 , n220014 );
not ( n220016 , n219718 );
not ( n220017 , n216065 );
or ( n220018 , n220016 , n220017 );
not ( n220019 , n215533 );
not ( n220020 , n216402 );
or ( n220021 , n220019 , n220020 );
not ( n220022 , n215533 );
nand ( n220023 , n216403 , n220022 );
nand ( n220024 , n220021 , n220023 );
nand ( n220025 , n216332 , n220024 );
nand ( n220026 , n220018 , n220025 );
xor ( n220027 , n220015 , n220026 );
xor ( n220028 , n220004 , n220014 );
and ( n220029 , n220028 , n220026 );
and ( n220030 , n220004 , n220014 );
or ( n220031 , n220029 , n220030 );
buf ( n220032 , n215761 );
not ( n220033 , n220032 );
not ( n220034 , n220033 );
not ( n220035 , n216281 );
not ( n220036 , n214820 );
or ( n220037 , n220035 , n220036 );
buf ( n220038 , n216277 );
nand ( n220039 , n215228 , n220038 );
nand ( n220040 , n220037 , n220039 );
not ( n220041 , n220040 );
or ( n220042 , n220034 , n220041 );
nand ( n220043 , n219668 , n217486 );
nand ( n220044 , n220042 , n220043 );
not ( n220045 , n219819 );
buf ( n220046 , n217089 );
not ( n220047 , n220046 );
or ( n220048 , n220045 , n220047 );
not ( n220049 , n216934 );
not ( n220050 , n216928 );
not ( n220051 , n220050 );
or ( n220052 , n220049 , n220051 );
nand ( n220053 , n216929 , n216940 );
nand ( n220054 , n220052 , n220053 );
nand ( n220055 , n220054 , n217388 );
nand ( n220056 , n220048 , n220055 );
xor ( n220057 , n220044 , n220056 );
not ( n220058 , n219829 );
not ( n220059 , n217630 );
not ( n220060 , n220059 );
or ( n220061 , n220058 , n220060 );
not ( n220062 , n215075 );
not ( n220063 , n218253 );
or ( n220064 , n220062 , n220063 );
nand ( n220065 , n218560 , n215899 );
nand ( n220066 , n220064 , n220065 );
buf ( n220067 , n217230 );
nand ( n220068 , n220066 , n220067 );
nand ( n220069 , n220061 , n220068 );
xor ( n220070 , n220057 , n220069 );
xor ( n220071 , n220044 , n220056 );
and ( n220072 , n220071 , n220069 );
and ( n220073 , n220044 , n220056 );
or ( n220074 , n220072 , n220073 );
not ( n220075 , n216239 );
not ( n220076 , n215113 );
not ( n220077 , n41164 );
not ( n220078 , n220077 );
or ( n220079 , n220076 , n220078 );
nand ( n220080 , n41165 , n217944 );
nand ( n220081 , n220079 , n220080 );
not ( n220082 , n220081 );
or ( n220083 , n220075 , n220082 );
nand ( n220084 , n219929 , n214717 );
nand ( n220085 , n220083 , n220084 );
xor ( n220086 , n219968 , n220085 );
not ( n220087 , n219843 );
not ( n220088 , n219836 );
or ( n220089 , n220087 , n220088 );
not ( n220090 , n216964 );
not ( n220091 , n218775 );
not ( n220092 , n220091 );
or ( n220093 , n220090 , n220092 );
not ( n220094 , n219475 );
nand ( n220095 , n220094 , n218208 );
nand ( n220096 , n220093 , n220095 );
nand ( n220097 , n220096 , n218231 );
nand ( n220098 , n220089 , n220097 );
xor ( n220099 , n220086 , n220098 );
not ( n220100 , n217023 );
not ( n220101 , n219904 );
or ( n220102 , n220100 , n220101 );
not ( n220103 , n219577 );
not ( n220104 , n217147 );
or ( n220105 , n220103 , n220104 );
not ( n220106 , n216519 );
not ( n220107 , n220106 );
nand ( n220108 , n220107 , n215971 );
nand ( n220109 , n220105 , n220108 );
nand ( n220110 , n220109 , n219175 );
nand ( n220111 , n220102 , n220110 );
xor ( n220112 , n220111 , n220027 );
xor ( n220113 , n220112 , n220070 );
xor ( n220114 , n220099 , n220113 );
xor ( n220115 , n220114 , n219984 );
xor ( n220116 , n220099 , n220113 );
and ( n220117 , n220116 , n219984 );
and ( n220118 , n220099 , n220113 );
or ( n220119 , n220117 , n220118 );
not ( n220120 , n219854 );
not ( n220121 , n218835 );
or ( n220122 , n220120 , n220121 );
not ( n220123 , n217044 );
not ( n220124 , n218876 );
or ( n220125 , n220123 , n220124 );
not ( n220126 , n218876 );
nand ( n220127 , n220126 , n215131 );
nand ( n220128 , n220125 , n220127 );
nand ( n220129 , n220128 , n218843 );
nand ( n220130 , n220122 , n220129 );
nor ( n220131 , n37546 , n37584 );
not ( n220132 , n220131 );
not ( n220133 , n36319 );
or ( n220134 , n220132 , n220133 );
nand ( n220135 , n220134 , n37555 );
not ( n220136 , n34056 );
not ( n220137 , n34061 );
or ( n220138 , n220136 , n220137 );
nand ( n220139 , n220138 , n34078 );
and ( n220140 , n220135 , n220139 );
not ( n220141 , n220135 );
not ( n220142 , n220139 );
and ( n220143 , n220141 , n220142 );
nor ( n220144 , n220140 , n220143 );
not ( n220145 , n220144 );
buf ( n220146 , n220145 );
not ( n220147 , n220146 );
and ( n220148 , n213751 , n220147 );
not ( n220149 , n213751 );
not ( n220150 , n220147 );
buf ( n220151 , n220150 );
and ( n220152 , n220149 , n220151 );
nor ( n220153 , n220148 , n220152 );
not ( n220154 , n220153 );
not ( n220155 , n220145 );
nand ( n220156 , n220155 , n219775 );
nand ( n220157 , n220145 , n219771 );
nand ( n220158 , n220156 , n220157 );
not ( n220159 , n220158 );
xor ( n220160 , n219416 , n219775 );
nand ( n220161 , n220159 , n220160 );
not ( n220162 , n220161 );
buf ( n220163 , n220162 );
buf ( n220164 , n220163 );
not ( n220165 , n220164 );
or ( n220166 , n220154 , n220165 );
and ( n220167 , n220151 , n216076 );
not ( n220168 , n220151 );
and ( n220169 , n220168 , n218224 );
or ( n220170 , n220167 , n220169 );
nand ( n220171 , n220170 , n219779 );
nand ( n220172 , n220166 , n220171 );
xor ( n220173 , n220130 , n220172 );
not ( n220174 , n219802 );
not ( n220175 , n219792 );
or ( n220176 , n220174 , n220175 );
not ( n220177 , n213583 );
not ( n220178 , n219440 );
or ( n220179 , n220177 , n220178 );
not ( n220180 , n219439 );
not ( n220181 , n220180 );
or ( n220182 , n220181 , n213583 );
nand ( n220183 , n220179 , n220182 );
nand ( n220184 , n220183 , n219076 );
nand ( n220185 , n220176 , n220184 );
xor ( n220186 , n220173 , n220185 );
xor ( n220187 , n219988 , n220186 );
xor ( n220188 , n220187 , n219992 );
xor ( n220189 , n219988 , n220186 );
and ( n220190 , n220189 , n219992 );
and ( n220191 , n219988 , n220186 );
or ( n220192 , n220190 , n220191 );
xor ( n220193 , n219972 , n219976 );
xor ( n220194 , n220193 , n219980 );
xor ( n220195 , n219996 , n220194 );
xor ( n220196 , n220195 , n219788 );
xor ( n220197 , n219996 , n220194 );
and ( n220198 , n220197 , n219788 );
and ( n220199 , n219996 , n220194 );
or ( n220200 , n220198 , n220199 );
not ( n220201 , n213498 );
not ( n220202 , n213735 );
buf ( n220203 , n208078 );
not ( n220204 , n220203 );
not ( n220205 , n220204 );
or ( n220206 , n220202 , n220205 );
nand ( n220207 , n220203 , n213732 );
nand ( n220208 , n220206 , n220207 );
not ( n220209 , n220208 );
or ( n220210 , n220201 , n220209 );
nand ( n220211 , n219756 , n213577 );
nand ( n220212 , n220210 , n220211 );
not ( n220213 , n217969 );
not ( n220214 , n219746 );
or ( n220215 , n220213 , n220214 );
not ( n220216 , n40668 );
not ( n220217 , n220216 );
not ( n220218 , n220217 );
nand ( n220219 , n220218 , n213381 );
not ( n220220 , n220216 );
nand ( n220221 , n220220 , n213382 );
nand ( n220222 , n220219 , n220221 , n211314 );
nand ( n220223 , n220215 , n220222 );
xor ( n220224 , n220212 , n220223 );
not ( n220225 , n214694 );
not ( n220226 , n217115 );
not ( n220227 , n220226 );
not ( n220228 , n220227 );
not ( n220229 , n216810 );
or ( n220230 , n220228 , n220229 );
or ( n220231 , n220227 , n216810 );
nand ( n220232 , n220230 , n220231 );
not ( n220233 , n220232 );
or ( n220234 , n220225 , n220233 );
nand ( n220235 , n219894 , n216562 );
nand ( n220236 , n220234 , n220235 );
xor ( n220237 , n220236 , n219701 );
xor ( n220238 , n220237 , n219738 );
xor ( n220239 , n220224 , n220238 );
not ( n220240 , n215383 );
not ( n220241 , n217573 );
not ( n220242 , n218268 );
or ( n220243 , n220241 , n220242 );
nand ( n220244 , n40710 , n217397 );
nand ( n220245 , n220243 , n220244 );
not ( n220246 , n220245 );
or ( n220247 , n220240 , n220246 );
nand ( n220248 , n219863 , n215605 );
nand ( n220249 , n220247 , n220248 );
not ( n220250 , n219680 );
not ( n220251 , n218647 );
or ( n220252 , n220250 , n220251 );
not ( n220253 , n219343 );
not ( n220254 , n216593 );
or ( n220255 , n220253 , n220254 );
nand ( n220256 , n216762 , n219348 );
nand ( n220257 , n220255 , n220256 );
nand ( n220258 , n219501 , n220257 );
nand ( n220259 , n220252 , n220258 );
not ( n220260 , n219314 );
not ( n220261 , n219687 );
not ( n220262 , n217066 );
or ( n220263 , n220261 , n220262 );
not ( n220264 , n219305 );
nand ( n220265 , n220264 , n216938 );
nand ( n220266 , n220263 , n220265 );
not ( n220267 , n220266 );
or ( n220268 , n220260 , n220267 );
nand ( n220269 , n219694 , n216204 );
nand ( n220270 , n220268 , n220269 );
xor ( n220271 , n220259 , n220270 );
not ( n220272 , n217549 );
not ( n220273 , n220272 );
and ( n220274 , n217130 , n215955 );
not ( n220275 , n217130 );
and ( n220276 , n220275 , n219358 );
or ( n220277 , n220274 , n220276 );
not ( n220278 , n220277 );
or ( n220279 , n220273 , n220278 );
not ( n220280 , n217551 );
nand ( n220281 , n219917 , n220280 );
nand ( n220282 , n220279 , n220281 );
xor ( n220283 , n220271 , n220282 );
not ( n220284 , n213750 );
not ( n220285 , n219771 );
or ( n220286 , n220284 , n220285 );
nand ( n220287 , n220286 , n220181 );
nand ( n220288 , n219775 , n213751 );
and ( n220289 , n220287 , n220288 );
not ( n220290 , n220151 );
nor ( n220291 , n220289 , n220290 );
xor ( n220292 , n220283 , n220291 );
xor ( n220293 , n220249 , n220292 );
not ( n220294 , n213874 );
not ( n220295 , n219884 );
or ( n220296 , n220294 , n220295 );
not ( n220297 , n214818 );
not ( n220298 , n219518 );
or ( n220299 , n220297 , n220298 );
not ( n220300 , n214818 );
nand ( n220301 , n219522 , n220300 );
nand ( n220302 , n220299 , n220301 );
not ( n220303 , n220302 );
or ( n220304 , n220303 , n218150 );
nand ( n220305 , n220296 , n220304 );
xor ( n220306 , n220293 , n220305 );
xor ( n220307 , n220239 , n220306 );
xor ( n220308 , n220307 , n219811 );
xor ( n220309 , n220239 , n220306 );
and ( n220310 , n220309 , n219811 );
and ( n220311 , n220239 , n220306 );
or ( n220312 , n220310 , n220311 );
xor ( n220313 , n220115 , n220188 );
xor ( n220314 , n220313 , n219875 );
xor ( n220315 , n220115 , n220188 );
and ( n220316 , n220315 , n219875 );
and ( n220317 , n220115 , n220188 );
or ( n220318 , n220316 , n220317 );
xor ( n220319 , n219940 , n220196 );
xor ( n220320 , n220319 , n220308 );
xor ( n220321 , n219940 , n220196 );
and ( n220322 , n220321 , n220308 );
and ( n220323 , n219940 , n220196 );
or ( n220324 , n220322 , n220323 );
xor ( n220325 , n219946 , n220314 );
xor ( n220326 , n220325 , n219952 );
xor ( n220327 , n219946 , n220314 );
and ( n220328 , n220327 , n219952 );
and ( n220329 , n219946 , n220314 );
or ( n220330 , n220328 , n220329 );
xor ( n220331 , n220320 , n219958 );
xor ( n220332 , n220331 , n220326 );
xor ( n220333 , n220320 , n219958 );
and ( n220334 , n220333 , n220326 );
and ( n220335 , n220320 , n219958 );
or ( n220336 , n220334 , n220335 );
xor ( n220337 , n220271 , n220282 );
and ( n220338 , n220337 , n220291 );
and ( n220339 , n220271 , n220282 );
or ( n220340 , n220338 , n220339 );
xor ( n220341 , n220236 , n219701 );
and ( n220342 , n220341 , n219738 );
and ( n220343 , n220236 , n219701 );
or ( n220344 , n220342 , n220343 );
xor ( n220345 , n220111 , n220027 );
and ( n220346 , n220345 , n220070 );
and ( n220347 , n220111 , n220027 );
or ( n220348 , n220346 , n220347 );
xor ( n220349 , n219968 , n220085 );
and ( n220350 , n220349 , n220098 );
and ( n220351 , n219968 , n220085 );
or ( n220352 , n220350 , n220351 );
xor ( n220353 , n220130 , n220172 );
and ( n220354 , n220353 , n220185 );
and ( n220355 , n220130 , n220172 );
or ( n220356 , n220354 , n220355 );
xor ( n220357 , n219972 , n219976 );
and ( n220358 , n220357 , n219980 );
and ( n220359 , n219972 , n219976 );
or ( n220360 , n220358 , n220359 );
xor ( n220361 , n220249 , n220292 );
and ( n220362 , n220361 , n220305 );
and ( n220363 , n220249 , n220292 );
or ( n220364 , n220362 , n220363 );
xor ( n220365 , n220212 , n220223 );
and ( n220366 , n220365 , n220238 );
and ( n220367 , n220212 , n220223 );
or ( n220368 , n220366 , n220367 );
not ( n220369 , n220257 );
not ( n220370 , n216586 );
or ( n220371 , n220369 , n220370 );
not ( n220372 , n218981 );
not ( n220373 , n216569 );
or ( n220374 , n220372 , n220373 );
nand ( n220375 , n216421 , n218980 );
nand ( n220376 , n220374 , n220375 );
nand ( n220377 , n220376 , n219501 );
nand ( n220378 , n220371 , n220377 );
not ( n220379 , n215550 );
not ( n220380 , n215165 );
not ( n220381 , n218503 );
or ( n220382 , n220380 , n220381 );
nand ( n220383 , n219326 , n208725 );
nand ( n220384 , n220382 , n220383 );
not ( n220385 , n220384 );
or ( n220386 , n220379 , n220385 );
nand ( n220387 , n220002 , n215183 );
nand ( n220388 , n220386 , n220387 );
xor ( n220389 , n220378 , n220388 );
not ( n220390 , n219314 );
not ( n220391 , n219687 );
not ( n220392 , n215428 );
or ( n220393 , n220391 , n220392 );
nand ( n220394 , n41701 , n219092 );
nand ( n220395 , n220393 , n220394 );
not ( n220396 , n220395 );
or ( n220397 , n220390 , n220396 );
nand ( n220398 , n220266 , n216426 );
nand ( n220399 , n220397 , n220398 );
xor ( n220400 , n220389 , n220399 );
xor ( n220401 , n220378 , n220388 );
and ( n220402 , n220401 , n220399 );
and ( n220403 , n220378 , n220388 );
or ( n220404 , n220402 , n220403 );
not ( n220405 , n220024 );
or ( n220406 , n216066 , n220405 );
and ( n220407 , n216068 , n214628 );
not ( n220408 , n216068 );
and ( n220409 , n220408 , n30997 );
or ( n220410 , n220407 , n220409 );
not ( n220411 , n220410 );
or ( n220412 , n220411 , n216795 );
nand ( n220413 , n220406 , n220412 );
not ( n220414 , n216730 );
not ( n220415 , n220414 );
not ( n220416 , n220040 );
or ( n220417 , n220415 , n220416 );
not ( n220418 , n215766 );
not ( n220419 , n215833 );
or ( n220420 , n220418 , n220419 );
not ( n220421 , n831 );
not ( n220422 , n186143 );
or ( n220423 , n220421 , n220422 );
nand ( n220424 , n220423 , n32112 );
nand ( n220425 , n220424 , n216277 );
nand ( n220426 , n220420 , n220425 );
nand ( n220427 , n220426 , n220033 );
nand ( n220428 , n220417 , n220427 );
xor ( n220429 , n220413 , n220428 );
not ( n220430 , n220054 );
not ( n220431 , n219368 );
or ( n220432 , n220430 , n220431 );
not ( n220433 , n219102 );
not ( n220434 , n220050 );
or ( n220435 , n220433 , n220434 );
not ( n220436 , n219102 );
nand ( n220437 , n216929 , n220436 );
nand ( n220438 , n220435 , n220437 );
nand ( n220439 , n220438 , n217388 );
nand ( n220440 , n220432 , n220439 );
xor ( n220441 , n220429 , n220440 );
xor ( n220442 , n220413 , n220428 );
and ( n220443 , n220442 , n220440 );
and ( n220444 , n220413 , n220428 );
or ( n220445 , n220443 , n220444 );
not ( n220446 , n217023 );
not ( n220447 , n220109 );
or ( n220448 , n220446 , n220447 );
not ( n220449 , n217017 );
not ( n220450 , n217317 );
or ( n220451 , n220449 , n220450 );
nand ( n220452 , n216859 , n219583 );
nand ( n220453 , n220451 , n220452 );
nand ( n220454 , n220453 , n219175 );
nand ( n220455 , n220448 , n220454 );
xor ( n220456 , n220031 , n220455 );
xor ( n220457 , n220456 , n220400 );
xor ( n220458 , n220348 , n220457 );
xor ( n220459 , n220441 , n220074 );
not ( n220460 , n220096 );
not ( n220461 , n219836 );
or ( n220462 , n220460 , n220461 );
not ( n220463 , n216208 );
not ( n220464 , n220091 );
or ( n220465 , n220463 , n220464 );
not ( n220466 , n218226 );
nand ( n220467 , n220466 , n216207 );
nand ( n220468 , n220465 , n220467 );
nand ( n220469 , n220468 , n218533 );
nand ( n220470 , n220462 , n220469 );
xor ( n220471 , n220459 , n220470 );
xor ( n220472 , n220458 , n220471 );
xor ( n220473 , n220348 , n220457 );
and ( n220474 , n220473 , n220471 );
and ( n220475 , n220348 , n220457 );
or ( n220476 , n220474 , n220475 );
xor ( n220477 , n220356 , n220352 );
not ( n220478 , n220128 );
not ( n220479 , n218834 );
buf ( n220480 , n220479 );
not ( n220481 , n220480 );
or ( n220482 , n220478 , n220481 );
not ( n220483 , n214537 );
not ( n220484 , n218876 );
or ( n220485 , n220483 , n220484 );
not ( n220486 , n214537 );
nand ( n220487 , n220486 , n218815 );
nand ( n220488 , n220485 , n220487 );
nand ( n220489 , n220488 , n218843 );
nand ( n220490 , n220482 , n220489 );
not ( n220491 , n220170 );
buf ( n220492 , n220163 );
not ( n220493 , n220492 );
or ( n220494 , n220491 , n220493 );
not ( n220495 , n213347 );
not ( n220496 , n220151 );
not ( n220497 , n220496 );
or ( n220498 , n220495 , n220497 );
buf ( n220499 , n220147 );
not ( n220500 , n220499 );
nand ( n220501 , n220500 , n214616 );
nand ( n220502 , n220498 , n220501 );
nand ( n220503 , n220502 , n219779 );
nand ( n220504 , n220494 , n220503 );
xor ( n220505 , n220490 , n220504 );
not ( n220506 , n220183 );
not ( n220507 , n219791 );
not ( n220508 , n220507 );
or ( n220509 , n220506 , n220508 );
not ( n220510 , n214956 );
not ( n220511 , n219797 );
or ( n220512 , n220510 , n220511 );
nand ( n220513 , n219800 , n214960 );
nand ( n220514 , n220512 , n220513 );
nand ( n220515 , n220514 , n219076 );
nand ( n220516 , n220509 , n220515 );
xor ( n220517 , n220505 , n220516 );
xor ( n220518 , n220477 , n220517 );
xor ( n220519 , n220356 , n220352 );
and ( n220520 , n220519 , n220517 );
and ( n220521 , n220356 , n220352 );
or ( n220522 , n220520 , n220521 );
xor ( n220523 , n220364 , n220368 );
not ( n220524 , n220066 );
not ( n220525 , n217890 );
or ( n220526 , n220524 , n220525 );
not ( n220527 , n218514 );
not ( n220528 , n217637 );
or ( n220529 , n220527 , n220528 );
nand ( n220530 , n217614 , n216170 );
nand ( n220531 , n220529 , n220530 );
nand ( n220532 , n220531 , n220067 );
nand ( n220533 , n220526 , n220532 );
not ( n220534 , n214458 );
not ( n220535 , n216166 );
not ( n220536 , n216261 );
or ( n220537 , n220535 , n220536 );
not ( n220538 , n214416 );
nand ( n220539 , n208717 , n220538 );
nand ( n220540 , n220537 , n220539 );
not ( n220541 , n220540 );
or ( n220542 , n220534 , n220541 );
nand ( n220543 , n220012 , n219731 );
nand ( n220544 , n220542 , n220543 );
xor ( n220545 , n220533 , n220544 );
and ( n220546 , n220259 , n220270 );
xor ( n220547 , n220545 , n220546 );
xor ( n220548 , n220547 , n220340 );
xor ( n220549 , n220548 , n220344 );
xor ( n220550 , n220523 , n220549 );
xor ( n220551 , n220364 , n220368 );
and ( n220552 , n220551 , n220549 );
and ( n220553 , n220364 , n220368 );
or ( n220554 , n220552 , n220553 );
xor ( n220555 , n220360 , n220472 );
not ( n220556 , n216239 );
not ( n220557 , n217944 );
not ( n220558 , n40724 );
or ( n220559 , n220557 , n220558 );
nand ( n220560 , n217964 , n215113 );
nand ( n220561 , n220559 , n220560 );
not ( n220562 , n220561 );
or ( n220563 , n220556 , n220562 );
nand ( n220564 , n220081 , n214717 );
nand ( n220565 , n220563 , n220564 );
not ( n220566 , n215137 );
not ( n220567 , n217573 );
not ( n220568 , n219238 );
not ( n220569 , n220568 );
not ( n220570 , n220569 );
or ( n220571 , n220567 , n220570 );
nand ( n220572 , n208044 , n215388 );
nand ( n220573 , n220571 , n220572 );
not ( n220574 , n220573 );
or ( n220575 , n220566 , n220574 );
nand ( n220576 , n220245 , n214086 );
nand ( n220577 , n220575 , n220576 );
xor ( n220578 , n220565 , n220577 );
not ( n220579 , n217142 );
not ( n220580 , n216262 );
not ( n220581 , n207936 );
not ( n220582 , n220581 );
or ( n220583 , n220580 , n220582 );
nand ( n220584 , n207938 , n220300 );
nand ( n220585 , n220583 , n220584 );
not ( n220586 , n220585 );
or ( n220587 , n220579 , n220586 );
nand ( n220588 , n220302 , n213874 );
nand ( n220589 , n220587 , n220588 );
xor ( n220590 , n220578 , n220589 );
xor ( n220591 , n220555 , n220590 );
xor ( n220592 , n220360 , n220472 );
and ( n220593 , n220592 , n220590 );
and ( n220594 , n220360 , n220472 );
or ( n220595 , n220593 , n220594 );
not ( n220596 , n40410 );
and ( n220597 , n213382 , n220596 );
not ( n220598 , n213382 );
not ( n220599 , n40409 );
not ( n220600 , n220599 );
and ( n220601 , n220598 , n220600 );
nor ( n220602 , n220597 , n220601 );
or ( n220603 , n220602 , n213171 );
nand ( n220604 , n220219 , n220221 , n217969 );
nand ( n220605 , n220603 , n220604 );
not ( n220606 , n219353 );
not ( n220607 , n215955 );
not ( n220608 , n219899 );
or ( n220609 , n220607 , n220608 );
nand ( n220610 , n216306 , n219358 );
nand ( n220611 , n220609 , n220610 );
not ( n220612 , n220611 );
or ( n220613 , n220606 , n220612 );
nand ( n220614 , n220277 , n217552 );
nand ( n220615 , n220613 , n220614 );
not ( n220616 , n36650 );
not ( n220617 , n36998 );
or ( n220618 , n220616 , n220617 );
nor ( n220619 , n36645 , n36316 );
nand ( n220620 , n220618 , n220619 );
not ( n220621 , n220620 );
buf ( n220622 , n35319 );
buf ( n220623 , n36316 );
nor ( n220624 , n220622 , n220623 );
nor ( n220625 , n220624 , n34124 );
not ( n220626 , n220625 );
or ( n220627 , n220621 , n220626 );
nand ( n220628 , n220627 , n37535 );
not ( n220629 , n37609 );
and ( n220630 , n220628 , n220629 );
not ( n220631 , n220628 );
and ( n220632 , n220631 , n37609 );
nor ( n220633 , n220630 , n220632 );
xnor ( n220634 , n220633 , n220145 );
not ( n220635 , n220634 );
buf ( n220636 , n220635 );
not ( n220637 , n220636 );
nor ( n220638 , n220637 , n213751 );
xor ( n220639 , n220615 , n220638 );
not ( n220640 , n216299 );
not ( n220641 , n220232 );
or ( n220642 , n220640 , n220641 );
not ( n220643 , n215290 );
not ( n220644 , n217977 );
or ( n220645 , n220643 , n220644 );
nand ( n220646 , n219201 , n215289 );
nand ( n220647 , n220645 , n220646 );
nand ( n220648 , n220647 , n214694 );
nand ( n220649 , n220642 , n220648 );
xor ( n220650 , n220639 , n220649 );
xor ( n220651 , n220605 , n220650 );
not ( n220652 , n220208 );
not ( n220653 , n213577 );
or ( n220654 , n220652 , n220653 );
and ( n220655 , n213735 , n40561 );
not ( n220656 , n213735 );
not ( n220657 , n219223 );
and ( n220658 , n220656 , n220657 );
or ( n220659 , n220655 , n220658 );
not ( n220660 , n220659 );
or ( n220661 , n220660 , n216335 );
nand ( n220662 , n220654 , n220661 );
xor ( n220663 , n220651 , n220662 );
xor ( n220664 , n220663 , n220119 );
xor ( n220665 , n220664 , n220518 );
xor ( n220666 , n220663 , n220119 );
and ( n220667 , n220666 , n220518 );
and ( n220668 , n220663 , n220119 );
or ( n220669 , n220667 , n220668 );
xor ( n220670 , n220192 , n220200 );
xor ( n220671 , n220670 , n220550 );
xor ( n220672 , n220192 , n220200 );
and ( n220673 , n220672 , n220550 );
and ( n220674 , n220192 , n220200 );
or ( n220675 , n220673 , n220674 );
xor ( n220676 , n220312 , n220665 );
xor ( n220677 , n220676 , n220591 );
xor ( n220678 , n220312 , n220665 );
and ( n220679 , n220678 , n220591 );
and ( n220680 , n220312 , n220665 );
or ( n220681 , n220679 , n220680 );
xor ( n220682 , n220318 , n220671 );
xor ( n220683 , n220682 , n220324 );
xor ( n220684 , n220318 , n220671 );
and ( n220685 , n220684 , n220324 );
and ( n220686 , n220318 , n220671 );
or ( n220687 , n220685 , n220686 );
xor ( n220688 , n220677 , n220683 );
xor ( n220689 , n220688 , n220330 );
xor ( n220690 , n220677 , n220683 );
and ( n220691 , n220690 , n220330 );
and ( n220692 , n220677 , n220683 );
or ( n220693 , n220691 , n220692 );
xor ( n220694 , n220533 , n220544 );
and ( n220695 , n220694 , n220546 );
and ( n220696 , n220533 , n220544 );
or ( n220697 , n220695 , n220696 );
xor ( n220698 , n220615 , n220638 );
and ( n220699 , n220698 , n220649 );
and ( n220700 , n220615 , n220638 );
or ( n220701 , n220699 , n220700 );
xor ( n220702 , n220031 , n220455 );
and ( n220703 , n220702 , n220400 );
and ( n220704 , n220031 , n220455 );
or ( n220705 , n220703 , n220704 );
xor ( n220706 , n220441 , n220074 );
and ( n220707 , n220706 , n220470 );
and ( n220708 , n220441 , n220074 );
or ( n220709 , n220707 , n220708 );
xor ( n220710 , n220490 , n220504 );
and ( n220711 , n220710 , n220516 );
and ( n220712 , n220490 , n220504 );
or ( n220713 , n220711 , n220712 );
xor ( n220714 , n220547 , n220340 );
and ( n220715 , n220714 , n220344 );
and ( n220716 , n220547 , n220340 );
or ( n220717 , n220715 , n220716 );
xor ( n220718 , n220565 , n220577 );
and ( n220719 , n220718 , n220589 );
and ( n220720 , n220565 , n220577 );
or ( n220721 , n220719 , n220720 );
xor ( n220722 , n220605 , n220650 );
and ( n220723 , n220722 , n220662 );
and ( n220724 , n220605 , n220650 );
or ( n220725 , n220723 , n220724 );
not ( n220726 , n216426 );
not ( n220727 , n220395 );
or ( n220728 , n220726 , n220727 );
not ( n220729 , n219687 );
not ( n220730 , n41563 );
or ( n220731 , n220729 , n220730 );
nand ( n220732 , n41564 , n216938 );
nand ( n220733 , n220731 , n220732 );
nand ( n220734 , n220733 , n214808 );
nand ( n220735 , n220728 , n220734 );
not ( n220736 , n217047 );
not ( n220737 , n216327 );
not ( n220738 , n216555 );
or ( n220739 , n220737 , n220738 );
not ( n220740 , n214821 );
nand ( n220741 , n220740 , n216014 );
nand ( n220742 , n220739 , n220741 );
not ( n220743 , n220742 );
or ( n220744 , n220736 , n220743 );
nand ( n220745 , n217864 , n220410 );
nand ( n220746 , n220744 , n220745 );
xor ( n220747 , n220735 , n220746 );
not ( n220748 , n220033 );
buf ( n220749 , n215572 );
not ( n220750 , n220749 );
not ( n220751 , n218670 );
or ( n220752 , n220750 , n220751 );
not ( n220753 , n220749 );
nand ( n220754 , n214837 , n220753 );
nand ( n220755 , n220752 , n220754 );
not ( n220756 , n220755 );
or ( n220757 , n220748 , n220756 );
nand ( n220758 , n220426 , n217486 );
nand ( n220759 , n220757 , n220758 );
xor ( n220760 , n220747 , n220759 );
xor ( n220761 , n220735 , n220746 );
and ( n220762 , n220761 , n220759 );
and ( n220763 , n220735 , n220746 );
or ( n220764 , n220762 , n220763 );
not ( n220765 , n220438 );
not ( n220766 , n220046 );
or ( n220767 , n220765 , n220766 );
not ( n220768 , n219343 );
not ( n220769 , n217602 );
or ( n220770 , n220768 , n220769 );
not ( n220771 , n217093 );
nand ( n220772 , n220771 , n219348 );
nand ( n220773 , n220770 , n220772 );
nand ( n220774 , n220773 , n217388 );
nand ( n220775 , n220767 , n220774 );
not ( n220776 , n220531 );
not ( n220777 , n217631 );
or ( n220778 , n220776 , n220777 );
not ( n220779 , n216934 );
not ( n220780 , n217611 );
or ( n220781 , n220779 , n220780 );
nand ( n220782 , n218560 , n216940 );
nand ( n220783 , n220781 , n220782 );
nand ( n220784 , n220783 , n218762 );
nand ( n220785 , n220778 , n220784 );
xor ( n220786 , n220775 , n220785 );
not ( n220787 , n215550 );
not ( n220788 , n215165 );
not ( n220789 , n219305 );
or ( n220790 , n220788 , n220789 );
nand ( n220791 , n41609 , n219326 );
nand ( n220792 , n220790 , n220791 );
not ( n220793 , n220792 );
or ( n220794 , n220787 , n220793 );
nand ( n220795 , n220384 , n219332 );
nand ( n220796 , n220794 , n220795 );
not ( n220797 , n220376 );
not ( n220798 , n217505 );
or ( n220799 , n220797 , n220798 );
not ( n220800 , n216200 );
not ( n220801 , n215533 );
not ( n220802 , n216572 );
not ( n220803 , n220802 );
or ( n220804 , n220801 , n220803 );
nand ( n220805 , n216762 , n214190 );
nand ( n220806 , n220804 , n220805 );
nand ( n220807 , n220800 , n220806 );
nand ( n220808 , n220799 , n220807 );
and ( n220809 , n220796 , n220808 );
not ( n220810 , n220796 );
not ( n220811 , n220808 );
and ( n220812 , n220810 , n220811 );
nor ( n220813 , n220809 , n220812 );
xor ( n220814 , n220786 , n220813 );
xor ( n220815 , n220775 , n220785 );
and ( n220816 , n220815 , n220813 );
and ( n220817 , n220775 , n220785 );
or ( n220818 , n220816 , n220817 );
not ( n220819 , n214694 );
not ( n220820 , n220819 );
not ( n220821 , n220820 );
not ( n220822 , n216810 );
not ( n220823 , n41165 );
not ( n220824 , n220823 );
or ( n220825 , n220822 , n220824 );
nand ( n220826 , n219389 , n215289 );
nand ( n220827 , n220825 , n220826 );
not ( n220828 , n220827 );
or ( n220829 , n220821 , n220828 );
nand ( n220830 , n220647 , n216299 );
nand ( n220831 , n220829 , n220830 );
xor ( n220832 , n220760 , n220831 );
not ( n220833 , n220468 );
not ( n220834 , n219461 );
or ( n220835 , n220833 , n220834 );
not ( n220836 , n215075 );
not ( n220837 , n218209 );
or ( n220838 , n220836 , n220837 );
nand ( n220839 , n218771 , n215899 );
nand ( n220840 , n220838 , n220839 );
nand ( n220841 , n220840 , n218533 );
nand ( n220842 , n220835 , n220841 );
xor ( n220843 , n220832 , n220842 );
xor ( n220844 , n220713 , n220843 );
xor ( n220845 , n220844 , n220709 );
xor ( n220846 , n220713 , n220843 );
and ( n220847 , n220846 , n220709 );
and ( n220848 , n220713 , n220843 );
or ( n220849 , n220847 , n220848 );
not ( n220850 , n220488 );
buf ( n220851 , n218832 );
buf ( n220852 , n218826 );
nor ( n220853 , n220851 , n220852 );
not ( n220854 , n220853 );
or ( n220855 , n220850 , n220854 );
not ( n220856 , n216964 );
not ( n220857 , n218876 );
or ( n220858 , n220856 , n220857 );
not ( n220859 , n218814 );
buf ( n220860 , n220859 );
nand ( n220861 , n220860 , n214678 );
nand ( n220862 , n220858 , n220861 );
nand ( n220863 , n218843 , n220862 );
nand ( n220864 , n220855 , n220863 );
xor ( n220865 , n220864 , n220814 );
not ( n220866 , n220514 );
not ( n220867 , n219435 );
or ( n220868 , n220866 , n220867 );
not ( n220869 , n217044 );
not ( n220870 , n220181 );
or ( n220871 , n220869 , n220870 );
nand ( n220872 , n219800 , n215131 );
nand ( n220873 , n220871 , n220872 );
nand ( n220874 , n219076 , n220873 );
nand ( n220875 , n220868 , n220874 );
xor ( n220876 , n220865 , n220875 );
xor ( n220877 , n220717 , n220876 );
not ( n220878 , n220502 );
not ( n220879 , n220492 );
or ( n220880 , n220878 , n220879 );
buf ( n220881 , n219778 );
not ( n220882 , n213583 );
not ( n220883 , n220499 );
or ( n220884 , n220882 , n220883 );
nand ( n220885 , n220150 , n214134 );
nand ( n220886 , n220884 , n220885 );
nand ( n220887 , n220881 , n220886 );
nand ( n220888 , n220880 , n220887 );
not ( n220889 , n37704 );
not ( n220890 , n219064 );
or ( n220891 , n220889 , n220890 );
nand ( n220892 , n220891 , n37458 );
nand ( n220893 , n33568 , n33573 );
not ( n220894 , n220893 );
and ( n220895 , n220892 , n220894 );
not ( n220896 , n220892 );
and ( n220897 , n220896 , n220893 );
nor ( n220898 , n220895 , n220897 );
buf ( n220899 , n220898 );
buf ( n220900 , n220899 );
not ( n220901 , n220900 );
and ( n220902 , n213750 , n220901 );
not ( n220903 , n213750 );
not ( n220904 , n220899 );
buf ( n220905 , n220904 );
not ( n220906 , n220905 );
and ( n220907 , n220903 , n220906 );
or ( n220908 , n220902 , n220907 );
not ( n220909 , n220908 );
not ( n220910 , n220899 );
not ( n220911 , n220633 );
not ( n220912 , n220911 );
not ( n220913 , n220912 );
and ( n220914 , n220910 , n220913 );
and ( n220915 , n220899 , n220912 );
nor ( n220916 , n220914 , n220915 );
not ( n220917 , n220635 );
nand ( n220918 , n220916 , n220917 );
not ( n220919 , n220918 );
not ( n220920 , n220919 );
or ( n220921 , n220909 , n220920 );
not ( n220922 , n218224 );
not ( n220923 , n220901 );
or ( n220924 , n220922 , n220923 );
not ( n220925 , n220901 );
nand ( n220926 , n220925 , n216076 );
nand ( n220927 , n220924 , n220926 );
buf ( n220928 , n220634 );
not ( n220929 , n220928 );
buf ( n220930 , n220929 );
nand ( n220931 , n220927 , n220930 );
nand ( n220932 , n220921 , n220931 );
xor ( n220933 , n220888 , n220932 );
xor ( n220934 , n220933 , n220697 );
xor ( n220935 , n220877 , n220934 );
xor ( n220936 , n220717 , n220876 );
and ( n220937 , n220936 , n220934 );
and ( n220938 , n220717 , n220876 );
or ( n220939 , n220937 , n220938 );
xor ( n220940 , n220721 , n220725 );
not ( n220941 , n214563 );
not ( n220942 , n220941 );
not ( n220943 , n217573 );
not ( n220944 , n218912 );
or ( n220945 , n220943 , n220944 );
nand ( n220946 , n218911 , n219390 );
nand ( n220947 , n220945 , n220946 );
not ( n220948 , n220947 );
or ( n220949 , n220942 , n220948 );
nand ( n220950 , n220573 , n218467 );
nand ( n220951 , n220949 , n220950 );
xor ( n220952 , n220701 , n220951 );
and ( n220953 , n220912 , n213750 );
nor ( n220954 , n220953 , n220150 );
nor ( n220955 , n220912 , n213750 );
or ( n220956 , n220954 , n220955 );
nand ( n220957 , n220956 , n220925 );
not ( n220958 , n220957 );
xor ( n220959 , n220958 , n220404 );
xor ( n220960 , n220959 , n220445 );
xor ( n220961 , n220952 , n220960 );
xor ( n220962 , n220940 , n220961 );
xor ( n220963 , n220721 , n220725 );
and ( n220964 , n220963 , n220961 );
and ( n220965 , n220721 , n220725 );
or ( n220966 , n220964 , n220965 );
not ( n220967 , n40258 );
not ( n220968 , n213382 );
and ( n220969 , n220967 , n220968 );
not ( n220970 , n40258 );
not ( n220971 , n220970 );
and ( n220972 , n220971 , n213382 );
nor ( n220973 , n220969 , n220972 );
or ( n220974 , n220973 , n213171 );
not ( n220975 , n220602 );
nand ( n220976 , n220975 , n217969 );
nand ( n220977 , n220974 , n220976 );
xor ( n220978 , n220705 , n220977 );
not ( n220979 , n215113 );
not ( n220980 , n218268 );
or ( n220981 , n220979 , n220980 );
nand ( n220982 , n40710 , n216037 );
nand ( n220983 , n220981 , n220982 );
not ( n220984 , n220983 );
buf ( n220985 , n216239 );
not ( n220986 , n220985 );
or ( n220987 , n220984 , n220986 );
nand ( n220988 , n214717 , n220561 );
nand ( n220989 , n220987 , n220988 );
xor ( n220990 , n220978 , n220989 );
not ( n220991 , n214458 );
not ( n220992 , n219033 );
not ( n220993 , n215989 );
or ( n220994 , n220992 , n220993 );
nand ( n220995 , n217133 , n220538 );
nand ( n220996 , n220994 , n220995 );
not ( n220997 , n220996 );
or ( n220998 , n220991 , n220997 );
nand ( n220999 , n220540 , n219731 );
nand ( n221000 , n220998 , n220999 );
not ( n221001 , n219175 );
not ( n221002 , n218661 );
not ( n221003 , n220226 );
or ( n221004 , n221002 , n221003 );
nand ( n221005 , n217017 , n217119 );
nand ( n221006 , n221004 , n221005 );
not ( n221007 , n221006 );
or ( n221008 , n221001 , n221007 );
nand ( n221009 , n220453 , n217023 );
nand ( n221010 , n221008 , n221009 );
xor ( n221011 , n221000 , n221010 );
not ( n221012 , n219353 );
not ( n221013 , n217542 );
not ( n221014 , n217147 );
or ( n221015 , n221013 , n221014 );
not ( n221016 , n217147 );
nand ( n221017 , n221016 , n219358 );
nand ( n221018 , n221015 , n221017 );
not ( n221019 , n221018 );
or ( n221020 , n221012 , n221019 );
nand ( n221021 , n220611 , n217552 );
nand ( n221022 , n221020 , n221021 );
xor ( n221023 , n221011 , n221022 );
not ( n221024 , n213874 );
not ( n221025 , n220585 );
or ( n221026 , n221024 , n221025 );
not ( n221027 , n216262 );
not ( n221028 , n40668 );
not ( n221029 , n221028 );
or ( n221030 , n221027 , n221029 );
not ( n221031 , n40668 );
not ( n221032 , n221031 );
nand ( n221033 , n221032 , n220300 );
nand ( n221034 , n221030 , n221033 );
nand ( n221035 , n221034 , n217142 );
nand ( n221036 , n221026 , n221035 );
xor ( n221037 , n221023 , n221036 );
not ( n221038 , n216336 );
not ( n221039 , n213735 );
not ( n221040 , n40623 );
not ( n221041 , n221040 );
or ( n221042 , n221039 , n221041 );
nand ( n221043 , n219522 , n213732 );
nand ( n221044 , n221042 , n221043 );
not ( n221045 , n221044 );
or ( n221046 , n221038 , n221045 );
nand ( n221047 , n220659 , n213577 );
nand ( n221048 , n221046 , n221047 );
xor ( n221049 , n221037 , n221048 );
xor ( n221050 , n220990 , n221049 );
xor ( n221051 , n221050 , n220476 );
xor ( n221052 , n220990 , n221049 );
and ( n221053 , n221052 , n220476 );
and ( n221054 , n220990 , n221049 );
or ( n221055 , n221053 , n221054 );
xor ( n221056 , n220845 , n220522 );
xor ( n221057 , n221056 , n220935 );
xor ( n221058 , n220845 , n220522 );
and ( n221059 , n221058 , n220935 );
and ( n221060 , n220845 , n220522 );
or ( n221061 , n221059 , n221060 );
xor ( n221062 , n220554 , n220962 );
xor ( n221063 , n221062 , n220595 );
xor ( n221064 , n220554 , n220962 );
and ( n221065 , n221064 , n220595 );
and ( n221066 , n220554 , n220962 );
or ( n221067 , n221065 , n221066 );
xor ( n221068 , n221051 , n220669 );
xor ( n221069 , n221068 , n221057 );
xor ( n221070 , n221051 , n220669 );
and ( n221071 , n221070 , n221057 );
and ( n221072 , n221051 , n220669 );
or ( n221073 , n221071 , n221072 );
xor ( n221074 , n220675 , n220681 );
xor ( n221075 , n221074 , n221063 );
xor ( n221076 , n220675 , n220681 );
and ( n221077 , n221076 , n221063 );
and ( n221078 , n220675 , n220681 );
or ( n221079 , n221077 , n221078 );
xor ( n221080 , n221069 , n220687 );
xor ( n221081 , n221080 , n221075 );
xor ( n221082 , n221069 , n220687 );
and ( n221083 , n221082 , n221075 );
and ( n221084 , n221069 , n220687 );
or ( n221085 , n221083 , n221084 );
xor ( n221086 , n221000 , n221010 );
and ( n221087 , n221086 , n221022 );
and ( n221088 , n221000 , n221010 );
or ( n221089 , n221087 , n221088 );
xor ( n221090 , n220958 , n220404 );
and ( n221091 , n221090 , n220445 );
and ( n221092 , n220958 , n220404 );
or ( n221093 , n221091 , n221092 );
xor ( n221094 , n220760 , n220831 );
and ( n221095 , n221094 , n220842 );
and ( n221096 , n220760 , n220831 );
or ( n221097 , n221095 , n221096 );
xor ( n221098 , n220864 , n220814 );
and ( n221099 , n221098 , n220875 );
and ( n221100 , n220864 , n220814 );
or ( n221101 , n221099 , n221100 );
xor ( n221102 , n220888 , n220932 );
and ( n221103 , n221102 , n220697 );
and ( n221104 , n220888 , n220932 );
or ( n221105 , n221103 , n221104 );
xor ( n221106 , n220701 , n220951 );
and ( n221107 , n221106 , n220960 );
and ( n221108 , n220701 , n220951 );
or ( n221109 , n221107 , n221108 );
xor ( n221110 , n221023 , n221036 );
and ( n221111 , n221110 , n221048 );
and ( n221112 , n221023 , n221036 );
or ( n221113 , n221111 , n221112 );
xor ( n221114 , n220705 , n220977 );
and ( n221115 , n221114 , n220989 );
and ( n221116 , n220705 , n220977 );
or ( n221117 , n221115 , n221116 );
not ( n221118 , n217824 );
not ( n221119 , n214628 );
not ( n221120 , n221119 );
not ( n221121 , n216420 );
or ( n221122 , n221120 , n221121 );
nand ( n221123 , n214628 , n216762 );
nand ( n221124 , n221122 , n221123 );
not ( n221125 , n221124 );
or ( n221126 , n221118 , n221125 );
nand ( n221127 , n220806 , n218647 );
nand ( n221128 , n221126 , n221127 );
not ( n221129 , n215550 );
not ( n221130 , n215165 );
not ( n221131 , n216339 );
or ( n221132 , n221130 , n221131 );
not ( n221133 , n219724 );
nand ( n221134 , n221133 , n219326 );
nand ( n221135 , n221132 , n221134 );
not ( n221136 , n221135 );
or ( n221137 , n221129 , n221136 );
nand ( n221138 , n220792 , n215183 );
nand ( n221139 , n221137 , n221138 );
xor ( n221140 , n221128 , n221139 );
not ( n221141 , n216324 );
not ( n221142 , n220742 );
or ( n221143 , n221141 , n221142 );
and ( n221144 , n216068 , n215833 );
not ( n221145 , n216068 );
and ( n221146 , n221145 , n41716 );
or ( n221147 , n221144 , n221146 );
nand ( n221148 , n221147 , n216630 );
nand ( n221149 , n221143 , n221148 );
xor ( n221150 , n221140 , n221149 );
xor ( n221151 , n221128 , n221139 );
and ( n221152 , n221151 , n221149 );
and ( n221153 , n221128 , n221139 );
or ( n221154 , n221152 , n221153 );
not ( n221155 , n217486 );
not ( n221156 , n220755 );
or ( n221157 , n221155 , n221156 );
and ( n221158 , n218503 , n220749 );
not ( n221159 , n218503 );
and ( n221160 , n221159 , n216280 );
or ( n221161 , n221158 , n221160 );
nand ( n221162 , n221161 , n215587 );
nand ( n221163 , n221157 , n221162 );
not ( n221164 , n220773 );
not ( n221165 , n217089 );
or ( n221166 , n221164 , n221165 );
not ( n221167 , n218981 );
not ( n221168 , n216929 );
not ( n221169 , n221168 );
or ( n221170 , n221167 , n221169 );
nand ( n221171 , n217080 , n218980 );
nand ( n221172 , n221170 , n221171 );
nand ( n221173 , n221172 , n219119 );
nand ( n221174 , n221166 , n221173 );
xor ( n221175 , n221163 , n221174 );
not ( n221176 , n220783 );
not ( n221177 , n220059 );
or ( n221178 , n221176 , n221177 );
and ( n221179 , n217473 , n219102 );
not ( n221180 , n217473 );
and ( n221181 , n221180 , n216139 );
or ( n221182 , n221179 , n221181 );
nand ( n221183 , n221182 , n220067 );
nand ( n221184 , n221178 , n221183 );
xor ( n221185 , n221175 , n221184 );
xor ( n221186 , n221163 , n221174 );
and ( n221187 , n221186 , n221184 );
and ( n221188 , n221163 , n221174 );
or ( n221189 , n221187 , n221188 );
not ( n221190 , n217969 );
not ( n221191 , n220973 );
not ( n221192 , n221191 );
or ( n221193 , n221190 , n221192 );
not ( n221194 , n40396 );
and ( n221195 , n213382 , n221194 );
not ( n221196 , n213382 );
and ( n221197 , n221196 , n40397 );
or ( n221198 , n221195 , n221197 );
nand ( n221199 , n221198 , n214319 );
nand ( n221200 , n221193 , n221199 );
xor ( n221201 , n220764 , n221185 );
xor ( n221202 , n221201 , n221150 );
xor ( n221203 , n221200 , n221202 );
xor ( n221204 , n221203 , n221101 );
xor ( n221205 , n221200 , n221202 );
and ( n221206 , n221205 , n221101 );
and ( n221207 , n221200 , n221202 );
or ( n221208 , n221206 , n221207 );
xor ( n221209 , n221097 , n221105 );
not ( n221210 , n220840 );
not ( n221211 , n218525 );
or ( n221212 , n221210 , n221211 );
not ( n221213 , n218514 );
not ( n221214 , n218208 );
not ( n221215 , n221214 );
or ( n221216 , n221213 , n221215 );
nand ( n221217 , n219141 , n216170 );
nand ( n221218 , n221216 , n221217 );
nand ( n221219 , n221218 , n218232 );
nand ( n221220 , n221212 , n221219 );
not ( n221221 , n220873 );
not ( n221222 , n219792 );
or ( n221223 , n221221 , n221222 );
not ( n221224 , n214537 );
not ( n221225 , n219440 );
or ( n221226 , n221224 , n221225 );
buf ( n221227 , n219416 );
buf ( n221228 , n221227 );
nand ( n221229 , n221228 , n214899 );
nand ( n221230 , n221226 , n221229 );
nand ( n221231 , n219076 , n221230 );
nand ( n221232 , n221223 , n221231 );
xor ( n221233 , n221220 , n221232 );
not ( n221234 , n219449 );
not ( n221235 , n220862 );
or ( n221236 , n221234 , n221235 );
not ( n221237 , n218843 );
not ( n221238 , n220860 );
and ( n221239 , n216208 , n221238 );
not ( n221240 , n216208 );
buf ( n221241 , n219128 );
and ( n221242 , n221240 , n221241 );
nor ( n221243 , n221239 , n221242 );
or ( n221244 , n221237 , n221243 );
nand ( n221245 , n221236 , n221244 );
xor ( n221246 , n221233 , n221245 );
xor ( n221247 , n221209 , n221246 );
xor ( n221248 , n221097 , n221105 );
and ( n221249 , n221248 , n221246 );
and ( n221250 , n221097 , n221105 );
or ( n221251 , n221249 , n221250 );
not ( n221252 , n220886 );
not ( n221253 , n220492 );
or ( n221254 , n221252 , n221253 );
not ( n221255 , n214956 );
not ( n221256 , n220146 );
buf ( n221257 , n221256 );
not ( n221258 , n221257 );
or ( n221259 , n221255 , n221258 );
nand ( n221260 , n220151 , n214960 );
nand ( n221261 , n221259 , n221260 );
nand ( n221262 , n220881 , n221261 );
nand ( n221263 , n221254 , n221262 );
not ( n221264 , n220927 );
not ( n221265 , n220918 );
buf ( n221266 , n221265 );
not ( n221267 , n221266 );
or ( n221268 , n221264 , n221267 );
not ( n221269 , n213347 );
not ( n221270 , n220905 );
or ( n221271 , n221269 , n221270 );
nand ( n221272 , n220925 , n214616 );
nand ( n221273 , n221271 , n221272 );
nand ( n221274 , n221273 , n220930 );
nand ( n221275 , n221268 , n221274 );
xor ( n221276 , n221263 , n221275 );
xor ( n221277 , n221276 , n220818 );
xor ( n221278 , n221277 , n221117 );
not ( n221279 , n219314 );
not ( n221280 , n219687 );
not ( n221281 , n217394 );
or ( n221282 , n221280 , n221281 );
not ( n221283 , n219687 );
nand ( n221284 , n208717 , n221283 );
nand ( n221285 , n221282 , n221284 );
not ( n221286 , n221285 );
or ( n221287 , n221279 , n221286 );
nand ( n221288 , n220733 , n216426 );
nand ( n221289 , n221287 , n221288 );
and ( n221290 , n220796 , n220808 );
xor ( n221291 , n221289 , n221290 );
not ( n221292 , n214458 );
not ( n221293 , n219033 );
not ( n221294 , n219899 );
or ( n221295 , n221293 , n221294 );
nand ( n221296 , n216311 , n220538 );
nand ( n221297 , n221295 , n221296 );
not ( n221298 , n221297 );
or ( n221299 , n221292 , n221298 );
nand ( n221300 , n220996 , n219731 );
nand ( n221301 , n221299 , n221300 );
xor ( n221302 , n221291 , n221301 );
not ( n221303 , n214694 );
not ( n221304 , n216810 );
not ( n221305 , n219151 );
or ( n221306 , n221304 , n221305 );
not ( n221307 , n216810 );
nand ( n221308 , n208002 , n221307 );
nand ( n221309 , n221306 , n221308 );
not ( n221310 , n221309 );
or ( n221311 , n221303 , n221310 );
nand ( n221312 , n220827 , n216562 );
nand ( n221313 , n221311 , n221312 );
xor ( n221314 , n221302 , n221313 );
xor ( n221315 , n221314 , n221089 );
xor ( n221316 , n221278 , n221315 );
xor ( n221317 , n221277 , n221117 );
and ( n221318 , n221317 , n221315 );
and ( n221319 , n221277 , n221117 );
or ( n221320 , n221318 , n221319 );
xor ( n221321 , n221113 , n221109 );
xor ( n221322 , n221321 , n220849 );
xor ( n221323 , n221113 , n221109 );
and ( n221324 , n221323 , n220849 );
and ( n221325 , n221113 , n221109 );
or ( n221326 , n221324 , n221325 );
not ( n221327 , n213874 );
not ( n221328 , n221034 );
or ( n221329 , n221327 , n221328 );
not ( n221330 , n40409 );
and ( n221331 , n221330 , n216262 );
not ( n221332 , n221330 );
and ( n221333 , n221332 , n214824 );
or ( n221334 , n221331 , n221333 );
nand ( n221335 , n221334 , n217142 );
nand ( n221336 , n221329 , n221335 );
not ( n221337 , n220985 );
not ( n221338 , n217944 );
not ( n221339 , n221338 );
not ( n221340 , n40768 );
or ( n221341 , n221339 , n221340 );
not ( n221342 , n219234 );
nand ( n221343 , n221342 , n217944 );
nand ( n221344 , n221341 , n221343 );
not ( n221345 , n221344 );
or ( n221346 , n221337 , n221345 );
nand ( n221347 , n220983 , n214717 );
nand ( n221348 , n221346 , n221347 );
xor ( n221349 , n221336 , n221348 );
not ( n221350 , n213577 );
not ( n221351 , n221044 );
or ( n221352 , n221350 , n221351 );
not ( n221353 , n213735 );
not ( n221354 , n219742 );
or ( n221355 , n221353 , n221354 );
not ( n221356 , n207936 );
or ( n221357 , n221356 , n213735 );
nand ( n221358 , n221355 , n221357 );
nand ( n221359 , n221358 , n216336 );
nand ( n221360 , n221352 , n221359 );
xor ( n221361 , n221349 , n221360 );
not ( n221362 , n214086 );
not ( n221363 , n220947 );
or ( n221364 , n221362 , n221363 );
and ( n221365 , n217397 , n219880 );
not ( n221366 , n217397 );
and ( n221367 , n221366 , n219226 );
nor ( n221368 , n221365 , n221367 );
nand ( n221369 , n221368 , n215137 );
nand ( n221370 , n221364 , n221369 );
xor ( n221371 , n221093 , n221370 );
not ( n221372 , n217023 );
not ( n221373 , n221006 );
or ( n221374 , n221372 , n221373 );
and ( n221375 , n218661 , n218420 );
not ( n221376 , n218661 );
and ( n221377 , n221376 , n41069 );
nor ( n221378 , n221375 , n221377 );
nand ( n221379 , n221378 , n219175 );
nand ( n221380 , n221374 , n221379 );
and ( n221381 , n36640 , n37598 );
not ( n221382 , n36640 );
and ( n221383 , n221382 , n37597 );
nor ( n221384 , n221381 , n221383 );
xor ( n221385 , n220898 , n221384 );
not ( n221386 , n221385 );
not ( n221387 , n221386 );
and ( n221388 , n221387 , n215999 );
xor ( n221389 , n221380 , n221388 );
not ( n221390 , n217552 );
not ( n221391 , n221018 );
or ( n221392 , n221390 , n221391 );
not ( n221393 , n215955 );
not ( n221394 , n217314 );
or ( n221395 , n221393 , n221394 );
nand ( n221396 , n216859 , n219358 );
nand ( n221397 , n221395 , n221396 );
nand ( n221398 , n221397 , n219353 );
nand ( n221399 , n221392 , n221398 );
xor ( n221400 , n221389 , n221399 );
xor ( n221401 , n221371 , n221400 );
xor ( n221402 , n221361 , n221401 );
xor ( n221403 , n221402 , n221247 );
xor ( n221404 , n221361 , n221401 );
and ( n221405 , n221404 , n221247 );
and ( n221406 , n221361 , n221401 );
or ( n221407 , n221405 , n221406 );
xor ( n221408 , n220939 , n221204 );
xor ( n221409 , n221408 , n221322 );
xor ( n221410 , n220939 , n221204 );
and ( n221411 , n221410 , n221322 );
and ( n221412 , n220939 , n221204 );
or ( n221413 , n221411 , n221412 );
xor ( n221414 , n220966 , n221316 );
xor ( n221415 , n221414 , n221055 );
xor ( n221416 , n220966 , n221316 );
and ( n221417 , n221416 , n221055 );
and ( n221418 , n220966 , n221316 );
or ( n221419 , n221417 , n221418 );
xor ( n221420 , n221403 , n221061 );
xor ( n221421 , n221420 , n221067 );
xor ( n221422 , n221403 , n221061 );
and ( n221423 , n221422 , n221067 );
and ( n221424 , n221403 , n221061 );
or ( n221425 , n221423 , n221424 );
xor ( n221426 , n221409 , n221415 );
xor ( n221427 , n221426 , n221073 );
xor ( n221428 , n221409 , n221415 );
and ( n221429 , n221428 , n221073 );
and ( n221430 , n221409 , n221415 );
or ( n221431 , n221429 , n221430 );
xor ( n221432 , n221421 , n221079 );
xor ( n221433 , n221432 , n221427 );
xor ( n221434 , n221421 , n221079 );
and ( n221435 , n221434 , n221427 );
and ( n221436 , n221421 , n221079 );
or ( n221437 , n221435 , n221436 );
xor ( n221438 , n221289 , n221290 );
and ( n221439 , n221438 , n221301 );
and ( n221440 , n221289 , n221290 );
or ( n221441 , n221439 , n221440 );
xor ( n221442 , n221380 , n221388 );
and ( n221443 , n221442 , n221399 );
and ( n221444 , n221380 , n221388 );
or ( n221445 , n221443 , n221444 );
xor ( n221446 , n220764 , n221185 );
and ( n221447 , n221446 , n221150 );
and ( n221448 , n220764 , n221185 );
or ( n221449 , n221447 , n221448 );
xor ( n221450 , n221220 , n221232 );
and ( n221451 , n221450 , n221245 );
and ( n221452 , n221220 , n221232 );
or ( n221453 , n221451 , n221452 );
xor ( n221454 , n221263 , n221275 );
and ( n221455 , n221454 , n220818 );
and ( n221456 , n221263 , n221275 );
or ( n221457 , n221455 , n221456 );
xor ( n221458 , n221302 , n221313 );
and ( n221459 , n221458 , n221089 );
and ( n221460 , n221302 , n221313 );
or ( n221461 , n221459 , n221460 );
xor ( n221462 , n221093 , n221370 );
and ( n221463 , n221462 , n221400 );
and ( n221464 , n221093 , n221370 );
or ( n221465 , n221463 , n221464 );
xor ( n221466 , n221336 , n221348 );
and ( n221467 , n221466 , n221360 );
and ( n221468 , n221336 , n221348 );
or ( n221469 , n221467 , n221468 );
not ( n221470 , n217047 );
not ( n221471 , n216327 );
not ( n221472 , n214834 );
or ( n221473 , n221471 , n221472 );
nand ( n221474 , n214837 , n216014 );
nand ( n221475 , n221473 , n221474 );
not ( n221476 , n221475 );
or ( n221477 , n221470 , n221476 );
nand ( n221478 , n217864 , n221147 );
nand ( n221479 , n221477 , n221478 );
not ( n221480 , n216598 );
not ( n221481 , n216594 );
not ( n221482 , n216555 );
or ( n221483 , n221481 , n221482 );
nand ( n221484 , n215228 , n220802 );
nand ( n221485 , n221483 , n221484 );
not ( n221486 , n221485 );
or ( n221487 , n221480 , n221486 );
nand ( n221488 , n216586 , n221124 );
nand ( n221489 , n221487 , n221488 );
xor ( n221490 , n221479 , n221489 );
not ( n221491 , n221172 );
not ( n221492 , n220046 );
or ( n221493 , n221491 , n221492 );
buf ( n221494 , n214190 );
not ( n221495 , n221494 );
not ( n221496 , n221495 );
not ( n221497 , n217076 );
or ( n221498 , n221496 , n221497 );
nand ( n221499 , n216929 , n221494 );
nand ( n221500 , n221498 , n221499 );
nand ( n221501 , n221500 , n217388 );
nand ( n221502 , n221493 , n221501 );
xor ( n221503 , n221490 , n221502 );
xor ( n221504 , n221479 , n221489 );
and ( n221505 , n221504 , n221502 );
and ( n221506 , n221479 , n221489 );
or ( n221507 , n221505 , n221506 );
not ( n221508 , n220059 );
not ( n221509 , n221182 );
or ( n221510 , n221508 , n221509 );
and ( n221511 , n217611 , n219343 );
and ( n221512 , n217634 , n219348 );
nor ( n221513 , n221511 , n221512 );
or ( n221514 , n221513 , n217640 );
nand ( n221515 , n221510 , n221514 );
not ( n221516 , n215550 );
not ( n221517 , n218990 );
not ( n221518 , n215613 );
or ( n221519 , n221517 , n221518 );
not ( n221520 , n216089 );
not ( n221521 , n221520 );
nand ( n221522 , n221521 , n219326 );
nand ( n221523 , n221519 , n221522 );
not ( n221524 , n221523 );
or ( n221525 , n221516 , n221524 );
nand ( n221526 , n221135 , n215183 );
nand ( n221527 , n221525 , n221526 );
not ( n221528 , n217486 );
not ( n221529 , n221161 );
or ( n221530 , n221528 , n221529 );
not ( n221531 , n215766 );
not ( n221532 , n216046 );
or ( n221533 , n221531 , n221532 );
nand ( n221534 , n216608 , n216277 );
nand ( n221535 , n221533 , n221534 );
nand ( n221536 , n221535 , n220033 );
nand ( n221537 , n221530 , n221536 );
xor ( n221538 , n221527 , n221537 );
xor ( n221539 , n221515 , n221538 );
not ( n221540 , n220272 );
not ( n221541 , n217542 );
not ( n221542 , n217119 );
or ( n221543 , n221541 , n221542 );
nand ( n221544 , n217564 , n219358 );
nand ( n221545 , n221543 , n221544 );
not ( n221546 , n221545 );
or ( n221547 , n221540 , n221546 );
nand ( n221548 , n221397 , n220280 );
nand ( n221549 , n221547 , n221548 );
xor ( n221550 , n221539 , n221549 );
xor ( n221551 , n221515 , n221538 );
and ( n221552 , n221551 , n221549 );
and ( n221553 , n221515 , n221538 );
or ( n221554 , n221552 , n221553 );
not ( n221555 , n219175 );
not ( n221556 , n219577 );
not ( n221557 , n220823 );
or ( n221558 , n221556 , n221557 );
not ( n221559 , n220077 );
nand ( n221560 , n221559 , n219583 );
nand ( n221561 , n221558 , n221560 );
not ( n221562 , n221561 );
or ( n221563 , n221555 , n221562 );
nand ( n221564 , n221378 , n217023 );
nand ( n221565 , n221563 , n221564 );
xor ( n221566 , n221154 , n221565 );
xor ( n221567 , n221566 , n221503 );
xor ( n221568 , n221567 , n221453 );
xor ( n221569 , n221568 , n221457 );
xor ( n221570 , n221567 , n221453 );
and ( n221571 , n221570 , n221457 );
and ( n221572 , n221567 , n221453 );
or ( n221573 , n221571 , n221572 );
not ( n221574 , n221230 );
not ( n221575 , n219433 );
buf ( n221576 , n221575 );
not ( n221577 , n221576 );
or ( n221578 , n221574 , n221577 );
not ( n221579 , n216964 );
not ( n221580 , n219440 );
or ( n221581 , n221579 , n221580 );
nand ( n221582 , n220180 , n214678 );
nand ( n221583 , n221581 , n221582 );
nand ( n221584 , n221583 , n219076 );
nand ( n221585 , n221578 , n221584 );
not ( n221586 , n221261 );
not ( n221587 , n220164 );
or ( n221588 , n221586 , n221587 );
not ( n221589 , n214357 );
not ( n221590 , n220496 );
or ( n221591 , n221589 , n221590 );
not ( n221592 , n217044 );
not ( n221593 , n221257 );
nand ( n221594 , n221592 , n221593 );
nand ( n221595 , n221591 , n221594 );
nand ( n221596 , n219779 , n221595 );
nand ( n221597 , n221588 , n221596 );
xor ( n221598 , n221585 , n221597 );
buf ( n221599 , n33454 );
nand ( n221600 , n221599 , n33582 );
not ( n221601 , n221600 );
and ( n221602 , n36708 , n221601 );
not ( n221603 , n36708 );
and ( n221604 , n221603 , n221600 );
nor ( n221605 , n221602 , n221604 );
buf ( n221606 , n221605 );
buf ( n221607 , n221606 );
buf ( n221608 , n221607 );
and ( n221609 , n215999 , n221608 );
not ( n221610 , n215999 );
not ( n221611 , n221606 );
buf ( n221612 , n221611 );
and ( n221613 , n221610 , n221612 );
nor ( n221614 , n221609 , n221613 );
not ( n221615 , n221614 );
not ( n221616 , n221384 );
not ( n221617 , n221616 );
not ( n221618 , n221606 );
not ( n221619 , n221618 );
or ( n221620 , n221617 , n221619 );
nand ( n221621 , n221606 , n221384 );
nand ( n221622 , n221620 , n221621 );
nor ( n221623 , n221622 , n221385 );
not ( n221624 , n221623 );
not ( n221625 , n221624 );
buf ( n221626 , n221625 );
not ( n221627 , n221626 );
or ( n221628 , n221615 , n221627 );
not ( n221629 , n218224 );
not ( n221630 , n221612 );
or ( n221631 , n221629 , n221630 );
not ( n221632 , n221607 );
not ( n221633 , n221632 );
nand ( n221634 , n221633 , n216076 );
nand ( n221635 , n221631 , n221634 );
not ( n221636 , n221387 );
not ( n221637 , n221636 );
nand ( n221638 , n221635 , n221637 );
nand ( n221639 , n221628 , n221638 );
xor ( n221640 , n221598 , n221639 );
not ( n221641 , n221218 );
not ( n221642 , n218221 );
or ( n221643 , n221641 , n221642 );
not ( n221644 , n216934 );
not ( n221645 , n218226 );
or ( n221646 , n221644 , n221645 );
nand ( n221647 , n218208 , n216940 );
nand ( n221648 , n221646 , n221647 );
nand ( n221649 , n221648 , n218231 );
nand ( n221650 , n221643 , n221649 );
xor ( n221651 , n221189 , n221650 );
or ( n221652 , n221234 , n221243 );
not ( n221653 , n218815 );
not ( n221654 , n215899 );
and ( n221655 , n221653 , n221654 );
and ( n221656 , n220860 , n215899 );
nor ( n221657 , n221655 , n221656 );
or ( n221658 , n218456 , n221657 );
nand ( n221659 , n221652 , n221658 );
xor ( n221660 , n221651 , n221659 );
xor ( n221661 , n221640 , n221660 );
xor ( n221662 , n221661 , n221461 );
xor ( n221663 , n221640 , n221660 );
and ( n221664 , n221663 , n221461 );
and ( n221665 , n221640 , n221660 );
or ( n221666 , n221664 , n221665 );
not ( n221667 , n221273 );
not ( n221668 , n221266 );
or ( n221669 , n221667 , n221668 );
and ( n221670 , n213583 , n220901 );
not ( n221671 , n213583 );
and ( n221672 , n221671 , n220925 );
or ( n221673 , n221670 , n221672 );
not ( n221674 , n220928 );
nand ( n221675 , n221673 , n221674 );
nand ( n221676 , n221669 , n221675 );
xor ( n221677 , n221676 , n221550 );
xor ( n221678 , n221677 , n221441 );
xor ( n221679 , n221469 , n221678 );
xor ( n221680 , n221679 , n221465 );
xor ( n221681 , n221469 , n221678 );
and ( n221682 , n221681 , n221465 );
and ( n221683 , n221469 , n221678 );
or ( n221684 , n221682 , n221683 );
not ( n221685 , n215137 );
not ( n221686 , n213960 );
not ( n221687 , n40624 );
not ( n221688 , n221687 );
or ( n221689 , n221686 , n221688 );
not ( n221690 , n221040 );
nand ( n221691 , n221690 , n217397 );
nand ( n221692 , n221689 , n221691 );
not ( n221693 , n221692 );
or ( n221694 , n221685 , n221693 );
nand ( n221695 , n221368 , n215605 );
nand ( n221696 , n221694 , n221695 );
xor ( n221697 , n221445 , n221696 );
not ( n221698 , n214717 );
not ( n221699 , n221344 );
or ( n221700 , n221698 , n221699 );
not ( n221701 , n215113 );
not ( n221702 , n220204 );
or ( n221703 , n221701 , n221702 );
nand ( n221704 , n218911 , n216037 );
nand ( n221705 , n221703 , n221704 );
nand ( n221706 , n221705 , n220985 );
nand ( n221707 , n221700 , n221706 );
xor ( n221708 , n221697 , n221707 );
not ( n221709 , n214319 );
not ( n221710 , n213382 );
not ( n221711 , n40180 );
buf ( n221712 , n221711 );
not ( n221713 , n221712 );
or ( n221714 , n221710 , n221713 );
not ( n221715 , n40180 );
not ( n221716 , n221715 );
nand ( n221717 , n221716 , n217715 );
nand ( n221718 , n221714 , n221717 );
not ( n221719 , n221718 );
or ( n221720 , n221709 , n221719 );
nand ( n221721 , n221198 , n217969 );
nand ( n221722 , n221720 , n221721 );
not ( n221723 , n213498 );
not ( n221724 , n213735 );
not ( n221725 , n40668 );
not ( n221726 , n221725 );
or ( n221727 , n221724 , n221726 );
not ( n221728 , n221028 );
nand ( n221729 , n221728 , n213732 );
nand ( n221730 , n221727 , n221729 );
not ( n221731 , n221730 );
or ( n221732 , n221723 , n221731 );
nand ( n221733 , n221358 , n213577 );
nand ( n221734 , n221732 , n221733 );
xor ( n221735 , n221722 , n221734 );
xor ( n221736 , n221735 , n221449 );
xor ( n221737 , n221708 , n221736 );
not ( n221738 , n217142 );
not ( n221739 , n214818 );
not ( n221740 , n220971 );
or ( n221741 , n221739 , n221740 );
not ( n221742 , n40257 );
buf ( n221743 , n221742 );
nand ( n221744 , n221743 , n218887 );
nand ( n221745 , n221741 , n221744 );
not ( n221746 , n221745 );
or ( n221747 , n221738 , n221746 );
nand ( n221748 , n221334 , n213874 );
nand ( n221749 , n221747 , n221748 );
not ( n221750 , n219731 );
not ( n221751 , n221297 );
or ( n221752 , n221750 , n221751 );
not ( n221753 , n219033 );
not ( n221754 , n41249 );
or ( n221755 , n221753 , n221754 );
nand ( n221756 , n221016 , n220538 );
nand ( n221757 , n221755 , n221756 );
nand ( n221758 , n221757 , n214458 );
nand ( n221759 , n221752 , n221758 );
not ( n221760 , n219314 );
not ( n221761 , n219687 );
not ( n221762 , n215989 );
or ( n221763 , n221761 , n221762 );
nand ( n221764 , n219582 , n221283 );
nand ( n221765 , n221763 , n221764 );
not ( n221766 , n221765 );
or ( n221767 , n221760 , n221766 );
nand ( n221768 , n221285 , n216426 );
nand ( n221769 , n221767 , n221768 );
xor ( n221770 , n221759 , n221769 );
not ( n221771 , n220925 );
not ( n221772 , n221616 );
nand ( n221773 , n221772 , n215999 );
nand ( n221774 , n221771 , n221773 );
nand ( n221775 , n221616 , n213751 );
and ( n221776 , n221774 , n221775 );
not ( n221777 , n221607 );
buf ( n221778 , n221777 );
nor ( n221779 , n221776 , n221778 );
xor ( n221780 , n221770 , n221779 );
xor ( n221781 , n221749 , n221780 );
not ( n221782 , n221309 );
not ( n221783 , n216299 );
or ( n221784 , n221782 , n221783 );
not ( n221785 , n216810 );
not ( n221786 , n218268 );
or ( n221787 , n221785 , n221786 );
nand ( n221788 , n219594 , n215289 );
nand ( n221789 , n221787 , n221788 );
not ( n221790 , n221789 );
or ( n221791 , n221790 , n220819 );
nand ( n221792 , n221784 , n221791 );
xor ( n221793 , n221781 , n221792 );
xor ( n221794 , n221737 , n221793 );
xor ( n221795 , n221708 , n221736 );
and ( n221796 , n221795 , n221793 );
and ( n221797 , n221708 , n221736 );
or ( n221798 , n221796 , n221797 );
xor ( n221799 , n221208 , n221251 );
xor ( n221800 , n221799 , n221569 );
xor ( n221801 , n221208 , n221251 );
and ( n221802 , n221801 , n221569 );
and ( n221803 , n221208 , n221251 );
or ( n221804 , n221802 , n221803 );
xor ( n221805 , n221320 , n221662 );
xor ( n221806 , n221805 , n221680 );
xor ( n221807 , n221320 , n221662 );
and ( n221808 , n221807 , n221680 );
and ( n221809 , n221320 , n221662 );
or ( n221810 , n221808 , n221809 );
xor ( n221811 , n221326 , n221407 );
xor ( n221812 , n221811 , n221794 );
xor ( n221813 , n221326 , n221407 );
and ( n221814 , n221813 , n221794 );
and ( n221815 , n221326 , n221407 );
or ( n221816 , n221814 , n221815 );
xor ( n221817 , n221800 , n221419 );
xor ( n221818 , n221817 , n221413 );
xor ( n221819 , n221800 , n221419 );
and ( n221820 , n221819 , n221413 );
and ( n221821 , n221800 , n221419 );
or ( n221822 , n221820 , n221821 );
xor ( n221823 , n221806 , n221812 );
xor ( n221824 , n221823 , n221425 );
xor ( n221825 , n221806 , n221812 );
and ( n221826 , n221825 , n221425 );
and ( n221827 , n221806 , n221812 );
or ( n221828 , n221826 , n221827 );
xor ( n221829 , n221818 , n221431 );
xor ( n221830 , n221829 , n221824 );
xor ( n221831 , n221818 , n221431 );
and ( n221832 , n221831 , n221824 );
and ( n221833 , n221818 , n221431 );
or ( n221834 , n221832 , n221833 );
xor ( n221835 , n221759 , n221769 );
and ( n221836 , n221835 , n221779 );
and ( n221837 , n221759 , n221769 );
or ( n221838 , n221836 , n221837 );
xor ( n221839 , n221154 , n221565 );
and ( n221840 , n221839 , n221503 );
and ( n221841 , n221154 , n221565 );
or ( n221842 , n221840 , n221841 );
xor ( n221843 , n221189 , n221650 );
and ( n221844 , n221843 , n221659 );
and ( n221845 , n221189 , n221650 );
or ( n221846 , n221844 , n221845 );
xor ( n221847 , n221585 , n221597 );
and ( n221848 , n221847 , n221639 );
and ( n221849 , n221585 , n221597 );
or ( n221850 , n221848 , n221849 );
xor ( n221851 , n221676 , n221550 );
and ( n221852 , n221851 , n221441 );
and ( n221853 , n221676 , n221550 );
or ( n221854 , n221852 , n221853 );
xor ( n221855 , n221445 , n221696 );
and ( n221856 , n221855 , n221707 );
and ( n221857 , n221445 , n221696 );
or ( n221858 , n221856 , n221857 );
xor ( n221859 , n221749 , n221780 );
and ( n221860 , n221859 , n221792 );
and ( n221861 , n221749 , n221780 );
or ( n221862 , n221860 , n221861 );
xor ( n221863 , n221722 , n221734 );
and ( n221864 , n221863 , n221449 );
and ( n221865 , n221722 , n221734 );
or ( n221866 , n221864 , n221865 );
not ( n221867 , n215587 );
not ( n221868 , n220749 );
not ( n221869 , n216339 );
or ( n221870 , n221868 , n221869 );
not ( n221871 , n215820 );
nand ( n221872 , n221871 , n216277 );
nand ( n221873 , n221870 , n221872 );
not ( n221874 , n221873 );
or ( n221875 , n221867 , n221874 );
not ( n221876 , n216730 );
nand ( n221877 , n221876 , n221535 );
nand ( n221878 , n221875 , n221877 );
not ( n221879 , n216324 );
not ( n221880 , n221475 );
or ( n221881 , n221879 , n221880 );
not ( n221882 , n216068 );
not ( n221883 , n218503 );
or ( n221884 , n221882 , n221883 );
nand ( n221885 , n208725 , n216014 );
nand ( n221886 , n221884 , n221885 );
nand ( n221887 , n221886 , n216332 );
nand ( n221888 , n221881 , n221887 );
xor ( n221889 , n221878 , n221888 );
not ( n221890 , n217505 );
not ( n221891 , n221485 );
or ( n221892 , n221890 , n221891 );
not ( n221893 , n217511 );
not ( n221894 , n220424 );
not ( n221895 , n221894 );
or ( n221896 , n221893 , n221895 );
not ( n221897 , n215833 );
nand ( n221898 , n221897 , n216593 );
nand ( n221899 , n221896 , n221898 );
nand ( n221900 , n221899 , n216201 );
nand ( n221901 , n221892 , n221900 );
xor ( n221902 , n221889 , n221901 );
xor ( n221903 , n221878 , n221888 );
and ( n221904 , n221903 , n221901 );
and ( n221905 , n221878 , n221888 );
or ( n221906 , n221904 , n221905 );
not ( n221907 , n221500 );
not ( n221908 , n219368 );
or ( n221909 , n221907 , n221908 );
not ( n221910 , n30997 );
not ( n221911 , n221168 );
or ( n221912 , n221910 , n221911 );
nand ( n221913 , n216929 , n214628 );
nand ( n221914 , n221912 , n221913 );
nand ( n221915 , n221914 , n217388 );
nand ( n221916 , n221909 , n221915 );
not ( n221917 , n221513 );
not ( n221918 , n221917 );
not ( n221919 , n217631 );
or ( n221920 , n221918 , n221919 );
not ( n221921 , n218980 );
not ( n221922 , n221921 );
buf ( n221923 , n217472 );
not ( n221924 , n221923 );
not ( n221925 , n221924 );
or ( n221926 , n221922 , n221925 );
nand ( n221927 , n217614 , n218980 );
nand ( n221928 , n221926 , n221927 );
nand ( n221929 , n221928 , n218762 );
nand ( n221930 , n221920 , n221929 );
xor ( n221931 , n221916 , n221930 );
not ( n221932 , n215550 );
not ( n221933 , n221932 );
not ( n221934 , n221933 );
buf ( n221935 , n215165 );
and ( n221936 , n216261 , n221935 );
not ( n221937 , n216261 );
buf ( n221938 , n219326 );
and ( n221939 , n221937 , n221938 );
or ( n221940 , n221936 , n221939 );
not ( n221941 , n221940 );
or ( n221942 , n221934 , n221941 );
nand ( n221943 , n221523 , n219332 );
nand ( n221944 , n221942 , n221943 );
xor ( n221945 , n221931 , n221944 );
xor ( n221946 , n221916 , n221930 );
and ( n221947 , n221946 , n221944 );
and ( n221948 , n221916 , n221930 );
or ( n221949 , n221947 , n221948 );
not ( n221950 , n213577 );
not ( n221951 , n221730 );
or ( n221952 , n221950 , n221951 );
not ( n221953 , n213735 );
not ( n221954 , n220599 );
or ( n221955 , n221953 , n221954 );
not ( n221956 , n221330 );
nand ( n221957 , n221956 , n213732 );
nand ( n221958 , n221955 , n221957 );
nand ( n221959 , n221958 , n216336 );
nand ( n221960 , n221952 , n221959 );
xor ( n221961 , n221960 , n221842 );
xor ( n221962 , n221961 , n221846 );
xor ( n221963 , n221960 , n221842 );
and ( n221964 , n221963 , n221846 );
and ( n221965 , n221960 , n221842 );
or ( n221966 , n221964 , n221965 );
not ( n221967 , n221657 );
not ( n221968 , n221967 );
not ( n221969 , n219449 );
or ( n221970 , n221968 , n221969 );
not ( n221971 , n218514 );
not ( n221972 , n218876 );
or ( n221973 , n221971 , n221972 );
nand ( n221974 , n218815 , n216170 );
nand ( n221975 , n221973 , n221974 );
nand ( n221976 , n218843 , n221975 );
nand ( n221977 , n221970 , n221976 );
not ( n221978 , n221583 );
not ( n221979 , n219792 );
or ( n221980 , n221978 , n221979 );
not ( n221981 , n216208 );
not ( n221982 , n220181 );
or ( n221983 , n221981 , n221982 );
nand ( n221984 , n221228 , n216207 );
nand ( n221985 , n221983 , n221984 );
nand ( n221986 , n219076 , n221985 );
nand ( n221987 , n221980 , n221986 );
xor ( n221988 , n221977 , n221987 );
xor ( n221989 , n221988 , n221945 );
xor ( n221990 , n221850 , n221989 );
not ( n221991 , n221673 );
not ( n221992 , n220919 );
or ( n221993 , n221991 , n221992 );
not ( n221994 , n214956 );
not ( n221995 , n220901 );
or ( n221996 , n221994 , n221995 );
nand ( n221997 , n220925 , n214960 );
nand ( n221998 , n221996 , n221997 );
nand ( n221999 , n221998 , n220930 );
nand ( n222000 , n221993 , n221999 );
xor ( n222001 , n221902 , n222000 );
not ( n222002 , n219461 );
not ( n222003 , n221648 );
or ( n222004 , n222002 , n222003 );
not ( n222005 , n219102 );
not ( n222006 , n218209 );
or ( n222007 , n222005 , n222006 );
or ( n222008 , n218226 , n219102 );
nand ( n222009 , n222007 , n222008 );
not ( n222010 , n222009 );
or ( n222011 , n222010 , n217936 );
nand ( n222012 , n222004 , n222011 );
xor ( n222013 , n222001 , n222012 );
xor ( n222014 , n221990 , n222013 );
xor ( n222015 , n221850 , n221989 );
and ( n222016 , n222015 , n222013 );
and ( n222017 , n221850 , n221989 );
or ( n222018 , n222016 , n222017 );
not ( n222019 , n221595 );
not ( n222020 , n220492 );
or ( n222021 , n222019 , n222020 );
and ( n222022 , n214537 , n220499 );
not ( n222023 , n214537 );
and ( n222024 , n222023 , n220151 );
or ( n222025 , n222022 , n222024 );
nand ( n222026 , n219779 , n222025 );
nand ( n222027 , n222021 , n222026 );
not ( n222028 , n221635 );
not ( n222029 , n221626 );
or ( n222030 , n222028 , n222029 );
buf ( n222031 , n214616 );
not ( n222032 , n222031 );
and ( n222033 , n222032 , n221612 );
not ( n222034 , n222032 );
not ( n222035 , n221612 );
and ( n222036 , n222034 , n222035 );
nor ( n222037 , n222033 , n222036 );
not ( n222038 , n222037 );
nand ( n222039 , n222038 , n221637 );
nand ( n222040 , n222030 , n222039 );
xor ( n222041 , n222027 , n222040 );
not ( n222042 , n219175 );
not ( n222043 , n219577 );
not ( n222044 , n219151 );
or ( n222045 , n222043 , n222044 );
nand ( n222046 , n208002 , n218661 );
nand ( n222047 , n222045 , n222046 );
not ( n222048 , n222047 );
or ( n222049 , n222042 , n222048 );
nand ( n222050 , n221561 , n217023 );
nand ( n222051 , n222049 , n222050 );
xor ( n222052 , n222041 , n222051 );
xor ( n222053 , n221854 , n222052 );
xor ( n222054 , n222053 , n221862 );
xor ( n222055 , n221854 , n222052 );
and ( n222056 , n222055 , n221862 );
and ( n222057 , n221854 , n222052 );
or ( n222058 , n222056 , n222057 );
xor ( n222059 , n221858 , n221866 );
xor ( n222060 , n221554 , n221838 );
not ( n222061 , n215383 );
not ( n222062 , n213960 );
not ( n222063 , n220581 );
or ( n222064 , n222062 , n222063 );
nand ( n222065 , n207936 , n217397 );
nand ( n222066 , n222064 , n222065 );
not ( n222067 , n222066 );
or ( n222068 , n222061 , n222067 );
nand ( n222069 , n221692 , n214086 );
nand ( n222070 , n222068 , n222069 );
xor ( n222071 , n222060 , n222070 );
xor ( n222072 , n222059 , n222071 );
xor ( n222073 , n221858 , n221866 );
and ( n222074 , n222073 , n222071 );
and ( n222075 , n221858 , n221866 );
or ( n222076 , n222074 , n222075 );
xor ( n222077 , n221962 , n221573 );
not ( n222078 , n214717 );
not ( n222079 , n221705 );
or ( n222080 , n222078 , n222079 );
not ( n222081 , n40559 );
and ( n222082 , n222081 , n215113 );
not ( n222083 , n222081 );
and ( n222084 , n222083 , n217944 );
or ( n222085 , n222082 , n222084 );
nand ( n222086 , n222085 , n216239 );
nand ( n222087 , n222080 , n222086 );
not ( n222088 , n216562 );
not ( n222089 , n221789 );
or ( n222090 , n222088 , n222089 );
not ( n222091 , n216810 );
not ( n222092 , n220569 );
or ( n222093 , n222091 , n222092 );
nand ( n222094 , n208044 , n215289 );
nand ( n222095 , n222093 , n222094 );
nand ( n222096 , n222095 , n214694 );
nand ( n222097 , n222090 , n222096 );
xor ( n222098 , n222087 , n222097 );
not ( n222099 , n214319 );
not ( n222100 , n40421 );
not ( n222101 , n222100 );
and ( n222102 , n222101 , n217715 );
not ( n222103 , n222101 );
and ( n222104 , n222103 , n213382 );
or ( n222105 , n222102 , n222104 );
not ( n222106 , n222105 );
or ( n222107 , n222099 , n222106 );
nand ( n222108 , n221718 , n217969 );
nand ( n222109 , n222107 , n222108 );
xor ( n222110 , n222098 , n222109 );
xor ( n222111 , n222077 , n222110 );
xor ( n222112 , n221962 , n221573 );
and ( n222113 , n222112 , n222110 );
and ( n222114 , n221962 , n221573 );
or ( n222115 , n222113 , n222114 );
not ( n222116 , n213874 );
not ( n222117 , n221745 );
or ( n222118 , n222116 , n222117 );
not ( n222119 , n214818 );
not ( n222120 , n40396 );
buf ( n222121 , n222120 );
not ( n222122 , n222121 );
or ( n222123 , n222119 , n222122 );
not ( n222124 , n221194 );
nand ( n222125 , n222124 , n214824 );
nand ( n222126 , n222123 , n222125 );
nand ( n222127 , n222126 , n217142 );
nand ( n222128 , n222118 , n222127 );
not ( n222129 , n219314 );
not ( n222130 , n219687 );
not ( n222131 , n219899 );
or ( n222132 , n222130 , n222131 );
nand ( n222133 , n41319 , n221283 );
nand ( n222134 , n222132 , n222133 );
not ( n222135 , n222134 );
or ( n222136 , n222129 , n222135 );
nand ( n222137 , n221765 , n216426 );
nand ( n222138 , n222136 , n222137 );
not ( n222139 , n36673 );
nor ( n222140 , n222139 , n36593 );
not ( n222141 , n222140 );
not ( n222142 , n36319 );
or ( n222143 , n222141 , n222142 );
nand ( n222144 , n222143 , n37433 );
nand ( n222145 , n36615 , n36617 );
and ( n222146 , n222144 , n222145 );
not ( n222147 , n222144 );
not ( n222148 , n222145 );
and ( n222149 , n222147 , n222148 );
nor ( n222150 , n222146 , n222149 );
not ( n222151 , n222150 );
not ( n222152 , n222151 );
and ( n222153 , n221606 , n222152 );
not ( n222154 , n221606 );
and ( n222155 , n222154 , n222151 );
nor ( n222156 , n222153 , n222155 );
not ( n222157 , n222156 );
buf ( n222158 , n222157 );
not ( n222159 , n222158 );
nor ( n222160 , n222159 , n213751 );
xor ( n222161 , n222138 , n222160 );
xor ( n222162 , n222161 , n221507 );
xor ( n222163 , n222128 , n222162 );
and ( n222164 , n221527 , n221537 );
not ( n222165 , n217552 );
not ( n222166 , n221545 );
or ( n222167 , n222165 , n222166 );
not ( n222168 , n215955 );
not ( n222169 , n217330 );
or ( n222170 , n222168 , n222169 );
nand ( n222171 , n219201 , n219358 );
nand ( n222172 , n222170 , n222171 );
nand ( n222173 , n222172 , n219353 );
nand ( n222174 , n222167 , n222173 );
xor ( n222175 , n222164 , n222174 );
not ( n222176 , n219731 );
not ( n222177 , n221757 );
or ( n222178 , n222176 , n222177 );
not ( n222179 , n216166 );
not ( n222180 , n216859 );
not ( n222181 , n222180 );
or ( n222182 , n222179 , n222181 );
nand ( n222183 , n219050 , n220538 );
nand ( n222184 , n222182 , n222183 );
buf ( n222185 , n218077 );
nand ( n222186 , n222184 , n222185 );
nand ( n222187 , n222178 , n222186 );
xor ( n222188 , n222175 , n222187 );
xor ( n222189 , n222163 , n222188 );
xor ( n222190 , n222189 , n221666 );
xor ( n222191 , n222190 , n221684 );
xor ( n222192 , n222189 , n221666 );
and ( n222193 , n222192 , n221684 );
and ( n222194 , n222189 , n221666 );
or ( n222195 , n222193 , n222194 );
xor ( n222196 , n222054 , n222014 );
xor ( n222197 , n222196 , n222072 );
xor ( n222198 , n222054 , n222014 );
and ( n222199 , n222198 , n222072 );
and ( n222200 , n222054 , n222014 );
or ( n222201 , n222199 , n222200 );
xor ( n222202 , n221798 , n221804 );
xor ( n222203 , n222202 , n222111 );
xor ( n222204 , n221798 , n221804 );
and ( n222205 , n222204 , n222111 );
and ( n222206 , n221798 , n221804 );
or ( n222207 , n222205 , n222206 );
xor ( n222208 , n222191 , n221810 );
xor ( n222209 , n222208 , n222197 );
xor ( n222210 , n222191 , n221810 );
and ( n222211 , n222210 , n222197 );
and ( n222212 , n222191 , n221810 );
or ( n222213 , n222211 , n222212 );
xor ( n222214 , n221816 , n222203 );
xor ( n222215 , n222214 , n221822 );
xor ( n222216 , n221816 , n222203 );
and ( n222217 , n222216 , n221822 );
and ( n222218 , n221816 , n222203 );
or ( n222219 , n222217 , n222218 );
xor ( n222220 , n222164 , n222174 );
and ( n222221 , n222220 , n222187 );
and ( n222222 , n222164 , n222174 );
or ( n222223 , n222221 , n222222 );
xor ( n222224 , n222209 , n222215 );
xor ( n222225 , n222224 , n221828 );
xor ( n222226 , n222209 , n222215 );
and ( n222227 , n222226 , n221828 );
and ( n222228 , n222209 , n222215 );
or ( n222229 , n222227 , n222228 );
xor ( n222230 , n222138 , n222160 );
and ( n222231 , n222230 , n221507 );
and ( n222232 , n222138 , n222160 );
or ( n222233 , n222231 , n222232 );
xor ( n222234 , n221902 , n222000 );
and ( n222235 , n222234 , n222012 );
and ( n222236 , n221902 , n222000 );
or ( n222237 , n222235 , n222236 );
xor ( n222238 , n221977 , n221987 );
and ( n222239 , n222238 , n221945 );
and ( n222240 , n221977 , n221987 );
or ( n222241 , n222239 , n222240 );
xor ( n222242 , n222027 , n222040 );
and ( n222243 , n222242 , n222051 );
and ( n222244 , n222027 , n222040 );
or ( n222245 , n222243 , n222244 );
xor ( n222246 , n221554 , n221838 );
and ( n222247 , n222246 , n222070 );
and ( n222248 , n221554 , n221838 );
or ( n222249 , n222247 , n222248 );
xor ( n222250 , n222128 , n222162 );
and ( n222251 , n222250 , n222188 );
and ( n222252 , n222128 , n222162 );
or ( n222253 , n222251 , n222252 );
xor ( n222254 , n222087 , n222097 );
and ( n222255 , n222254 , n222109 );
and ( n222256 , n222087 , n222097 );
or ( n222257 , n222255 , n222256 );
not ( n222258 , n219501 );
not ( n222259 , n216594 );
not ( n222260 , n214834 );
or ( n222261 , n222259 , n222260 );
nand ( n222262 , n215642 , n216593 );
nand ( n222263 , n222261 , n222262 );
not ( n222264 , n222263 );
or ( n222265 , n222258 , n222264 );
nand ( n222266 , n217289 , n221899 );
nand ( n222267 , n222265 , n222266 );
not ( n222268 , n221914 );
not ( n222269 , n218544 );
not ( n222270 , n222269 );
not ( n222271 , n222270 );
or ( n222272 , n222268 , n222271 );
not ( n222273 , n41725 );
not ( n222274 , n217076 );
and ( n222275 , n222273 , n222274 );
and ( n222276 , n215228 , n217076 );
nor ( n222277 , n222275 , n222276 );
not ( n222278 , n222277 );
nand ( n222279 , n222278 , n217099 );
nand ( n222280 , n222272 , n222279 );
xor ( n222281 , n222267 , n222280 );
not ( n222282 , n221928 );
not ( n222283 , n220059 );
or ( n222284 , n222282 , n222283 );
not ( n222285 , n215533 );
not ( n222286 , n217615 );
or ( n222287 , n222285 , n222286 );
nand ( n222288 , n221923 , n220022 );
nand ( n222289 , n222287 , n222288 );
nand ( n222290 , n222289 , n220067 );
nand ( n222291 , n222284 , n222290 );
xor ( n222292 , n222281 , n222291 );
xor ( n222293 , n222267 , n222280 );
and ( n222294 , n222293 , n222291 );
and ( n222295 , n222267 , n222280 );
or ( n222296 , n222294 , n222295 );
not ( n222297 , n215587 );
and ( n222298 , n41563 , n220749 );
not ( n222299 , n41563 );
and ( n222300 , n222299 , n216277 );
or ( n222301 , n222298 , n222300 );
not ( n222302 , n222301 );
or ( n222303 , n222297 , n222302 );
nand ( n222304 , n221873 , n216731 );
nand ( n222305 , n222303 , n222304 );
not ( n222306 , n216065 );
not ( n222307 , n221886 );
or ( n222308 , n222306 , n222307 );
not ( n222309 , n216623 );
not ( n222310 , n216607 );
or ( n222311 , n222309 , n222310 );
nand ( n222312 , n41608 , n216014 );
nand ( n222313 , n222311 , n222312 );
nand ( n222314 , n222313 , n217047 );
nand ( n222315 , n222308 , n222314 );
xor ( n222316 , n222305 , n222315 );
not ( n222317 , n216204 );
not ( n222318 , n222134 );
or ( n222319 , n222317 , n222318 );
not ( n222320 , n219687 );
not ( n222321 , n41249 );
or ( n222322 , n222320 , n222321 );
not ( n222323 , n219687 );
nand ( n222324 , n216519 , n222323 );
nand ( n222325 , n222322 , n222324 );
nand ( n222326 , n222325 , n219314 );
nand ( n222327 , n222319 , n222326 );
xor ( n222328 , n222316 , n222327 );
not ( n222329 , n221933 );
not ( n222330 , n221935 );
not ( n222331 , n216500 );
or ( n222332 , n222330 , n222331 );
not ( n222333 , n221935 );
nand ( n222334 , n218786 , n222333 );
nand ( n222335 , n222332 , n222334 );
not ( n222336 , n222335 );
or ( n222337 , n222329 , n222336 );
nand ( n222338 , n221940 , n219332 );
nand ( n222339 , n222337 , n222338 );
xor ( n222340 , n222328 , n222339 );
xor ( n222341 , n222316 , n222327 );
and ( n222342 , n222341 , n222339 );
and ( n222343 , n222316 , n222327 );
or ( n222344 , n222342 , n222343 );
not ( n222345 , n219353 );
not ( n222346 , n215955 );
not ( n222347 , n219386 );
or ( n222348 , n222346 , n222347 );
nand ( n222349 , n41165 , n216989 );
nand ( n222350 , n222348 , n222349 );
not ( n222351 , n222350 );
or ( n222352 , n222345 , n222351 );
nand ( n222353 , n222172 , n220280 );
nand ( n222354 , n222352 , n222353 );
xor ( n222355 , n222292 , n222354 );
not ( n222356 , n222009 );
not ( n222357 , n218221 );
or ( n222358 , n222356 , n222357 );
not ( n222359 , n219343 );
not ( n222360 , n218226 );
or ( n222361 , n222359 , n222360 );
nand ( n222362 , n219141 , n219348 );
nand ( n222363 , n222361 , n222362 );
nand ( n222364 , n222363 , n218232 );
nand ( n222365 , n222358 , n222364 );
xor ( n222366 , n222355 , n222365 );
xor ( n222367 , n222366 , n222237 );
xor ( n222368 , n222367 , n222241 );
xor ( n222369 , n222366 , n222237 );
and ( n222370 , n222369 , n222241 );
and ( n222371 , n222366 , n222237 );
or ( n222372 , n222370 , n222371 );
not ( n222373 , n221975 );
not ( n222374 , n220853 );
or ( n222375 , n222373 , n222374 );
not ( n222376 , n218456 );
not ( n222377 , n216934 );
not ( n222378 , n218876 );
or ( n222379 , n222377 , n222378 );
nand ( n222380 , n220859 , n216940 );
nand ( n222381 , n222379 , n222380 );
nand ( n222382 , n222376 , n222381 );
nand ( n222383 , n222375 , n222382 );
not ( n222384 , n221985 );
not ( n222385 , n219792 );
or ( n222386 , n222384 , n222385 );
not ( n222387 , n215075 );
not ( n222388 , n220181 );
or ( n222389 , n222387 , n222388 );
nand ( n222390 , n221228 , n215899 );
nand ( n222391 , n222389 , n222390 );
nand ( n222392 , n219076 , n222391 );
nand ( n222393 , n222386 , n222392 );
xor ( n222394 , n222383 , n222393 );
not ( n222395 , n221998 );
not ( n222396 , n221266 );
or ( n222397 , n222395 , n222396 );
not ( n222398 , n217044 );
buf ( n222399 , n220900 );
not ( n222400 , n222399 );
not ( n222401 , n222400 );
or ( n222402 , n222398 , n222401 );
nand ( n222403 , n222399 , n215131 );
nand ( n222404 , n222402 , n222403 );
nand ( n222405 , n222404 , n220930 );
nand ( n222406 , n222397 , n222405 );
xor ( n222407 , n222394 , n222406 );
not ( n222408 , n222025 );
not ( n222409 , n220492 );
or ( n222410 , n222408 , n222409 );
not ( n222411 , n219475 );
not ( n222412 , n220145 );
not ( n222413 , n222412 );
not ( n222414 , n222413 );
not ( n222415 , n222414 );
or ( n222416 , n222411 , n222415 );
nand ( n222417 , n220150 , n214678 );
nand ( n222418 , n222416 , n222417 );
nand ( n222419 , n219779 , n222418 );
nand ( n222420 , n222410 , n222419 );
not ( n222421 , n37702 );
not ( n222422 , n222421 );
not ( n222423 , n36622 );
not ( n222424 , n222423 );
or ( n222425 , n222422 , n222424 );
nand ( n222426 , n36622 , n37702 );
nand ( n222427 , n222425 , n222426 );
buf ( n222428 , n222427 );
not ( n222429 , n222428 );
not ( n222430 , n222429 );
and ( n222431 , n215999 , n222430 );
not ( n222432 , n215999 );
buf ( n222433 , n222428 );
buf ( n222434 , n222433 );
not ( n222435 , n222434 );
and ( n222436 , n222432 , n222435 );
nor ( n222437 , n222431 , n222436 );
not ( n222438 , n222437 );
not ( n222439 , n222151 );
not ( n222440 , n222421 );
not ( n222441 , n222423 );
or ( n222442 , n222440 , n222441 );
nand ( n222443 , n222442 , n222426 );
not ( n222444 , n222443 );
and ( n222445 , n222439 , n222444 );
and ( n222446 , n222443 , n222151 );
nor ( n222447 , n222445 , n222446 );
not ( n222448 , n221606 );
or ( n222449 , n222448 , n222150 );
nand ( n222450 , n221618 , n222150 );
nand ( n222451 , n222449 , n222450 );
nand ( n222452 , n222447 , n222451 );
not ( n222453 , n222452 );
buf ( n222454 , n222453 );
not ( n222455 , n222454 );
or ( n222456 , n222438 , n222455 );
not ( n222457 , n218224 );
not ( n222458 , n222428 );
not ( n222459 , n222458 );
or ( n222460 , n222457 , n222459 );
not ( n222461 , n222433 );
not ( n222462 , n222461 );
nand ( n222463 , n222462 , n216076 );
nand ( n222464 , n222460 , n222463 );
not ( n222465 , n222156 );
not ( n222466 , n222465 );
not ( n222467 , n222466 );
nand ( n222468 , n222464 , n222467 );
nand ( n222469 , n222456 , n222468 );
xor ( n222470 , n222420 , n222469 );
not ( n222471 , n221626 );
or ( n222472 , n222471 , n222037 );
not ( n222473 , n213583 );
not ( n222474 , n221778 );
or ( n222475 , n222473 , n222474 );
nand ( n222476 , n221608 , n214134 );
nand ( n222477 , n222475 , n222476 );
not ( n222478 , n222477 );
or ( n222479 , n222478 , n221636 );
nand ( n222480 , n222472 , n222479 );
xor ( n222481 , n222470 , n222480 );
xor ( n222482 , n222407 , n222481 );
xor ( n222483 , n222482 , n222245 );
xor ( n222484 , n222407 , n222481 );
and ( n222485 , n222484 , n222245 );
and ( n222486 , n222407 , n222481 );
or ( n222487 , n222485 , n222486 );
xor ( n222488 , n222257 , n222249 );
xor ( n222489 , n221949 , n222223 );
xor ( n222490 , n222489 , n222233 );
xor ( n222491 , n222488 , n222490 );
xor ( n222492 , n222257 , n222249 );
and ( n222493 , n222492 , n222490 );
and ( n222494 , n222257 , n222249 );
or ( n222495 , n222493 , n222494 );
not ( n222496 , n215605 );
not ( n222497 , n222066 );
or ( n222498 , n222496 , n222497 );
not ( n222499 , n213960 );
not ( n222500 , n40668 );
not ( n222501 , n222500 );
or ( n222502 , n222499 , n222501 );
nand ( n222503 , n40668 , n215388 );
nand ( n222504 , n222502 , n222503 );
nand ( n222505 , n222504 , n215137 );
nand ( n222506 , n222498 , n222505 );
not ( n222507 , n211314 );
not ( n222508 , n213382 );
not ( n222509 , n40413 );
not ( n222510 , n222509 );
or ( n222511 , n222508 , n222510 );
not ( n222512 , n40413 );
not ( n222513 , n222512 );
nand ( n222514 , n222513 , n213381 );
nand ( n222515 , n222511 , n222514 );
not ( n222516 , n222515 );
or ( n222517 , n222507 , n222516 );
nand ( n222518 , n222105 , n217969 );
nand ( n222519 , n222517 , n222518 );
xor ( n222520 , n222506 , n222519 );
not ( n222521 , n213874 );
not ( n222522 , n222126 );
or ( n222523 , n222521 , n222522 );
not ( n222524 , n214818 );
not ( n222525 , n40181 );
or ( n222526 , n222524 , n222525 );
nand ( n222527 , n221716 , n214824 );
nand ( n222528 , n222526 , n222527 );
not ( n222529 , n222528 );
or ( n222530 , n222529 , n218150 );
nand ( n222531 , n222523 , n222530 );
xor ( n222532 , n222520 , n222531 );
xor ( n222533 , n222253 , n222532 );
xor ( n222534 , n222533 , n221966 );
xor ( n222535 , n222253 , n222532 );
and ( n222536 , n222535 , n221966 );
and ( n222537 , n222253 , n222532 );
or ( n222538 , n222536 , n222537 );
not ( n222539 , n220820 );
not ( n222540 , n216810 );
not ( n222541 , n219532 );
or ( n222542 , n222540 , n222541 );
not ( n222543 , n220204 );
nand ( n222544 , n222543 , n215289 );
nand ( n222545 , n222542 , n222544 );
not ( n222546 , n222545 );
or ( n222547 , n222539 , n222546 );
nand ( n222548 , n222095 , n216299 );
nand ( n222549 , n222547 , n222548 );
not ( n222550 , n216336 );
not ( n222551 , n213735 );
not ( n222552 , n221743 );
not ( n222553 , n222552 );
or ( n222554 , n222551 , n222553 );
nand ( n222555 , n220970 , n213732 );
nand ( n222556 , n222554 , n222555 );
not ( n222557 , n222556 );
or ( n222558 , n222550 , n222557 );
nand ( n222559 , n221958 , n213577 );
nand ( n222560 , n222558 , n222559 );
xor ( n222561 , n222549 , n222560 );
not ( n222562 , n219175 );
not ( n222563 , n219577 );
not ( n222564 , n218884 );
or ( n222565 , n222563 , n222564 );
nand ( n222566 , n219599 , n219583 );
nand ( n222567 , n222565 , n222566 );
not ( n222568 , n222567 );
or ( n222569 , n222562 , n222568 );
nand ( n222570 , n222047 , n217023 );
nand ( n222571 , n222569 , n222570 );
xor ( n222572 , n222561 , n222571 );
not ( n222573 , n214458 );
not ( n222574 , n216166 );
not ( n222575 , n220227 );
or ( n222576 , n222574 , n222575 );
nand ( n222577 , n220538 , n220226 );
nand ( n222578 , n222576 , n222577 );
not ( n222579 , n222578 );
or ( n222580 , n222573 , n222579 );
nand ( n222581 , n222184 , n219731 );
nand ( n222582 , n222580 , n222581 );
buf ( n222583 , n222151 );
nand ( n222584 , n222583 , n215999 );
not ( n222585 , n222584 );
not ( n222586 , n221608 );
not ( n222587 , n222586 );
or ( n222588 , n222585 , n222587 );
not ( n222589 , n222583 );
nand ( n222590 , n222589 , n213751 );
nand ( n222591 , n222588 , n222590 );
and ( n222592 , n222591 , n222462 );
xor ( n222593 , n222582 , n222592 );
xor ( n222594 , n222593 , n221906 );
not ( n222595 , n220985 );
not ( n222596 , n215113 );
not ( n222597 , n221687 );
or ( n222598 , n222596 , n222597 );
nand ( n222599 , n221690 , n216037 );
nand ( n222600 , n222598 , n222599 );
not ( n222601 , n222600 );
or ( n222602 , n222595 , n222601 );
nand ( n222603 , n222085 , n214717 );
nand ( n222604 , n222602 , n222603 );
xor ( n222605 , n222594 , n222604 );
xor ( n222606 , n222605 , n222340 );
xor ( n222607 , n222572 , n222606 );
xor ( n222608 , n222607 , n222018 );
xor ( n222609 , n222572 , n222606 );
and ( n222610 , n222609 , n222018 );
and ( n222611 , n222572 , n222606 );
or ( n222612 , n222610 , n222611 );
xor ( n222613 , n222368 , n222483 );
xor ( n222614 , n222613 , n222058 );
xor ( n222615 , n222368 , n222483 );
and ( n222616 , n222615 , n222058 );
and ( n222617 , n222368 , n222483 );
or ( n222618 , n222616 , n222617 );
xor ( n222619 , n222076 , n222491 );
xor ( n222620 , n222619 , n222115 );
xor ( n222621 , n222076 , n222491 );
and ( n222622 , n222621 , n222115 );
and ( n222623 , n222076 , n222491 );
or ( n222624 , n222622 , n222623 );
xor ( n222625 , n222608 , n222534 );
xor ( n222626 , n222625 , n222195 );
xor ( n222627 , n222608 , n222534 );
and ( n222628 , n222627 , n222195 );
and ( n222629 , n222608 , n222534 );
or ( n222630 , n222628 , n222629 );
xor ( n222631 , n222614 , n222201 );
xor ( n222632 , n222631 , n222620 );
xor ( n222633 , n222614 , n222201 );
and ( n222634 , n222633 , n222620 );
and ( n222635 , n222614 , n222201 );
or ( n222636 , n222634 , n222635 );
xor ( n222637 , n222207 , n222626 );
xor ( n222638 , n222637 , n222213 );
xor ( n222639 , n222207 , n222626 );
and ( n222640 , n222639 , n222213 );
and ( n222641 , n222207 , n222626 );
or ( n222642 , n222640 , n222641 );
xor ( n222643 , n222582 , n222592 );
and ( n222644 , n222643 , n221906 );
and ( n222645 , n222582 , n222592 );
or ( n222646 , n222644 , n222645 );
xor ( n222647 , n222632 , n222638 );
xor ( n222648 , n222647 , n222219 );
xor ( n222649 , n222632 , n222638 );
and ( n222650 , n222649 , n222219 );
and ( n222651 , n222632 , n222638 );
or ( n222652 , n222650 , n222651 );
xor ( n222653 , n222292 , n222354 );
and ( n222654 , n222653 , n222365 );
and ( n222655 , n222292 , n222354 );
or ( n222656 , n222654 , n222655 );
xor ( n222657 , n222383 , n222393 );
and ( n222658 , n222657 , n222406 );
and ( n222659 , n222383 , n222393 );
or ( n222660 , n222658 , n222659 );
xor ( n222661 , n222420 , n222469 );
and ( n222662 , n222661 , n222480 );
and ( n222663 , n222420 , n222469 );
or ( n222664 , n222662 , n222663 );
xor ( n222665 , n221949 , n222223 );
and ( n222666 , n222665 , n222233 );
and ( n222667 , n221949 , n222223 );
or ( n222668 , n222666 , n222667 );
xor ( n222669 , n222506 , n222519 );
and ( n222670 , n222669 , n222531 );
and ( n222671 , n222506 , n222519 );
or ( n222672 , n222670 , n222671 );
xor ( n222673 , n222594 , n222604 );
and ( n222674 , n222673 , n222340 );
and ( n222675 , n222594 , n222604 );
or ( n222676 , n222674 , n222675 );
xor ( n222677 , n222549 , n222560 );
and ( n222678 , n222677 , n222571 );
and ( n222679 , n222549 , n222560 );
or ( n222680 , n222678 , n222679 );
not ( n222681 , n217864 );
not ( n222682 , n222313 );
or ( n222683 , n222681 , n222682 );
not ( n222684 , n216068 );
not ( n222685 , n215820 );
or ( n222686 , n222684 , n222685 );
nand ( n222687 , n211451 , n216402 );
nand ( n222688 , n222686 , n222687 );
nand ( n222689 , n222688 , n216630 );
nand ( n222690 , n222683 , n222689 );
not ( n222691 , n217289 );
not ( n222692 , n222263 );
or ( n222693 , n222691 , n222692 );
not ( n222694 , n217511 );
not ( n222695 , n218503 );
or ( n222696 , n222694 , n222695 );
nand ( n222697 , n208725 , n216592 );
nand ( n222698 , n222696 , n222697 );
nand ( n222699 , n222698 , n216598 );
nand ( n222700 , n222693 , n222699 );
xor ( n222701 , n222690 , n222700 );
or ( n222702 , n222269 , n222277 );
not ( n222703 , n216928 );
not ( n222704 , n215833 );
or ( n222705 , n222703 , n222704 );
nand ( n222706 , n41716 , n217079 );
nand ( n222707 , n222705 , n222706 );
not ( n222708 , n222707 );
or ( n222709 , n222708 , n217098 );
nand ( n222710 , n222702 , n222709 );
xor ( n222711 , n222701 , n222710 );
xor ( n222712 , n222690 , n222700 );
and ( n222713 , n222712 , n222710 );
and ( n222714 , n222690 , n222700 );
or ( n222715 , n222713 , n222714 );
not ( n222716 , n222289 );
not ( n222717 , n217631 );
or ( n222718 , n222716 , n222717 );
not ( n222719 , n221119 );
not ( n222720 , n217473 );
or ( n222721 , n222719 , n222720 );
nand ( n222722 , n217614 , n217278 );
nand ( n222723 , n222721 , n222722 );
nand ( n222724 , n222723 , n218762 );
nand ( n222725 , n222718 , n222724 );
and ( n222726 , n222305 , n222315 );
xor ( n222727 , n222725 , n222726 );
not ( n222728 , n220033 );
not ( n222729 , n215766 );
not ( n222730 , n215793 );
or ( n222731 , n222729 , n222730 );
nand ( n222732 , n220753 , n215796 );
nand ( n222733 , n222731 , n222732 );
not ( n222734 , n222733 );
or ( n222735 , n222728 , n222734 );
nand ( n222736 , n222301 , n220414 );
nand ( n222737 , n222735 , n222736 );
xor ( n222738 , n222727 , n222737 );
xor ( n222739 , n222725 , n222726 );
and ( n222740 , n222739 , n222737 );
and ( n222741 , n222725 , n222726 );
or ( n222742 , n222740 , n222741 );
not ( n222743 , n219175 );
not ( n222744 , n219577 );
not ( n222745 , n219235 );
or ( n222746 , n222744 , n222745 );
nand ( n222747 , n220568 , n215971 );
nand ( n222748 , n222746 , n222747 );
not ( n222749 , n222748 );
or ( n222750 , n222743 , n222749 );
nand ( n222751 , n222567 , n217023 );
nand ( n222752 , n222750 , n222751 );
not ( n222753 , n222443 );
not ( n222754 , n222753 );
and ( n222755 , n36688 , n37596 );
not ( n222756 , n36688 );
and ( n222757 , n222756 , n37595 );
nor ( n222758 , n222755 , n222757 );
not ( n222759 , n222758 );
or ( n222760 , n222754 , n222759 );
and ( n222761 , n36688 , n37596 );
not ( n222762 , n36688 );
and ( n222763 , n222762 , n37595 );
nor ( n222764 , n222761 , n222763 );
not ( n222765 , n222764 );
nand ( n222766 , n222765 , n222443 );
nand ( n222767 , n222760 , n222766 );
buf ( n222768 , n222767 );
buf ( n222769 , n222768 );
and ( n222770 , n222769 , n215999 );
xor ( n222771 , n222770 , n222711 );
xor ( n222772 , n222771 , n222296 );
xor ( n222773 , n222752 , n222772 );
xor ( n222774 , n222773 , n222664 );
xor ( n222775 , n222752 , n222772 );
and ( n222776 , n222775 , n222664 );
and ( n222777 , n222752 , n222772 );
or ( n222778 , n222776 , n222777 );
xor ( n222779 , n222656 , n222660 );
xor ( n222780 , n222779 , n222668 );
xor ( n222781 , n222656 , n222660 );
and ( n222782 , n222781 , n222668 );
and ( n222783 , n222656 , n222660 );
or ( n222784 , n222782 , n222783 );
not ( n222785 , n222418 );
not ( n222786 , n220163 );
or ( n222787 , n222785 , n222786 );
not ( n222788 , n216208 );
not ( n222789 , n221256 );
or ( n222790 , n222788 , n222789 );
not ( n222791 , n220147 );
nand ( n222792 , n222791 , n216207 );
nand ( n222793 , n222790 , n222792 );
nand ( n222794 , n219779 , n222793 );
nand ( n222795 , n222787 , n222794 );
not ( n222796 , n222404 );
not ( n222797 , n220919 );
or ( n222798 , n222796 , n222797 );
not ( n222799 , n214537 );
not ( n222800 , n220905 );
or ( n222801 , n222799 , n222800 );
nand ( n222802 , n220900 , n214899 );
nand ( n222803 , n222801 , n222802 );
nand ( n222804 , n222803 , n220636 );
nand ( n222805 , n222798 , n222804 );
xor ( n222806 , n222795 , n222805 );
not ( n222807 , n222477 );
not ( n222808 , n221626 );
or ( n222809 , n222807 , n222808 );
not ( n222810 , n214956 );
not ( n222811 , n221777 );
or ( n222812 , n222810 , n222811 );
nand ( n222813 , n221607 , n214960 );
nand ( n222814 , n222812 , n222813 );
nand ( n222815 , n221387 , n222814 );
nand ( n222816 , n222809 , n222815 );
xor ( n222817 , n222806 , n222816 );
not ( n222818 , n222363 );
not ( n222819 , n218525 );
or ( n222820 , n222818 , n222819 );
not ( n222821 , n218980 );
not ( n222822 , n222821 );
not ( n222823 , n218226 );
or ( n222824 , n222822 , n222823 );
nand ( n222825 , n218208 , n218980 );
nand ( n222826 , n222824 , n222825 );
nand ( n222827 , n222826 , n218533 );
nand ( n222828 , n222820 , n222827 );
not ( n222829 , n222381 );
not ( n222830 , n219449 );
or ( n222831 , n222829 , n222830 );
and ( n222832 , n219102 , n218814 );
not ( n222833 , n219102 );
and ( n222834 , n222833 , n219128 );
or ( n222835 , n222832 , n222834 );
nand ( n222836 , n218843 , n222835 );
nand ( n222837 , n222831 , n222836 );
xor ( n222838 , n222828 , n222837 );
not ( n222839 , n222391 );
not ( n222840 , n219792 );
or ( n222841 , n222839 , n222840 );
not ( n222842 , n218514 );
not ( n222843 , n219440 );
or ( n222844 , n222842 , n222843 );
nand ( n222845 , n221228 , n216170 );
nand ( n222846 , n222844 , n222845 );
nand ( n222847 , n219076 , n222846 );
nand ( n222848 , n222841 , n222847 );
xor ( n222849 , n222838 , n222848 );
xor ( n222850 , n222817 , n222849 );
not ( n222851 , n220272 );
not ( n222852 , n217542 );
not ( n222853 , n219151 );
or ( n222854 , n222852 , n222853 );
nand ( n222855 , n40724 , n219358 );
nand ( n222856 , n222854 , n222855 );
not ( n222857 , n222856 );
or ( n222858 , n222851 , n222857 );
nand ( n222859 , n222350 , n220280 );
nand ( n222860 , n222858 , n222859 );
xor ( n222861 , n222860 , n222646 );
not ( n222862 , n214086 );
not ( n222863 , n222504 );
or ( n222864 , n222862 , n222863 );
not ( n222865 , n213960 );
not ( n222866 , n220596 );
or ( n222867 , n222865 , n222866 );
nand ( n222868 , n40410 , n217397 );
nand ( n222869 , n222867 , n222868 );
nand ( n222870 , n222869 , n220941 );
nand ( n222871 , n222864 , n222870 );
xor ( n222872 , n222861 , n222871 );
xor ( n222873 , n222850 , n222872 );
xor ( n222874 , n222817 , n222849 );
and ( n222875 , n222874 , n222872 );
and ( n222876 , n222817 , n222849 );
or ( n222877 , n222875 , n222876 );
xor ( n222878 , n222672 , n222676 );
xor ( n222879 , n222878 , n222680 );
xor ( n222880 , n222672 , n222676 );
and ( n222881 , n222880 , n222680 );
and ( n222882 , n222672 , n222676 );
or ( n222883 , n222881 , n222882 );
not ( n222884 , n222464 );
buf ( n222885 , n222452 );
not ( n222886 , n222885 );
not ( n222887 , n222886 );
or ( n222888 , n222884 , n222887 );
not ( n222889 , n222032 );
not ( n222890 , n222458 );
or ( n222891 , n222889 , n222890 );
not ( n222892 , n222458 );
nand ( n222893 , n222892 , n222031 );
nand ( n222894 , n222891 , n222893 );
nand ( n222895 , n222894 , n222467 );
nand ( n222896 , n222888 , n222895 );
xor ( n222897 , n222896 , n222738 );
xor ( n222898 , n222897 , n222344 );
not ( n222899 , n214717 );
not ( n222900 , n222600 );
or ( n222901 , n222899 , n222900 );
not ( n222902 , n215113 );
not ( n222903 , n221356 );
or ( n222904 , n222902 , n222903 );
nand ( n222905 , n207936 , n216037 );
nand ( n222906 , n222904 , n222905 );
nand ( n222907 , n222906 , n220985 );
nand ( n222908 , n222901 , n222907 );
not ( n222909 , n216562 );
not ( n222910 , n222545 );
or ( n222911 , n222909 , n222910 );
not ( n222912 , n215290 );
not ( n222913 , n40560 );
or ( n222914 , n222912 , n222913 );
nand ( n222915 , n40559 , n215289 );
nand ( n222916 , n222914 , n222915 );
nand ( n222917 , n222916 , n214694 );
nand ( n222918 , n222911 , n222917 );
xor ( n222919 , n222908 , n222918 );
not ( n222920 , n213577 );
not ( n222921 , n222556 );
or ( n222922 , n222920 , n222921 );
not ( n222923 , n213735 );
not ( n222924 , n222121 );
or ( n222925 , n222923 , n222924 );
nand ( n222926 , n40397 , n213732 );
nand ( n222927 , n222925 , n222926 );
nand ( n222928 , n222927 , n216336 );
nand ( n222929 , n222922 , n222928 );
xor ( n222930 , n222919 , n222929 );
xor ( n222931 , n222898 , n222930 );
xor ( n222932 , n222931 , n222372 );
xor ( n222933 , n222898 , n222930 );
and ( n222934 , n222933 , n222372 );
and ( n222935 , n222898 , n222930 );
or ( n222936 , n222934 , n222935 );
not ( n222937 , n217969 );
not ( n222938 , n222515 );
or ( n222939 , n222937 , n222938 );
not ( n222940 , n40484 );
and ( n222941 , n213382 , n222940 );
not ( n222942 , n213382 );
and ( n222943 , n222942 , n40485 );
or ( n222944 , n222941 , n222943 );
nand ( n222945 , n222944 , n213912 );
nand ( n222946 , n222939 , n222945 );
not ( n222947 , n213874 );
not ( n222948 , n222528 );
or ( n222949 , n222947 , n222948 );
not ( n222950 , n214824 );
not ( n222951 , n40421 );
not ( n222952 , n222951 );
not ( n222953 , n222952 );
or ( n222954 , n222950 , n222953 );
not ( n222955 , n222100 );
not ( n222956 , n222955 );
nand ( n222957 , n222956 , n216262 );
nand ( n222958 , n222954 , n222957 );
nand ( n222959 , n222958 , n217142 );
nand ( n222960 , n222949 , n222959 );
xor ( n222961 , n222946 , n222960 );
not ( n222962 , n216426 );
not ( n222963 , n222325 );
or ( n222964 , n222962 , n222963 );
not ( n222965 , n219687 );
not ( n222966 , n217856 );
or ( n222967 , n222965 , n222966 );
nand ( n222968 , n208164 , n222323 );
nand ( n222969 , n222967 , n222968 );
nand ( n222970 , n222969 , n219314 );
nand ( n222971 , n222964 , n222970 );
not ( n222972 , n219332 );
not ( n222973 , n222335 );
or ( n222974 , n222972 , n222973 );
not ( n222975 , n215165 );
not ( n222976 , n208594 );
or ( n222977 , n222975 , n222976 );
nand ( n222978 , n216306 , n219326 );
nand ( n222979 , n222977 , n222978 );
nand ( n222980 , n222979 , n221933 );
nand ( n222981 , n222974 , n222980 );
xor ( n222982 , n222971 , n222981 );
not ( n222983 , n214458 );
not ( n222984 , n219201 );
and ( n222985 , n222984 , n219033 );
not ( n222986 , n222984 );
and ( n222987 , n222986 , n219034 );
or ( n222988 , n222985 , n222987 );
not ( n222989 , n222988 );
or ( n222990 , n222983 , n222989 );
nand ( n222991 , n222578 , n219731 );
nand ( n222992 , n222990 , n222991 );
xor ( n222993 , n222982 , n222992 );
xor ( n222994 , n222961 , n222993 );
xor ( n222995 , n222994 , n222487 );
xor ( n222996 , n222995 , n222780 );
xor ( n222997 , n222994 , n222487 );
and ( n222998 , n222997 , n222780 );
and ( n222999 , n222994 , n222487 );
or ( n223000 , n222998 , n222999 );
xor ( n223001 , n222774 , n222873 );
xor ( n223002 , n223001 , n222495 );
xor ( n223003 , n222774 , n222873 );
and ( n223004 , n223003 , n222495 );
and ( n223005 , n222774 , n222873 );
or ( n223006 , n223004 , n223005 );
xor ( n223007 , n222879 , n222538 );
xor ( n223008 , n223007 , n222932 );
xor ( n223009 , n222879 , n222538 );
and ( n223010 , n223009 , n222932 );
and ( n223011 , n222879 , n222538 );
or ( n223012 , n223010 , n223011 );
xor ( n223013 , n222612 , n222996 );
xor ( n223014 , n223013 , n222618 );
xor ( n223015 , n222612 , n222996 );
and ( n223016 , n223015 , n222618 );
and ( n223017 , n222612 , n222996 );
or ( n223018 , n223016 , n223017 );
xor ( n223019 , n222624 , n223002 );
xor ( n223020 , n223019 , n223008 );
xor ( n223021 , n222624 , n223002 );
and ( n223022 , n223021 , n223008 );
and ( n223023 , n222624 , n223002 );
or ( n223024 , n223022 , n223023 );
xor ( n223025 , n222971 , n222981 );
and ( n223026 , n223025 , n222992 );
and ( n223027 , n222971 , n222981 );
or ( n223028 , n223026 , n223027 );
xor ( n223029 , n222630 , n223014 );
xor ( n223030 , n223029 , n222636 );
xor ( n223031 , n222630 , n223014 );
and ( n223032 , n223031 , n222636 );
and ( n223033 , n222630 , n223014 );
or ( n223034 , n223032 , n223033 );
xor ( n223035 , n223020 , n222642 );
xor ( n223036 , n223035 , n223030 );
xor ( n223037 , n223020 , n222642 );
and ( n223038 , n223037 , n223030 );
and ( n223039 , n223020 , n222642 );
or ( n223040 , n223038 , n223039 );
xor ( n223041 , n222770 , n222711 );
and ( n223042 , n223041 , n222296 );
and ( n223043 , n222770 , n222711 );
or ( n223044 , n223042 , n223043 );
xor ( n223045 , n222828 , n222837 );
and ( n223046 , n223045 , n222848 );
and ( n223047 , n222828 , n222837 );
or ( n223048 , n223046 , n223047 );
xor ( n223049 , n222795 , n222805 );
and ( n223050 , n223049 , n222816 );
and ( n223051 , n222795 , n222805 );
or ( n223052 , n223050 , n223051 );
xor ( n223053 , n222896 , n222738 );
and ( n223054 , n223053 , n222344 );
and ( n223055 , n222896 , n222738 );
or ( n223056 , n223054 , n223055 );
xor ( n223057 , n222860 , n222646 );
and ( n223058 , n223057 , n222871 );
and ( n223059 , n222860 , n222646 );
or ( n223060 , n223058 , n223059 );
xor ( n223061 , n222946 , n222960 );
and ( n223062 , n223061 , n222993 );
and ( n223063 , n222946 , n222960 );
or ( n223064 , n223062 , n223063 );
xor ( n223065 , n222908 , n222918 );
and ( n223066 , n223065 , n222929 );
and ( n223067 , n222908 , n222918 );
or ( n223068 , n223066 , n223067 );
not ( n223069 , n222707 );
not ( n223070 , n217875 );
or ( n223071 , n223069 , n223070 );
not ( n223072 , n216928 );
not ( n223073 , n216530 );
or ( n223074 , n223072 , n223073 );
nand ( n223075 , n30962 , n217079 );
nand ( n223076 , n223074 , n223075 );
nand ( n223077 , n223076 , n219119 );
nand ( n223078 , n223071 , n223077 );
not ( n223079 , n222723 );
not ( n223080 , n218239 );
or ( n223081 , n223079 , n223080 );
not ( n223082 , n217614 );
not ( n223083 , n214488 );
or ( n223084 , n223082 , n223083 );
nand ( n223085 , n217637 , n41725 );
nand ( n223086 , n223084 , n223085 );
nand ( n223087 , n223086 , n217230 );
nand ( n223088 , n223081 , n223087 );
xor ( n223089 , n223078 , n223088 );
not ( n223090 , n217864 );
not ( n223091 , n222688 );
or ( n223092 , n223090 , n223091 );
not ( n223093 , n216623 );
not ( n223094 , n41563 );
or ( n223095 , n223093 , n223094 );
nand ( n223096 , n216542 , n216402 );
nand ( n223097 , n223095 , n223096 );
nand ( n223098 , n223097 , n216630 );
nand ( n223099 , n223092 , n223098 );
not ( n223100 , n216762 );
not ( n223101 , n217066 );
or ( n223102 , n223100 , n223101 );
nand ( n223103 , n216420 , n41608 );
nand ( n223104 , n223102 , n223103 );
not ( n223105 , n223104 );
not ( n223106 , n216598 );
or ( n223107 , n223105 , n223106 );
nand ( n223108 , n222698 , n218647 );
nand ( n223109 , n223107 , n223108 );
xor ( n223110 , n223099 , n223109 );
xor ( n223111 , n223089 , n223110 );
xor ( n223112 , n223078 , n223088 );
and ( n223113 , n223112 , n223110 );
and ( n223114 , n223078 , n223088 );
or ( n223115 , n223113 , n223114 );
not ( n223116 , n215550 );
not ( n223117 , n218990 );
not ( n223118 , n41249 );
or ( n223119 , n223117 , n223118 );
nand ( n223120 , n218283 , n219326 );
nand ( n223121 , n223119 , n223120 );
not ( n223122 , n223121 );
or ( n223123 , n223116 , n223122 );
nand ( n223124 , n222979 , n215183 );
nand ( n223125 , n223123 , n223124 );
not ( n223126 , n220033 );
not ( n223127 , n215766 );
not ( n223128 , n215989 );
or ( n223129 , n223127 , n223128 );
nand ( n223130 , n41397 , n220038 );
nand ( n223131 , n223129 , n223130 );
not ( n223132 , n223131 );
or ( n223133 , n223126 , n223132 );
nand ( n223134 , n222733 , n217486 );
nand ( n223135 , n223133 , n223134 );
xor ( n223136 , n223125 , n223135 );
not ( n223137 , n213750 );
not ( n223138 , n222764 );
or ( n223139 , n223137 , n223138 );
nand ( n223140 , n223139 , n222461 );
not ( n223141 , n222764 );
nand ( n223142 , n223141 , n213751 );
and ( n223143 , n223140 , n223142 );
not ( n223144 , n37572 );
not ( n223145 , n36374 );
or ( n223146 , n223144 , n223145 );
nand ( n223147 , n223146 , n37476 );
nand ( n223148 , n33601 , n33426 );
not ( n223149 , n223148 );
and ( n223150 , n223147 , n223149 );
not ( n223151 , n223147 );
and ( n223152 , n223151 , n223148 );
nor ( n223153 , n223150 , n223152 );
buf ( n223154 , n223153 );
buf ( n223155 , n223154 );
not ( n223156 , n223155 );
nor ( n223157 , n223143 , n223156 );
xor ( n223158 , n223136 , n223157 );
xor ( n223159 , n223125 , n223135 );
and ( n223160 , n223159 , n223157 );
and ( n223161 , n223125 , n223135 );
or ( n223162 , n223160 , n223161 );
xor ( n223163 , n223044 , n223052 );
xor ( n223164 , n223163 , n223048 );
xor ( n223165 , n223044 , n223052 );
and ( n223166 , n223165 , n223048 );
and ( n223167 , n223044 , n223052 );
or ( n223168 , n223166 , n223167 );
not ( n223169 , n222814 );
not ( n223170 , n221625 );
or ( n223171 , n223169 , n223170 );
and ( n223172 , n217044 , n221607 );
not ( n223173 , n217044 );
and ( n223174 , n223173 , n221611 );
nor ( n223175 , n223172 , n223174 );
buf ( n223176 , n221386 );
not ( n223177 , n223176 );
nand ( n223178 , n223175 , n223177 );
nand ( n223179 , n223171 , n223178 );
xor ( n223180 , n223111 , n223179 );
not ( n223181 , n215999 );
buf ( n223182 , n223155 );
not ( n223183 , n223182 );
not ( n223184 , n223183 );
or ( n223185 , n223181 , n223184 );
not ( n223186 , n223155 );
not ( n223187 , n223186 );
nand ( n223188 , n223187 , n213751 );
nand ( n223189 , n223185 , n223188 );
not ( n223190 , n223189 );
and ( n223191 , n222427 , n222765 );
not ( n223192 , n222427 );
and ( n223193 , n223192 , n222764 );
nor ( n223194 , n223191 , n223193 );
xor ( n223195 , n223154 , n222764 );
nand ( n223196 , n223194 , n223195 );
not ( n223197 , n223196 );
not ( n223198 , n223197 );
or ( n223199 , n223190 , n223198 );
not ( n223200 , n218224 );
buf ( n223201 , n223154 );
buf ( n223202 , n223201 );
not ( n223203 , n223202 );
not ( n223204 , n223203 );
or ( n223205 , n223200 , n223204 );
nand ( n223206 , n223201 , n213077 );
nand ( n223207 , n223205 , n223206 );
nand ( n223208 , n222768 , n223207 );
nand ( n223209 , n223199 , n223208 );
xor ( n223210 , n223180 , n223209 );
xor ( n223211 , n223056 , n223210 );
not ( n223212 , n222793 );
not ( n223213 , n220163 );
or ( n223214 , n223212 , n223213 );
not ( n223215 , n215075 );
not ( n223216 , n220147 );
or ( n223217 , n223215 , n223216 );
nand ( n223218 , n222791 , n215899 );
nand ( n223219 , n223217 , n223218 );
nand ( n223220 , n223219 , n220881 );
nand ( n223221 , n223214 , n223220 );
not ( n223222 , n222803 );
and ( n223223 , n220916 , n220917 );
not ( n223224 , n223223 );
or ( n223225 , n223222 , n223224 );
not ( n223226 , n216964 );
not ( n223227 , n220900 );
buf ( n223228 , n223227 );
not ( n223229 , n223228 );
or ( n223230 , n223226 , n223229 );
nand ( n223231 , n220900 , n214678 );
nand ( n223232 , n223230 , n223231 );
nand ( n223233 , n223232 , n220636 );
nand ( n223234 , n223225 , n223233 );
xor ( n223235 , n223221 , n223234 );
not ( n223236 , n222894 );
not ( n223237 , n222886 );
or ( n223238 , n223236 , n223237 );
and ( n223239 , n213583 , n222458 );
not ( n223240 , n213583 );
and ( n223241 , n223240 , n222434 );
or ( n223242 , n223239 , n223241 );
not ( n223243 , n222156 );
buf ( n223244 , n223243 );
nand ( n223245 , n223242 , n223244 );
nand ( n223246 , n223238 , n223245 );
xor ( n223247 , n223235 , n223246 );
xor ( n223248 , n223211 , n223247 );
xor ( n223249 , n223056 , n223210 );
and ( n223250 , n223249 , n223247 );
and ( n223251 , n223056 , n223210 );
or ( n223252 , n223250 , n223251 );
not ( n223253 , n222826 );
not ( n223254 , n218525 );
or ( n223255 , n223253 , n223254 );
not ( n223256 , n215533 );
not ( n223257 , n218226 );
or ( n223258 , n223256 , n223257 );
nand ( n223259 , n218208 , n221494 );
nand ( n223260 , n223258 , n223259 );
nand ( n223261 , n223260 , n218533 );
nand ( n223262 , n223255 , n223261 );
not ( n223263 , n222835 );
not ( n223264 , n219449 );
or ( n223265 , n223263 , n223264 );
not ( n223266 , n219343 );
not ( n223267 , n218818 );
or ( n223268 , n223266 , n223267 );
not ( n223269 , n219343 );
nand ( n223270 , n219128 , n223269 );
nand ( n223271 , n223268 , n223270 );
nand ( n223272 , n223271 , n218843 );
nand ( n223273 , n223265 , n223272 );
xor ( n223274 , n223262 , n223273 );
not ( n223275 , n222846 );
not ( n223276 , n219435 );
or ( n223277 , n223275 , n223276 );
not ( n223278 , n216934 );
not ( n223279 , n219440 );
or ( n223280 , n223278 , n223279 );
nand ( n223281 , n220180 , n216940 );
nand ( n223282 , n223280 , n223281 );
nand ( n223283 , n219076 , n223282 );
nand ( n223284 , n223277 , n223283 );
xor ( n223285 , n223274 , n223284 );
xor ( n223286 , n223285 , n223060 );
xor ( n223287 , n222742 , n223028 );
not ( n223288 , n219314 );
and ( n223289 , n219687 , n217116 );
not ( n223290 , n219687 );
and ( n223291 , n223290 , n218137 );
or ( n223292 , n223289 , n223291 );
not ( n223293 , n223292 );
or ( n223294 , n223288 , n223293 );
nand ( n223295 , n222969 , n216426 );
nand ( n223296 , n223294 , n223295 );
xor ( n223297 , n222715 , n223296 );
not ( n223298 , n222185 );
not ( n223299 , n219033 );
not ( n223300 , n217710 );
or ( n223301 , n223299 , n223300 );
nand ( n223302 , n41165 , n220538 );
nand ( n223303 , n223301 , n223302 );
not ( n223304 , n223303 );
or ( n223305 , n223298 , n223304 );
nand ( n223306 , n222988 , n219731 );
nand ( n223307 , n223305 , n223306 );
xor ( n223308 , n223297 , n223307 );
xor ( n223309 , n223287 , n223308 );
xor ( n223310 , n223286 , n223309 );
xor ( n223311 , n223285 , n223060 );
and ( n223312 , n223311 , n223309 );
and ( n223313 , n223285 , n223060 );
or ( n223314 , n223312 , n223313 );
xor ( n223315 , n223068 , n223064 );
not ( n223316 , n213577 );
not ( n223317 , n222927 );
or ( n223318 , n223316 , n223317 );
not ( n223319 , n213735 );
buf ( n223320 , n40180 );
not ( n223321 , n223320 );
not ( n223322 , n223321 );
or ( n223323 , n223319 , n223322 );
nand ( n223324 , n40182 , n213732 );
nand ( n223325 , n223323 , n223324 );
nand ( n223326 , n223325 , n216336 );
nand ( n223327 , n223318 , n223326 );
not ( n223328 , n214319 );
not ( n223329 , n213382 );
not ( n223330 , n40545 );
not ( n223331 , n223330 );
or ( n223332 , n223329 , n223331 );
not ( n223333 , n223330 );
nand ( n223334 , n223333 , n217715 );
nand ( n223335 , n223332 , n223334 );
not ( n223336 , n223335 );
or ( n223337 , n223328 , n223336 );
nand ( n223338 , n222944 , n217969 );
nand ( n223339 , n223337 , n223338 );
xor ( n223340 , n223327 , n223339 );
not ( n223341 , n217023 );
not ( n223342 , n222748 );
or ( n223343 , n223341 , n223342 );
not ( n223344 , n219577 );
not ( n223345 , n220204 );
or ( n223346 , n223344 , n223345 );
nand ( n223347 , n219533 , n218661 );
nand ( n223348 , n223346 , n223347 );
nand ( n223349 , n223348 , n219175 );
nand ( n223350 , n223343 , n223349 );
xor ( n223351 , n223340 , n223350 );
xor ( n223352 , n223315 , n223351 );
xor ( n223353 , n223068 , n223064 );
and ( n223354 , n223353 , n223351 );
and ( n223355 , n223068 , n223064 );
or ( n223356 , n223354 , n223355 );
not ( n223357 , n222856 );
not ( n223358 , n220280 );
or ( n223359 , n223357 , n223358 );
and ( n223360 , n215955 , n218268 );
not ( n223361 , n215955 );
and ( n223362 , n223361 , n40710 );
nor ( n223363 , n223360 , n223362 );
or ( n223364 , n223363 , n217549 );
nand ( n223365 , n223359 , n223364 );
not ( n223366 , n217142 );
not ( n223367 , n214818 );
not ( n223368 , n40414 );
not ( n223369 , n223368 );
or ( n223370 , n223367 , n223369 );
nand ( n223371 , n222513 , n218887 );
nand ( n223372 , n223370 , n223371 );
not ( n223373 , n223372 );
or ( n223374 , n223366 , n223373 );
nand ( n223375 , n222958 , n213874 );
nand ( n223376 , n223374 , n223375 );
xor ( n223377 , n223365 , n223376 );
not ( n223378 , n222869 );
not ( n223379 , n215605 );
or ( n223380 , n223378 , n223379 );
not ( n223381 , n213960 );
not ( n223382 , n221742 );
not ( n223383 , n223382 );
not ( n223384 , n223383 );
not ( n223385 , n223384 );
or ( n223386 , n223381 , n223385 );
nand ( n223387 , n220970 , n217397 );
nand ( n223388 , n223386 , n223387 );
not ( n223389 , n223388 );
not ( n223390 , n217571 );
or ( n223391 , n223389 , n223390 );
nand ( n223392 , n223380 , n223391 );
xor ( n223393 , n223377 , n223392 );
not ( n223394 , n216239 );
not ( n223395 , n215113 );
not ( n223396 , n222500 );
or ( n223397 , n223395 , n223396 );
nand ( n223398 , n217944 , n40668 );
nand ( n223399 , n223397 , n223398 );
not ( n223400 , n223399 );
or ( n223401 , n223394 , n223400 );
nand ( n223402 , n222906 , n214717 );
nand ( n223403 , n223401 , n223402 );
xor ( n223404 , n223403 , n223158 );
not ( n223405 , n214694 );
not ( n223406 , n215290 );
not ( n223407 , n221040 );
or ( n223408 , n223406 , n223407 );
nand ( n223409 , n219522 , n215289 );
nand ( n223410 , n223408 , n223409 );
not ( n223411 , n223410 );
or ( n223412 , n223405 , n223411 );
nand ( n223413 , n222916 , n216562 );
nand ( n223414 , n223412 , n223413 );
xor ( n223415 , n223404 , n223414 );
xor ( n223416 , n223393 , n223415 );
xor ( n223417 , n223416 , n222778 );
xor ( n223418 , n223393 , n223415 );
and ( n223419 , n223418 , n222778 );
and ( n223420 , n223393 , n223415 );
or ( n223421 , n223419 , n223420 );
xor ( n223422 , n222784 , n223164 );
xor ( n223423 , n223422 , n223248 );
xor ( n223424 , n222784 , n223164 );
and ( n223425 , n223424 , n223248 );
and ( n223426 , n222784 , n223164 );
or ( n223427 , n223425 , n223426 );
xor ( n223428 , n222877 , n222883 );
xor ( n223429 , n223428 , n223352 );
xor ( n223430 , n222877 , n222883 );
and ( n223431 , n223430 , n223352 );
and ( n223432 , n222877 , n222883 );
or ( n223433 , n223431 , n223432 );
xor ( n223434 , n222936 , n223310 );
xor ( n223435 , n223434 , n223000 );
xor ( n223436 , n222936 , n223310 );
and ( n223437 , n223436 , n223000 );
and ( n223438 , n222936 , n223310 );
or ( n223439 , n223437 , n223438 );
xor ( n223440 , n223417 , n223423 );
xor ( n223441 , n223440 , n223006 );
xor ( n223442 , n223417 , n223423 );
and ( n223443 , n223442 , n223006 );
and ( n223444 , n223417 , n223423 );
or ( n223445 , n223443 , n223444 );
xor ( n223446 , n223429 , n223012 );
xor ( n223447 , n223446 , n223435 );
xor ( n223448 , n223429 , n223012 );
and ( n223449 , n223448 , n223435 );
and ( n223450 , n223429 , n223012 );
or ( n223451 , n223449 , n223450 );
xor ( n223452 , n222715 , n223296 );
and ( n223453 , n223452 , n223307 );
and ( n223454 , n222715 , n223296 );
or ( n223455 , n223453 , n223454 );
xor ( n223456 , n223018 , n223441 );
xor ( n223457 , n223456 , n223024 );
xor ( n223458 , n223018 , n223441 );
and ( n223459 , n223458 , n223024 );
and ( n223460 , n223018 , n223441 );
or ( n223461 , n223459 , n223460 );
xor ( n223462 , n223447 , n223457 );
xor ( n223463 , n223462 , n223034 );
xor ( n223464 , n223447 , n223457 );
and ( n223465 , n223464 , n223034 );
and ( n223466 , n223447 , n223457 );
or ( n223467 , n223465 , n223466 );
xor ( n223468 , n223262 , n223273 );
and ( n223469 , n223468 , n223284 );
and ( n223470 , n223262 , n223273 );
or ( n223471 , n223469 , n223470 );
xor ( n223472 , n223221 , n223234 );
and ( n223473 , n223472 , n223246 );
and ( n223474 , n223221 , n223234 );
or ( n223475 , n223473 , n223474 );
xor ( n223476 , n223111 , n223179 );
and ( n223477 , n223476 , n223209 );
and ( n223478 , n223111 , n223179 );
or ( n223479 , n223477 , n223478 );
xor ( n223480 , n222742 , n223028 );
and ( n223481 , n223480 , n223308 );
and ( n223482 , n222742 , n223028 );
or ( n223483 , n223481 , n223482 );
xor ( n223484 , n223365 , n223376 );
and ( n223485 , n223484 , n223392 );
and ( n223486 , n223365 , n223376 );
or ( n223487 , n223485 , n223486 );
xor ( n223488 , n223403 , n223158 );
and ( n223489 , n223488 , n223414 );
and ( n223490 , n223403 , n223158 );
or ( n223491 , n223489 , n223490 );
xor ( n223492 , n223327 , n223339 );
and ( n223493 , n223492 , n223350 );
and ( n223494 , n223327 , n223339 );
or ( n223495 , n223493 , n223494 );
not ( n223496 , n216201 );
not ( n223497 , n216762 );
not ( n223498 , n215820 );
or ( n223499 , n223497 , n223498 );
nand ( n223500 , n211451 , n216593 );
nand ( n223501 , n223499 , n223500 );
not ( n223502 , n223501 );
or ( n223503 , n223496 , n223502 );
nand ( n223504 , n223104 , n217289 );
nand ( n223505 , n223503 , n223504 );
not ( n223506 , n223076 );
not ( n223507 , n217089 );
or ( n223508 , n223506 , n223507 );
not ( n223509 , n216928 );
not ( n223510 , n218503 );
or ( n223511 , n223509 , n223510 );
nand ( n223512 , n219689 , n217602 );
nand ( n223513 , n223511 , n223512 );
nand ( n223514 , n223513 , n219119 );
nand ( n223515 , n223508 , n223514 );
xor ( n223516 , n223505 , n223515 );
not ( n223517 , n223086 );
not ( n223518 , n220059 );
or ( n223519 , n223517 , n223518 );
not ( n223520 , n218560 );
not ( n223521 , n215833 );
or ( n223522 , n223520 , n223521 );
nand ( n223523 , n221924 , n220424 );
nand ( n223524 , n223522 , n223523 );
nand ( n223525 , n223524 , n217641 );
nand ( n223526 , n223519 , n223525 );
xor ( n223527 , n223516 , n223526 );
xor ( n223528 , n223505 , n223515 );
and ( n223529 , n223528 , n223526 );
and ( n223530 , n223505 , n223515 );
or ( n223531 , n223529 , n223530 );
and ( n223532 , n223099 , n223109 );
not ( n223533 , n217047 );
not ( n223534 , n216015 );
not ( n223535 , n217941 );
or ( n223536 , n223534 , n223535 );
buf ( n223537 , n216059 );
nand ( n223538 , n218433 , n223537 );
nand ( n223539 , n223536 , n223538 );
not ( n223540 , n223539 );
or ( n223541 , n223533 , n223540 );
nand ( n223542 , n216619 , n223097 );
nand ( n223543 , n223541 , n223542 );
xor ( n223544 , n223532 , n223543 );
not ( n223545 , n221933 );
not ( n223546 , n215165 );
not ( n223547 , n217314 );
or ( n223548 , n223546 , n223547 );
not ( n223549 , n217856 );
nand ( n223550 , n223549 , n219326 );
nand ( n223551 , n223548 , n223550 );
not ( n223552 , n223551 );
or ( n223553 , n223545 , n223552 );
nand ( n223554 , n223121 , n215183 );
nand ( n223555 , n223553 , n223554 );
xor ( n223556 , n223544 , n223555 );
xor ( n223557 , n223532 , n223543 );
and ( n223558 , n223557 , n223555 );
and ( n223559 , n223532 , n223543 );
or ( n223560 , n223558 , n223559 );
not ( n223561 , n217023 );
not ( n223562 , n223348 );
or ( n223563 , n223561 , n223562 );
not ( n223564 , n219577 );
not ( n223565 , n222081 );
or ( n223566 , n223564 , n223565 );
nand ( n223567 , n40559 , n215971 );
nand ( n223568 , n223566 , n223567 );
nand ( n223569 , n223568 , n219175 );
nand ( n223570 , n223563 , n223569 );
xor ( n223571 , n223570 , n223455 );
xor ( n223572 , n223571 , n223475 );
xor ( n223573 , n223570 , n223455 );
and ( n223574 , n223573 , n223475 );
and ( n223575 , n223570 , n223455 );
or ( n223576 , n223574 , n223575 );
xor ( n223577 , n223479 , n223471 );
not ( n223578 , n223175 );
not ( n223579 , n221624 );
not ( n223580 , n223579 );
or ( n223581 , n223578 , n223580 );
and ( n223582 , n214899 , n221611 );
not ( n223583 , n214899 );
not ( n223584 , n221611 );
and ( n223585 , n223583 , n223584 );
nor ( n223586 , n223582 , n223585 );
not ( n223587 , n221386 );
nand ( n223588 , n223586 , n223587 );
nand ( n223589 , n223581 , n223588 );
not ( n223590 , n223207 );
not ( n223591 , n223196 );
not ( n223592 , n223591 );
or ( n223593 , n223590 , n223592 );
not ( n223594 , n222032 );
not ( n223595 , n223155 );
not ( n223596 , n223595 );
or ( n223597 , n223594 , n223596 );
nand ( n223598 , n223202 , n214616 );
nand ( n223599 , n223597 , n223598 );
nand ( n223600 , n223599 , n222769 );
nand ( n223601 , n223593 , n223600 );
xor ( n223602 , n223589 , n223601 );
not ( n223603 , n223242 );
not ( n223604 , n222886 );
or ( n223605 , n223603 , n223604 );
not ( n223606 , n214956 );
not ( n223607 , n222435 );
or ( n223608 , n223606 , n223607 );
nand ( n223609 , n222434 , n214960 );
nand ( n223610 , n223608 , n223609 );
nand ( n223611 , n223610 , n223244 );
nand ( n223612 , n223605 , n223611 );
xor ( n223613 , n223602 , n223612 );
xor ( n223614 , n223577 , n223613 );
xor ( n223615 , n223479 , n223471 );
and ( n223616 , n223615 , n223613 );
and ( n223617 , n223479 , n223471 );
or ( n223618 , n223616 , n223617 );
not ( n223619 , n223282 );
not ( n223620 , n219434 );
not ( n223621 , n223620 );
or ( n223622 , n223619 , n223621 );
not ( n223623 , n219102 );
not ( n223624 , n219440 );
or ( n223625 , n223623 , n223624 );
nand ( n223626 , n220180 , n216139 );
nand ( n223627 , n223625 , n223626 );
nand ( n223628 , n223627 , n219076 );
nand ( n223629 , n223622 , n223628 );
not ( n223630 , n223232 );
not ( n223631 , n223223 );
or ( n223632 , n223630 , n223631 );
not ( n223633 , n216208 );
not ( n223634 , n223227 );
or ( n223635 , n223633 , n223634 );
nand ( n223636 , n220900 , n216207 );
nand ( n223637 , n223635 , n223636 );
nand ( n223638 , n223637 , n221674 );
nand ( n223639 , n223632 , n223638 );
xor ( n223640 , n223629 , n223639 );
not ( n223641 , n223219 );
not ( n223642 , n220163 );
or ( n223643 , n223641 , n223642 );
not ( n223644 , n218514 );
not ( n223645 , n220147 );
or ( n223646 , n223644 , n223645 );
nand ( n223647 , n220150 , n216170 );
nand ( n223648 , n223646 , n223647 );
nand ( n223649 , n219779 , n223648 );
nand ( n223650 , n223643 , n223649 );
xor ( n223651 , n223640 , n223650 );
not ( n223652 , n223260 );
not ( n223653 , n219836 );
or ( n223654 , n223652 , n223653 );
not ( n223655 , n216293 );
not ( n223656 , n221214 );
or ( n223657 , n223655 , n223656 );
not ( n223658 , n216293 );
nand ( n223659 , n218208 , n223658 );
nand ( n223660 , n223657 , n223659 );
nand ( n223661 , n223660 , n218533 );
nand ( n223662 , n223654 , n223661 );
xor ( n223663 , n223527 , n223662 );
not ( n223664 , n223271 );
buf ( n223665 , n218835 );
not ( n223666 , n223665 );
or ( n223667 , n223664 , n223666 );
not ( n223668 , n221921 );
not ( n223669 , n218814 );
or ( n223670 , n223668 , n223669 );
buf ( n223671 , n218813 );
nand ( n223672 , n223671 , n218980 );
nand ( n223673 , n223670 , n223672 );
nand ( n223674 , n218843 , n223673 );
nand ( n223675 , n223667 , n223674 );
xor ( n223676 , n223663 , n223675 );
xor ( n223677 , n223651 , n223676 );
xor ( n223678 , n223677 , n223483 );
xor ( n223679 , n223651 , n223676 );
and ( n223680 , n223679 , n223483 );
and ( n223681 , n223651 , n223676 );
or ( n223682 , n223680 , n223681 );
xor ( n223683 , n223491 , n223487 );
not ( n223684 , n222185 );
not ( n223685 , n219033 );
not ( n223686 , n217964 );
or ( n223687 , n223685 , n223686 );
nand ( n223688 , n219034 , n40724 );
nand ( n223689 , n223687 , n223688 );
not ( n223690 , n223689 );
or ( n223691 , n223684 , n223690 );
nand ( n223692 , n223303 , n219731 );
nand ( n223693 , n223691 , n223692 );
xor ( n223694 , n223115 , n223693 );
xor ( n223695 , n223694 , n223556 );
xor ( n223696 , n223683 , n223695 );
xor ( n223697 , n223491 , n223487 );
and ( n223698 , n223697 , n223695 );
and ( n223699 , n223491 , n223487 );
or ( n223700 , n223698 , n223699 );
not ( n223701 , n220272 );
not ( n223702 , n215955 );
not ( n223703 , n219234 );
or ( n223704 , n223702 , n223703 );
nand ( n223705 , n208044 , n219358 );
nand ( n223706 , n223704 , n223705 );
not ( n223707 , n223706 );
or ( n223708 , n223701 , n223707 );
not ( n223709 , n223363 );
nand ( n223710 , n223709 , n217552 );
nand ( n223711 , n223708 , n223710 );
xor ( n223712 , n223162 , n223711 );
not ( n223713 , n213874 );
not ( n223714 , n223372 );
or ( n223715 , n223713 , n223714 );
not ( n223716 , n216262 );
not ( n223717 , n40485 );
not ( n223718 , n223717 );
or ( n223719 , n223716 , n223718 );
not ( n223720 , n214818 );
not ( n223721 , n40484 );
not ( n223722 , n223721 );
nand ( n223723 , n223720 , n223722 );
nand ( n223724 , n223719 , n223723 );
nand ( n223725 , n223724 , n217142 );
nand ( n223726 , n223715 , n223725 );
xor ( n223727 , n223712 , n223726 );
xor ( n223728 , n223495 , n223727 );
xor ( n223729 , n223728 , n223168 );
xor ( n223730 , n223495 , n223727 );
and ( n223731 , n223730 , n223168 );
and ( n223732 , n223495 , n223727 );
or ( n223733 , n223731 , n223732 );
not ( n223734 , n216562 );
not ( n223735 , n223410 );
or ( n223736 , n223734 , n223735 );
not ( n223737 , n215290 );
not ( n223738 , n221356 );
or ( n223739 , n223737 , n223738 );
nand ( n223740 , n207936 , n215289 );
nand ( n223741 , n223739 , n223740 );
nand ( n223742 , n223741 , n214694 );
nand ( n223743 , n223736 , n223742 );
not ( n223744 , n213577 );
not ( n223745 , n223325 );
or ( n223746 , n223744 , n223745 );
not ( n223747 , n213735 );
not ( n223748 , n40421 );
not ( n223749 , n223748 );
or ( n223750 , n223747 , n223749 );
not ( n223751 , n223748 );
nand ( n223752 , n223751 , n213732 );
nand ( n223753 , n223750 , n223752 );
nand ( n223754 , n216336 , n223753 );
nand ( n223755 , n223746 , n223754 );
xor ( n223756 , n223743 , n223755 );
not ( n223757 , n217969 );
not ( n223758 , n223335 );
or ( n223759 , n223757 , n223758 );
not ( n223760 , n213382 );
not ( n223761 , n40045 );
not ( n223762 , n223761 );
or ( n223763 , n223760 , n223762 );
not ( n223764 , n40044 );
not ( n223765 , n223764 );
nand ( n223766 , n223765 , n213381 );
nand ( n223767 , n223763 , n223766 );
nand ( n223768 , n223767 , n214319 );
nand ( n223769 , n223759 , n223768 );
xor ( n223770 , n223756 , n223769 );
xor ( n223771 , n223572 , n223770 );
not ( n223772 , n218467 );
not ( n223773 , n223388 );
or ( n223774 , n223772 , n223773 );
not ( n223775 , n217573 );
not ( n223776 , n221194 );
or ( n223777 , n223775 , n223776 );
nand ( n223778 , n40397 , n217397 );
nand ( n223779 , n223777 , n223778 );
nand ( n223780 , n223779 , n215137 );
nand ( n223781 , n223774 , n223780 );
not ( n223782 , n214717 );
not ( n223783 , n223399 );
or ( n223784 , n223782 , n223783 );
not ( n223785 , n215113 );
not ( n223786 , n40410 );
not ( n223787 , n223786 );
or ( n223788 , n223785 , n223787 );
nand ( n223789 , n221956 , n217944 );
nand ( n223790 , n223788 , n223789 );
nand ( n223791 , n223790 , n220985 );
nand ( n223792 , n223784 , n223791 );
xor ( n223793 , n223781 , n223792 );
not ( n223794 , n36319 );
not ( n223795 , n34127 );
or ( n223796 , n223794 , n223795 );
nand ( n223797 , n223796 , n37427 );
nand ( n223798 , n32541 , n36326 );
not ( n223799 , n223798 );
not ( n223800 , n223799 );
and ( n223801 , n223797 , n223800 );
not ( n223802 , n223797 );
and ( n223803 , n223802 , n223799 );
nor ( n223804 , n223801 , n223803 );
and ( n223805 , n223153 , n223804 );
not ( n223806 , n223153 );
not ( n223807 , n223804 );
and ( n223808 , n223806 , n223807 );
nor ( n223809 , n223805 , n223808 );
not ( n223810 , n223809 );
not ( n223811 , n223810 );
nor ( n223812 , n223811 , n213751 );
not ( n223813 , n220033 );
not ( n223814 , n220749 );
not ( n223815 , n216307 );
or ( n223816 , n223814 , n223815 );
nand ( n223817 , n41319 , n216277 );
nand ( n223818 , n223816 , n223817 );
not ( n223819 , n223818 );
or ( n223820 , n223813 , n223819 );
nand ( n223821 , n223131 , n220414 );
nand ( n223822 , n223820 , n223821 );
xor ( n223823 , n223812 , n223822 );
not ( n223824 , n223292 );
not ( n223825 , n216204 );
or ( n223826 , n223824 , n223825 );
not ( n223827 , n219687 );
not ( n223828 , n217977 );
or ( n223829 , n223827 , n223828 );
nand ( n223830 , n41069 , n221283 );
nand ( n223831 , n223829 , n223830 );
not ( n223832 , n223831 );
buf ( n223833 , n214793 );
or ( n223834 , n223832 , n223833 );
nand ( n223835 , n223826 , n223834 );
xor ( n223836 , n223823 , n223835 );
xor ( n223837 , n223793 , n223836 );
xor ( n223838 , n223771 , n223837 );
xor ( n223839 , n223572 , n223770 );
and ( n223840 , n223839 , n223837 );
and ( n223841 , n223572 , n223770 );
or ( n223842 , n223840 , n223841 );
xor ( n223843 , n223614 , n223252 );
xor ( n223844 , n223843 , n223678 );
xor ( n223845 , n223614 , n223252 );
and ( n223846 , n223845 , n223678 );
and ( n223847 , n223614 , n223252 );
or ( n223848 , n223846 , n223847 );
xor ( n223849 , n223314 , n223356 );
xor ( n223850 , n223849 , n223421 );
xor ( n223851 , n223314 , n223356 );
and ( n223852 , n223851 , n223421 );
and ( n223853 , n223314 , n223356 );
or ( n223854 , n223852 , n223853 );
xor ( n223855 , n223696 , n223838 );
xor ( n223856 , n223855 , n223729 );
xor ( n223857 , n223696 , n223838 );
and ( n223858 , n223857 , n223729 );
and ( n223859 , n223696 , n223838 );
or ( n223860 , n223858 , n223859 );
xor ( n223861 , n223844 , n223427 );
xor ( n223862 , n223861 , n223433 );
xor ( n223863 , n223844 , n223427 );
and ( n223864 , n223863 , n223433 );
and ( n223865 , n223844 , n223427 );
or ( n223866 , n223864 , n223865 );
xor ( n223867 , n223812 , n223822 );
and ( n223868 , n223867 , n223835 );
and ( n223869 , n223812 , n223822 );
or ( n223870 , n223868 , n223869 );
xor ( n223871 , n223850 , n223439 );
xor ( n223872 , n223871 , n223445 );
xor ( n223873 , n223850 , n223439 );
and ( n223874 , n223873 , n223445 );
and ( n223875 , n223850 , n223439 );
or ( n223876 , n223874 , n223875 );
xor ( n223877 , n223856 , n223862 );
xor ( n223878 , n223877 , n223451 );
xor ( n223879 , n223856 , n223862 );
and ( n223880 , n223879 , n223451 );
and ( n223881 , n223856 , n223862 );
or ( n223882 , n223880 , n223881 );
xor ( n223883 , n223872 , n223878 );
xor ( n223884 , n223883 , n223461 );
xor ( n223885 , n223872 , n223878 );
and ( n223886 , n223885 , n223461 );
and ( n223887 , n223872 , n223878 );
or ( n223888 , n223886 , n223887 );
xor ( n223889 , n223527 , n223662 );
and ( n223890 , n223889 , n223675 );
and ( n223891 , n223527 , n223662 );
or ( n223892 , n223890 , n223891 );
xor ( n223893 , n223629 , n223639 );
and ( n223894 , n223893 , n223650 );
and ( n223895 , n223629 , n223639 );
or ( n223896 , n223894 , n223895 );
xor ( n223897 , n223589 , n223601 );
and ( n223898 , n223897 , n223612 );
and ( n223899 , n223589 , n223601 );
or ( n223900 , n223898 , n223899 );
xor ( n223901 , n223115 , n223693 );
and ( n223902 , n223901 , n223556 );
and ( n223903 , n223115 , n223693 );
or ( n223904 , n223902 , n223903 );
xor ( n223905 , n223162 , n223711 );
and ( n223906 , n223905 , n223726 );
and ( n223907 , n223162 , n223711 );
or ( n223908 , n223906 , n223907 );
xor ( n223909 , n223781 , n223792 );
and ( n223910 , n223909 , n223836 );
and ( n223911 , n223781 , n223792 );
or ( n223912 , n223910 , n223911 );
xor ( n223913 , n223743 , n223755 );
and ( n223914 , n223913 , n223769 );
and ( n223915 , n223743 , n223755 );
or ( n223916 , n223914 , n223915 );
not ( n223917 , n223524 );
not ( n223918 , n220059 );
or ( n223919 , n223917 , n223918 );
and ( n223920 , n221924 , n30962 );
not ( n223921 , n221924 );
and ( n223922 , n223921 , n216530 );
or ( n223923 , n223920 , n223922 );
nand ( n223924 , n223923 , n220067 );
nand ( n223925 , n223919 , n223924 );
not ( n223926 , n216598 );
not ( n223927 , n216542 );
and ( n223928 , n217511 , n223927 );
not ( n223929 , n217511 );
and ( n223930 , n223929 , n41564 );
or ( n223931 , n223928 , n223930 );
not ( n223932 , n223931 );
or ( n223933 , n223926 , n223932 );
nand ( n223934 , n223501 , n218647 );
nand ( n223935 , n223933 , n223934 );
not ( n223936 , n223513 );
not ( n223937 , n217088 );
not ( n223938 , n223937 );
or ( n223939 , n223936 , n223938 );
not ( n223940 , n216928 );
not ( n223941 , n216607 );
or ( n223942 , n223940 , n223941 );
nand ( n223943 , n216608 , n217079 );
nand ( n223944 , n223942 , n223943 );
nand ( n223945 , n223944 , n217885 );
nand ( n223946 , n223939 , n223945 );
xor ( n223947 , n223935 , n223946 );
xor ( n223948 , n223925 , n223947 );
buf ( n223949 , n217047 );
not ( n223950 , n223949 );
not ( n223951 , n216015 );
not ( n223952 , n216500 );
or ( n223953 , n223951 , n223952 );
nand ( n223954 , n41397 , n216404 );
nand ( n223955 , n223953 , n223954 );
not ( n223956 , n223955 );
or ( n223957 , n223950 , n223956 );
nand ( n223958 , n223539 , n216619 );
nand ( n223959 , n223957 , n223958 );
xor ( n223960 , n223948 , n223959 );
xor ( n223961 , n223925 , n223947 );
and ( n223962 , n223961 , n223959 );
and ( n223963 , n223925 , n223947 );
or ( n223964 , n223962 , n223963 );
not ( n223965 , n223182 );
buf ( n223966 , n32549 );
nand ( n223967 , n223966 , n36329 );
not ( n223968 , n223967 );
not ( n223969 , n223968 );
and ( n223970 , n34100 , n32541 );
not ( n223971 , n223970 );
not ( n223972 , n220628 );
or ( n223973 , n223971 , n223972 );
not ( n223974 , n32541 );
not ( n223975 , n33604 );
or ( n223976 , n223974 , n223975 );
nand ( n223977 , n223976 , n36326 );
not ( n223978 , n223977 );
nand ( n223979 , n223973 , n223978 );
not ( n223980 , n223979 );
not ( n223981 , n223980 );
or ( n223982 , n223969 , n223981 );
not ( n223983 , n223970 );
not ( n223984 , n220628 );
or ( n223985 , n223983 , n223984 );
nand ( n223986 , n223985 , n223978 );
nand ( n223987 , n223986 , n223967 );
nand ( n223988 , n223982 , n223987 );
buf ( n223989 , n223988 );
nand ( n223990 , n223965 , n223989 );
buf ( n223991 , n223807 );
and ( n223992 , n223991 , n213750 );
or ( n223993 , n223990 , n223992 );
not ( n223994 , n213750 );
not ( n223995 , n223991 );
nand ( n223996 , n223994 , n223995 , n223989 );
nand ( n223997 , n223993 , n223996 );
not ( n223998 , n221933 );
not ( n223999 , n221935 );
not ( n224000 , n217116 );
or ( n224001 , n223999 , n224000 );
nand ( n224002 , n218137 , n218994 );
nand ( n224003 , n224001 , n224002 );
not ( n224004 , n224003 );
or ( n224005 , n223998 , n224004 );
nand ( n224006 , n223551 , n215183 );
nand ( n224007 , n224005 , n224006 );
xor ( n224008 , n223997 , n224007 );
not ( n224009 , n220033 );
not ( n224010 , n215766 );
not ( n224011 , n41249 );
or ( n224012 , n224010 , n224011 );
nand ( n224013 , n41250 , n220038 );
nand ( n224014 , n224012 , n224013 );
not ( n224015 , n224014 );
or ( n224016 , n224009 , n224015 );
nand ( n224017 , n223818 , n217486 );
nand ( n224018 , n224016 , n224017 );
xor ( n224019 , n224008 , n224018 );
xor ( n224020 , n223997 , n224007 );
and ( n224021 , n224020 , n224018 );
and ( n224022 , n223997 , n224007 );
or ( n224023 , n224021 , n224022 );
not ( n224024 , n219314 );
and ( n224025 , n219687 , n220077 );
not ( n224026 , n219687 );
and ( n224027 , n224026 , n41165 );
or ( n224028 , n224025 , n224027 );
not ( n224029 , n224028 );
or ( n224030 , n224024 , n224029 );
nand ( n224031 , n223831 , n216204 );
nand ( n224032 , n224030 , n224031 );
xor ( n224033 , n224032 , n223531 );
not ( n224034 , n223660 );
not ( n224035 , n218221 );
or ( n224036 , n224034 , n224035 );
buf ( n224037 , n215228 );
not ( n224038 , n224037 );
not ( n224039 , n221214 );
or ( n224040 , n224038 , n224039 );
not ( n224041 , n224037 );
nand ( n224042 , n218208 , n224041 );
nand ( n224043 , n224040 , n224042 );
nand ( n224044 , n224043 , n218232 );
nand ( n224045 , n224036 , n224044 );
xor ( n224046 , n224033 , n224045 );
xor ( n224047 , n223900 , n224046 );
xor ( n224048 , n224047 , n223896 );
xor ( n224049 , n223900 , n224046 );
and ( n224050 , n224049 , n223896 );
and ( n224051 , n223900 , n224046 );
or ( n224052 , n224050 , n224051 );
xor ( n224053 , n223892 , n223904 );
not ( n224054 , n223599 );
not ( n224055 , n223591 );
or ( n224056 , n224054 , n224055 );
and ( n224057 , n213583 , n223186 );
not ( n224058 , n213583 );
not ( n224059 , n223156 );
and ( n224060 , n224058 , n224059 );
or ( n224061 , n224057 , n224060 );
nand ( n224062 , n222769 , n224061 );
nand ( n224063 , n224056 , n224062 );
and ( n224064 , n223979 , n223968 );
not ( n224065 , n223979 );
and ( n224066 , n224065 , n223967 );
nor ( n224067 , n224064 , n224066 );
buf ( n224068 , n224067 );
not ( n224069 , n224068 );
and ( n224070 , n213751 , n224069 );
not ( n224071 , n213751 );
and ( n224072 , n224071 , n223989 );
nor ( n224073 , n224070 , n224072 );
not ( n224074 , n224073 );
not ( n224075 , n223968 );
not ( n224076 , n223980 );
or ( n224077 , n224075 , n224076 );
nand ( n224078 , n224077 , n223987 );
not ( n224079 , n223804 );
and ( n224080 , n224078 , n224079 );
not ( n224081 , n224078 );
not ( n224082 , n224079 );
and ( n224083 , n224081 , n224082 );
nor ( n224084 , n224080 , n224083 );
and ( n224085 , n224084 , n223809 );
buf ( n224086 , n224085 );
buf ( n224087 , n224086 );
not ( n224088 , n224087 );
or ( n224089 , n224074 , n224088 );
buf ( n224090 , n223810 );
not ( n224091 , n218224 );
not ( n224092 , n224069 );
or ( n224093 , n224091 , n224092 );
not ( n224094 , n224078 );
buf ( n224095 , n224094 );
not ( n224096 , n224095 );
nand ( n224097 , n224096 , n216076 );
nand ( n224098 , n224093 , n224097 );
nand ( n224099 , n224090 , n224098 );
nand ( n224100 , n224089 , n224099 );
xor ( n224101 , n224063 , n224100 );
xor ( n224102 , n224101 , n223960 );
xor ( n224103 , n224053 , n224102 );
xor ( n224104 , n223892 , n223904 );
and ( n224105 , n224104 , n224102 );
and ( n224106 , n223892 , n223904 );
or ( n224107 , n224105 , n224106 );
not ( n224108 , n223637 );
not ( n224109 , n220919 );
or ( n224110 , n224108 , n224109 );
not ( n224111 , n215075 );
not ( n224112 , n220900 );
not ( n224113 , n224112 );
or ( n224114 , n224111 , n224113 );
nand ( n224115 , n220900 , n215899 );
nand ( n224116 , n224114 , n224115 );
nand ( n224117 , n224116 , n221674 );
nand ( n224118 , n224110 , n224117 );
not ( n224119 , n223586 );
not ( n224120 , n221624 );
not ( n224121 , n224120 );
or ( n224122 , n224119 , n224121 );
not ( n224123 , n216964 );
not ( n224124 , n221612 );
or ( n224125 , n224123 , n224124 );
nand ( n224126 , n223584 , n214678 );
nand ( n224127 , n224125 , n224126 );
nand ( n224128 , n224127 , n223177 );
nand ( n224129 , n224122 , n224128 );
xor ( n224130 , n224118 , n224129 );
not ( n224131 , n223610 );
not ( n224132 , n222886 );
or ( n224133 , n224131 , n224132 );
not ( n224134 , n217044 );
not ( n224135 , n222429 );
or ( n224136 , n224134 , n224135 );
nand ( n224137 , n222462 , n215131 );
nand ( n224138 , n224136 , n224137 );
nand ( n224139 , n224138 , n222158 );
nand ( n224140 , n224133 , n224139 );
xor ( n224141 , n224130 , n224140 );
not ( n224142 , n223673 );
not ( n224143 , n220853 );
or ( n224144 , n224142 , n224143 );
not ( n224145 , n221495 );
not ( n224146 , n218876 );
or ( n224147 , n224145 , n224146 );
nand ( n224148 , n218815 , n221494 );
nand ( n224149 , n224147 , n224148 );
nand ( n224150 , n218843 , n224149 );
nand ( n224151 , n224144 , n224150 );
not ( n224152 , n223627 );
not ( n224153 , n219435 );
or ( n224154 , n224152 , n224153 );
not ( n224155 , n219343 );
not ( n224156 , n219420 );
or ( n224157 , n224155 , n224156 );
nand ( n224158 , n220180 , n223269 );
nand ( n224159 , n224157 , n224158 );
nand ( n224160 , n224159 , n219076 );
nand ( n224161 , n224154 , n224160 );
xor ( n224162 , n224151 , n224161 );
not ( n224163 , n220492 );
not ( n224164 , n223648 );
or ( n224165 , n224163 , n224164 );
and ( n224166 , n216940 , n220150 );
not ( n224167 , n216940 );
and ( n224168 , n224167 , n221257 );
nor ( n224169 , n224166 , n224168 );
buf ( n224170 , n220160 );
buf ( n224171 , n224170 );
or ( n224172 , n224169 , n224171 );
nand ( n224173 , n224165 , n224172 );
xor ( n224174 , n224162 , n224173 );
xor ( n224175 , n224141 , n224174 );
xor ( n224176 , n224175 , n223908 );
xor ( n224177 , n224141 , n224174 );
and ( n224178 , n224177 , n223908 );
and ( n224179 , n224141 , n224174 );
or ( n224180 , n224178 , n224179 );
xor ( n224181 , n223560 , n223870 );
not ( n224182 , n220272 );
not ( n224183 , n215955 );
not ( n224184 , n219532 );
or ( n224185 , n224183 , n224184 );
nand ( n224186 , n220203 , n219358 );
nand ( n224187 , n224185 , n224186 );
not ( n224188 , n224187 );
or ( n224189 , n224182 , n224188 );
nand ( n224190 , n223706 , n220280 );
nand ( n224191 , n224189 , n224190 );
xor ( n224192 , n224181 , n224191 );
xor ( n224193 , n223912 , n224192 );
xor ( n224194 , n224193 , n223916 );
xor ( n224195 , n223912 , n224192 );
and ( n224196 , n224195 , n223916 );
and ( n224197 , n223912 , n224192 );
or ( n224198 , n224196 , n224197 );
not ( n224199 , n215137 );
not ( n224200 , n217573 );
not ( n224201 , n40181 );
or ( n224202 , n224200 , n224201 );
nand ( n224203 , n223320 , n219390 );
nand ( n224204 , n224202 , n224203 );
not ( n224205 , n224204 );
or ( n224206 , n224199 , n224205 );
nand ( n224207 , n223779 , n215605 );
nand ( n224208 , n224206 , n224207 );
not ( n224209 , n222185 );
not ( n224210 , n219033 );
not ( n224211 , n218268 );
or ( n224212 , n224210 , n224211 );
nand ( n224213 , n219594 , n219034 );
nand ( n224214 , n224212 , n224213 );
not ( n224215 , n224214 );
or ( n224216 , n224209 , n224215 );
nand ( n224217 , n223689 , n219731 );
nand ( n224218 , n224216 , n224217 );
xor ( n224219 , n224208 , n224218 );
not ( n224220 , n220985 );
not ( n224221 , n215113 );
not ( n224222 , n40258 );
or ( n224223 , n224221 , n224222 );
nand ( n224224 , n220970 , n216037 );
nand ( n224225 , n224223 , n224224 );
not ( n224226 , n224225 );
or ( n224227 , n224220 , n224226 );
nand ( n224228 , n223790 , n214717 );
nand ( n224229 , n224227 , n224228 );
xor ( n224230 , n224219 , n224229 );
not ( n224231 , n220820 );
not ( n224232 , n216810 );
not ( n224233 , n221028 );
or ( n224234 , n224232 , n224233 );
nand ( n224235 , n40668 , n215289 );
nand ( n224236 , n224234 , n224235 );
not ( n224237 , n224236 );
or ( n224238 , n224231 , n224237 );
nand ( n224239 , n223741 , n216562 );
nand ( n224240 , n224238 , n224239 );
not ( n224241 , n216336 );
not ( n224242 , n213735 );
not ( n224243 , n223368 );
or ( n224244 , n224242 , n224243 );
nand ( n224245 , n222513 , n213732 );
nand ( n224246 , n224244 , n224245 );
not ( n224247 , n224246 );
or ( n224248 , n224241 , n224247 );
nand ( n224249 , n223753 , n213577 );
nand ( n224250 , n224248 , n224249 );
xor ( n224251 , n224240 , n224250 );
not ( n224252 , n219175 );
not ( n224253 , n219577 );
not ( n224254 , n219521 );
or ( n224255 , n224253 , n224254 );
nand ( n224256 , n40625 , n218661 );
nand ( n224257 , n224255 , n224256 );
not ( n224258 , n224257 );
or ( n224259 , n224252 , n224258 );
nand ( n224260 , n223568 , n217023 );
nand ( n224261 , n224259 , n224260 );
xor ( n224262 , n224251 , n224261 );
xor ( n224263 , n224230 , n224262 );
xor ( n224264 , n224263 , n223576 );
xor ( n224265 , n224230 , n224262 );
and ( n224266 , n224265 , n223576 );
and ( n224267 , n224230 , n224262 );
or ( n224268 , n224266 , n224267 );
not ( n224269 , n217969 );
not ( n224270 , n223767 );
or ( n224271 , n224269 , n224270 );
not ( n224272 , n39995 );
and ( n224273 , n224272 , n213381 );
not ( n224274 , n224272 );
and ( n224275 , n224274 , n213382 );
nor ( n224276 , n224273 , n224275 );
nand ( n224277 , n224276 , n213912 );
nand ( n224278 , n224271 , n224277 );
not ( n224279 , n213874 );
not ( n224280 , n223724 );
or ( n224281 , n224279 , n224280 );
not ( n224282 , n216262 );
not ( n224283 , n223330 );
or ( n224284 , n224282 , n224283 );
not ( n224285 , n40545 );
not ( n224286 , n224285 );
nand ( n224287 , n224286 , n220300 );
nand ( n224288 , n224284 , n224287 );
nand ( n224289 , n224288 , n217142 );
nand ( n224290 , n224281 , n224289 );
xor ( n224291 , n224278 , n224290 );
xor ( n224292 , n224291 , n224019 );
xor ( n224293 , n224292 , n223618 );
xor ( n224294 , n224293 , n224048 );
xor ( n224295 , n224292 , n223618 );
and ( n224296 , n224295 , n224048 );
and ( n224297 , n224292 , n223618 );
or ( n224298 , n224296 , n224297 );
xor ( n224299 , n223682 , n223700 );
xor ( n224300 , n224299 , n224176 );
xor ( n224301 , n223682 , n223700 );
and ( n224302 , n224301 , n224176 );
and ( n224303 , n223682 , n223700 );
or ( n224304 , n224302 , n224303 );
xor ( n224305 , n224103 , n223733 );
xor ( n224306 , n224305 , n223842 );
xor ( n224307 , n224103 , n223733 );
and ( n224308 , n224307 , n223842 );
and ( n224309 , n224103 , n223733 );
or ( n224310 , n224308 , n224309 );
xor ( n224311 , n224194 , n224264 );
xor ( n224312 , n224311 , n223848 );
xor ( n224313 , n224194 , n224264 );
and ( n224314 , n224313 , n223848 );
and ( n224315 , n224194 , n224264 );
or ( n224316 , n224314 , n224315 );
xor ( n224317 , n224294 , n224300 );
xor ( n224318 , n224317 , n223854 );
xor ( n224319 , n224294 , n224300 );
and ( n224320 , n224319 , n223854 );
and ( n224321 , n224294 , n224300 );
or ( n224322 , n224320 , n224321 );
xor ( n224323 , n224032 , n223531 );
and ( n224324 , n224323 , n224045 );
and ( n224325 , n224032 , n223531 );
or ( n224326 , n224324 , n224325 );
xor ( n224327 , n223860 , n224306 );
xor ( n224328 , n224327 , n224312 );
xor ( n224329 , n223860 , n224306 );
and ( n224330 , n224329 , n224312 );
and ( n224331 , n223860 , n224306 );
or ( n224332 , n224330 , n224331 );
xor ( n224333 , n223866 , n224318 );
xor ( n224334 , n224333 , n223876 );
xor ( n224335 , n223866 , n224318 );
and ( n224336 , n224335 , n223876 );
and ( n224337 , n223866 , n224318 );
or ( n224338 , n224336 , n224337 );
xor ( n224339 , n224328 , n223882 );
xor ( n224340 , n224339 , n224334 );
xor ( n224341 , n224328 , n223882 );
and ( n224342 , n224341 , n224334 );
and ( n224343 , n224328 , n223882 );
or ( n224344 , n224342 , n224343 );
xor ( n224345 , n224151 , n224161 );
and ( n224346 , n224345 , n224173 );
and ( n224347 , n224151 , n224161 );
or ( n224348 , n224346 , n224347 );
xor ( n224349 , n224118 , n224129 );
and ( n224350 , n224349 , n224140 );
and ( n224351 , n224118 , n224129 );
or ( n224352 , n224350 , n224351 );
xor ( n224353 , n224063 , n224100 );
and ( n224354 , n224353 , n223960 );
and ( n224355 , n224063 , n224100 );
or ( n224356 , n224354 , n224355 );
xor ( n224357 , n223560 , n223870 );
and ( n224358 , n224357 , n224191 );
and ( n224359 , n223560 , n223870 );
or ( n224360 , n224358 , n224359 );
xor ( n224361 , n224208 , n224218 );
and ( n224362 , n224361 , n224229 );
and ( n224363 , n224208 , n224218 );
or ( n224364 , n224362 , n224363 );
xor ( n224365 , n224278 , n224290 );
and ( n224366 , n224365 , n224019 );
and ( n224367 , n224278 , n224290 );
or ( n224368 , n224366 , n224367 );
xor ( n224369 , n224240 , n224250 );
and ( n224370 , n224369 , n224261 );
and ( n224371 , n224240 , n224250 );
or ( n224372 , n224370 , n224371 );
not ( n224373 , n223944 );
not ( n224374 , n217089 );
or ( n224375 , n224373 , n224374 );
not ( n224376 , n217080 );
not ( n224377 , n216339 );
or ( n224378 , n224376 , n224377 );
nand ( n224379 , n41701 , n217602 );
nand ( n224380 , n224378 , n224379 );
nand ( n224381 , n224380 , n219119 );
nand ( n224382 , n224375 , n224381 );
not ( n224383 , n223923 );
not ( n224384 , n217631 );
or ( n224385 , n224383 , n224384 );
not ( n224386 , n219689 );
not ( n224387 , n217611 );
or ( n224388 , n224386 , n224387 );
or ( n224389 , n219689 , n217473 );
nand ( n224390 , n224388 , n224389 );
nand ( n224391 , n224390 , n218762 );
nand ( n224392 , n224385 , n224391 );
xor ( n224393 , n224382 , n224392 );
not ( n224394 , n219501 );
not ( n224395 , n216762 );
not ( n224396 , n216261 );
or ( n224397 , n224395 , n224396 );
not ( n224398 , n216422 );
nand ( n224399 , n215796 , n224398 );
nand ( n224400 , n224397 , n224399 );
not ( n224401 , n224400 );
or ( n224402 , n224394 , n224401 );
nand ( n224403 , n223931 , n216586 );
nand ( n224404 , n224402 , n224403 );
xor ( n224405 , n224393 , n224404 );
xor ( n224406 , n224382 , n224392 );
and ( n224407 , n224406 , n224404 );
and ( n224408 , n224382 , n224392 );
or ( n224409 , n224407 , n224408 );
not ( n224410 , n223513 );
not ( n224411 , n223937 );
or ( n224412 , n224410 , n224411 );
nand ( n224413 , n224412 , n223945 );
and ( n224414 , n223935 , n224413 );
not ( n224415 , n217047 );
and ( n224416 , n216015 , n216307 );
not ( n224417 , n216015 );
and ( n224418 , n224417 , n216306 );
or ( n224419 , n224416 , n224418 );
not ( n224420 , n224419 );
or ( n224421 , n224415 , n224420 );
not ( n224422 , n216066 );
nand ( n224423 , n224422 , n223955 );
nand ( n224424 , n224421 , n224423 );
xor ( n224425 , n224414 , n224424 );
not ( n224426 , n224067 );
not ( n224427 , n36413 );
not ( n224428 , n224427 );
not ( n224429 , n34127 );
nor ( n224430 , n224429 , n37563 );
not ( n224431 , n224430 );
or ( n224432 , n224428 , n224431 );
and ( n224433 , n36380 , n37629 );
nor ( n224434 , n224433 , n36330 );
nand ( n224435 , n224432 , n224434 );
nand ( n224436 , n37581 , n32723 );
not ( n224437 , n224436 );
not ( n224438 , n224437 );
and ( n224439 , n224435 , n224438 );
not ( n224440 , n224435 );
and ( n224441 , n224440 , n224437 );
nor ( n224442 , n224439 , n224441 );
and ( n224443 , n224426 , n224442 );
not ( n224444 , n224426 );
not ( n224445 , n224442 );
and ( n224446 , n224444 , n224445 );
nor ( n224447 , n224443 , n224446 );
not ( n224448 , n224447 );
not ( n224449 , n224448 );
and ( n224450 , n224449 , n215999 );
xor ( n224451 , n224425 , n224450 );
xor ( n224452 , n224414 , n224424 );
and ( n224453 , n224452 , n224450 );
and ( n224454 , n224414 , n224424 );
or ( n224455 , n224453 , n224454 );
not ( n224456 , n211314 );
not ( n224457 , n213382 );
not ( n224458 , n39877 );
or ( n224459 , n224457 , n224458 );
nand ( n224460 , n39878 , n213381 );
nand ( n224461 , n224459 , n224460 );
not ( n224462 , n224461 );
or ( n224463 , n224456 , n224462 );
nand ( n224464 , n224276 , n217969 );
nand ( n224465 , n224463 , n224464 );
xor ( n224466 , n224465 , n224352 );
not ( n224467 , n221933 );
not ( n224468 , n221935 );
not ( n224469 , n217330 );
or ( n224470 , n224468 , n224469 );
nand ( n224471 , n41071 , n222333 );
nand ( n224472 , n224470 , n224471 );
not ( n224473 , n224472 );
or ( n224474 , n224467 , n224473 );
nand ( n224475 , n224003 , n219332 );
nand ( n224476 , n224474 , n224475 );
not ( n224477 , n220414 );
not ( n224478 , n224014 );
or ( n224479 , n224477 , n224478 );
not ( n224480 , n215766 );
not ( n224481 , n217317 );
or ( n224482 , n224480 , n224481 );
not ( n224483 , n216281 );
nand ( n224484 , n208164 , n224483 );
nand ( n224485 , n224482 , n224484 );
nand ( n224486 , n224485 , n220033 );
nand ( n224487 , n224479 , n224486 );
xor ( n224488 , n224476 , n224487 );
not ( n224489 , n224043 );
not ( n224490 , n218221 );
or ( n224491 , n224489 , n224490 );
not ( n224492 , n214642 );
not ( n224493 , n224492 );
not ( n224494 , n220091 );
or ( n224495 , n224493 , n224494 );
not ( n224496 , n224492 );
not ( n224497 , n218256 );
nand ( n224498 , n224496 , n224497 );
nand ( n224499 , n224495 , n224498 );
nand ( n224500 , n224499 , n218232 );
nand ( n224501 , n224491 , n224500 );
xor ( n224502 , n224488 , n224501 );
xor ( n224503 , n224466 , n224502 );
xor ( n224504 , n224465 , n224352 );
and ( n224505 , n224504 , n224502 );
and ( n224506 , n224465 , n224352 );
or ( n224507 , n224505 , n224506 );
xor ( n224508 , n224326 , n224348 );
xor ( n224509 , n224508 , n224356 );
xor ( n224510 , n224326 , n224348 );
and ( n224511 , n224510 , n224356 );
and ( n224512 , n224326 , n224348 );
or ( n224513 , n224511 , n224512 );
not ( n224514 , n224061 );
not ( n224515 , n223591 );
or ( n224516 , n224514 , n224515 );
not ( n224517 , n214956 );
not ( n224518 , n223203 );
or ( n224519 , n224517 , n224518 );
nand ( n224520 , n223202 , n214960 );
nand ( n224521 , n224519 , n224520 );
nand ( n224522 , n224521 , n222769 );
nand ( n224523 , n224516 , n224522 );
xor ( n224524 , n224523 , n224405 );
not ( n224525 , n224098 );
not ( n224526 , n224087 );
or ( n224527 , n224525 , n224526 );
not ( n224528 , n213347 );
not ( n224529 , n224095 );
or ( n224530 , n224528 , n224529 );
nand ( n224531 , n224068 , n214616 );
nand ( n224532 , n224530 , n224531 );
nand ( n224533 , n224090 , n224532 );
nand ( n224534 , n224527 , n224533 );
xor ( n224535 , n224524 , n224534 );
not ( n224536 , n224149 );
not ( n224537 , n220480 );
or ( n224538 , n224536 , n224537 );
not ( n224539 , n216293 );
not ( n224540 , n218814 );
or ( n224541 , n224539 , n224540 );
nand ( n224542 , n218815 , n223658 );
nand ( n224543 , n224541 , n224542 );
nand ( n224544 , n222376 , n224543 );
nand ( n224545 , n224538 , n224544 );
not ( n224546 , n224159 );
not ( n224547 , n221576 );
or ( n224548 , n224546 , n224547 );
not ( n224549 , n221921 );
not ( n224550 , n219440 );
or ( n224551 , n224549 , n224550 );
nand ( n224552 , n221228 , n218980 );
nand ( n224553 , n224551 , n224552 );
nand ( n224554 , n224553 , n219076 );
nand ( n224555 , n224548 , n224554 );
xor ( n224556 , n224545 , n224555 );
not ( n224557 , n224169 );
not ( n224558 , n224557 );
not ( n224559 , n220164 );
or ( n224560 , n224558 , n224559 );
not ( n224561 , n219102 );
not ( n224562 , n220146 );
buf ( n224563 , n224562 );
not ( n224564 , n224563 );
or ( n224565 , n224561 , n224564 );
nand ( n224566 , n222791 , n216139 );
nand ( n224567 , n224565 , n224566 );
nand ( n224568 , n219779 , n224567 );
nand ( n224569 , n224560 , n224568 );
xor ( n224570 , n224556 , n224569 );
xor ( n224571 , n224535 , n224570 );
not ( n224572 , n224116 );
not ( n224573 , n220919 );
or ( n224574 , n224572 , n224573 );
not ( n224575 , n218514 );
not ( n224576 , n223227 );
or ( n224577 , n224575 , n224576 );
nand ( n224578 , n220900 , n216170 );
nand ( n224579 , n224577 , n224578 );
nand ( n224580 , n224579 , n220636 );
nand ( n224581 , n224574 , n224580 );
not ( n224582 , n224127 );
not ( n224583 , n224120 );
or ( n224584 , n224582 , n224583 );
not ( n224585 , n216208 );
not ( n224586 , n222586 );
or ( n224587 , n224585 , n224586 );
nand ( n224588 , n221607 , n216207 );
nand ( n224589 , n224587 , n224588 );
nand ( n224590 , n224589 , n221387 );
nand ( n224591 , n224584 , n224590 );
xor ( n224592 , n224581 , n224591 );
not ( n224593 , n224138 );
not ( n224594 , n222454 );
or ( n224595 , n224593 , n224594 );
not ( n224596 , n214537 );
not ( n224597 , n222429 );
or ( n224598 , n224596 , n224597 );
nand ( n224599 , n222433 , n214899 );
nand ( n224600 , n224598 , n224599 );
nand ( n224601 , n223244 , n224600 );
nand ( n224602 , n224595 , n224601 );
xor ( n224603 , n224592 , n224602 );
xor ( n224604 , n224571 , n224603 );
xor ( n224605 , n224535 , n224570 );
and ( n224606 , n224605 , n224603 );
and ( n224607 , n224535 , n224570 );
or ( n224608 , n224606 , n224607 );
xor ( n224609 , n224360 , n224372 );
xor ( n224610 , n224609 , n224368 );
xor ( n224611 , n224360 , n224372 );
and ( n224612 , n224611 , n224368 );
and ( n224613 , n224360 , n224372 );
or ( n224614 , n224612 , n224613 );
not ( n224615 , n219314 );
not ( n224616 , n219687 );
not ( n224617 , n40724 );
not ( n224618 , n224617 );
or ( n224619 , n224616 , n224618 );
nand ( n224620 , n40724 , n221283 );
nand ( n224621 , n224619 , n224620 );
not ( n224622 , n224621 );
or ( n224623 , n224615 , n224622 );
not ( n224624 , n223825 );
nand ( n224625 , n224028 , n224624 );
nand ( n224626 , n224623 , n224625 );
xor ( n224627 , n224626 , n223964 );
xor ( n224628 , n224627 , n224023 );
xor ( n224629 , n224628 , n224364 );
not ( n224630 , n220280 );
not ( n224631 , n224187 );
or ( n224632 , n224630 , n224631 );
and ( n224633 , n215955 , n219226 );
not ( n224634 , n215955 );
and ( n224635 , n224634 , n219223 );
nor ( n224636 , n224633 , n224635 );
nand ( n224637 , n224636 , n219353 );
nand ( n224638 , n224632 , n224637 );
not ( n224639 , n222185 );
and ( n224640 , n219033 , n221342 );
not ( n224641 , n219033 );
not ( n224642 , n219238 );
not ( n224643 , n224642 );
and ( n224644 , n224641 , n224643 );
nor ( n224645 , n224640 , n224644 );
not ( n224646 , n224645 );
or ( n224647 , n224639 , n224646 );
nand ( n224648 , n224214 , n219731 );
nand ( n224649 , n224647 , n224648 );
xor ( n224650 , n224638 , n224649 );
not ( n224651 , n214717 );
not ( n224652 , n224225 );
or ( n224653 , n224651 , n224652 );
not ( n224654 , n218855 );
not ( n224655 , n222121 );
or ( n224656 , n224654 , n224655 );
nand ( n224657 , n40397 , n216037 );
nand ( n224658 , n224656 , n224657 );
nand ( n224659 , n224658 , n220985 );
nand ( n224660 , n224653 , n224659 );
xor ( n224661 , n224650 , n224660 );
xor ( n224662 , n224629 , n224661 );
xor ( n224663 , n224628 , n224364 );
and ( n224664 , n224663 , n224661 );
and ( n224665 , n224628 , n224364 );
or ( n224666 , n224664 , n224665 );
not ( n224667 , n213577 );
not ( n224668 , n224246 );
or ( n224669 , n224667 , n224668 );
not ( n224670 , n213735 );
not ( n224671 , n222940 );
or ( n224672 , n224670 , n224671 );
nand ( n224673 , n223722 , n213732 );
nand ( n224674 , n224672 , n224673 );
nand ( n224675 , n224674 , n216336 );
nand ( n224676 , n224669 , n224675 );
xor ( n224677 , n224451 , n224676 );
not ( n224678 , n217023 );
not ( n224679 , n224257 );
or ( n224680 , n224678 , n224679 );
not ( n224681 , n219577 );
not ( n224682 , n220581 );
or ( n224683 , n224681 , n224682 );
nand ( n224684 , n207936 , n218661 );
nand ( n224685 , n224683 , n224684 );
nand ( n224686 , n224685 , n219175 );
nand ( n224687 , n224680 , n224686 );
xor ( n224688 , n224677 , n224687 );
xor ( n224689 , n224688 , n224052 );
not ( n224690 , n217142 );
nand ( n224691 , n223765 , n214824 );
nand ( n224692 , n214818 , n223764 );
nand ( n224693 , n224691 , n224692 );
not ( n224694 , n224693 );
or ( n224695 , n224690 , n224694 );
nand ( n224696 , n224288 , n213874 );
nand ( n224697 , n224695 , n224696 );
not ( n224698 , n215137 );
not ( n224699 , n217573 );
not ( n224700 , n222101 );
not ( n224701 , n224700 );
or ( n224702 , n224699 , n224701 );
nand ( n224703 , n40422 , n217397 );
nand ( n224704 , n224702 , n224703 );
not ( n224705 , n224704 );
or ( n224706 , n224698 , n224705 );
nand ( n224707 , n224204 , n214086 );
nand ( n224708 , n224706 , n224707 );
xor ( n224709 , n224697 , n224708 );
not ( n224710 , n216810 );
not ( n224711 , n221330 );
or ( n224712 , n224710 , n224711 );
nand ( n224713 , n40410 , n221307 );
nand ( n224714 , n224712 , n224713 );
not ( n224715 , n224714 );
not ( n224716 , n220820 );
or ( n224717 , n224715 , n224716 );
not ( n224718 , n224236 );
or ( n224719 , n224718 , n216298 );
nand ( n224720 , n224717 , n224719 );
xor ( n224721 , n224709 , n224720 );
xor ( n224722 , n224689 , n224721 );
xor ( n224723 , n224688 , n224052 );
and ( n224724 , n224723 , n224721 );
and ( n224725 , n224688 , n224052 );
or ( n224726 , n224724 , n224725 );
xor ( n224727 , n224503 , n224509 );
xor ( n224728 , n224727 , n224107 );
xor ( n224729 , n224503 , n224509 );
and ( n224730 , n224729 , n224107 );
and ( n224731 , n224503 , n224509 );
or ( n224732 , n224730 , n224731 );
xor ( n224733 , n224604 , n224180 );
xor ( n224734 , n224733 , n224198 );
xor ( n224735 , n224604 , n224180 );
and ( n224736 , n224735 , n224198 );
and ( n224737 , n224604 , n224180 );
or ( n224738 , n224736 , n224737 );
xor ( n224739 , n224610 , n224268 );
xor ( n224740 , n224739 , n224662 );
xor ( n224741 , n224610 , n224268 );
and ( n224742 , n224741 , n224662 );
and ( n224743 , n224610 , n224268 );
or ( n224744 , n224742 , n224743 );
xor ( n224745 , n224722 , n224298 );
xor ( n224746 , n224745 , n224728 );
xor ( n224747 , n224722 , n224298 );
and ( n224748 , n224747 , n224728 );
and ( n224749 , n224722 , n224298 );
or ( n224750 , n224748 , n224749 );
xor ( n224751 , n224476 , n224487 );
and ( n224752 , n224751 , n224501 );
and ( n224753 , n224476 , n224487 );
or ( n224754 , n224752 , n224753 );
xor ( n224755 , n224304 , n224734 );
xor ( n224756 , n224755 , n224310 );
xor ( n224757 , n224304 , n224734 );
and ( n224758 , n224757 , n224310 );
and ( n224759 , n224304 , n224734 );
or ( n224760 , n224758 , n224759 );
xor ( n224761 , n224740 , n224746 );
xor ( n224762 , n224761 , n224316 );
xor ( n224763 , n224740 , n224746 );
and ( n224764 , n224763 , n224316 );
and ( n224765 , n224740 , n224746 );
or ( n224766 , n224764 , n224765 );
xor ( n224767 , n224322 , n224756 );
xor ( n224768 , n224767 , n224332 );
xor ( n224769 , n224322 , n224756 );
and ( n224770 , n224769 , n224332 );
and ( n224771 , n224322 , n224756 );
or ( n224772 , n224770 , n224771 );
xor ( n224773 , n224762 , n224768 );
xor ( n224774 , n224773 , n224338 );
xor ( n224775 , n224762 , n224768 );
and ( n224776 , n224775 , n224338 );
and ( n224777 , n224762 , n224768 );
or ( n224778 , n224776 , n224777 );
xor ( n224779 , n224545 , n224555 );
and ( n224780 , n224779 , n224569 );
and ( n224781 , n224545 , n224555 );
or ( n224782 , n224780 , n224781 );
xor ( n224783 , n224581 , n224591 );
and ( n224784 , n224783 , n224602 );
and ( n224785 , n224581 , n224591 );
or ( n224786 , n224784 , n224785 );
xor ( n224787 , n224523 , n224405 );
and ( n224788 , n224787 , n224534 );
and ( n224789 , n224523 , n224405 );
or ( n224790 , n224788 , n224789 );
xor ( n224791 , n224626 , n223964 );
and ( n224792 , n224791 , n224023 );
and ( n224793 , n224626 , n223964 );
or ( n224794 , n224792 , n224793 );
xor ( n224795 , n224638 , n224649 );
and ( n224796 , n224795 , n224660 );
and ( n224797 , n224638 , n224649 );
or ( n224798 , n224796 , n224797 );
xor ( n224799 , n224697 , n224708 );
and ( n224800 , n224799 , n224720 );
and ( n224801 , n224697 , n224708 );
or ( n224802 , n224800 , n224801 );
xor ( n224803 , n224451 , n224676 );
and ( n224804 , n224803 , n224687 );
and ( n224805 , n224451 , n224676 );
or ( n224806 , n224804 , n224805 );
not ( n224807 , n220033 );
not ( n224808 , n215766 );
not ( n224809 , n217119 );
or ( n224810 , n224808 , n224809 );
nand ( n224811 , n220226 , n224483 );
nand ( n224812 , n224810 , n224811 );
not ( n224813 , n224812 );
or ( n224814 , n224807 , n224813 );
nand ( n224815 , n224485 , n217486 );
nand ( n224816 , n224814 , n224815 );
and ( n224817 , n224435 , n224437 );
not ( n224818 , n224435 );
and ( n224819 , n224818 , n224436 );
nor ( n224820 , n224817 , n224819 );
not ( n224821 , n224820 );
nand ( n224822 , n224821 , n213751 );
not ( n224823 , n213750 );
not ( n224824 , n224820 );
or ( n224825 , n224823 , n224824 );
nand ( n224826 , n224825 , n224095 );
and ( n224827 , n224822 , n224826 );
not ( n224828 , n37564 );
not ( n224829 , n34102 );
or ( n224830 , n224828 , n224829 );
and ( n224831 , n37565 , n219064 );
nor ( n224832 , n224831 , n37582 );
nand ( n224833 , n224830 , n224832 );
not ( n224834 , n36336 );
nand ( n224835 , n224834 , n32805 );
not ( n224836 , n224835 );
and ( n224837 , n224833 , n224836 );
not ( n224838 , n224833 );
and ( n224839 , n224838 , n224835 );
nor ( n224840 , n224837 , n224839 );
not ( n224841 , n224840 );
not ( n224842 , n224841 );
buf ( n224843 , n224842 );
not ( n224844 , n224843 );
nor ( n224845 , n224827 , n224844 );
xor ( n224846 , n224816 , n224845 );
not ( n224847 , n224390 );
not ( n224848 , n217631 );
or ( n224849 , n224847 , n224848 );
not ( n224850 , n217473 );
not ( n224851 , n224850 );
not ( n224852 , n216607 );
or ( n224853 , n224851 , n224852 );
nand ( n224854 , n216608 , n217473 );
nand ( n224855 , n224853 , n224854 );
nand ( n224856 , n224855 , n217641 );
nand ( n224857 , n224849 , n224856 );
not ( n224858 , n224380 );
not ( n224859 , n219367 );
or ( n224860 , n224858 , n224859 );
not ( n224861 , n215616 );
not ( n224862 , n217602 );
and ( n224863 , n224861 , n224862 );
not ( n224864 , n221520 );
and ( n224865 , n224864 , n217079 );
nor ( n224866 , n224863 , n224865 );
not ( n224867 , n224866 );
nand ( n224868 , n224867 , n217885 );
nand ( n224869 , n224860 , n224868 );
xor ( n224870 , n224857 , n224869 );
xor ( n224871 , n224846 , n224870 );
xor ( n224872 , n224816 , n224845 );
and ( n224873 , n224872 , n224870 );
and ( n224874 , n224816 , n224845 );
or ( n224875 , n224873 , n224874 );
not ( n224876 , n216619 );
not ( n224877 , n224419 );
or ( n224878 , n224876 , n224877 );
and ( n224879 , n223537 , n41249 );
not ( n224880 , n223537 );
not ( n224881 , n41249 );
and ( n224882 , n224880 , n224881 );
or ( n224883 , n224879 , n224882 );
not ( n224884 , n224883 );
nand ( n224885 , n224884 , n223949 );
nand ( n224886 , n224878 , n224885 );
not ( n224887 , n216598 );
not ( n224888 , n216422 );
not ( n224889 , n217130 );
or ( n224890 , n224888 , n224889 );
nand ( n224891 , n219582 , n224398 );
nand ( n224892 , n224890 , n224891 );
not ( n224893 , n224892 );
or ( n224894 , n224887 , n224893 );
buf ( n224895 , n216585 );
not ( n224896 , n224895 );
nand ( n224897 , n224400 , n224896 );
nand ( n224898 , n224894 , n224897 );
xor ( n224899 , n224886 , n224898 );
not ( n224900 , n221933 );
not ( n224901 , n221935 );
not ( n224902 , n217710 );
or ( n224903 , n224901 , n224902 );
nand ( n224904 , n217714 , n218994 );
nand ( n224905 , n224903 , n224904 );
not ( n224906 , n224905 );
or ( n224907 , n224900 , n224906 );
nand ( n224908 , n224472 , n215183 );
nand ( n224909 , n224907 , n224908 );
xor ( n224910 , n224899 , n224909 );
xor ( n224911 , n224886 , n224898 );
and ( n224912 , n224911 , n224909 );
and ( n224913 , n224886 , n224898 );
or ( n224914 , n224912 , n224913 );
xor ( n224915 , n224786 , n224790 );
xor ( n224916 , n224915 , n224754 );
xor ( n224917 , n224786 , n224790 );
and ( n224918 , n224917 , n224754 );
and ( n224919 , n224786 , n224790 );
or ( n224920 , n224918 , n224919 );
xor ( n224921 , n224782 , n224794 );
not ( n224922 , n213750 );
buf ( n224923 , n224840 );
buf ( n224924 , n224923 );
not ( n224925 , n224924 );
not ( n224926 , n224925 );
or ( n224927 , n224922 , n224926 );
not ( n224928 , n215999 );
buf ( n224929 , n224923 );
nand ( n224930 , n224928 , n224929 );
nand ( n224931 , n224927 , n224930 );
not ( n224932 , n224931 );
and ( n224933 , n224923 , n224820 );
not ( n224934 , n224923 );
and ( n224935 , n224934 , n224821 );
nor ( n224936 , n224933 , n224935 );
nand ( n224937 , n224448 , n224936 );
not ( n224938 , n224937 );
not ( n224939 , n224938 );
or ( n224940 , n224932 , n224939 );
buf ( n224941 , n224449 );
not ( n224942 , n213077 );
buf ( n224943 , n224841 );
not ( n224944 , n224943 );
not ( n224945 , n224944 );
or ( n224946 , n224942 , n224945 );
not ( n224947 , n224929 );
nand ( n224948 , n224947 , n218224 );
nand ( n224949 , n224946 , n224948 );
nand ( n224950 , n224941 , n224949 );
nand ( n224951 , n224940 , n224950 );
xor ( n224952 , n224951 , n224409 );
xor ( n224953 , n224952 , n224455 );
xor ( n224954 , n224921 , n224953 );
xor ( n224955 , n224782 , n224794 );
and ( n224956 , n224955 , n224953 );
and ( n224957 , n224782 , n224794 );
or ( n224958 , n224956 , n224957 );
not ( n224959 , n224600 );
not ( n224960 , n222453 );
or ( n224961 , n224959 , n224960 );
not ( n224962 , n219475 );
not ( n224963 , n222458 );
or ( n224964 , n224962 , n224963 );
not ( n224965 , n222429 );
nand ( n224966 , n224965 , n214678 );
nand ( n224967 , n224964 , n224966 );
nand ( n224968 , n224967 , n222465 );
nand ( n224969 , n224961 , n224968 );
not ( n224970 , n224532 );
not ( n224971 , n224086 );
or ( n224972 , n224970 , n224971 );
not ( n224973 , n213583 );
not ( n224974 , n224094 );
not ( n224975 , n224974 );
not ( n224976 , n224975 );
or ( n224977 , n224973 , n224976 );
nand ( n224978 , n224068 , n214134 );
nand ( n224979 , n224977 , n224978 );
nand ( n224980 , n224090 , n224979 );
nand ( n224981 , n224972 , n224980 );
xor ( n224982 , n224969 , n224981 );
not ( n224983 , n224521 );
not ( n224984 , n223197 );
or ( n224985 , n224983 , n224984 );
not ( n224986 , n223155 );
and ( n224987 , n215131 , n224986 );
not ( n224988 , n215131 );
and ( n224989 , n224988 , n223155 );
or ( n224990 , n224987 , n224989 );
not ( n224991 , n224990 );
nand ( n224992 , n224991 , n222769 );
nand ( n224993 , n224985 , n224992 );
xor ( n224994 , n224982 , n224993 );
not ( n224995 , n224567 );
not ( n224996 , n220163 );
or ( n224997 , n224995 , n224996 );
not ( n224998 , n219343 );
not ( n224999 , n224563 );
or ( n225000 , n224998 , n224999 );
nand ( n225001 , n222791 , n219348 );
nand ( n225002 , n225000 , n225001 );
nand ( n225003 , n225002 , n220881 );
nand ( n225004 , n224997 , n225003 );
not ( n225005 , n224579 );
not ( n225006 , n223223 );
or ( n225007 , n225005 , n225006 );
not ( n225008 , n216934 );
not ( n225009 , n223228 );
or ( n225010 , n225008 , n225009 );
nand ( n225011 , n220900 , n216940 );
nand ( n225012 , n225010 , n225011 );
nand ( n225013 , n225012 , n220929 );
nand ( n225014 , n225007 , n225013 );
xor ( n225015 , n225004 , n225014 );
not ( n225016 , n224589 );
not ( n225017 , n224120 );
or ( n225018 , n225016 , n225017 );
and ( n225019 , n221607 , n215899 );
not ( n225020 , n221607 );
and ( n225021 , n225020 , n215075 );
nor ( n225022 , n225019 , n225021 );
not ( n225023 , n225022 );
nand ( n225024 , n225023 , n221387 );
nand ( n225025 , n225018 , n225024 );
xor ( n225026 , n225015 , n225025 );
xor ( n225027 , n224994 , n225026 );
not ( n225028 , n224499 );
not ( n225029 , n218221 );
or ( n225030 , n225028 , n225029 );
and ( n225031 , n214837 , n218771 );
not ( n225032 , n214837 );
and ( n225033 , n225032 , n221214 );
nor ( n225034 , n225031 , n225033 );
nand ( n225035 , n225034 , n218231 );
nand ( n225036 , n225030 , n225035 );
not ( n225037 , n224543 );
not ( n225038 , n218835 );
or ( n225039 , n225037 , n225038 );
not ( n225040 , n224037 );
not ( n225041 , n218814 );
or ( n225042 , n225040 , n225041 );
nand ( n225043 , n219128 , n224041 );
nand ( n225044 , n225042 , n225043 );
nand ( n225045 , n225044 , n218843 );
nand ( n225046 , n225039 , n225045 );
xor ( n225047 , n225036 , n225046 );
not ( n225048 , n224553 );
not ( n225049 , n221576 );
or ( n225050 , n225048 , n225049 );
not ( n225051 , n221495 );
not ( n225052 , n219440 );
or ( n225053 , n225051 , n225052 );
nand ( n225054 , n221228 , n221494 );
nand ( n225055 , n225053 , n225054 );
nand ( n225056 , n219076 , n225055 );
nand ( n225057 , n225050 , n225056 );
xor ( n225058 , n225047 , n225057 );
xor ( n225059 , n225027 , n225058 );
xor ( n225060 , n224994 , n225026 );
and ( n225061 , n225060 , n225058 );
and ( n225062 , n224994 , n225026 );
or ( n225063 , n225061 , n225062 );
xor ( n225064 , n224806 , n224802 );
xor ( n225065 , n225064 , n224798 );
xor ( n225066 , n224806 , n224802 );
and ( n225067 , n225066 , n224798 );
and ( n225068 , n224806 , n224802 );
or ( n225069 , n225067 , n225068 );
not ( n225070 , n213577 );
not ( n225071 , n224674 );
or ( n225072 , n225070 , n225071 );
not ( n225073 , n213735 );
not ( n225074 , n223330 );
or ( n225075 , n225073 , n225074 );
nand ( n225076 , n224286 , n213732 );
nand ( n225077 , n225075 , n225076 );
nand ( n225078 , n225077 , n216336 );
nand ( n225079 , n225072 , n225078 );
not ( n225080 , n219175 );
not ( n225081 , n219577 );
not ( n225082 , n221028 );
or ( n225083 , n225081 , n225082 );
nand ( n225084 , n40668 , n218661 );
nand ( n225085 , n225083 , n225084 );
not ( n225086 , n225085 );
or ( n225087 , n225080 , n225086 );
nand ( n225088 , n224685 , n217023 );
nand ( n225089 , n225087 , n225088 );
xor ( n225090 , n225079 , n225089 );
not ( n225091 , n217969 );
not ( n225092 , n224461 );
or ( n225093 , n225091 , n225092 );
not ( n225094 , n213382 );
not ( n225095 , n39926 );
or ( n225096 , n225094 , n225095 );
not ( n225097 , n39926 );
nand ( n225098 , n225097 , n217715 );
nand ( n225099 , n225096 , n225098 );
nand ( n225100 , n225099 , n211314 );
nand ( n225101 , n225093 , n225100 );
xor ( n225102 , n225090 , n225101 );
xor ( n225103 , n225102 , n224507 );
not ( n225104 , n213874 );
not ( n225105 , n224693 );
or ( n225106 , n225104 , n225105 );
not ( n225107 , n214818 );
not ( n225108 , n39995 );
not ( n225109 , n225108 );
or ( n225110 , n225107 , n225109 );
not ( n225111 , n225108 );
nand ( n225112 , n225111 , n218887 );
nand ( n225113 , n225110 , n225112 );
nand ( n225114 , n225113 , n217142 );
nand ( n225115 , n225106 , n225114 );
xor ( n225116 , n224910 , n225115 );
not ( n225117 , n220280 );
not ( n225118 , n224636 );
or ( n225119 , n225117 , n225118 );
not ( n225120 , n219358 );
not ( n225121 , n225120 );
not ( n225122 , n221040 );
or ( n225123 , n225121 , n225122 );
nand ( n225124 , n40624 , n216989 );
nand ( n225125 , n225123 , n225124 );
nand ( n225126 , n225125 , n219353 );
nand ( n225127 , n225119 , n225126 );
xor ( n225128 , n225116 , n225127 );
xor ( n225129 , n225103 , n225128 );
xor ( n225130 , n225102 , n224507 );
and ( n225131 , n225130 , n225128 );
and ( n225132 , n225102 , n224507 );
or ( n225133 , n225131 , n225132 );
not ( n225134 , n219731 );
not ( n225135 , n224645 );
or ( n225136 , n225134 , n225135 );
not ( n225137 , n216166 );
not ( n225138 , n220204 );
or ( n225139 , n225137 , n225138 );
not ( n225140 , n219532 );
nand ( n225141 , n225140 , n220538 );
nand ( n225142 , n225139 , n225141 );
nand ( n225143 , n225142 , n222185 );
nand ( n225144 , n225136 , n225143 );
not ( n225145 , n219314 );
not ( n225146 , n219687 );
not ( n225147 , n219595 );
or ( n225148 , n225146 , n225147 );
nand ( n225149 , n219599 , n221283 );
nand ( n225150 , n225148 , n225149 );
not ( n225151 , n225150 );
or ( n225152 , n225145 , n225151 );
nand ( n225153 , n224621 , n224624 );
nand ( n225154 , n225152 , n225153 );
xor ( n225155 , n225144 , n225154 );
not ( n225156 , n214086 );
not ( n225157 , n224704 );
or ( n225158 , n225156 , n225157 );
not ( n225159 , n217573 );
not ( n225160 , n222512 );
or ( n225161 , n225159 , n225160 );
nand ( n225162 , n40413 , n217397 );
nand ( n225163 , n225161 , n225162 );
nand ( n225164 , n225163 , n220941 );
nand ( n225165 , n225158 , n225164 );
xor ( n225166 , n225155 , n225165 );
not ( n225167 , n214717 );
not ( n225168 , n224658 );
or ( n225169 , n225167 , n225168 );
not ( n225170 , n221338 );
not ( n225171 , n40181 );
or ( n225172 , n225170 , n225171 );
not ( n225173 , n215113 );
nand ( n225174 , n225173 , n221716 );
nand ( n225175 , n225172 , n225174 );
nand ( n225176 , n225175 , n220985 );
nand ( n225177 , n225169 , n225176 );
not ( n225178 , n220820 );
not ( n225179 , n216810 );
not ( n225180 , n40258 );
or ( n225181 , n225179 , n225180 );
not ( n225182 , n215290 );
nand ( n225183 , n225182 , n223383 );
nand ( n225184 , n225181 , n225183 );
not ( n225185 , n225184 );
or ( n225186 , n225178 , n225185 );
nand ( n225187 , n224714 , n216299 );
nand ( n225188 , n225186 , n225187 );
xor ( n225189 , n225177 , n225188 );
xor ( n225190 , n225189 , n224871 );
xor ( n225191 , n225166 , n225190 );
xor ( n225192 , n225191 , n224916 );
xor ( n225193 , n225166 , n225190 );
and ( n225194 , n225193 , n224916 );
and ( n225195 , n225166 , n225190 );
or ( n225196 , n225194 , n225195 );
xor ( n225197 , n224513 , n224608 );
xor ( n225198 , n225197 , n225059 );
xor ( n225199 , n224513 , n224608 );
and ( n225200 , n225199 , n225059 );
and ( n225201 , n224513 , n224608 );
or ( n225202 , n225200 , n225201 );
xor ( n225203 , n224614 , n224954 );
xor ( n225204 , n225203 , n224726 );
xor ( n225205 , n224614 , n224954 );
and ( n225206 , n225205 , n224726 );
and ( n225207 , n224614 , n224954 );
or ( n225208 , n225206 , n225207 );
xor ( n225209 , n224666 , n225065 );
xor ( n225210 , n225209 , n224732 );
xor ( n225211 , n224666 , n225065 );
and ( n225212 , n225211 , n224732 );
and ( n225213 , n224666 , n225065 );
or ( n225214 , n225212 , n225213 );
xor ( n225215 , n225129 , n225192 );
xor ( n225216 , n225215 , n225198 );
xor ( n225217 , n225129 , n225192 );
and ( n225218 , n225217 , n225198 );
and ( n225219 , n225129 , n225192 );
or ( n225220 , n225218 , n225219 );
xor ( n225221 , n225036 , n225046 );
and ( n225222 , n225221 , n225057 );
and ( n225223 , n225036 , n225046 );
or ( n225224 , n225222 , n225223 );
xor ( n225225 , n224738 , n225204 );
xor ( n225226 , n225225 , n224744 );
xor ( n225227 , n224738 , n225204 );
and ( n225228 , n225227 , n224744 );
and ( n225229 , n224738 , n225204 );
or ( n225230 , n225228 , n225229 );
xor ( n225231 , n225210 , n225216 );
xor ( n225232 , n225231 , n224750 );
xor ( n225233 , n225210 , n225216 );
and ( n225234 , n225233 , n224750 );
and ( n225235 , n225210 , n225216 );
or ( n225236 , n225234 , n225235 );
xor ( n225237 , n224760 , n225226 );
xor ( n225238 , n225237 , n224766 );
xor ( n225239 , n224760 , n225226 );
and ( n225240 , n225239 , n224766 );
and ( n225241 , n224760 , n225226 );
or ( n225242 , n225240 , n225241 );
xor ( n225243 , n225232 , n225238 );
xor ( n225244 , n225243 , n224772 );
xor ( n225245 , n225232 , n225238 );
and ( n225246 , n225245 , n224772 );
and ( n225247 , n225232 , n225238 );
or ( n225248 , n225246 , n225247 );
xor ( n225249 , n225004 , n225014 );
and ( n225250 , n225249 , n225025 );
and ( n225251 , n225004 , n225014 );
or ( n225252 , n225250 , n225251 );
xor ( n225253 , n224969 , n224981 );
and ( n225254 , n225253 , n224993 );
and ( n225255 , n224969 , n224981 );
or ( n225256 , n225254 , n225255 );
xor ( n225257 , n224951 , n224409 );
and ( n225258 , n225257 , n224455 );
and ( n225259 , n224951 , n224409 );
or ( n225260 , n225258 , n225259 );
xor ( n225261 , n224910 , n225115 );
and ( n225262 , n225261 , n225127 );
and ( n225263 , n224910 , n225115 );
or ( n225264 , n225262 , n225263 );
xor ( n225265 , n225144 , n225154 );
and ( n225266 , n225265 , n225165 );
and ( n225267 , n225144 , n225154 );
or ( n225268 , n225266 , n225267 );
xor ( n225269 , n225177 , n225188 );
and ( n225270 , n225269 , n224871 );
and ( n225271 , n225177 , n225188 );
or ( n225272 , n225270 , n225271 );
xor ( n225273 , n225079 , n225089 );
and ( n225274 , n225273 , n225101 );
and ( n225275 , n225079 , n225089 );
or ( n225276 , n225274 , n225275 );
not ( n225277 , n224855 );
not ( n225278 , n218239 );
or ( n225279 , n225277 , n225278 );
and ( n225280 , n41701 , n217473 );
not ( n225281 , n41701 );
and ( n225282 , n225281 , n221923 );
or ( n225283 , n225280 , n225282 );
nand ( n225284 , n225283 , n217230 );
nand ( n225285 , n225279 , n225284 );
and ( n225286 , n208717 , n217602 );
not ( n225287 , n208717 );
and ( n225288 , n225287 , n216928 );
or ( n225289 , n225286 , n225288 );
not ( n225290 , n225289 );
or ( n225291 , n225290 , n217098 );
or ( n225292 , n217876 , n224866 );
nand ( n225293 , n225291 , n225292 );
xor ( n225294 , n225285 , n225293 );
not ( n225295 , n220414 );
not ( n225296 , n224812 );
or ( n225297 , n225295 , n225296 );
not ( n225298 , n215766 );
not ( n225299 , n41070 );
or ( n225300 , n225298 , n225299 );
nand ( n225301 , n41069 , n216277 );
nand ( n225302 , n225300 , n225301 );
nand ( n225303 , n225302 , n220033 );
nand ( n225304 , n225297 , n225303 );
xor ( n225305 , n225294 , n225304 );
xor ( n225306 , n225285 , n225293 );
and ( n225307 , n225306 , n225304 );
and ( n225308 , n225285 , n225293 );
or ( n225309 , n225307 , n225308 );
not ( n225310 , n224842 );
not ( n225311 , n36389 );
not ( n225312 , n225311 );
or ( n225313 , n225310 , n225312 );
nand ( n225314 , n224841 , n36389 );
nand ( n225315 , n225313 , n225314 );
not ( n225316 , n225315 );
nor ( n225317 , n225316 , n213751 );
not ( n225318 , n216619 );
not ( n225319 , n224883 );
not ( n225320 , n225319 );
or ( n225321 , n225318 , n225320 );
not ( n225322 , n223537 );
not ( n225323 , n40886 );
not ( n225324 , n225323 );
or ( n225325 , n225322 , n225324 );
or ( n225326 , n223537 , n225323 );
nand ( n225327 , n225325 , n225326 );
not ( n225328 , n217047 );
or ( n225329 , n225327 , n225328 );
nand ( n225330 , n225321 , n225329 );
xor ( n225331 , n225317 , n225330 );
and ( n225332 , n224857 , n224869 );
xor ( n225333 , n225331 , n225332 );
xor ( n225334 , n225317 , n225330 );
and ( n225335 , n225334 , n225332 );
and ( n225336 , n225317 , n225330 );
or ( n225337 , n225335 , n225336 );
not ( n225338 , n213874 );
not ( n225339 , n225113 );
or ( n225340 , n225338 , n225339 );
not ( n225341 , n216262 );
not ( n225342 , n39877 );
or ( n225343 , n225341 , n225342 );
not ( n225344 , n39877 );
nand ( n225345 , n225344 , n214824 );
nand ( n225346 , n225343 , n225345 );
nand ( n225347 , n225346 , n217142 );
nand ( n225348 , n225340 , n225347 );
xor ( n225349 , n225348 , n225252 );
xor ( n225350 , n225349 , n225256 );
xor ( n225351 , n225348 , n225252 );
and ( n225352 , n225351 , n225256 );
and ( n225353 , n225348 , n225252 );
or ( n225354 , n225352 , n225353 );
not ( n225355 , n213912 );
not ( n225356 , n213382 );
not ( n225357 , n39812 );
not ( n225358 , n225357 );
or ( n225359 , n225356 , n225358 );
nand ( n225360 , n39812 , n217715 );
nand ( n225361 , n225359 , n225360 );
not ( n225362 , n225361 );
or ( n225363 , n225355 , n225362 );
nand ( n225364 , n225099 , n217969 );
nand ( n225365 , n225363 , n225364 );
xor ( n225366 , n225365 , n225224 );
xor ( n225367 , n225366 , n225260 );
xor ( n225368 , n225365 , n225224 );
and ( n225369 , n225368 , n225260 );
and ( n225370 , n225365 , n225224 );
or ( n225371 , n225369 , n225370 );
and ( n225372 , n214899 , n223595 );
not ( n225373 , n214899 );
and ( n225374 , n225373 , n223201 );
or ( n225375 , n225372 , n225374 );
not ( n225376 , n222768 );
or ( n225377 , n225375 , n225376 );
not ( n225378 , n224990 );
nand ( n225379 , n223195 , n223194 );
not ( n225380 , n225379 );
nand ( n225381 , n225378 , n225380 );
nand ( n225382 , n225377 , n225381 );
not ( n225383 , n224949 );
not ( n225384 , n224938 );
or ( n225385 , n225383 , n225384 );
not ( n225386 , n222031 );
not ( n225387 , n224843 );
or ( n225388 , n225386 , n225387 );
not ( n225389 , n224929 );
nand ( n225390 , n225389 , n213347 );
nand ( n225391 , n225388 , n225390 );
nand ( n225392 , n225391 , n224449 );
nand ( n225393 , n225385 , n225392 );
xor ( n225394 , n225382 , n225393 );
not ( n225395 , n224905 );
not ( n225396 , n215183 );
or ( n225397 , n225395 , n225396 );
not ( n225398 , n40724 );
not ( n225399 , n221938 );
and ( n225400 , n225398 , n225399 );
and ( n225401 , n40724 , n218994 );
nor ( n225402 , n225400 , n225401 );
or ( n225403 , n225402 , n221932 );
nand ( n225404 , n225397 , n225403 );
xor ( n225405 , n225394 , n225404 );
or ( n225406 , n221624 , n225022 );
and ( n225407 , n218514 , n221607 );
not ( n225408 , n218514 );
and ( n225409 , n225408 , n221611 );
nor ( n225410 , n225407 , n225409 );
not ( n225411 , n225410 );
or ( n225412 , n225411 , n221386 );
nand ( n225413 , n225406 , n225412 );
not ( n225414 , n224967 );
not ( n225415 , n222453 );
or ( n225416 , n225414 , n225415 );
not ( n225417 , n216208 );
not ( n225418 , n222428 );
not ( n225419 , n225418 );
or ( n225420 , n225417 , n225419 );
nand ( n225421 , n222428 , n216207 );
nand ( n225422 , n225420 , n225421 );
nand ( n225423 , n225422 , n222158 );
nand ( n225424 , n225416 , n225423 );
xor ( n225425 , n225413 , n225424 );
not ( n225426 , n224979 );
not ( n225427 , n224086 );
or ( n225428 , n225426 , n225427 );
not ( n225429 , n214956 );
not ( n225430 , n224094 );
or ( n225431 , n225429 , n225430 );
nand ( n225432 , n224068 , n214960 );
nand ( n225433 , n225431 , n225432 );
nand ( n225434 , n224090 , n225433 );
nand ( n225435 , n225428 , n225434 );
xor ( n225436 , n225425 , n225435 );
xor ( n225437 , n225405 , n225436 );
not ( n225438 , n225055 );
not ( n225439 , n221576 );
or ( n225440 , n225438 , n225439 );
not ( n225441 , n216293 );
not ( n225442 , n219439 );
or ( n225443 , n225441 , n225442 );
nand ( n225444 , n219418 , n216290 );
nand ( n225445 , n225443 , n225444 );
nand ( n225446 , n219076 , n225445 );
nand ( n225447 , n225440 , n225446 );
not ( n225448 , n225002 );
not ( n225449 , n220163 );
or ( n225450 , n225448 , n225449 );
not ( n225451 , n221921 );
not ( n225452 , n220147 );
or ( n225453 , n225451 , n225452 );
not ( n225454 , n221256 );
nand ( n225455 , n225454 , n218980 );
nand ( n225456 , n225453 , n225455 );
nand ( n225457 , n220881 , n225456 );
nand ( n225458 , n225450 , n225457 );
xor ( n225459 , n225447 , n225458 );
not ( n225460 , n225012 );
not ( n225461 , n221266 );
or ( n225462 , n225460 , n225461 );
not ( n225463 , n219102 );
not ( n225464 , n220904 );
or ( n225465 , n225463 , n225464 );
nand ( n225466 , n220900 , n216139 );
nand ( n225467 , n225465 , n225466 );
not ( n225468 , n225467 );
or ( n225469 , n225468 , n220928 );
nand ( n225470 , n225462 , n225469 );
xor ( n225471 , n225459 , n225470 );
xor ( n225472 , n225437 , n225471 );
xor ( n225473 , n225405 , n225436 );
and ( n225474 , n225473 , n225471 );
and ( n225475 , n225405 , n225436 );
or ( n225476 , n225474 , n225475 );
not ( n225477 , n217505 );
not ( n225478 , n225477 );
not ( n225479 , n225478 );
not ( n225480 , n224892 );
or ( n225481 , n225479 , n225480 );
not ( n225482 , n208594 );
xor ( n225483 , n216419 , n225482 );
nand ( n225484 , n225483 , n219501 );
nand ( n225485 , n225481 , n225484 );
not ( n225486 , n225034 );
not ( n225487 , n219461 );
or ( n225488 , n225486 , n225487 );
buf ( n225489 , n218503 );
not ( n225490 , n225489 );
not ( n225491 , n225490 );
not ( n225492 , n218226 );
or ( n225493 , n225491 , n225492 );
nand ( n225494 , n218771 , n208726 );
nand ( n225495 , n225493 , n225494 );
nand ( n225496 , n225495 , n218231 );
nand ( n225497 , n225488 , n225496 );
xor ( n225498 , n225485 , n225497 );
not ( n225499 , n220853 );
not ( n225500 , n225044 );
or ( n225501 , n225499 , n225500 );
not ( n225502 , n224492 );
not ( n225503 , n218818 );
or ( n225504 , n225502 , n225503 );
buf ( n225505 , n214642 );
nand ( n225506 , n220859 , n225505 );
nand ( n225507 , n225504 , n225506 );
not ( n225508 , n225507 );
or ( n225509 , n221237 , n225508 );
nand ( n225510 , n225501 , n225509 );
xor ( n225511 , n225498 , n225510 );
xor ( n225512 , n225511 , n225268 );
xor ( n225513 , n225305 , n224875 );
not ( n225514 , n213577 );
not ( n225515 , n225077 );
or ( n225516 , n225514 , n225515 );
and ( n225517 , n40044 , n213732 );
not ( n225518 , n40044 );
and ( n225519 , n225518 , n213735 );
or ( n225520 , n225517 , n225519 );
nand ( n225521 , n225520 , n216336 );
nand ( n225522 , n225516 , n225521 );
xor ( n225523 , n225513 , n225522 );
xor ( n225524 , n225512 , n225523 );
xor ( n225525 , n225511 , n225268 );
and ( n225526 , n225525 , n225523 );
and ( n225527 , n225511 , n225268 );
or ( n225528 , n225526 , n225527 );
xor ( n225529 , n225272 , n225264 );
not ( n225530 , n219353 );
not ( n225531 , n215955 );
not ( n225532 , n221356 );
or ( n225533 , n225531 , n225532 );
nand ( n225534 , n207936 , n216989 );
nand ( n225535 , n225533 , n225534 );
not ( n225536 , n225535 );
or ( n225537 , n225530 , n225536 );
nand ( n225538 , n225125 , n217552 );
nand ( n225539 , n225537 , n225538 );
not ( n225540 , n219731 );
not ( n225541 , n225142 );
or ( n225542 , n225540 , n225541 );
not ( n225543 , n216166 );
not ( n225544 , n219880 );
or ( n225545 , n225543 , n225544 );
not ( n225546 , n222081 );
nand ( n225547 , n225546 , n219034 );
nand ( n225548 , n225545 , n225547 );
nand ( n225549 , n225548 , n222185 );
nand ( n225550 , n225542 , n225549 );
xor ( n225551 , n225539 , n225550 );
not ( n225552 , n219314 );
not ( n225553 , n219687 );
not ( n225554 , n219238 );
or ( n225555 , n225553 , n225554 );
not ( n225556 , n208042 );
nand ( n225557 , n225556 , n221283 );
nand ( n225558 , n225555 , n225557 );
not ( n225559 , n225558 );
or ( n225560 , n225552 , n225559 );
not ( n225561 , n225150 );
or ( n225562 , n225561 , n223825 );
nand ( n225563 , n225560 , n225562 );
xor ( n225564 , n225551 , n225563 );
xor ( n225565 , n225529 , n225564 );
xor ( n225566 , n225272 , n225264 );
and ( n225567 , n225566 , n225564 );
and ( n225568 , n225272 , n225264 );
or ( n225569 , n225567 , n225568 );
not ( n225570 , n216562 );
not ( n225571 , n225184 );
or ( n225572 , n225570 , n225571 );
not ( n225573 , n216810 );
not ( n225574 , n222120 );
or ( n225575 , n225573 , n225574 );
nand ( n225576 , n40396 , n215289 );
nand ( n225577 , n225575 , n225576 );
nand ( n225578 , n225577 , n220820 );
nand ( n225579 , n225572 , n225578 );
not ( n225580 , n217023 );
not ( n225581 , n225085 );
or ( n225582 , n225580 , n225581 );
not ( n225583 , n219577 );
not ( n225584 , n220599 );
or ( n225585 , n225583 , n225584 );
nand ( n225586 , n40410 , n219583 );
nand ( n225587 , n225585 , n225586 );
nand ( n225588 , n225587 , n219175 );
nand ( n225589 , n225582 , n225588 );
xor ( n225590 , n225579 , n225589 );
xor ( n225591 , n225590 , n224914 );
xor ( n225592 , n225591 , n225276 );
xor ( n225593 , n225592 , n224920 );
xor ( n225594 , n225591 , n225276 );
and ( n225595 , n225594 , n224920 );
and ( n225596 , n225591 , n225276 );
or ( n225597 , n225595 , n225596 );
not ( n225598 , n215137 );
and ( n225599 , n40484 , n217397 );
not ( n225600 , n40484 );
and ( n225601 , n225600 , n217573 );
or ( n225602 , n225599 , n225601 );
not ( n225603 , n225602 );
or ( n225604 , n225598 , n225603 );
nand ( n225605 , n225163 , n214086 );
nand ( n225606 , n225604 , n225605 );
not ( n225607 , n214717 );
not ( n225608 , n225175 );
or ( n225609 , n225607 , n225608 );
not ( n225610 , n221338 );
not ( n225611 , n222100 );
or ( n225612 , n225610 , n225611 );
nand ( n225613 , n40421 , n216037 );
nand ( n225614 , n225612 , n225613 );
nand ( n225615 , n225614 , n220985 );
nand ( n225616 , n225609 , n225615 );
xor ( n225617 , n225606 , n225616 );
xor ( n225618 , n225617 , n225333 );
xor ( n225619 , n225618 , n225063 );
xor ( n225620 , n225619 , n224958 );
xor ( n225621 , n225618 , n225063 );
and ( n225622 , n225621 , n224958 );
and ( n225623 , n225618 , n225063 );
or ( n225624 , n225622 , n225623 );
xor ( n225625 , n225367 , n225350 );
xor ( n225626 , n225625 , n225472 );
xor ( n225627 , n225367 , n225350 );
and ( n225628 , n225627 , n225472 );
and ( n225629 , n225367 , n225350 );
or ( n225630 , n225628 , n225629 );
xor ( n225631 , n225069 , n225133 );
xor ( n225632 , n225631 , n225565 );
xor ( n225633 , n225069 , n225133 );
and ( n225634 , n225633 , n225565 );
and ( n225635 , n225069 , n225133 );
or ( n225636 , n225634 , n225635 );
xor ( n225637 , n225524 , n225196 );
xor ( n225638 , n225637 , n225593 );
xor ( n225639 , n225524 , n225196 );
and ( n225640 , n225639 , n225593 );
and ( n225641 , n225524 , n225196 );
or ( n225642 , n225640 , n225641 );
xor ( n225643 , n225485 , n225497 );
and ( n225644 , n225643 , n225510 );
and ( n225645 , n225485 , n225497 );
or ( n225646 , n225644 , n225645 );
xor ( n225647 , n225626 , n225620 );
xor ( n225648 , n225647 , n225202 );
xor ( n225649 , n225626 , n225620 );
and ( n225650 , n225649 , n225202 );
and ( n225651 , n225626 , n225620 );
or ( n225652 , n225650 , n225651 );
xor ( n225653 , n225208 , n225214 );
xor ( n225654 , n225653 , n225632 );
xor ( n225655 , n225208 , n225214 );
and ( n225656 , n225655 , n225632 );
and ( n225657 , n225208 , n225214 );
or ( n225658 , n225656 , n225657 );
xor ( n225659 , n225638 , n225220 );
xor ( n225660 , n225659 , n225230 );
xor ( n225661 , n225638 , n225220 );
and ( n225662 , n225661 , n225230 );
and ( n225663 , n225638 , n225220 );
or ( n225664 , n225662 , n225663 );
xor ( n225665 , n225648 , n225654 );
xor ( n225666 , n225665 , n225236 );
xor ( n225667 , n225648 , n225654 );
and ( n225668 , n225667 , n225236 );
and ( n225669 , n225648 , n225654 );
or ( n225670 , n225668 , n225669 );
xor ( n225671 , n225660 , n225242 );
xor ( n225672 , n225671 , n225666 );
xor ( n225673 , n225660 , n225242 );
and ( n225674 , n225673 , n225666 );
and ( n225675 , n225660 , n225242 );
or ( n225676 , n225674 , n225675 );
xor ( n225677 , n225447 , n225458 );
and ( n225678 , n225677 , n225470 );
and ( n225679 , n225447 , n225458 );
or ( n225680 , n225678 , n225679 );
xor ( n225681 , n225413 , n225424 );
and ( n225682 , n225681 , n225435 );
and ( n225683 , n225413 , n225424 );
or ( n225684 , n225682 , n225683 );
xor ( n225685 , n225382 , n225393 );
and ( n225686 , n225685 , n225404 );
and ( n225687 , n225382 , n225393 );
or ( n225688 , n225686 , n225687 );
xor ( n225689 , n225305 , n224875 );
and ( n225690 , n225689 , n225522 );
and ( n225691 , n225305 , n224875 );
or ( n225692 , n225690 , n225691 );
xor ( n225693 , n225539 , n225550 );
and ( n225694 , n225693 , n225563 );
and ( n225695 , n225539 , n225550 );
or ( n225696 , n225694 , n225695 );
xor ( n225697 , n225606 , n225616 );
and ( n225698 , n225697 , n225333 );
and ( n225699 , n225606 , n225616 );
or ( n225700 , n225698 , n225699 );
xor ( n225701 , n225579 , n225589 );
and ( n225702 , n225701 , n224914 );
and ( n225703 , n225579 , n225589 );
or ( n225704 , n225702 , n225703 );
not ( n225705 , n217289 );
not ( n225706 , n225483 );
or ( n225707 , n225705 , n225706 );
not ( n225708 , n216593 );
and ( n225709 , n831 , n41246 );
not ( n225710 , n831 );
and ( n225711 , n225710 , n208484 );
nor ( n225712 , n225709 , n225711 );
or ( n225713 , n225708 , n225712 );
nand ( n225714 , n225712 , n217511 );
nand ( n225715 , n225713 , n225714 );
nand ( n225716 , n225715 , n217824 );
nand ( n225717 , n225707 , n225716 );
not ( n225718 , n217099 );
not ( n225719 , n216929 );
not ( n225720 , n218290 );
or ( n225721 , n225719 , n225720 );
nand ( n225722 , n41396 , n217076 );
nand ( n225723 , n225721 , n225722 );
not ( n225724 , n225723 );
or ( n225725 , n225718 , n225724 );
nand ( n225726 , n225289 , n218544 );
nand ( n225727 , n225725 , n225726 );
xor ( n225728 , n225717 , n225727 );
not ( n225729 , n213750 );
not ( n225730 , n36389 );
not ( n225731 , n225730 );
not ( n225732 , n225731 );
or ( n225733 , n225729 , n225732 );
nand ( n225734 , n225733 , n224943 );
nand ( n225735 , n225730 , n213751 );
and ( n225736 , n225734 , n225735 );
and ( n225737 , n36422 , n37605 );
not ( n225738 , n36422 );
not ( n225739 , n37605 );
and ( n225740 , n225738 , n225739 );
nor ( n225741 , n225737 , n225740 );
not ( n225742 , n225741 );
not ( n225743 , n225742 );
nor ( n225744 , n225736 , n225743 );
xor ( n225745 , n225728 , n225744 );
xor ( n225746 , n225717 , n225727 );
and ( n225747 , n225746 , n225744 );
and ( n225748 , n225717 , n225727 );
or ( n225749 , n225747 , n225748 );
not ( n225750 , n225302 );
not ( n225751 , n217486 );
or ( n225752 , n225750 , n225751 );
not ( n225753 , n220032 );
and ( n225754 , n41165 , n215766 );
not ( n225755 , n41165 );
and ( n225756 , n225755 , n220038 );
nor ( n225757 , n225754 , n225756 );
nand ( n225758 , n225753 , n225757 );
nand ( n225759 , n225752 , n225758 );
not ( n225760 , n225495 );
not ( n225761 , n218221 );
or ( n225762 , n225760 , n225761 );
not ( n225763 , n220264 );
not ( n225764 , n225763 );
not ( n225765 , n225764 );
not ( n225766 , n221214 );
or ( n225767 , n225765 , n225766 );
not ( n225768 , n216607 );
not ( n225769 , n225768 );
nand ( n225770 , n218208 , n225769 );
nand ( n225771 , n225767 , n225770 );
nand ( n225772 , n225771 , n218231 );
nand ( n225773 , n225762 , n225772 );
xor ( n225774 , n225759 , n225773 );
not ( n225775 , n225507 );
not ( n225776 , n218835 );
or ( n225777 , n225775 , n225776 );
not ( n225778 , n214837 );
not ( n225779 , n218814 );
or ( n225780 , n225778 , n225779 );
nand ( n225781 , n223671 , n218670 );
nand ( n225782 , n225780 , n225781 );
nand ( n225783 , n218843 , n225782 );
nand ( n225784 , n225777 , n225783 );
xor ( n225785 , n225774 , n225784 );
xor ( n225786 , n225759 , n225773 );
and ( n225787 , n225786 , n225784 );
and ( n225788 , n225759 , n225773 );
or ( n225789 , n225787 , n225788 );
not ( n225790 , n214319 );
not ( n225791 , n213382 );
not ( n225792 , n39711 );
not ( n225793 , n225792 );
or ( n225794 , n225791 , n225793 );
not ( n225795 , n39712 );
nand ( n225796 , n225795 , n213381 );
nand ( n225797 , n225794 , n225796 );
not ( n225798 , n225797 );
or ( n225799 , n225790 , n225798 );
nand ( n225800 , n225361 , n217969 );
nand ( n225801 , n225799 , n225800 );
xor ( n225802 , n225684 , n225801 );
xor ( n225803 , n225802 , n225646 );
xor ( n225804 , n225684 , n225801 );
and ( n225805 , n225804 , n225646 );
and ( n225806 , n225684 , n225801 );
or ( n225807 , n225805 , n225806 );
not ( n225808 , n225445 );
not ( n225809 , n221575 );
or ( n225810 , n225808 , n225809 );
xor ( n225811 , n214820 , n219439 );
nand ( n225812 , n225811 , n219075 );
nand ( n225813 , n225810 , n225812 );
not ( n225814 , n225456 );
not ( n225815 , n220162 );
or ( n225816 , n225814 , n225815 );
not ( n225817 , n221495 );
not ( n225818 , n224562 );
or ( n225819 , n225817 , n225818 );
nand ( n225820 , n225454 , n220022 );
nand ( n225821 , n225819 , n225820 );
nand ( n225822 , n225821 , n219778 );
nand ( n225823 , n225816 , n225822 );
xor ( n225824 , n225813 , n225823 );
not ( n225825 , n225467 );
not ( n225826 , n223223 );
or ( n225827 , n225825 , n225826 );
not ( n225828 , n219343 );
not ( n225829 , n224112 );
or ( n225830 , n225828 , n225829 );
nand ( n225831 , n220900 , n223269 );
nand ( n225832 , n225830 , n225831 );
nand ( n225833 , n225832 , n220929 );
nand ( n225834 , n225827 , n225833 );
xor ( n225835 , n225824 , n225834 );
xor ( n225836 , n225835 , n225688 );
not ( n225837 , n225433 );
not ( n225838 , n224084 );
nor ( n225839 , n225838 , n223810 );
not ( n225840 , n225839 );
or ( n225841 , n225837 , n225840 );
and ( n225842 , n217044 , n224974 );
not ( n225843 , n217044 );
not ( n225844 , n224974 );
and ( n225845 , n225843 , n225844 );
nor ( n225846 , n225842 , n225845 );
nand ( n225847 , n225846 , n223810 );
nand ( n225848 , n225841 , n225847 );
not ( n225849 , n225391 );
nand ( n225850 , n224448 , n224936 );
not ( n225851 , n225850 );
not ( n225852 , n225851 );
or ( n225853 , n225849 , n225852 );
not ( n225854 , n213583 );
not ( n225855 , n224943 );
or ( n225856 , n225854 , n225855 );
nand ( n225857 , n224929 , n214134 );
nand ( n225858 , n225856 , n225857 );
nand ( n225859 , n225858 , n224449 );
nand ( n225860 , n225853 , n225859 );
xor ( n225861 , n225848 , n225860 );
not ( n225862 , n225283 );
not ( n225863 , n217631 );
or ( n225864 , n225862 , n225863 );
not ( n225865 , n217614 );
buf ( n225866 , n41563 );
not ( n225867 , n225866 );
or ( n225868 , n225865 , n225867 );
nand ( n225869 , n217611 , n41564 );
nand ( n225870 , n225868 , n225869 );
nand ( n225871 , n225870 , n217641 );
nand ( n225872 , n225864 , n225871 );
not ( n225873 , n216630 );
and ( n225874 , n217119 , n216074 );
not ( n225875 , n217119 );
and ( n225876 , n225875 , n216624 );
or ( n225877 , n225874 , n225876 );
not ( n225878 , n225877 );
or ( n225879 , n225873 , n225878 );
not ( n225880 , n225327 );
nand ( n225881 , n225880 , n216619 );
nand ( n225882 , n225879 , n225881 );
xor ( n225883 , n225872 , n225882 );
xor ( n225884 , n225861 , n225883 );
xor ( n225885 , n225836 , n225884 );
xor ( n225886 , n225835 , n225688 );
and ( n225887 , n225886 , n225884 );
and ( n225888 , n225835 , n225688 );
or ( n225889 , n225887 , n225888 );
not ( n225890 , n223587 );
not ( n225891 , n216934 );
not ( n225892 , n221611 );
or ( n225893 , n225891 , n225892 );
nand ( n225894 , n221607 , n216940 );
nand ( n225895 , n225893 , n225894 );
not ( n225896 , n225895 );
or ( n225897 , n225890 , n225896 );
nand ( n225898 , n225410 , n221623 );
nand ( n225899 , n225897 , n225898 );
not ( n225900 , n225422 );
nand ( n225901 , n222447 , n222451 );
not ( n225902 , n225901 );
not ( n225903 , n225902 );
or ( n225904 , n225900 , n225903 );
not ( n225905 , n215075 );
not ( n225906 , n225418 );
or ( n225907 , n225905 , n225906 );
nand ( n225908 , n222428 , n215899 );
nand ( n225909 , n225907 , n225908 );
nand ( n225910 , n222157 , n225909 );
nand ( n225911 , n225904 , n225910 );
xor ( n225912 , n225899 , n225911 );
not ( n225913 , n216964 );
not ( n225914 , n223201 );
not ( n225915 , n225914 );
or ( n225916 , n225913 , n225915 );
nand ( n225917 , n223201 , n214678 );
nand ( n225918 , n225916 , n225917 );
not ( n225919 , n225918 );
not ( n225920 , n222768 );
or ( n225921 , n225919 , n225920 );
not ( n225922 , n225375 );
nand ( n225923 , n225922 , n223197 );
nand ( n225924 , n225921 , n225923 );
xor ( n225925 , n225912 , n225924 );
xor ( n225926 , n225925 , n225785 );
xor ( n225927 , n225926 , n225696 );
xor ( n225928 , n225925 , n225785 );
and ( n225929 , n225928 , n225696 );
and ( n225930 , n225925 , n225785 );
or ( n225931 , n225929 , n225930 );
xor ( n225932 , n225700 , n225704 );
not ( n225933 , n215999 );
not ( n225934 , n225743 );
or ( n225935 , n225933 , n225934 );
not ( n225936 , n225743 );
nand ( n225937 , n225936 , n213751 );
nand ( n225938 , n225935 , n225937 );
not ( n225939 , n225938 );
buf ( n225940 , n225741 );
and ( n225941 , n225940 , n225730 );
not ( n225942 , n225940 );
and ( n225943 , n225942 , n36389 );
nor ( n225944 , n225941 , n225943 );
and ( n225945 , n225316 , n225944 );
not ( n225946 , n225945 );
or ( n225947 , n225939 , n225946 );
not ( n225948 , n225316 );
not ( n225949 , n213126 );
not ( n225950 , n225940 );
or ( n225951 , n225949 , n225950 );
buf ( n225952 , n225742 );
nand ( n225953 , n225952 , n216076 );
nand ( n225954 , n225951 , n225953 );
nand ( n225955 , n225948 , n225954 );
nand ( n225956 , n225947 , n225955 );
xor ( n225957 , n225956 , n225309 );
xor ( n225958 , n225957 , n225337 );
xor ( n225959 , n225932 , n225958 );
xor ( n225960 , n225700 , n225704 );
and ( n225961 , n225960 , n225958 );
and ( n225962 , n225700 , n225704 );
or ( n225963 , n225961 , n225962 );
not ( n225964 , n213498 );
xnor ( n225965 , n213732 , n39995 );
not ( n225966 , n225965 );
or ( n225967 , n225964 , n225966 );
nand ( n225968 , n225520 , n213577 );
nand ( n225969 , n225967 , n225968 );
xor ( n225970 , n225969 , n225745 );
not ( n225971 , n219175 );
not ( n225972 , n217017 );
not ( n225973 , n223384 );
or ( n225974 , n225972 , n225973 );
nand ( n225975 , n221743 , n218661 );
nand ( n225976 , n225974 , n225975 );
not ( n225977 , n225976 );
or ( n225978 , n225971 , n225977 );
nand ( n225979 , n225587 , n217023 );
nand ( n225980 , n225978 , n225979 );
xor ( n225981 , n225970 , n225980 );
xor ( n225982 , n225692 , n225981 );
not ( n225983 , n225602 );
or ( n225984 , n225983 , n214085 );
not ( n225985 , n40545 );
not ( n225986 , n215388 );
and ( n225987 , n225985 , n225986 );
and ( n225988 , n40545 , n217397 );
nor ( n225989 , n225987 , n225988 );
or ( n225990 , n223390 , n225989 );
nand ( n225991 , n225984 , n225990 );
not ( n225992 , n225535 );
or ( n225993 , n225992 , n217551 );
and ( n225994 , n40668 , n215955 );
not ( n225995 , n40668 );
and ( n225996 , n225995 , n219358 );
or ( n225997 , n225994 , n225996 );
or ( n225998 , n217549 , n225997 );
nand ( n225999 , n225993 , n225998 );
xor ( n226000 , n225991 , n225999 );
not ( n226001 , n222185 );
not ( n226002 , n216166 );
and ( n226003 , n40623 , n226002 );
not ( n226004 , n40623 );
and ( n226005 , n226004 , n219033 );
or ( n226006 , n226003 , n226005 );
not ( n226007 , n226006 );
or ( n226008 , n226001 , n226007 );
not ( n226009 , n225548 );
not ( n226010 , n219731 );
or ( n226011 , n226009 , n226010 );
nand ( n226012 , n226008 , n226011 );
xor ( n226013 , n226000 , n226012 );
xor ( n226014 , n225982 , n226013 );
xor ( n226015 , n225692 , n225981 );
and ( n226016 , n226015 , n226013 );
and ( n226017 , n225692 , n225981 );
or ( n226018 , n226016 , n226017 );
not ( n226019 , n216204 );
not ( n226020 , n225558 );
or ( n226021 , n226019 , n226020 );
and ( n226022 , n221283 , n219532 );
not ( n226023 , n221283 );
and ( n226024 , n226023 , n40802 );
nor ( n226025 , n226022 , n226024 );
nand ( n226026 , n226025 , n219314 );
nand ( n226027 , n226021 , n226026 );
not ( n226028 , n214717 );
not ( n226029 , n225614 );
or ( n226030 , n226028 , n226029 );
and ( n226031 , n40413 , n216037 );
not ( n226032 , n40413 );
and ( n226033 , n226032 , n215113 );
or ( n226034 , n226031 , n226033 );
nand ( n226035 , n226034 , n220985 );
nand ( n226036 , n226030 , n226035 );
xor ( n226037 , n226027 , n226036 );
not ( n226038 , n218990 );
not ( n226039 , n218883 );
or ( n226040 , n226038 , n226039 );
nand ( n226041 , n40710 , n218994 );
nand ( n226042 , n226040 , n226041 );
not ( n226043 , n226042 );
or ( n226044 , n226043 , n221932 );
not ( n226045 , n225402 );
nand ( n226046 , n226045 , n219332 );
nand ( n226047 , n226044 , n226046 );
xor ( n226048 , n226037 , n226047 );
xor ( n226049 , n225354 , n226048 );
not ( n226050 , n220820 );
not ( n226051 , n216810 );
not ( n226052 , n40181 );
or ( n226053 , n226051 , n226052 );
nand ( n226054 , n223320 , n215289 );
nand ( n226055 , n226053 , n226054 );
not ( n226056 , n226055 );
or ( n226057 , n226050 , n226056 );
nand ( n226058 , n225577 , n216299 );
nand ( n226059 , n226057 , n226058 );
not ( n226060 , n213874 );
not ( n226061 , n225346 );
or ( n226062 , n226060 , n226061 );
not ( n226063 , n220300 );
not ( n226064 , n225097 );
or ( n226065 , n226063 , n226064 );
nand ( n226066 , n39926 , n216262 );
nand ( n226067 , n226065 , n226066 );
nand ( n226068 , n226067 , n217142 );
nand ( n226069 , n226062 , n226068 );
xor ( n226070 , n226059 , n226069 );
xor ( n226071 , n226070 , n225680 );
xor ( n226072 , n226049 , n226071 );
xor ( n226073 , n225354 , n226048 );
and ( n226074 , n226073 , n226071 );
and ( n226075 , n225354 , n226048 );
or ( n226076 , n226074 , n226075 );
xor ( n226077 , n225371 , n225476 );
xor ( n226078 , n226077 , n225803 );
xor ( n226079 , n225371 , n225476 );
and ( n226080 , n226079 , n225803 );
and ( n226081 , n225371 , n225476 );
or ( n226082 , n226080 , n226081 );
xor ( n226083 , n225885 , n225927 );
xor ( n226084 , n226083 , n225528 );
xor ( n226085 , n225885 , n225927 );
and ( n226086 , n226085 , n225528 );
and ( n226087 , n225885 , n225927 );
or ( n226088 , n226086 , n226087 );
xor ( n226089 , n225959 , n225597 );
xor ( n226090 , n226089 , n225569 );
xor ( n226091 , n225959 , n225597 );
and ( n226092 , n226091 , n225569 );
and ( n226093 , n225959 , n225597 );
or ( n226094 , n226092 , n226093 );
xor ( n226095 , n225624 , n226014 );
xor ( n226096 , n226095 , n226072 );
xor ( n226097 , n225624 , n226014 );
and ( n226098 , n226097 , n226072 );
and ( n226099 , n225624 , n226014 );
or ( n226100 , n226098 , n226099 );
xor ( n226101 , n225813 , n225823 );
and ( n226102 , n226101 , n225834 );
and ( n226103 , n225813 , n225823 );
or ( n226104 , n226102 , n226103 );
xor ( n226105 , n226078 , n225630 );
xor ( n226106 , n226105 , n226084 );
xor ( n226107 , n226078 , n225630 );
and ( n226108 , n226107 , n226084 );
and ( n226109 , n226078 , n225630 );
or ( n226110 , n226108 , n226109 );
xor ( n226111 , n225636 , n226090 );
xor ( n226112 , n226111 , n225642 );
xor ( n226113 , n225636 , n226090 );
and ( n226114 , n226113 , n225642 );
and ( n226115 , n225636 , n226090 );
or ( n226116 , n226114 , n226115 );
xor ( n226117 , n225652 , n226096 );
xor ( n226118 , n226117 , n226106 );
xor ( n226119 , n225652 , n226096 );
and ( n226120 , n226119 , n226106 );
and ( n226121 , n225652 , n226096 );
or ( n226122 , n226120 , n226121 );
xor ( n226123 , n225658 , n226112 );
xor ( n226124 , n226123 , n225664 );
xor ( n226125 , n225658 , n226112 );
and ( n226126 , n226125 , n225664 );
and ( n226127 , n225658 , n226112 );
or ( n226128 , n226126 , n226127 );
xor ( n226129 , n226118 , n225670 );
xor ( n226130 , n226129 , n226124 );
xor ( n226131 , n226118 , n225670 );
and ( n226132 , n226131 , n226124 );
and ( n226133 , n226118 , n225670 );
or ( n226134 , n226132 , n226133 );
xor ( n226135 , n225899 , n225911 );
and ( n226136 , n226135 , n225924 );
and ( n226137 , n225899 , n225911 );
or ( n226138 , n226136 , n226137 );
xor ( n226139 , n225848 , n225860 );
and ( n226140 , n226139 , n225883 );
and ( n226141 , n225848 , n225860 );
or ( n226142 , n226140 , n226141 );
xor ( n226143 , n225956 , n225309 );
and ( n226144 , n226143 , n225337 );
and ( n226145 , n225956 , n225309 );
or ( n226146 , n226144 , n226145 );
xor ( n226147 , n225991 , n225999 );
and ( n226148 , n226147 , n226012 );
and ( n226149 , n225991 , n225999 );
or ( n226150 , n226148 , n226149 );
xor ( n226151 , n226027 , n226036 );
and ( n226152 , n226151 , n226047 );
and ( n226153 , n226027 , n226036 );
or ( n226154 , n226152 , n226153 );
xor ( n226155 , n225969 , n225745 );
and ( n226156 , n226155 , n225980 );
and ( n226157 , n225969 , n225745 );
or ( n226158 , n226156 , n226157 );
xor ( n226159 , n226059 , n226069 );
and ( n226160 , n226159 , n225680 );
and ( n226161 , n226059 , n226069 );
or ( n226162 , n226160 , n226161 );
not ( n226163 , n218762 );
not ( n226164 , n218560 );
not ( n226165 , n215793 );
or ( n226166 , n226164 , n226165 );
not ( n226167 , n221923 );
nand ( n226168 , n226167 , n208717 );
nand ( n226169 , n226166 , n226168 );
not ( n226170 , n226169 );
or ( n226171 , n226163 , n226170 );
not ( n226172 , n217629 );
nand ( n226173 , n226172 , n225870 );
nand ( n226174 , n226171 , n226173 );
not ( n226175 , n216619 );
not ( n226176 , n225877 );
or ( n226177 , n226175 , n226176 );
not ( n226178 , n216015 );
not ( n226179 , n218420 );
or ( n226180 , n226178 , n226179 );
nand ( n226181 , n41069 , n216404 );
nand ( n226182 , n226180 , n226181 );
nand ( n226183 , n226182 , n223949 );
nand ( n226184 , n226177 , n226183 );
xor ( n226185 , n226174 , n226184 );
not ( n226186 , n216598 );
not ( n226187 , n216762 );
not ( n226188 , n219051 );
or ( n226189 , n226187 , n226188 );
nand ( n226190 , n219050 , n224398 );
nand ( n226191 , n226189 , n226190 );
not ( n226192 , n226191 );
or ( n226193 , n226186 , n226192 );
buf ( n226194 , n225715 );
nand ( n226195 , n217505 , n226194 );
nand ( n226196 , n226193 , n226195 );
xor ( n226197 , n226185 , n226196 );
xor ( n226198 , n226174 , n226184 );
and ( n226199 , n226198 , n226196 );
and ( n226200 , n226174 , n226184 );
or ( n226201 , n226199 , n226200 );
not ( n226202 , n217388 );
not ( n226203 , n216929 );
not ( n226204 , n41318 );
or ( n226205 , n226203 , n226204 );
nand ( n226206 , n216311 , n220050 );
nand ( n226207 , n226205 , n226206 );
not ( n226208 , n226207 );
or ( n226209 , n226202 , n226208 );
nand ( n226210 , n225723 , n219368 );
nand ( n226211 , n226209 , n226210 );
not ( n226212 , n36370 );
and ( n226213 , n225742 , n226212 );
not ( n226214 , n225742 );
and ( n226215 , n226214 , n36370 );
nor ( n226216 , n226213 , n226215 );
buf ( n226217 , n226216 );
not ( n226218 , n226217 );
and ( n226219 , n226218 , n213750 );
xor ( n226220 , n226211 , n226219 );
not ( n226221 , n225771 );
not ( n226222 , n218221 );
or ( n226223 , n226221 , n226222 );
buf ( n226224 , n216339 );
not ( n226225 , n226224 );
not ( n226226 , n226225 );
not ( n226227 , n218772 );
or ( n226228 , n226226 , n226227 );
nand ( n226229 , n218208 , n226224 );
nand ( n226230 , n226228 , n226229 );
nand ( n226231 , n226230 , n218231 );
nand ( n226232 , n226223 , n226231 );
xor ( n226233 , n226220 , n226232 );
xor ( n226234 , n226211 , n226219 );
and ( n226235 , n226234 , n226232 );
and ( n226236 , n226211 , n226219 );
or ( n226237 , n226235 , n226236 );
xor ( n226238 , n226138 , n226142 );
not ( n226239 , n217969 );
not ( n226240 , n225797 );
or ( n226241 , n226239 , n226240 );
not ( n226242 , n213382 );
not ( n226243 , n39747 );
not ( n226244 , n226243 );
or ( n226245 , n226242 , n226244 );
nand ( n226246 , n39747 , n217715 );
nand ( n226247 , n226245 , n226246 );
nand ( n226248 , n226247 , n211314 );
nand ( n226249 , n226241 , n226248 );
xor ( n226250 , n226238 , n226249 );
xor ( n226251 , n226138 , n226142 );
and ( n226252 , n226251 , n226249 );
and ( n226253 , n226138 , n226142 );
or ( n226254 , n226252 , n226253 );
not ( n226255 , n225965 );
not ( n226256 , n213577 );
or ( n226257 , n226255 , n226256 );
and ( n226258 , n213735 , n39877 );
not ( n226259 , n213735 );
and ( n226260 , n226259 , n39878 );
nor ( n226261 , n226258 , n226260 );
or ( n226262 , n226261 , n216335 );
nand ( n226263 , n226257 , n226262 );
xor ( n226264 , n226233 , n226263 );
xor ( n226265 , n226264 , n225789 );
xor ( n226266 , n226233 , n226263 );
and ( n226267 , n226266 , n225789 );
and ( n226268 , n226233 , n226263 );
or ( n226269 , n226267 , n226268 );
not ( n226270 , n225954 );
nand ( n226271 , n225316 , n225944 );
not ( n226272 , n226271 );
not ( n226273 , n226272 );
or ( n226274 , n226270 , n226273 );
not ( n226275 , n222032 );
not ( n226276 , n225952 );
not ( n226277 , n226276 );
or ( n226278 , n226275 , n226277 );
not ( n226279 , n213347 );
nand ( n226280 , n226279 , n225952 );
nand ( n226281 , n226278 , n226280 );
nand ( n226282 , n226281 , n225948 );
nand ( n226283 , n226274 , n226282 );
and ( n226284 , n225882 , n225872 );
xor ( n226285 , n226283 , n226284 );
not ( n226286 , n220033 );
not ( n226287 , n226286 );
not ( n226288 , n226287 );
not ( n226289 , n220038 );
not ( n226290 , n40724 );
or ( n226291 , n226289 , n226290 );
buf ( n226292 , n220749 );
nand ( n226293 , n224617 , n226292 );
nand ( n226294 , n226291 , n226293 );
not ( n226295 , n226294 );
or ( n226296 , n226288 , n226295 );
nand ( n226297 , n225757 , n220414 );
nand ( n226298 , n226296 , n226297 );
xor ( n226299 , n226285 , n226298 );
xor ( n226300 , n226146 , n226299 );
not ( n226301 , n225782 );
not ( n226302 , n220479 );
or ( n226303 , n226301 , n226302 );
buf ( n226304 , n219689 );
not ( n226305 , n226304 );
not ( n226306 , n218814 );
or ( n226307 , n226305 , n226306 );
nand ( n226308 , n220126 , n225489 );
nand ( n226309 , n226307 , n226308 );
nand ( n226310 , n226309 , n218455 );
nand ( n226311 , n226303 , n226310 );
not ( n226312 , n225811 );
not ( n226313 , n223620 );
or ( n226314 , n226312 , n226313 );
not ( n226315 , n224492 );
not ( n226316 , n219423 );
or ( n226317 , n226315 , n226316 );
nand ( n226318 , n219443 , n214642 );
nand ( n226319 , n226317 , n226318 );
nand ( n226320 , n226319 , n219076 );
nand ( n226321 , n226314 , n226320 );
xor ( n226322 , n226311 , n226321 );
not ( n226323 , n225821 );
not ( n226324 , n220492 );
or ( n226325 , n226323 , n226324 );
not ( n226326 , n216293 );
not ( n226327 , n222412 );
or ( n226328 , n226326 , n226327 );
nand ( n226329 , n225454 , n223658 );
nand ( n226330 , n226328 , n226329 );
nand ( n226331 , n219779 , n226330 );
nand ( n226332 , n226325 , n226331 );
xor ( n226333 , n226322 , n226332 );
xor ( n226334 , n226300 , n226333 );
xor ( n226335 , n226146 , n226299 );
and ( n226336 , n226335 , n226333 );
and ( n226337 , n226146 , n226299 );
or ( n226338 , n226336 , n226337 );
not ( n226339 , n225380 );
not ( n226340 , n225918 );
or ( n226341 , n226339 , n226340 );
not ( n226342 , n216208 );
not ( n226343 , n223595 );
or ( n226344 , n226342 , n226343 );
nand ( n226345 , n223155 , n216207 );
nand ( n226346 , n226344 , n226345 );
nand ( n226347 , n226346 , n222768 );
nand ( n226348 , n226341 , n226347 );
not ( n226349 , n225846 );
not ( n226350 , n224086 );
or ( n226351 , n226349 , n226350 );
not ( n226352 , n214537 );
not ( n226353 , n224069 );
or ( n226354 , n226352 , n226353 );
not ( n226355 , n224069 );
nand ( n226356 , n226355 , n214899 );
nand ( n226357 , n226354 , n226356 );
nand ( n226358 , n224090 , n226357 );
nand ( n226359 , n226351 , n226358 );
xor ( n226360 , n226348 , n226359 );
not ( n226361 , n225858 );
not ( n226362 , n224938 );
or ( n226363 , n226361 , n226362 );
and ( n226364 , n224843 , n214960 );
not ( n226365 , n224843 );
and ( n226366 , n226365 , n214956 );
or ( n226367 , n226364 , n226366 );
nand ( n226368 , n226367 , n224941 );
nand ( n226369 , n226363 , n226368 );
xor ( n226370 , n226360 , n226369 );
not ( n226371 , n225832 );
not ( n226372 , n223223 );
or ( n226373 , n226371 , n226372 );
not ( n226374 , n222821 );
not ( n226375 , n223227 );
or ( n226376 , n226374 , n226375 );
not ( n226377 , n220904 );
nand ( n226378 , n226377 , n218980 );
nand ( n226379 , n226376 , n226378 );
nand ( n226380 , n226379 , n221674 );
nand ( n226381 , n226373 , n226380 );
not ( n226382 , n225895 );
not ( n226383 , n224120 );
or ( n226384 , n226382 , n226383 );
not ( n226385 , n219102 );
not ( n226386 , n221777 );
or ( n226387 , n226385 , n226386 );
not ( n226388 , n221612 );
nand ( n226389 , n226388 , n216139 );
nand ( n226390 , n226387 , n226389 );
nand ( n226391 , n226390 , n221387 );
nand ( n226392 , n226384 , n226391 );
xor ( n226393 , n226381 , n226392 );
not ( n226394 , n225909 );
not ( n226395 , n222454 );
or ( n226396 , n226394 , n226395 );
not ( n226397 , n218514 );
not ( n226398 , n222429 );
or ( n226399 , n226397 , n226398 );
nand ( n226400 , n222428 , n216170 );
nand ( n226401 , n226399 , n226400 );
nand ( n226402 , n222467 , n226401 );
nand ( n226403 , n226396 , n226402 );
xor ( n226404 , n226393 , n226403 );
xor ( n226405 , n226370 , n226404 );
xor ( n226406 , n226405 , n226150 );
xor ( n226407 , n226370 , n226404 );
and ( n226408 , n226407 , n226150 );
and ( n226409 , n226370 , n226404 );
or ( n226410 , n226408 , n226409 );
xor ( n226411 , n226158 , n226154 );
xor ( n226412 , n226411 , n226162 );
xor ( n226413 , n226158 , n226154 );
and ( n226414 , n226413 , n226162 );
and ( n226415 , n226158 , n226154 );
or ( n226416 , n226414 , n226415 );
not ( n226417 , n215137 );
not ( n226418 , n217573 );
not ( n226419 , n223761 );
or ( n226420 , n226418 , n226419 );
nand ( n226421 , n40045 , n217397 );
nand ( n226422 , n226420 , n226421 );
not ( n226423 , n226422 );
or ( n226424 , n226417 , n226423 );
not ( n226425 , n225989 );
nand ( n226426 , n226425 , n215605 );
nand ( n226427 , n226424 , n226426 );
xor ( n226428 , n226197 , n226427 );
not ( n226429 , n214694 );
not ( n226430 , n216810 );
not ( n226431 , n223748 );
or ( n226432 , n226430 , n226431 );
nand ( n226433 , n40422 , n215289 );
nand ( n226434 , n226432 , n226433 );
not ( n226435 , n226434 );
or ( n226436 , n226429 , n226435 );
nand ( n226437 , n226055 , n216562 );
nand ( n226438 , n226436 , n226437 );
xor ( n226439 , n226428 , n226438 );
not ( n226440 , n214717 );
not ( n226441 , n226034 );
or ( n226442 , n226440 , n226441 );
not ( n226443 , n215113 );
not ( n226444 , n40484 );
not ( n226445 , n226444 );
or ( n226446 , n226443 , n226445 );
nand ( n226447 , n40484 , n217944 );
nand ( n226448 , n226446 , n226447 );
nand ( n226449 , n226448 , n216239 );
nand ( n226450 , n226442 , n226449 );
xor ( n226451 , n225749 , n226450 );
or ( n226452 , n225997 , n217551 );
xor ( n226453 , n219358 , n40409 );
or ( n226454 , n226453 , n217549 );
nand ( n226455 , n226452 , n226454 );
xor ( n226456 , n226451 , n226455 );
xor ( n226457 , n226439 , n226456 );
xor ( n226458 , n226457 , n225807 );
xor ( n226459 , n226439 , n226456 );
and ( n226460 , n226459 , n225807 );
and ( n226461 , n226439 , n226456 );
or ( n226462 , n226460 , n226461 );
not ( n226463 , n219731 );
not ( n226464 , n226006 );
or ( n226465 , n226463 , n226464 );
and ( n226466 , n40658 , n220538 );
not ( n226467 , n40658 );
and ( n226468 , n226467 , n219033 );
or ( n226469 , n226466 , n226468 );
nand ( n226470 , n226469 , n214458 );
nand ( n226471 , n226465 , n226470 );
not ( n226472 , n224624 );
not ( n226473 , n226025 );
or ( n226474 , n226472 , n226473 );
not ( n226475 , n219687 );
not ( n226476 , n222081 );
or ( n226477 , n226475 , n226476 );
nand ( n226478 , n40559 , n221283 );
nand ( n226479 , n226477 , n226478 );
nand ( n226480 , n226479 , n219314 );
nand ( n226481 , n226474 , n226480 );
xor ( n226482 , n226471 , n226481 );
not ( n226483 , n221933 );
not ( n226484 , n221938 );
not ( n226485 , n226484 );
buf ( n226486 , n219238 );
not ( n226487 , n226486 );
or ( n226488 , n226485 , n226487 );
buf ( n226489 , n225556 );
nand ( n226490 , n226489 , n218994 );
nand ( n226491 , n226488 , n226490 );
not ( n226492 , n226491 );
or ( n226493 , n226483 , n226492 );
nand ( n226494 , n226042 , n215183 );
nand ( n226495 , n226493 , n226494 );
xor ( n226496 , n226482 , n226495 );
xor ( n226497 , n226496 , n225889 );
not ( n226498 , n217023 );
not ( n226499 , n225976 );
or ( n226500 , n226498 , n226499 );
not ( n226501 , n219577 );
not ( n226502 , n222121 );
or ( n226503 , n226501 , n226502 );
not ( n226504 , n40396 );
not ( n226505 , n226504 );
nand ( n226506 , n226505 , n218661 );
nand ( n226507 , n226503 , n226506 );
nand ( n226508 , n226507 , n219175 );
nand ( n226509 , n226500 , n226508 );
not ( n226510 , n213874 );
not ( n226511 , n226067 );
or ( n226512 , n226510 , n226511 );
not ( n226513 , n214818 );
not ( n226514 , n225357 );
or ( n226515 , n226513 , n226514 );
nand ( n226516 , n39812 , n216265 );
nand ( n226517 , n226515 , n226516 );
nand ( n226518 , n226517 , n217142 );
nand ( n226519 , n226512 , n226518 );
xor ( n226520 , n226509 , n226519 );
xor ( n226521 , n226520 , n226104 );
xor ( n226522 , n226497 , n226521 );
xor ( n226523 , n226496 , n225889 );
and ( n226524 , n226523 , n226521 );
and ( n226525 , n226496 , n225889 );
or ( n226526 , n226524 , n226525 );
xor ( n226527 , n226250 , n226265 );
xor ( n226528 , n226527 , n226334 );
xor ( n226529 , n226250 , n226265 );
and ( n226530 , n226529 , n226334 );
and ( n226531 , n226250 , n226265 );
or ( n226532 , n226530 , n226531 );
xor ( n226533 , n225931 , n226406 );
xor ( n226534 , n226533 , n225963 );
xor ( n226535 , n225931 , n226406 );
and ( n226536 , n226535 , n225963 );
and ( n226537 , n225931 , n226406 );
or ( n226538 , n226536 , n226537 );
xor ( n226539 , n226018 , n226412 );
xor ( n226540 , n226539 , n226076 );
xor ( n226541 , n226018 , n226412 );
and ( n226542 , n226541 , n226076 );
and ( n226543 , n226018 , n226412 );
or ( n226544 , n226542 , n226543 );
xor ( n226545 , n226311 , n226321 );
and ( n226546 , n226545 , n226332 );
and ( n226547 , n226311 , n226321 );
or ( n226548 , n226546 , n226547 );
xor ( n226549 , n226082 , n226458 );
xor ( n226550 , n226549 , n226088 );
xor ( n226551 , n226082 , n226458 );
and ( n226552 , n226551 , n226088 );
and ( n226553 , n226082 , n226458 );
or ( n226554 , n226552 , n226553 );
xor ( n226555 , n226522 , n226528 );
xor ( n226556 , n226555 , n226534 );
xor ( n226557 , n226522 , n226528 );
and ( n226558 , n226557 , n226534 );
and ( n226559 , n226522 , n226528 );
or ( n226560 , n226558 , n226559 );
xor ( n226561 , n226094 , n226540 );
xor ( n226562 , n226561 , n226100 );
xor ( n226563 , n226094 , n226540 );
and ( n226564 , n226563 , n226100 );
and ( n226565 , n226094 , n226540 );
or ( n226566 , n226564 , n226565 );
xor ( n226567 , n226550 , n226110 );
xor ( n226568 , n226567 , n226556 );
xor ( n226569 , n226550 , n226110 );
and ( n226570 , n226569 , n226556 );
and ( n226571 , n226550 , n226110 );
or ( n226572 , n226570 , n226571 );
xor ( n226573 , n226116 , n226562 );
xor ( n226574 , n226573 , n226122 );
xor ( n226575 , n226116 , n226562 );
and ( n226576 , n226575 , n226122 );
and ( n226577 , n226116 , n226562 );
or ( n226578 , n226576 , n226577 );
xor ( n226579 , n226568 , n226574 );
xor ( n226580 , n226579 , n226128 );
xor ( n226581 , n226568 , n226574 );
and ( n226582 , n226581 , n226128 );
and ( n226583 , n226568 , n226574 );
or ( n226584 , n226582 , n226583 );
xor ( n226585 , n226381 , n226392 );
and ( n226586 , n226585 , n226403 );
and ( n226587 , n226381 , n226392 );
or ( n226588 , n226586 , n226587 );
xor ( n226589 , n226348 , n226359 );
and ( n226590 , n226589 , n226369 );
and ( n226591 , n226348 , n226359 );
or ( n226592 , n226590 , n226591 );
xor ( n226593 , n226283 , n226284 );
and ( n226594 , n226593 , n226298 );
and ( n226595 , n226283 , n226284 );
or ( n226596 , n226594 , n226595 );
xor ( n226597 , n225749 , n226450 );
and ( n226598 , n226597 , n226455 );
and ( n226599 , n225749 , n226450 );
or ( n226600 , n226598 , n226599 );
xor ( n226601 , n226471 , n226481 );
and ( n226602 , n226601 , n226495 );
and ( n226603 , n226471 , n226481 );
or ( n226604 , n226602 , n226603 );
xor ( n226605 , n226197 , n226427 );
and ( n226606 , n226605 , n226438 );
and ( n226607 , n226197 , n226427 );
or ( n226608 , n226606 , n226607 );
xor ( n226609 , n226509 , n226519 );
and ( n226610 , n226609 , n226104 );
and ( n226611 , n226509 , n226519 );
or ( n226612 , n226610 , n226611 );
not ( n226613 , n220046 );
not ( n226614 , n226207 );
or ( n226615 , n226613 , n226614 );
not ( n226616 , n216929 );
not ( n226617 , n217147 );
or ( n226618 , n226616 , n226617 );
nand ( n226619 , n224881 , n217076 );
nand ( n226620 , n226618 , n226619 );
nand ( n226621 , n226620 , n217388 );
nand ( n226622 , n226615 , n226621 );
not ( n226623 , n225743 );
not ( n226624 , n226212 );
nand ( n226625 , n226624 , n213750 );
not ( n226626 , n226625 );
or ( n226627 , n226623 , n226626 );
nand ( n226628 , n226212 , n213751 );
nand ( n226629 , n226627 , n226628 );
not ( n226630 , n36575 );
nand ( n226631 , n226630 , n36557 );
not ( n226632 , n226631 );
nand ( n226633 , n37561 , n36320 );
and ( n226634 , n37559 , n36340 );
not ( n226635 , n36361 );
not ( n226636 , n36349 );
or ( n226637 , n226635 , n226636 );
nand ( n226638 , n226637 , n36364 );
nor ( n226639 , n226634 , n226638 );
nand ( n226640 , n37695 , n226633 , n226639 );
not ( n226641 , n226640 );
or ( n226642 , n226632 , n226641 );
not ( n226643 , n226631 );
and ( n226644 , n226639 , n226643 );
nand ( n226645 , n226644 , n37695 , n226633 );
nand ( n226646 , n226642 , n226645 );
buf ( n226647 , n226646 );
buf ( n226648 , n226647 );
not ( n226649 , n226648 );
buf ( n226650 , n226649 );
not ( n226651 , n226650 );
and ( n226652 , n226629 , n226651 );
xor ( n226653 , n226622 , n226652 );
not ( n226654 , n223949 );
buf ( n226655 , n216015 );
not ( n226656 , n226655 );
not ( n226657 , n219386 );
or ( n226658 , n226656 , n226657 );
nand ( n226659 , n41165 , n218736 );
nand ( n226660 , n226658 , n226659 );
not ( n226661 , n226660 );
or ( n226662 , n226654 , n226661 );
nand ( n226663 , n226182 , n216619 );
nand ( n226664 , n226662 , n226663 );
xor ( n226665 , n226653 , n226664 );
xor ( n226666 , n226622 , n226652 );
and ( n226667 , n226666 , n226664 );
and ( n226668 , n226622 , n226652 );
or ( n226669 , n226667 , n226668 );
not ( n226670 , n226230 );
not ( n226671 , n218221 );
or ( n226672 , n226670 , n226671 );
not ( n226673 , n41565 );
not ( n226674 , n221214 );
or ( n226675 , n226673 , n226674 );
nand ( n226676 , n218771 , n216543 );
nand ( n226677 , n226675 , n226676 );
nand ( n226678 , n226677 , n218231 );
nand ( n226679 , n226672 , n226678 );
not ( n226680 , n226309 );
not ( n226681 , n219449 );
or ( n226682 , n226680 , n226681 );
not ( n226683 , n225764 );
not ( n226684 , n218876 );
or ( n226685 , n226683 , n226684 );
nand ( n226686 , n220859 , n225769 );
nand ( n226687 , n226685 , n226686 );
nand ( n226688 , n226687 , n218455 );
nand ( n226689 , n226682 , n226688 );
xor ( n226690 , n226679 , n226689 );
not ( n226691 , n226319 );
not ( n226692 , n219435 );
or ( n226693 , n226691 , n226692 );
not ( n226694 , n214837 );
not ( n226695 , n219419 );
or ( n226696 , n226694 , n226695 );
not ( n226697 , n219439 );
not ( n226698 , n214837 );
nand ( n226699 , n226697 , n226698 );
nand ( n226700 , n226696 , n226699 );
nand ( n226701 , n219076 , n226700 );
nand ( n226702 , n226693 , n226701 );
xor ( n226703 , n226690 , n226702 );
xor ( n226704 , n226679 , n226689 );
and ( n226705 , n226704 , n226702 );
and ( n226706 , n226679 , n226689 );
or ( n226707 , n226705 , n226706 );
not ( n226708 , n213912 );
not ( n226709 , n39607 );
and ( n226710 , n213382 , n226709 );
not ( n226711 , n213382 );
not ( n226712 , n39606 );
not ( n226713 , n226712 );
and ( n226714 , n226711 , n226713 );
or ( n226715 , n226710 , n226714 );
not ( n226716 , n226715 );
or ( n226717 , n226708 , n226716 );
nand ( n226718 , n226247 , n217969 );
nand ( n226719 , n226717 , n226718 );
xor ( n226720 , n226592 , n226719 );
not ( n226721 , n216336 );
not ( n226722 , n213735 );
not ( n226723 , n39926 );
not ( n226724 , n226723 );
not ( n226725 , n226724 );
or ( n226726 , n226722 , n226725 );
not ( n226727 , n39927 );
nand ( n226728 , n226727 , n213732 );
nand ( n226729 , n226726 , n226728 );
not ( n226730 , n226729 );
or ( n226731 , n226721 , n226730 );
not ( n226732 , n226261 );
nand ( n226733 , n226732 , n213577 );
nand ( n226734 , n226731 , n226733 );
xor ( n226735 , n226720 , n226734 );
xor ( n226736 , n226592 , n226719 );
and ( n226737 , n226736 , n226734 );
and ( n226738 , n226592 , n226719 );
or ( n226739 , n226737 , n226738 );
xor ( n226740 , n226237 , n226596 );
not ( n226741 , n226367 );
not ( n226742 , n224937 );
not ( n226743 , n226742 );
or ( n226744 , n226741 , n226743 );
not ( n226745 , n224448 );
not ( n226746 , n217044 );
not ( n226747 , n224923 );
not ( n226748 , n226747 );
or ( n226749 , n226746 , n226748 );
nand ( n226750 , n224924 , n215131 );
nand ( n226751 , n226749 , n226750 );
nand ( n226752 , n226745 , n226751 );
nand ( n226753 , n226744 , n226752 );
not ( n226754 , n226281 );
not ( n226755 , n226271 );
not ( n226756 , n226755 );
or ( n226757 , n226754 , n226756 );
and ( n226758 , n225952 , n214134 );
not ( n226759 , n225952 );
and ( n226760 , n226759 , n213583 );
or ( n226761 , n226758 , n226760 );
nand ( n226762 , n225948 , n226761 );
nand ( n226763 , n226757 , n226762 );
xor ( n226764 , n226753 , n226763 );
not ( n226765 , n218762 );
not ( n226766 , n217614 );
not ( n226767 , n215989 );
or ( n226768 , n226766 , n226767 );
nand ( n226769 , n41397 , n221924 );
nand ( n226770 , n226768 , n226769 );
not ( n226771 , n226770 );
or ( n226772 , n226765 , n226771 );
nand ( n226773 , n226169 , n217890 );
nand ( n226774 , n226772 , n226773 );
not ( n226775 , n219501 );
not ( n226776 , n216594 );
not ( n226777 , n217115 );
or ( n226778 , n226776 , n226777 );
nand ( n226779 , n224398 , n220226 );
nand ( n226780 , n226778 , n226779 );
not ( n226781 , n226780 );
or ( n226782 , n226775 , n226781 );
nand ( n226783 , n226191 , n218647 );
nand ( n226784 , n226782 , n226783 );
xor ( n226785 , n226774 , n226784 );
xor ( n226786 , n226764 , n226785 );
xor ( n226787 , n226740 , n226786 );
xor ( n226788 , n226237 , n226596 );
and ( n226789 , n226788 , n226786 );
and ( n226790 , n226237 , n226596 );
or ( n226791 , n226789 , n226790 );
not ( n226792 , n226401 );
not ( n226793 , n222453 );
or ( n226794 , n226792 , n226793 );
not ( n226795 , n216934 );
not ( n226796 , n225418 );
or ( n226797 , n226795 , n226796 );
nand ( n226798 , n222428 , n216940 );
nand ( n226799 , n226797 , n226798 );
nand ( n226800 , n222157 , n226799 );
nand ( n226801 , n226794 , n226800 );
not ( n226802 , n226346 );
not ( n226803 , n225380 );
or ( n226804 , n226802 , n226803 );
not ( n226805 , n215075 );
not ( n226806 , n223182 );
not ( n226807 , n226806 );
or ( n226808 , n226805 , n226807 );
not ( n226809 , n224986 );
nand ( n226810 , n226809 , n215899 );
nand ( n226811 , n226808 , n226810 );
nand ( n226812 , n226811 , n222768 );
nand ( n226813 , n226804 , n226812 );
xor ( n226814 , n226801 , n226813 );
not ( n226815 , n226357 );
not ( n226816 , n224086 );
or ( n226817 , n226815 , n226816 );
and ( n226818 , n224068 , n214678 );
not ( n226819 , n224068 );
and ( n226820 , n226819 , n219475 );
or ( n226821 , n226818 , n226820 );
nand ( n226822 , n224090 , n226821 );
nand ( n226823 , n226817 , n226822 );
xor ( n226824 , n226814 , n226823 );
xor ( n226825 , n226824 , n226703 );
not ( n226826 , n226330 );
not ( n226827 , n220162 );
or ( n226828 , n226826 , n226827 );
not ( n226829 , n215228 );
not ( n226830 , n220147 );
or ( n226831 , n226829 , n226830 );
nand ( n226832 , n225454 , n214820 );
nand ( n226833 , n226831 , n226832 );
nand ( n226834 , n226833 , n219778 );
nand ( n226835 , n226828 , n226834 );
not ( n226836 , n226379 );
not ( n226837 , n223223 );
or ( n226838 , n226836 , n226837 );
not ( n226839 , n41835 );
not ( n226840 , n223227 );
or ( n226841 , n226839 , n226840 );
nand ( n226842 , n220900 , n221494 );
nand ( n226843 , n226841 , n226842 );
nand ( n226844 , n226843 , n220929 );
nand ( n226845 , n226838 , n226844 );
xor ( n226846 , n226835 , n226845 );
not ( n226847 , n226390 );
not ( n226848 , n221625 );
or ( n226849 , n226847 , n226848 );
not ( n226850 , n219343 );
not ( n226851 , n221777 );
or ( n226852 , n226850 , n226851 );
nand ( n226853 , n221608 , n219348 );
nand ( n226854 , n226852 , n226853 );
nand ( n226855 , n226854 , n223587 );
nand ( n226856 , n226849 , n226855 );
xor ( n226857 , n226846 , n226856 );
xor ( n226858 , n226825 , n226857 );
xor ( n226859 , n226824 , n226703 );
and ( n226860 , n226859 , n226857 );
and ( n226861 , n226824 , n226703 );
or ( n226862 , n226860 , n226861 );
xor ( n226863 , n226600 , n226604 );
xor ( n226864 , n226863 , n226608 );
xor ( n226865 , n226600 , n226604 );
and ( n226866 , n226865 , n226608 );
and ( n226867 , n226600 , n226604 );
or ( n226868 , n226866 , n226867 );
not ( n226869 , n215999 );
not ( n226870 , n226649 );
or ( n226871 , n226869 , n226870 );
nand ( n226872 , n226648 , n213751 );
nand ( n226873 , n226871 , n226872 );
not ( n226874 , n226873 );
and ( n226875 , n226647 , n36370 );
not ( n226876 , n226647 );
and ( n226877 , n226876 , n226212 );
nor ( n226878 , n226875 , n226877 );
nand ( n226879 , n226216 , n226878 );
not ( n226880 , n226879 );
buf ( n226881 , n226880 );
not ( n226882 , n226881 );
or ( n226883 , n226874 , n226882 );
buf ( n226884 , n226217 );
not ( n226885 , n226884 );
not ( n226886 , n218224 );
not ( n226887 , n226646 );
buf ( n226888 , n226887 );
not ( n226889 , n226888 );
or ( n226890 , n226886 , n226889 );
nand ( n226891 , n226648 , n216076 );
nand ( n226892 , n226890 , n226891 );
nand ( n226893 , n226885 , n226892 );
nand ( n226894 , n226883 , n226893 );
xor ( n226895 , n226894 , n226201 );
xor ( n226896 , n226895 , n226665 );
not ( n226897 , n216239 );
not ( n226898 , n215113 );
not ( n226899 , n224285 );
or ( n226900 , n226898 , n226899 );
nand ( n226901 , n40545 , n217944 );
nand ( n226902 , n226900 , n226901 );
not ( n226903 , n226902 );
or ( n226904 , n226897 , n226903 );
nand ( n226905 , n226448 , n214717 );
nand ( n226906 , n226904 , n226905 );
not ( n226907 , n219353 );
not ( n226908 , n215955 );
not ( n226909 , n223384 );
or ( n226910 , n226908 , n226909 );
not ( n226911 , n40258 );
nand ( n226912 , n226911 , n216989 );
nand ( n226913 , n226910 , n226912 );
not ( n226914 , n226913 );
or ( n226915 , n226907 , n226914 );
not ( n226916 , n226453 );
nand ( n226917 , n226916 , n217552 );
nand ( n226918 , n226915 , n226917 );
xor ( n226919 , n226906 , n226918 );
not ( n226920 , n222185 );
not ( n226921 , n40668 );
not ( n226922 , n226921 );
not ( n226923 , n226922 );
not ( n226924 , n220538 );
or ( n226925 , n226923 , n226924 );
nand ( n226926 , n221725 , n219033 );
nand ( n226927 , n226925 , n226926 );
not ( n226928 , n226927 );
or ( n226929 , n226920 , n226928 );
nand ( n226930 , n226469 , n219731 );
nand ( n226931 , n226929 , n226930 );
xor ( n226932 , n226919 , n226931 );
xor ( n226933 , n226896 , n226932 );
not ( n226934 , n226292 );
not ( n226935 , n218883 );
or ( n226936 , n226934 , n226935 );
nand ( n226937 , n40710 , n220038 );
nand ( n226938 , n226936 , n226937 );
not ( n226939 , n226938 );
buf ( n226940 , n220032 );
or ( n226941 , n226939 , n226940 );
not ( n226942 , n217486 );
not ( n226943 , n226942 );
nand ( n226944 , n226294 , n226943 );
nand ( n226945 , n226941 , n226944 );
not ( n226946 , n217023 );
not ( n226947 , n226507 );
or ( n226948 , n226946 , n226947 );
not ( n226949 , n219577 );
not ( n226950 , n223321 );
or ( n226951 , n226949 , n226950 );
nand ( n226952 , n221716 , n218661 );
nand ( n226953 , n226951 , n226952 );
nand ( n226954 , n226953 , n219175 );
nand ( n226955 , n226948 , n226954 );
xor ( n226956 , n226945 , n226955 );
not ( n226957 , n218467 );
not ( n226958 , n226422 );
or ( n226959 , n226957 , n226958 );
not ( n226960 , n217573 );
buf ( n226961 , n224272 );
not ( n226962 , n226961 );
or ( n226963 , n226960 , n226962 );
buf ( n226964 , n225111 );
nand ( n226965 , n226964 , n219390 );
nand ( n226966 , n226963 , n226965 );
nand ( n226967 , n226966 , n215137 );
nand ( n226968 , n226959 , n226967 );
xor ( n226969 , n226956 , n226968 );
xor ( n226970 , n226933 , n226969 );
xor ( n226971 , n226896 , n226932 );
and ( n226972 , n226971 , n226969 );
and ( n226973 , n226896 , n226932 );
or ( n226974 , n226972 , n226973 );
xor ( n226975 , n226254 , n226269 );
xor ( n226976 , n226975 , n226612 );
xor ( n226977 , n226254 , n226269 );
and ( n226978 , n226977 , n226612 );
and ( n226979 , n226254 , n226269 );
or ( n226980 , n226978 , n226979 );
not ( n226981 , n216204 );
not ( n226982 , n226479 );
or ( n226983 , n226981 , n226982 );
not ( n226984 , n40624 );
not ( n226985 , n221283 );
and ( n226986 , n226984 , n226985 );
and ( n226987 , n219522 , n221283 );
nor ( n226988 , n226986 , n226987 );
or ( n226989 , n226988 , n223833 );
nand ( n226990 , n226983 , n226989 );
not ( n226991 , n221933 );
not ( n226992 , n221935 );
not ( n226993 , n220204 );
or ( n226994 , n226992 , n226993 );
nand ( n226995 , n218911 , n221938 );
nand ( n226996 , n226994 , n226995 );
not ( n226997 , n226996 );
or ( n226998 , n226991 , n226997 );
nand ( n226999 , n226491 , n215183 );
nand ( n227000 , n226998 , n226999 );
xor ( n227001 , n226990 , n227000 );
not ( n227002 , n214694 );
not ( n227003 , n216810 );
buf ( n227004 , n222512 );
not ( n227005 , n227004 );
or ( n227006 , n227003 , n227005 );
not ( n227007 , n222509 );
nand ( n227008 , n227007 , n221307 );
nand ( n227009 , n227006 , n227008 );
not ( n227010 , n227009 );
or ( n227011 , n227002 , n227010 );
nand ( n227012 , n226434 , n216299 );
nand ( n227013 , n227011 , n227012 );
xor ( n227014 , n227001 , n227013 );
xor ( n227015 , n227014 , n226338 );
not ( n227016 , n217142 );
not ( n227017 , n216262 );
not ( n227018 , n225792 );
or ( n227019 , n227017 , n227018 );
nand ( n227020 , n39713 , n214824 );
nand ( n227021 , n227019 , n227020 );
not ( n227022 , n227021 );
or ( n227023 , n227016 , n227022 );
nand ( n227024 , n226517 , n213874 );
nand ( n227025 , n227023 , n227024 );
xor ( n227026 , n227025 , n226548 );
xor ( n227027 , n227026 , n226588 );
xor ( n227028 , n227015 , n227027 );
xor ( n227029 , n227014 , n226338 );
and ( n227030 , n227029 , n227027 );
and ( n227031 , n227014 , n226338 );
or ( n227032 , n227030 , n227031 );
xor ( n227033 , n226735 , n226410 );
xor ( n227034 , n227033 , n226858 );
xor ( n227035 , n226735 , n226410 );
and ( n227036 , n227035 , n226858 );
and ( n227037 , n226735 , n226410 );
or ( n227038 , n227036 , n227037 );
xor ( n227039 , n226787 , n226864 );
xor ( n227040 , n227039 , n226462 );
xor ( n227041 , n226787 , n226864 );
and ( n227042 , n227041 , n226462 );
and ( n227043 , n226787 , n226864 );
or ( n227044 , n227042 , n227043 );
xor ( n227045 , n226416 , n226526 );
xor ( n227046 , n227045 , n226970 );
xor ( n227047 , n226416 , n226526 );
and ( n227048 , n227047 , n226970 );
and ( n227049 , n226416 , n226526 );
or ( n227050 , n227048 , n227049 );
xor ( n227051 , n226835 , n226845 );
and ( n227052 , n227051 , n226856 );
and ( n227053 , n226835 , n226845 );
or ( n227054 , n227052 , n227053 );
xor ( n227055 , n226976 , n226532 );
xor ( n227056 , n227055 , n227028 );
xor ( n227057 , n226976 , n226532 );
and ( n227058 , n227057 , n227028 );
and ( n227059 , n226976 , n226532 );
or ( n227060 , n227058 , n227059 );
xor ( n227061 , n226538 , n227034 );
xor ( n227062 , n227061 , n227040 );
xor ( n227063 , n226538 , n227034 );
and ( n227064 , n227063 , n227040 );
and ( n227065 , n226538 , n227034 );
or ( n227066 , n227064 , n227065 );
xor ( n227067 , n226544 , n227046 );
xor ( n227068 , n227067 , n226554 );
xor ( n227069 , n226544 , n227046 );
and ( n227070 , n227069 , n226554 );
and ( n227071 , n226544 , n227046 );
or ( n227072 , n227070 , n227071 );
xor ( n227073 , n227056 , n226560 );
xor ( n227074 , n227073 , n227062 );
xor ( n227075 , n227056 , n226560 );
and ( n227076 , n227075 , n227062 );
and ( n227077 , n227056 , n226560 );
or ( n227078 , n227076 , n227077 );
xor ( n227079 , n226566 , n227068 );
xor ( n227080 , n227079 , n226572 );
xor ( n227081 , n226566 , n227068 );
and ( n227082 , n227081 , n226572 );
and ( n227083 , n226566 , n227068 );
or ( n227084 , n227082 , n227083 );
xor ( n227085 , n227074 , n226578 );
xor ( n227086 , n227085 , n227080 );
xor ( n227087 , n227074 , n226578 );
and ( n227088 , n227087 , n227080 );
and ( n227089 , n227074 , n226578 );
or ( n227090 , n227088 , n227089 );
xor ( n227091 , n226801 , n226813 );
and ( n227092 , n227091 , n226823 );
and ( n227093 , n226801 , n226813 );
or ( n227094 , n227092 , n227093 );
xor ( n227095 , n226753 , n226763 );
and ( n227096 , n227095 , n226785 );
and ( n227097 , n226753 , n226763 );
or ( n227098 , n227096 , n227097 );
xor ( n227099 , n226894 , n226201 );
and ( n227100 , n227099 , n226665 );
and ( n227101 , n226894 , n226201 );
or ( n227102 , n227100 , n227101 );
xor ( n227103 , n226906 , n226918 );
and ( n227104 , n227103 , n226931 );
and ( n227105 , n226906 , n226918 );
or ( n227106 , n227104 , n227105 );
xor ( n227107 , n226990 , n227000 );
and ( n227108 , n227107 , n227013 );
and ( n227109 , n226990 , n227000 );
or ( n227110 , n227108 , n227109 );
xor ( n227111 , n226945 , n226955 );
and ( n227112 , n227111 , n226968 );
and ( n227113 , n226945 , n226955 );
or ( n227114 , n227112 , n227113 );
xor ( n227115 , n227025 , n226548 );
and ( n227116 , n227115 , n226588 );
and ( n227117 , n227025 , n226548 );
or ( n227118 , n227116 , n227117 );
not ( n227119 , n226780 );
or ( n227120 , n227119 , n224895 );
not ( n227121 , n219501 );
not ( n227122 , n41069 );
not ( n227123 , n216569 );
and ( n227124 , n227122 , n227123 );
and ( n227125 , n219201 , n216593 );
nor ( n227126 , n227124 , n227125 );
or ( n227127 , n227121 , n227126 );
nand ( n227128 , n227120 , n227127 );
not ( n227129 , n226770 );
not ( n227130 , n220059 );
or ( n227131 , n227129 , n227130 );
not ( n227132 , n218560 );
not ( n227133 , n41318 );
or ( n227134 , n227132 , n227133 );
nand ( n227135 , n217637 , n216306 );
nand ( n227136 , n227134 , n227135 );
not ( n227137 , n227136 );
not ( n227138 , n220067 );
or ( n227139 , n227137 , n227138 );
nand ( n227140 , n227131 , n227139 );
xor ( n227141 , n227128 , n227140 );
not ( n227142 , n217388 );
not ( n227143 , n216929 );
not ( n227144 , n222180 );
or ( n227145 , n227143 , n227144 );
nand ( n227146 , n208164 , n217076 );
nand ( n227147 , n227145 , n227146 );
not ( n227148 , n227147 );
or ( n227149 , n227142 , n227148 );
nand ( n227150 , n226620 , n219368 );
nand ( n227151 , n227149 , n227150 );
xor ( n227152 , n227141 , n227151 );
xor ( n227153 , n227128 , n227140 );
and ( n227154 , n227153 , n227151 );
and ( n227155 , n227128 , n227140 );
or ( n227156 , n227154 , n227155 );
not ( n227157 , n37602 );
not ( n227158 , n227157 );
not ( n227159 , n36582 );
not ( n227160 , n227159 );
or ( n227161 , n227158 , n227160 );
nand ( n227162 , n36582 , n37602 );
nand ( n227163 , n227161 , n227162 );
xor ( n227164 , n226887 , n227163 );
not ( n227165 , n227164 );
and ( n227166 , n227165 , n215999 );
not ( n227167 , n226677 );
not ( n227168 , n219836 );
or ( n227169 , n227167 , n227168 );
not ( n227170 , n215796 );
not ( n227171 , n218226 );
or ( n227172 , n227170 , n227171 );
nand ( n227173 , n218771 , n216261 );
nand ( n227174 , n227172 , n227173 );
nand ( n227175 , n227174 , n218231 );
nand ( n227176 , n227169 , n227175 );
xor ( n227177 , n227166 , n227176 );
not ( n227178 , n226687 );
not ( n227179 , n219449 );
or ( n227180 , n227178 , n227179 );
not ( n227181 , n41701 );
not ( n227182 , n218876 );
or ( n227183 , n227181 , n227182 );
nand ( n227184 , n223671 , n226224 );
nand ( n227185 , n227183 , n227184 );
nand ( n227186 , n218455 , n227185 );
nand ( n227187 , n227180 , n227186 );
xor ( n227188 , n227177 , n227187 );
xor ( n227189 , n227166 , n227176 );
and ( n227190 , n227189 , n227187 );
and ( n227191 , n227166 , n227176 );
or ( n227192 , n227190 , n227191 );
xor ( n227193 , n227054 , n227094 );
xor ( n227194 , n227193 , n227098 );
xor ( n227195 , n227054 , n227094 );
and ( n227196 , n227195 , n227098 );
and ( n227197 , n227054 , n227094 );
or ( n227198 , n227196 , n227197 );
not ( n227199 , n211314 );
not ( n227200 , n213382 );
not ( n227201 , n39088 );
not ( n227202 , n227201 );
or ( n227203 , n227200 , n227202 );
nand ( n227204 , n39088 , n217715 );
nand ( n227205 , n227203 , n227204 );
not ( n227206 , n227205 );
or ( n227207 , n227199 , n227206 );
nand ( n227208 , n226715 , n217969 );
nand ( n227209 , n227207 , n227208 );
not ( n227210 , n217142 );
not ( n227211 , n216262 );
not ( n227212 , n39748 );
or ( n227213 , n227211 , n227212 );
nand ( n227214 , n39747 , n214824 );
nand ( n227215 , n227213 , n227214 );
not ( n227216 , n227215 );
or ( n227217 , n227210 , n227216 );
nand ( n227218 , n227021 , n213874 );
nand ( n227219 , n227217 , n227218 );
xor ( n227220 , n227209 , n227219 );
not ( n227221 , n216336 );
not ( n227222 , n213735 );
buf ( n227223 , n39812 );
not ( n227224 , n227223 );
not ( n227225 , n227224 );
or ( n227226 , n227222 , n227225 );
nand ( n227227 , n227223 , n213732 );
nand ( n227228 , n227226 , n227227 );
not ( n227229 , n227228 );
or ( n227230 , n227221 , n227229 );
nand ( n227231 , n226729 , n213577 );
nand ( n227232 , n227230 , n227231 );
xor ( n227233 , n227220 , n227232 );
xor ( n227234 , n227209 , n227219 );
and ( n227235 , n227234 , n227232 );
and ( n227236 , n227209 , n227219 );
or ( n227237 , n227235 , n227236 );
not ( n227238 , n226892 );
not ( n227239 , n226880 );
or ( n227240 , n227238 , n227239 );
not ( n227241 , n226217 );
not ( n227242 , n213347 );
not ( n227243 , n226649 );
or ( n227244 , n227242 , n227243 );
not ( n227245 , n226888 );
nand ( n227246 , n227245 , n222031 );
nand ( n227247 , n227244 , n227246 );
nand ( n227248 , n227241 , n227247 );
nand ( n227249 , n227240 , n227248 );
and ( n227250 , n226784 , n226774 );
xor ( n227251 , n227249 , n227250 );
not ( n227252 , n223949 );
not ( n227253 , n226655 );
not ( n227254 , n224617 );
or ( n227255 , n227253 , n227254 );
nand ( n227256 , n40724 , n218736 );
nand ( n227257 , n227255 , n227256 );
not ( n227258 , n227257 );
or ( n227259 , n227252 , n227258 );
buf ( n227260 , n216619 );
nand ( n227261 , n226660 , n227260 );
nand ( n227262 , n227259 , n227261 );
xor ( n227263 , n227251 , n227262 );
xor ( n227264 , n227263 , n227188 );
not ( n227265 , n226854 );
not ( n227266 , n221625 );
or ( n227267 , n227265 , n227266 );
not ( n227268 , n221921 );
not ( n227269 , n221777 );
or ( n227270 , n227268 , n227269 );
nand ( n227271 , n221608 , n218980 );
nand ( n227272 , n227270 , n227271 );
nand ( n227273 , n227272 , n221387 );
nand ( n227274 , n227267 , n227273 );
not ( n227275 , n226799 );
not ( n227276 , n222453 );
or ( n227277 , n227275 , n227276 );
not ( n227278 , n219102 );
not ( n227279 , n222458 );
or ( n227280 , n227278 , n227279 );
nand ( n227281 , n222462 , n216139 );
nand ( n227282 , n227280 , n227281 );
nand ( n227283 , n227282 , n222158 );
nand ( n227284 , n227277 , n227283 );
xor ( n227285 , n227274 , n227284 );
not ( n227286 , n223197 );
not ( n227287 , n226811 );
or ( n227288 , n227286 , n227287 );
not ( n227289 , n218514 );
not ( n227290 , n223186 );
or ( n227291 , n227289 , n227290 );
nand ( n227292 , n223182 , n216170 );
nand ( n227293 , n227291 , n227292 );
buf ( n227294 , n222767 );
nand ( n227295 , n227293 , n227294 );
nand ( n227296 , n227288 , n227295 );
xor ( n227297 , n227285 , n227296 );
xor ( n227298 , n227264 , n227297 );
xor ( n227299 , n227263 , n227188 );
and ( n227300 , n227299 , n227297 );
and ( n227301 , n227263 , n227188 );
or ( n227302 , n227300 , n227301 );
not ( n227303 , n226700 );
not ( n227304 , n221575 );
or ( n227305 , n227303 , n227304 );
not ( n227306 , n219689 );
not ( n227307 , n219423 );
or ( n227308 , n227306 , n227307 );
not ( n227309 , n219423 );
nand ( n227310 , n227309 , n208726 );
nand ( n227311 , n227308 , n227310 );
nand ( n227312 , n227311 , n219075 );
nand ( n227313 , n227305 , n227312 );
not ( n227314 , n226833 );
not ( n227315 , n220163 );
or ( n227316 , n227314 , n227315 );
not ( n227317 , n224492 );
not ( n227318 , n222412 );
or ( n227319 , n227317 , n227318 );
not ( n227320 , n220147 );
nand ( n227321 , n227320 , n214642 );
nand ( n227322 , n227319 , n227321 );
nand ( n227323 , n227322 , n220881 );
nand ( n227324 , n227316 , n227323 );
xor ( n227325 , n227313 , n227324 );
not ( n227326 , n223223 );
not ( n227327 , n226843 );
or ( n227328 , n227326 , n227327 );
xor ( n227329 , n220900 , n223658 );
or ( n227330 , n227329 , n220928 );
nand ( n227331 , n227328 , n227330 );
xor ( n227332 , n227325 , n227331 );
not ( n227333 , n226821 );
not ( n227334 , n225839 );
or ( n227335 , n227333 , n227334 );
not ( n227336 , n216208 );
not ( n227337 , n224094 );
or ( n227338 , n227336 , n227337 );
nand ( n227339 , n224067 , n216207 );
nand ( n227340 , n227338 , n227339 );
nand ( n227341 , n223810 , n227340 );
nand ( n227342 , n227335 , n227341 );
not ( n227343 , n226751 );
not ( n227344 , n225851 );
or ( n227345 , n227343 , n227344 );
not ( n227346 , n214537 );
not ( n227347 , n224943 );
or ( n227348 , n227346 , n227347 );
nand ( n227349 , n224924 , n214899 );
nand ( n227350 , n227348 , n227349 );
nand ( n227351 , n227350 , n224449 );
nand ( n227352 , n227345 , n227351 );
xor ( n227353 , n227342 , n227352 );
not ( n227354 , n226761 );
not ( n227355 , n226755 );
or ( n227356 , n227354 , n227355 );
and ( n227357 , n225952 , n214960 );
not ( n227358 , n225952 );
and ( n227359 , n227358 , n214956 );
or ( n227360 , n227357 , n227359 );
nand ( n227361 , n225948 , n227360 );
nand ( n227362 , n227356 , n227361 );
xor ( n227363 , n227353 , n227362 );
xor ( n227364 , n227332 , n227363 );
xor ( n227365 , n227364 , n227106 );
xor ( n227366 , n227332 , n227363 );
and ( n227367 , n227366 , n227106 );
and ( n227368 , n227332 , n227363 );
or ( n227369 , n227367 , n227368 );
xor ( n227370 , n227102 , n227110 );
xor ( n227371 , n227370 , n227114 );
xor ( n227372 , n227102 , n227110 );
and ( n227373 , n227372 , n227114 );
and ( n227374 , n227102 , n227110 );
or ( n227375 , n227373 , n227374 );
not ( n227376 , n220414 );
not ( n227377 , n226938 );
or ( n227378 , n227376 , n227377 );
not ( n227379 , n226292 );
not ( n227380 , n40766 );
or ( n227381 , n227379 , n227380 );
nand ( n227382 , n219239 , n220038 );
nand ( n227383 , n227381 , n227382 );
nand ( n227384 , n227383 , n220033 );
nand ( n227385 , n227378 , n227384 );
not ( n227386 , n217023 );
not ( n227387 , n226953 );
or ( n227388 , n227386 , n227387 );
not ( n227389 , n219577 );
not ( n227390 , n222951 );
or ( n227391 , n227389 , n227390 );
nand ( n227392 , n222955 , n218661 );
nand ( n227393 , n227391 , n227392 );
nand ( n227394 , n227393 , n219175 );
nand ( n227395 , n227388 , n227394 );
xor ( n227396 , n227385 , n227395 );
not ( n227397 , n220985 );
and ( n227398 , n223764 , n221338 );
not ( n227399 , n223764 );
and ( n227400 , n227399 , n216037 );
or ( n227401 , n227398 , n227400 );
not ( n227402 , n227401 );
or ( n227403 , n227397 , n227402 );
nand ( n227404 , n226902 , n214717 );
nand ( n227405 , n227403 , n227404 );
xor ( n227406 , n227396 , n227405 );
xor ( n227407 , n227406 , n227118 );
xor ( n227408 , n227407 , n226739 );
xor ( n227409 , n227406 , n227118 );
and ( n227410 , n227409 , n226739 );
and ( n227411 , n227406 , n227118 );
or ( n227412 , n227410 , n227411 );
not ( n227413 , n220272 );
not ( n227414 , n217542 );
not ( n227415 , n222121 );
or ( n227416 , n227414 , n227415 );
nand ( n227417 , n40397 , n219358 );
nand ( n227418 , n227416 , n227417 );
not ( n227419 , n227418 );
or ( n227420 , n227413 , n227419 );
nand ( n227421 , n226913 , n220280 );
nand ( n227422 , n227420 , n227421 );
not ( n227423 , n218678 );
not ( n227424 , n226927 );
or ( n227425 , n227423 , n227424 );
not ( n227426 , n216166 );
not ( n227427 , n220599 );
or ( n227428 , n227426 , n227427 );
nand ( n227429 , n40409 , n220538 );
nand ( n227430 , n227428 , n227429 );
nand ( n227431 , n227430 , n222185 );
nand ( n227432 , n227425 , n227431 );
xor ( n227433 , n227422 , n227432 );
xor ( n227434 , n227433 , n227152 );
not ( n227435 , n219314 );
not ( n227436 , n219687 );
not ( n227437 , n220581 );
or ( n227438 , n227436 , n227437 );
nand ( n227439 , n207936 , n222323 );
nand ( n227440 , n227438 , n227439 );
not ( n227441 , n227440 );
or ( n227442 , n227435 , n227441 );
not ( n227443 , n226988 );
nand ( n227444 , n227443 , n224624 );
nand ( n227445 , n227442 , n227444 );
not ( n227446 , n221933 );
not ( n227447 , n221935 );
not ( n227448 , n219226 );
not ( n227449 , n227448 );
or ( n227450 , n227447 , n227449 );
nand ( n227451 , n219222 , n221938 );
nand ( n227452 , n227450 , n227451 );
not ( n227453 , n227452 );
or ( n227454 , n227446 , n227453 );
nand ( n227455 , n226996 , n215183 );
nand ( n227456 , n227454 , n227455 );
xor ( n227457 , n227445 , n227456 );
not ( n227458 , n216562 );
not ( n227459 , n227009 );
or ( n227460 , n227458 , n227459 );
not ( n227461 , n216810 );
not ( n227462 , n222940 );
or ( n227463 , n227461 , n227462 );
nand ( n227464 , n40485 , n215289 );
nand ( n227465 , n227463 , n227464 );
nand ( n227466 , n227465 , n214694 );
nand ( n227467 , n227460 , n227466 );
xor ( n227468 , n227457 , n227467 );
xor ( n227469 , n227434 , n227468 );
xor ( n227470 , n227469 , n226791 );
xor ( n227471 , n227434 , n227468 );
and ( n227472 , n227471 , n226791 );
and ( n227473 , n227434 , n227468 );
or ( n227474 , n227472 , n227473 );
not ( n227475 , n215137 );
not ( n227476 , n213960 );
not ( n227477 , n39878 );
not ( n227478 , n227477 );
or ( n227479 , n227476 , n227478 );
nand ( n227480 , n225344 , n215388 );
nand ( n227481 , n227479 , n227480 );
not ( n227482 , n227481 );
or ( n227483 , n227475 , n227482 );
nand ( n227484 , n226966 , n214086 );
nand ( n227485 , n227483 , n227484 );
xor ( n227486 , n226669 , n227485 );
xor ( n227487 , n227486 , n226707 );
xor ( n227488 , n227194 , n227487 );
xor ( n227489 , n227488 , n227233 );
xor ( n227490 , n227194 , n227487 );
and ( n227491 , n227490 , n227233 );
and ( n227492 , n227194 , n227487 );
or ( n227493 , n227491 , n227492 );
xor ( n227494 , n226862 , n226868 );
xor ( n227495 , n227494 , n227365 );
xor ( n227496 , n226862 , n226868 );
and ( n227497 , n227496 , n227365 );
and ( n227498 , n226862 , n226868 );
or ( n227499 , n227497 , n227498 );
xor ( n227500 , n227298 , n226980 );
xor ( n227501 , n227500 , n227371 );
xor ( n227502 , n227298 , n226980 );
and ( n227503 , n227502 , n227371 );
and ( n227504 , n227298 , n226980 );
or ( n227505 , n227503 , n227504 );
xor ( n227506 , n227313 , n227324 );
and ( n227507 , n227506 , n227331 );
and ( n227508 , n227313 , n227324 );
or ( n227509 , n227507 , n227508 );
xor ( n227510 , n226974 , n227032 );
xor ( n227511 , n227510 , n227470 );
xor ( n227512 , n226974 , n227032 );
and ( n227513 , n227512 , n227470 );
and ( n227514 , n226974 , n227032 );
or ( n227515 , n227513 , n227514 );
xor ( n227516 , n227408 , n227038 );
xor ( n227517 , n227516 , n227489 );
xor ( n227518 , n227408 , n227038 );
and ( n227519 , n227518 , n227489 );
and ( n227520 , n227408 , n227038 );
or ( n227521 , n227519 , n227520 );
xor ( n227522 , n227495 , n227044 );
xor ( n227523 , n227522 , n227050 );
xor ( n227524 , n227495 , n227044 );
and ( n227525 , n227524 , n227050 );
and ( n227526 , n227495 , n227044 );
or ( n227527 , n227525 , n227526 );
xor ( n227528 , n227501 , n227511 );
xor ( n227529 , n227528 , n227060 );
xor ( n227530 , n227501 , n227511 );
and ( n227531 , n227530 , n227060 );
and ( n227532 , n227501 , n227511 );
or ( n227533 , n227531 , n227532 );
xor ( n227534 , n227517 , n227523 );
xor ( n227535 , n227534 , n227066 );
xor ( n227536 , n227517 , n227523 );
and ( n227537 , n227536 , n227066 );
and ( n227538 , n227517 , n227523 );
or ( n227539 , n227537 , n227538 );
xor ( n227540 , n227072 , n227529 );
xor ( n227541 , n227540 , n227078 );
xor ( n227542 , n227072 , n227529 );
and ( n227543 , n227542 , n227078 );
and ( n227544 , n227072 , n227529 );
or ( n227545 , n227543 , n227544 );
xor ( n227546 , n227535 , n227084 );
xor ( n227547 , n227546 , n227541 );
xor ( n227548 , n227535 , n227084 );
and ( n227549 , n227548 , n227541 );
and ( n227550 , n227535 , n227084 );
or ( n227551 , n227549 , n227550 );
xor ( n227552 , n227274 , n227284 );
and ( n227553 , n227552 , n227296 );
and ( n227554 , n227274 , n227284 );
or ( n227555 , n227553 , n227554 );
xor ( n227556 , n227342 , n227352 );
and ( n227557 , n227556 , n227362 );
and ( n227558 , n227342 , n227352 );
or ( n227559 , n227557 , n227558 );
xor ( n227560 , n227249 , n227250 );
and ( n227561 , n227560 , n227262 );
and ( n227562 , n227249 , n227250 );
or ( n227563 , n227561 , n227562 );
xor ( n227564 , n227422 , n227432 );
and ( n227565 , n227564 , n227152 );
and ( n227566 , n227422 , n227432 );
or ( n227567 , n227565 , n227566 );
xor ( n227568 , n227445 , n227456 );
and ( n227569 , n227568 , n227467 );
and ( n227570 , n227445 , n227456 );
or ( n227571 , n227569 , n227570 );
xor ( n227572 , n227385 , n227395 );
and ( n227573 , n227572 , n227405 );
and ( n227574 , n227385 , n227395 );
or ( n227575 , n227573 , n227574 );
xor ( n227576 , n226669 , n227485 );
and ( n227577 , n227576 , n226707 );
and ( n227578 , n226669 , n227485 );
or ( n227579 , n227577 , n227578 );
not ( n227580 , n226648 );
not ( n227581 , n227157 );
not ( n227582 , n227159 );
or ( n227583 , n227581 , n227582 );
nand ( n227584 , n227583 , n227162 );
buf ( n227585 , n227584 );
nand ( n227586 , n227585 , n213750 );
nand ( n227587 , n227580 , n227586 );
not ( n227588 , n227585 );
nand ( n227589 , n227588 , n213751 );
and ( n227590 , n227587 , n227589 );
and ( n227591 , n36946 , n37441 );
nand ( n227592 , n37557 , n224427 );
nand ( n227593 , n227592 , n37099 , n37451 );
xor ( n227594 , n227591 , n227593 );
buf ( n227595 , n227594 );
not ( n227596 , n227595 );
nor ( n227597 , n227590 , n227596 );
not ( n227598 , n221559 );
not ( n227599 , n216422 );
not ( n227600 , n227599 );
and ( n227601 , n227598 , n227600 );
not ( n227602 , n216422 );
and ( n227603 , n41165 , n227602 );
nor ( n227604 , n227601 , n227603 );
not ( n227605 , n216598 );
or ( n227606 , n227604 , n227605 );
not ( n227607 , n227126 );
nand ( n227608 , n227607 , n224896 );
nand ( n227609 , n227606 , n227608 );
xor ( n227610 , n227597 , n227609 );
not ( n227611 , n227174 );
or ( n227612 , n218220 , n227611 );
and ( n227613 , n41396 , n218204 );
not ( n227614 , n41396 );
and ( n227615 , n227614 , n218217 );
or ( n227616 , n227613 , n227615 );
not ( n227617 , n227616 );
or ( n227618 , n227617 , n217936 );
nand ( n227619 , n227612 , n227618 );
xor ( n227620 , n227610 , n227619 );
xor ( n227621 , n227597 , n227609 );
and ( n227622 , n227621 , n227619 );
and ( n227623 , n227597 , n227609 );
or ( n227624 , n227622 , n227623 );
not ( n227625 , n227185 );
not ( n227626 , n218835 );
or ( n227627 , n227625 , n227626 );
not ( n227628 , n41564 );
not ( n227629 , n218814 );
or ( n227630 , n227628 , n227629 );
not ( n227631 , n218875 );
nand ( n227632 , n227631 , n216543 );
nand ( n227633 , n227630 , n227632 );
nand ( n227634 , n218455 , n227633 );
nand ( n227635 , n227627 , n227634 );
not ( n227636 , n227311 );
not ( n227637 , n223620 );
or ( n227638 , n227636 , n227637 );
not ( n227639 , n217066 );
not ( n227640 , n227639 );
not ( n227641 , n219440 );
or ( n227642 , n227640 , n227641 );
nand ( n227643 , n221227 , n225763 );
nand ( n227644 , n227642 , n227643 );
nand ( n227645 , n219076 , n227644 );
nand ( n227646 , n227638 , n227645 );
xor ( n227647 , n227635 , n227646 );
not ( n227648 , n227322 );
not ( n227649 , n220163 );
or ( n227650 , n227648 , n227649 );
and ( n227651 , n214834 , n224562 );
not ( n227652 , n214834 );
and ( n227653 , n227652 , n220146 );
or ( n227654 , n227651 , n227653 );
not ( n227655 , n227654 );
nand ( n227656 , n227655 , n219779 );
nand ( n227657 , n227650 , n227656 );
xor ( n227658 , n227647 , n227657 );
xor ( n227659 , n227635 , n227646 );
and ( n227660 , n227659 , n227657 );
and ( n227661 , n227635 , n227646 );
or ( n227662 , n227660 , n227661 );
not ( n227663 , n213784 );
not ( n227664 , n227205 );
or ( n227665 , n227663 , n227664 );
not ( n227666 , n213382 );
not ( n227667 , n38531 );
not ( n227668 , n227667 );
or ( n227669 , n227666 , n227668 );
nand ( n227670 , n38531 , n217715 );
nand ( n227671 , n227669 , n227670 );
nand ( n227672 , n227671 , n213912 );
nand ( n227673 , n227665 , n227672 );
xor ( n227674 , n227559 , n227673 );
not ( n227675 , n213874 );
not ( n227676 , n227215 );
or ( n227677 , n227675 , n227676 );
and ( n227678 , n39606 , n214824 );
not ( n227679 , n39606 );
and ( n227680 , n227679 , n216262 );
or ( n227681 , n227678 , n227680 );
nand ( n227682 , n227681 , n217142 );
nand ( n227683 , n227677 , n227682 );
xor ( n227684 , n227674 , n227683 );
xor ( n227685 , n227559 , n227673 );
and ( n227686 , n227685 , n227683 );
and ( n227687 , n227559 , n227673 );
or ( n227688 , n227686 , n227687 );
not ( n227689 , n213577 );
not ( n227690 , n227228 );
or ( n227691 , n227689 , n227690 );
not ( n227692 , n213735 );
not ( n227693 , n39713 );
not ( n227694 , n227693 );
or ( n227695 , n227692 , n227694 );
not ( n227696 , n225792 );
nand ( n227697 , n227696 , n213732 );
nand ( n227698 , n227695 , n227697 );
nand ( n227699 , n227698 , n216336 );
nand ( n227700 , n227691 , n227699 );
xor ( n227701 , n227620 , n227700 );
xor ( n227702 , n227701 , n227563 );
xor ( n227703 , n227620 , n227700 );
and ( n227704 , n227703 , n227563 );
and ( n227705 , n227620 , n227700 );
or ( n227706 , n227704 , n227705 );
not ( n227707 , n227360 );
not ( n227708 , n225945 );
or ( n227709 , n227707 , n227708 );
not ( n227710 , n225316 );
and ( n227711 , n225952 , n215131 );
not ( n227712 , n225952 );
and ( n227713 , n227712 , n217044 );
or ( n227714 , n227711 , n227713 );
nand ( n227715 , n227710 , n227714 );
nand ( n227716 , n227709 , n227715 );
not ( n227717 , n213751 );
not ( n227718 , n227595 );
or ( n227719 , n227717 , n227718 );
nand ( n227720 , n227596 , n213750 );
nand ( n227721 , n227719 , n227720 );
not ( n227722 , n227721 );
not ( n227723 , n227594 );
not ( n227724 , n227584 );
and ( n227725 , n227723 , n227724 );
not ( n227726 , n227723 );
and ( n227727 , n227726 , n227584 );
nor ( n227728 , n227725 , n227727 );
and ( n227729 , n226647 , n227724 );
not ( n227730 , n226647 );
and ( n227731 , n227730 , n227163 );
nor ( n227732 , n227729 , n227731 );
nand ( n227733 , n227728 , n227732 );
not ( n227734 , n227733 );
not ( n227735 , n227734 );
or ( n227736 , n227722 , n227735 );
not ( n227737 , n227164 );
and ( n227738 , n227595 , n213077 );
not ( n227739 , n227595 );
and ( n227740 , n227739 , n218224 );
or ( n227741 , n227738 , n227740 );
nand ( n227742 , n227737 , n227741 );
nand ( n227743 , n227736 , n227742 );
xor ( n227744 , n227716 , n227743 );
not ( n227745 , n217388 );
not ( n227746 , n217080 );
not ( n227747 , n208259 );
not ( n227748 , n227747 );
or ( n227749 , n227746 , n227748 );
nand ( n227750 , n208259 , n217602 );
nand ( n227751 , n227749 , n227750 );
not ( n227752 , n227751 );
or ( n227753 , n227745 , n227752 );
nand ( n227754 , n227147 , n219368 );
nand ( n227755 , n227753 , n227754 );
not ( n227756 , n217890 );
not ( n227757 , n227136 );
or ( n227758 , n227756 , n227757 );
not ( n227759 , n221923 );
not ( n227760 , n41249 );
or ( n227761 , n227759 , n227760 );
nand ( n227762 , n218283 , n217611 );
nand ( n227763 , n227761 , n227762 );
nand ( n227764 , n227763 , n217641 );
nand ( n227765 , n227758 , n227764 );
xor ( n227766 , n227755 , n227765 );
xor ( n227767 , n227744 , n227766 );
xor ( n227768 , n227658 , n227767 );
not ( n227769 , n227293 );
not ( n227770 , n223197 );
or ( n227771 , n227769 , n227770 );
not ( n227772 , n216934 );
not ( n227773 , n225914 );
or ( n227774 , n227772 , n227773 );
nand ( n227775 , n223182 , n216940 );
nand ( n227776 , n227774 , n227775 );
nand ( n227777 , n222769 , n227776 );
nand ( n227778 , n227771 , n227777 );
not ( n227779 , n227340 );
not ( n227780 , n224087 );
or ( n227781 , n227779 , n227780 );
buf ( n227782 , n224090 );
not ( n227783 , n215075 );
not ( n227784 , n224069 );
or ( n227785 , n227783 , n227784 );
nand ( n227786 , n224974 , n215899 );
nand ( n227787 , n227785 , n227786 );
nand ( n227788 , n227782 , n227787 );
nand ( n227789 , n227781 , n227788 );
xor ( n227790 , n227778 , n227789 );
not ( n227791 , n227350 );
buf ( n227792 , n226742 );
not ( n227793 , n227792 );
or ( n227794 , n227791 , n227793 );
not ( n227795 , n219475 );
not ( n227796 , n224844 );
or ( n227797 , n227795 , n227796 );
nand ( n227798 , n224843 , n214678 );
nand ( n227799 , n227797 , n227798 );
nand ( n227800 , n224941 , n227799 );
nand ( n227801 , n227794 , n227800 );
xor ( n227802 , n227790 , n227801 );
xor ( n227803 , n227768 , n227802 );
xor ( n227804 , n227658 , n227767 );
and ( n227805 , n227804 , n227802 );
and ( n227806 , n227658 , n227767 );
or ( n227807 , n227805 , n227806 );
not ( n227808 , n220929 );
not ( n227809 , n215228 );
not ( n227810 , n220904 );
or ( n227811 , n227809 , n227810 );
nand ( n227812 , n226377 , n214820 );
nand ( n227813 , n227811 , n227812 );
not ( n227814 , n227813 );
or ( n227815 , n227808 , n227814 );
not ( n227816 , n227329 );
nand ( n227817 , n227816 , n223223 );
nand ( n227818 , n227815 , n227817 );
not ( n227819 , n221626 );
not ( n227820 , n227272 );
or ( n227821 , n227819 , n227820 );
not ( n227822 , n221495 );
not ( n227823 , n221777 );
or ( n227824 , n227822 , n227823 );
nand ( n227825 , n221608 , n220022 );
nand ( n227826 , n227824 , n227825 );
nand ( n227827 , n221387 , n227826 );
nand ( n227828 , n227821 , n227827 );
xor ( n227829 , n227818 , n227828 );
not ( n227830 , n227282 );
not ( n227831 , n222454 );
or ( n227832 , n227830 , n227831 );
not ( n227833 , n219343 );
not ( n227834 , n222429 );
or ( n227835 , n227833 , n227834 );
nand ( n227836 , n222428 , n223269 );
nand ( n227837 , n227835 , n227836 );
nand ( n227838 , n222467 , n227837 );
nand ( n227839 , n227832 , n227838 );
xor ( n227840 , n227829 , n227839 );
xor ( n227841 , n227840 , n227575 );
xor ( n227842 , n227841 , n227567 );
xor ( n227843 , n227840 , n227575 );
and ( n227844 , n227843 , n227567 );
and ( n227845 , n227840 , n227575 );
or ( n227846 , n227844 , n227845 );
not ( n227847 , n227247 );
buf ( n227848 , n226879 );
not ( n227849 , n227848 );
not ( n227850 , n227849 );
or ( n227851 , n227847 , n227850 );
buf ( n227852 , n226218 );
not ( n227853 , n213583 );
not ( n227854 , n226650 );
or ( n227855 , n227853 , n227854 );
nand ( n227856 , n226648 , n214134 );
nand ( n227857 , n227855 , n227856 );
nand ( n227858 , n227852 , n227857 );
nand ( n227859 , n227851 , n227858 );
xor ( n227860 , n227859 , n227156 );
not ( n227861 , n227418 );
or ( n227862 , n227861 , n217551 );
not ( n227863 , n217542 );
not ( n227864 , n221711 );
or ( n227865 , n227863 , n227864 );
nand ( n227866 , n40180 , n219358 );
nand ( n227867 , n227865 , n227866 );
not ( n227868 , n227867 );
or ( n227869 , n227868 , n217549 );
nand ( n227870 , n227862 , n227869 );
xor ( n227871 , n227860 , n227870 );
xor ( n227872 , n227571 , n227871 );
not ( n227873 , n214717 );
not ( n227874 , n227401 );
or ( n227875 , n227873 , n227874 );
not ( n227876 , n221338 );
not ( n227877 , n224272 );
or ( n227878 , n227876 , n227877 );
nand ( n227879 , n39995 , n216037 );
nand ( n227880 , n227878 , n227879 );
nand ( n227881 , n227880 , n216239 );
nand ( n227882 , n227875 , n227881 );
not ( n227883 , n216299 );
not ( n227884 , n227465 );
or ( n227885 , n227883 , n227884 );
not ( n227886 , n215290 );
not ( n227887 , n40546 );
or ( n227888 , n227886 , n227887 );
nand ( n227889 , n40545 , n215289 );
nand ( n227890 , n227888 , n227889 );
nand ( n227891 , n227890 , n220820 );
nand ( n227892 , n227885 , n227891 );
xor ( n227893 , n227882 , n227892 );
not ( n227894 , n218467 );
not ( n227895 , n227481 );
or ( n227896 , n227894 , n227895 );
not ( n227897 , n217573 );
not ( n227898 , n39927 );
or ( n227899 , n227897 , n227898 );
not ( n227900 , n39926 );
nand ( n227901 , n227900 , n217397 );
nand ( n227902 , n227899 , n227901 );
nand ( n227903 , n227902 , n215383 );
nand ( n227904 , n227896 , n227903 );
xor ( n227905 , n227893 , n227904 );
xor ( n227906 , n227872 , n227905 );
xor ( n227907 , n227571 , n227871 );
and ( n227908 , n227907 , n227905 );
and ( n227909 , n227571 , n227871 );
or ( n227910 , n227908 , n227909 );
not ( n227911 , n226287 );
not ( n227912 , n220038 );
not ( n227913 , n227912 );
not ( n227914 , n219532 );
or ( n227915 , n227913 , n227914 );
buf ( n227916 , n208078 );
nand ( n227917 , n227916 , n220038 );
nand ( n227918 , n227915 , n227917 );
not ( n227919 , n227918 );
or ( n227920 , n227911 , n227919 );
nand ( n227921 , n227383 , n226943 );
nand ( n227922 , n227920 , n227921 );
not ( n227923 , n223949 );
not ( n227924 , n226655 );
not ( n227925 , n218268 );
or ( n227926 , n227924 , n227925 );
not ( n227927 , n226655 );
nand ( n227928 , n218882 , n227927 );
nand ( n227929 , n227926 , n227928 );
not ( n227930 , n227929 );
or ( n227931 , n227923 , n227930 );
nand ( n227932 , n227257 , n227260 );
nand ( n227933 , n227931 , n227932 );
xor ( n227934 , n227922 , n227933 );
not ( n227935 , n227393 );
or ( n227936 , n227935 , n217367 );
not ( n227937 , n217017 );
not ( n227938 , n222512 );
or ( n227939 , n227937 , n227938 );
nand ( n227940 , n40414 , n215971 );
nand ( n227941 , n227939 , n227940 );
not ( n227942 , n227941 );
not ( n227943 , n219175 );
or ( n227944 , n227942 , n227943 );
nand ( n227945 , n227936 , n227944 );
xor ( n227946 , n227934 , n227945 );
xor ( n227947 , n227237 , n227946 );
xor ( n227948 , n227947 , n227579 );
xor ( n227949 , n227237 , n227946 );
and ( n227950 , n227949 , n227579 );
and ( n227951 , n227237 , n227946 );
or ( n227952 , n227950 , n227951 );
not ( n227953 , n222185 );
and ( n227954 , n40258 , n219033 );
not ( n227955 , n40258 );
and ( n227956 , n227955 , n220538 );
or ( n227957 , n227954 , n227956 );
not ( n227958 , n227957 );
or ( n227959 , n227953 , n227958 );
nand ( n227960 , n227430 , n219731 );
nand ( n227961 , n227959 , n227960 );
not ( n227962 , n216204 );
not ( n227963 , n227440 );
or ( n227964 , n227962 , n227963 );
not ( n227965 , n219687 );
not ( n227966 , n222500 );
or ( n227967 , n227965 , n227966 );
nand ( n227968 , n40668 , n222323 );
nand ( n227969 , n227967 , n227968 );
nand ( n227970 , n227969 , n219314 );
nand ( n227971 , n227964 , n227970 );
xor ( n227972 , n227961 , n227971 );
not ( n227973 , n221933 );
not ( n227974 , n221935 );
not ( n227975 , n219521 );
or ( n227976 , n227974 , n227975 );
nand ( n227977 , n40624 , n222333 );
nand ( n227978 , n227976 , n227977 );
not ( n227979 , n227978 );
or ( n227980 , n227973 , n227979 );
nand ( n227981 , n227452 , n215183 );
nand ( n227982 , n227980 , n227981 );
xor ( n227983 , n227972 , n227982 );
xor ( n227984 , n227983 , n227198 );
xor ( n227985 , n227984 , n227302 );
xor ( n227986 , n227983 , n227198 );
and ( n227987 , n227986 , n227302 );
and ( n227988 , n227983 , n227198 );
or ( n227989 , n227987 , n227988 );
xor ( n227990 , n227192 , n227509 );
xor ( n227991 , n227990 , n227555 );
xor ( n227992 , n227684 , n227991 );
xor ( n227993 , n227992 , n227702 );
xor ( n227994 , n227684 , n227991 );
and ( n227995 , n227994 , n227702 );
and ( n227996 , n227684 , n227991 );
or ( n227997 , n227995 , n227996 );
xor ( n227998 , n227803 , n227375 );
xor ( n227999 , n227998 , n227369 );
xor ( n228000 , n227803 , n227375 );
and ( n228001 , n228000 , n227369 );
and ( n228002 , n227803 , n227375 );
or ( n228003 , n228001 , n228002 );
xor ( n228004 , n227842 , n227412 );
xor ( n228005 , n228004 , n227906 );
xor ( n228006 , n227842 , n227412 );
and ( n228007 , n228006 , n227906 );
and ( n228008 , n227842 , n227412 );
or ( n228009 , n228007 , n228008 );
xor ( n228010 , n227818 , n227828 );
and ( n228011 , n228010 , n227839 );
and ( n228012 , n227818 , n227828 );
or ( n228013 , n228011 , n228012 );
xor ( n228014 , n227985 , n227474 );
xor ( n228015 , n228014 , n227948 );
xor ( n228016 , n227985 , n227474 );
and ( n228017 , n228016 , n227948 );
and ( n228018 , n227985 , n227474 );
or ( n228019 , n228017 , n228018 );
xor ( n228020 , n227493 , n227993 );
xor ( n228021 , n228020 , n227499 );
xor ( n228022 , n227493 , n227993 );
and ( n228023 , n228022 , n227499 );
and ( n228024 , n227493 , n227993 );
or ( n228025 , n228023 , n228024 );
xor ( n228026 , n227505 , n227999 );
xor ( n228027 , n228026 , n228005 );
xor ( n228028 , n227505 , n227999 );
and ( n228029 , n228028 , n228005 );
and ( n228030 , n227505 , n227999 );
or ( n228031 , n228029 , n228030 );
xor ( n228032 , n227515 , n227521 );
xor ( n228033 , n228032 , n228015 );
xor ( n228034 , n227515 , n227521 );
and ( n228035 , n228034 , n228015 );
and ( n228036 , n227515 , n227521 );
or ( n228037 , n228035 , n228036 );
xor ( n228038 , n228021 , n227527 );
xor ( n228039 , n228038 , n228027 );
xor ( n228040 , n228021 , n227527 );
and ( n228041 , n228040 , n228027 );
and ( n228042 , n228021 , n227527 );
or ( n228043 , n228041 , n228042 );
xor ( n228044 , n227533 , n228033 );
xor ( n228045 , n228044 , n227539 );
xor ( n228046 , n227533 , n228033 );
and ( n228047 , n228046 , n227539 );
and ( n228048 , n227533 , n228033 );
or ( n228049 , n228047 , n228048 );
xor ( n228050 , n228039 , n228045 );
xor ( n228051 , n228050 , n227545 );
xor ( n228052 , n228039 , n228045 );
and ( n228053 , n228052 , n227545 );
and ( n228054 , n228039 , n228045 );
or ( n228055 , n228053 , n228054 );
xor ( n228056 , n227778 , n227789 );
and ( n228057 , n228056 , n227801 );
and ( n228058 , n227778 , n227789 );
or ( n228059 , n228057 , n228058 );
xor ( n228060 , n227716 , n227743 );
and ( n228061 , n228060 , n227766 );
and ( n228062 , n227716 , n227743 );
or ( n228063 , n228061 , n228062 );
xor ( n228064 , n227859 , n227156 );
and ( n228065 , n228064 , n227870 );
and ( n228066 , n227859 , n227156 );
or ( n228067 , n228065 , n228066 );
xor ( n228068 , n227961 , n227971 );
and ( n228069 , n228068 , n227982 );
and ( n228070 , n227961 , n227971 );
or ( n228071 , n228069 , n228070 );
xor ( n228072 , n227922 , n227933 );
and ( n228073 , n228072 , n227945 );
and ( n228074 , n227922 , n227933 );
or ( n228075 , n228073 , n228074 );
xor ( n228076 , n227882 , n227892 );
and ( n228077 , n228076 , n227904 );
and ( n228078 , n227882 , n227892 );
or ( n228079 , n228077 , n228078 );
xor ( n228080 , n227192 , n227509 );
and ( n228081 , n228080 , n227555 );
and ( n228082 , n227192 , n227509 );
or ( n228083 , n228081 , n228082 );
not ( n228084 , n218544 );
not ( n228085 , n227751 );
or ( n228086 , n228084 , n228085 );
and ( n228087 , n41068 , n217602 );
not ( n228088 , n41068 );
and ( n228089 , n228088 , n216929 );
or ( n228090 , n228087 , n228089 );
nand ( n228091 , n228090 , n217099 );
nand ( n228092 , n228086 , n228091 );
not ( n228093 , n217890 );
not ( n228094 , n227763 );
or ( n228095 , n228093 , n228094 );
not ( n228096 , n221923 );
not ( n228097 , n216858 );
or ( n228098 , n228096 , n228097 );
or ( n228099 , n225323 , n224850 );
nand ( n228100 , n228098 , n228099 );
nand ( n228101 , n228100 , n218762 );
nand ( n228102 , n228095 , n228101 );
xor ( n228103 , n228092 , n228102 );
not ( n228104 , n37603 );
nand ( n228105 , n36960 , n37691 , n37445 );
not ( n228106 , n228105 );
or ( n228107 , n228104 , n228106 );
not ( n228108 , n37603 );
nand ( n228109 , n228108 , n36960 , n37691 , n37445 );
nand ( n228110 , n228107 , n228109 );
not ( n228111 , n228110 );
and ( n228112 , n227594 , n228111 );
not ( n228113 , n227594 );
and ( n228114 , n228113 , n228110 );
nor ( n228115 , n228112 , n228114 );
buf ( n228116 , n228115 );
nor ( n228117 , n228116 , n213751 );
xor ( n228118 , n228103 , n228117 );
xor ( n228119 , n228092 , n228102 );
and ( n228120 , n228119 , n228117 );
and ( n228121 , n228092 , n228102 );
or ( n228122 , n228120 , n228121 );
not ( n228123 , n227616 );
not ( n228124 , n218219 );
not ( n228125 , n228124 );
or ( n228126 , n228123 , n228125 );
not ( n228127 , n217935 );
not ( n228128 , n216310 );
not ( n228129 , n218204 );
or ( n228130 , n228128 , n228129 );
nand ( n228131 , n208594 , n218217 );
nand ( n228132 , n228130 , n228131 );
nand ( n228133 , n228127 , n228132 );
nand ( n228134 , n228126 , n228133 );
not ( n228135 , n227633 );
nor ( n228136 , n218832 , n218826 );
not ( n228137 , n228136 );
or ( n228138 , n228135 , n228137 );
not ( n228139 , n208717 );
not ( n228140 , n218814 );
or ( n228141 , n228139 , n228140 );
nand ( n228142 , n223671 , n217941 );
nand ( n228143 , n228141 , n228142 );
nand ( n228144 , n228143 , n218454 );
nand ( n228145 , n228138 , n228144 );
xor ( n228146 , n228134 , n228145 );
not ( n228147 , n227644 );
not ( n228148 , n221575 );
or ( n228149 , n228147 , n228148 );
not ( n228150 , n41701 );
not ( n228151 , n219419 );
or ( n228152 , n228150 , n228151 );
nand ( n228153 , n221227 , n226224 );
nand ( n228154 , n228152 , n228153 );
nand ( n228155 , n228154 , n219075 );
nand ( n228156 , n228149 , n228155 );
xor ( n228157 , n228146 , n228156 );
xor ( n228158 , n228134 , n228145 );
and ( n228159 , n228158 , n228156 );
and ( n228160 , n228134 , n228145 );
or ( n228161 , n228159 , n228160 );
not ( n228162 , n214319 );
not ( n228163 , n213382 );
buf ( n228164 , n39363 );
not ( n228165 , n228164 );
not ( n228166 , n228165 );
or ( n228167 , n228163 , n228166 );
nand ( n228168 , n39365 , n213381 );
nand ( n228169 , n228167 , n228168 );
not ( n228170 , n228169 );
or ( n228171 , n228162 , n228170 );
nand ( n228172 , n227671 , n217969 );
nand ( n228173 , n228171 , n228172 );
xor ( n228174 , n228173 , n228013 );
xor ( n228175 , n228174 , n228059 );
xor ( n228176 , n228173 , n228013 );
and ( n228177 , n228176 , n228059 );
and ( n228178 , n228173 , n228013 );
or ( n228179 , n228177 , n228178 );
not ( n228180 , n213874 );
not ( n228181 , n227681 );
or ( n228182 , n228180 , n228181 );
not ( n228183 , n216262 );
not ( n228184 , n39088 );
not ( n228185 , n228184 );
or ( n228186 , n228183 , n228185 );
nand ( n228187 , n39088 , n216265 );
nand ( n228188 , n228186 , n228187 );
nand ( n228189 , n228188 , n217142 );
nand ( n228190 , n228182 , n228189 );
xor ( n228191 , n228190 , n228063 );
not ( n228192 , n227880 );
not ( n228193 , n214717 );
or ( n228194 , n228192 , n228193 );
buf ( n228195 , n39878 );
and ( n228196 , n217944 , n228195 );
not ( n228197 , n217944 );
and ( n228198 , n228197 , n39879 );
nor ( n228199 , n228196 , n228198 );
or ( n228200 , n228199 , n220986 );
nand ( n228201 , n228194 , n228200 );
xor ( n228202 , n228191 , n228201 );
xor ( n228203 , n228190 , n228063 );
and ( n228204 , n228203 , n228201 );
and ( n228205 , n228190 , n228063 );
or ( n228206 , n228204 , n228205 );
not ( n228207 , n213577 );
not ( n228208 , n227698 );
or ( n228209 , n228207 , n228208 );
not ( n228210 , n213735 );
and ( n228211 , n831 , n18376 );
not ( n228212 , n831 );
and ( n228213 , n228212 , n39743 );
nor ( n228214 , n228211 , n228213 );
not ( n228215 , n228214 );
not ( n228216 , n228215 );
not ( n228217 , n228216 );
or ( n228218 , n228210 , n228217 );
nand ( n228219 , n39747 , n213732 );
nand ( n228220 , n228218 , n228219 );
nand ( n228221 , n228220 , n216336 );
nand ( n228222 , n228209 , n228221 );
not ( n228223 , n227857 );
not ( n228224 , n227849 );
or ( n228225 , n228223 , n228224 );
and ( n228226 , n214960 , n226648 );
not ( n228227 , n214960 );
and ( n228228 , n228227 , n226649 );
nor ( n228229 , n228226 , n228228 );
not ( n228230 , n228229 );
nand ( n228231 , n228230 , n227241 );
nand ( n228232 , n228225 , n228231 );
and ( n228233 , n227755 , n227765 );
xor ( n228234 , n228232 , n228233 );
not ( n228235 , n227604 );
nand ( n228236 , n228235 , n225478 );
not ( n228237 , n227121 );
not ( n228238 , n216422 );
not ( n228239 , n224617 );
or ( n228240 , n228238 , n228239 );
nand ( n228241 , n40724 , n227602 );
nand ( n228242 , n228240 , n228241 );
nand ( n228243 , n228237 , n228242 );
nand ( n228244 , n228236 , n228243 );
xor ( n228245 , n228234 , n228244 );
xor ( n228246 , n228222 , n228245 );
not ( n228247 , n227714 );
not ( n228248 , n225945 );
or ( n228249 , n228247 , n228248 );
not ( n228250 , n214899 );
not ( n228251 , n225952 );
or ( n228252 , n228250 , n228251 );
not ( n228253 , n225936 );
nand ( n228254 , n228253 , n214537 );
nand ( n228255 , n228252 , n228254 );
nand ( n228256 , n227710 , n228255 );
nand ( n228257 , n228249 , n228256 );
not ( n228258 , n227776 );
not ( n228259 , n223591 );
or ( n228260 , n228258 , n228259 );
not ( n228261 , n223155 );
not ( n228262 , n220436 );
and ( n228263 , n228261 , n228262 );
and ( n228264 , n223201 , n220436 );
nor ( n228265 , n228263 , n228264 );
not ( n228266 , n228265 );
nand ( n228267 , n228266 , n222769 );
nand ( n228268 , n228260 , n228267 );
xor ( n228269 , n228257 , n228268 );
buf ( n228270 , n227733 );
not ( n228271 , n227741 );
or ( n228272 , n228270 , n228271 );
not ( n228273 , n227737 );
not ( n228274 , n227723 );
not ( n228275 , n228274 );
not ( n228276 , n214616 );
and ( n228277 , n228275 , n228276 );
not ( n228278 , n227595 );
not ( n228279 , n228278 );
and ( n228280 , n228279 , n222031 );
nor ( n228281 , n228277 , n228280 );
or ( n228282 , n228273 , n228281 );
nand ( n228283 , n228272 , n228282 );
xor ( n228284 , n228269 , n228283 );
xor ( n228285 , n228246 , n228284 );
xor ( n228286 , n228222 , n228245 );
and ( n228287 , n228286 , n228284 );
and ( n228288 , n228222 , n228245 );
or ( n228289 , n228287 , n228288 );
not ( n228290 , n227837 );
not ( n228291 , n225902 );
or ( n228292 , n228290 , n228291 );
and ( n228293 , n222821 , n222428 );
not ( n228294 , n222821 );
not ( n228295 , n222428 );
and ( n228296 , n228294 , n228295 );
nor ( n228297 , n228293 , n228296 );
nand ( n228298 , n228297 , n222157 );
nand ( n228299 , n228292 , n228298 );
not ( n228300 , n227787 );
not ( n228301 , n224086 );
or ( n228302 , n228300 , n228301 );
not ( n228303 , n218514 );
not ( n228304 , n224069 );
or ( n228305 , n228303 , n228304 );
not ( n228306 , n224094 );
nand ( n228307 , n228306 , n216170 );
nand ( n228308 , n228305 , n228307 );
nand ( n228309 , n224090 , n228308 );
nand ( n228310 , n228302 , n228309 );
xor ( n228311 , n228299 , n228310 );
not ( n228312 , n227799 );
not ( n228313 , n226742 );
or ( n228314 , n228312 , n228313 );
not ( n228315 , n216208 );
not ( n228316 , n224844 );
or ( n228317 , n228315 , n228316 );
nand ( n228318 , n224944 , n216207 );
nand ( n228319 , n228317 , n228318 );
nand ( n228320 , n226745 , n228319 );
nand ( n228321 , n228314 , n228320 );
xor ( n228322 , n228311 , n228321 );
not ( n228323 , n227654 );
not ( n228324 , n228323 );
nand ( n228325 , n220156 , n220157 );
nor ( n228326 , n219777 , n228325 );
not ( n228327 , n228326 );
or ( n228328 , n228324 , n228327 );
not ( n228329 , n224170 );
not ( n228330 , n221256 );
not ( n228331 , n208725 );
or ( n228332 , n228330 , n228331 );
not ( n228333 , n220146 );
or ( n228334 , n228333 , n208727 );
nand ( n228335 , n228332 , n228334 );
nand ( n228336 , n228329 , n228335 );
nand ( n228337 , n228328 , n228336 );
not ( n228338 , n227813 );
not ( n228339 , n220899 );
nand ( n228340 , n228339 , n220911 );
nand ( n228341 , n220899 , n220912 );
and ( n228342 , n228340 , n220634 , n228341 );
not ( n228343 , n228342 );
or ( n228344 , n228338 , n228343 );
not ( n228345 , n224492 );
not ( n228346 , n220904 );
or ( n228347 , n228345 , n228346 );
nand ( n228348 , n226377 , n215833 );
nand ( n228349 , n228347 , n228348 );
nand ( n228350 , n228349 , n220929 );
nand ( n228351 , n228344 , n228350 );
xor ( n228352 , n228337 , n228351 );
not ( n228353 , n227826 );
not ( n228354 , n221625 );
or ( n228355 , n228353 , n228354 );
not ( n228356 , n216293 );
not ( n228357 , n221777 );
or ( n228358 , n228356 , n228357 );
nand ( n228359 , n221608 , n223658 );
nand ( n228360 , n228358 , n228359 );
nand ( n228361 , n228360 , n221387 );
nand ( n228362 , n228355 , n228361 );
xor ( n228363 , n228352 , n228362 );
xor ( n228364 , n228322 , n228363 );
xor ( n228365 , n228364 , n228157 );
xor ( n228366 , n228322 , n228363 );
and ( n228367 , n228366 , n228157 );
and ( n228368 , n228322 , n228363 );
or ( n228369 , n228367 , n228368 );
xor ( n228370 , n228075 , n228067 );
xor ( n228371 , n228370 , n228071 );
xor ( n228372 , n228075 , n228067 );
and ( n228373 , n228372 , n228071 );
and ( n228374 , n228075 , n228067 );
or ( n228375 , n228373 , n228374 );
not ( n228376 , n216562 );
not ( n228377 , n227890 );
or ( n228378 , n228376 , n228377 );
not ( n228379 , n215290 );
not ( n228380 , n223764 );
or ( n228381 , n228379 , n228380 );
nand ( n228382 , n40045 , n215289 );
nand ( n228383 , n228381 , n228382 );
nand ( n228384 , n228383 , n214694 );
nand ( n228385 , n228378 , n228384 );
xor ( n228386 , n228118 , n228385 );
not ( n228387 , n217023 );
not ( n228388 , n227941 );
or ( n228389 , n228387 , n228388 );
and ( n228390 , n40484 , n218661 );
not ( n228391 , n40484 );
and ( n228392 , n228391 , n219577 );
or ( n228393 , n228390 , n228392 );
nand ( n228394 , n228393 , n219175 );
nand ( n228395 , n228389 , n228394 );
xor ( n228396 , n228386 , n228395 );
xor ( n228397 , n228396 , n228079 );
xor ( n228398 , n228397 , n228083 );
xor ( n228399 , n228396 , n228079 );
and ( n228400 , n228399 , n228083 );
and ( n228401 , n228396 , n228079 );
or ( n228402 , n228400 , n228401 );
not ( n228403 , n220280 );
not ( n228404 , n227867 );
or ( n228405 , n228403 , n228404 );
not ( n228406 , n217542 );
not ( n228407 , n223748 );
or ( n228408 , n228406 , n228407 );
nand ( n228409 , n40421 , n216989 );
nand ( n228410 , n228408 , n228409 );
nand ( n228411 , n228410 , n220272 );
nand ( n228412 , n228405 , n228411 );
not ( n228413 , n219731 );
not ( n228414 , n227957 );
or ( n228415 , n228413 , n228414 );
and ( n228416 , n40396 , n219034 );
not ( n228417 , n40396 );
and ( n228418 , n228417 , n219033 );
or ( n228419 , n228416 , n228418 );
nand ( n228420 , n228419 , n222185 );
nand ( n228421 , n228415 , n228420 );
xor ( n228422 , n228412 , n228421 );
not ( n228423 , n224624 );
not ( n228424 , n227969 );
or ( n228425 , n228423 , n228424 );
not ( n228426 , n219687 );
not ( n228427 , n220599 );
or ( n228428 , n228426 , n228427 );
nand ( n228429 , n40410 , n222323 );
nand ( n228430 , n228428 , n228429 );
nand ( n228431 , n228430 , n219314 );
nand ( n228432 , n228425 , n228431 );
xor ( n228433 , n228422 , n228432 );
xor ( n228434 , n227688 , n228433 );
not ( n228435 , n219332 );
not ( n228436 , n227978 );
or ( n228437 , n228435 , n228436 );
not ( n228438 , n226484 );
not ( n228439 , n221356 );
or ( n228440 , n228438 , n228439 );
nand ( n228441 , n207936 , n221938 );
nand ( n228442 , n228440 , n228441 );
nand ( n228443 , n228442 , n221933 );
nand ( n228444 , n228437 , n228443 );
not ( n228445 , n226943 );
not ( n228446 , n227918 );
or ( n228447 , n228445 , n228446 );
not ( n228448 , n227912 );
not ( n228449 , n219226 );
not ( n228450 , n228449 );
or ( n228451 , n228448 , n228450 );
not ( n228452 , n219226 );
or ( n228453 , n228452 , n227912 );
nand ( n228454 , n228451 , n228453 );
nand ( n228455 , n228454 , n226287 );
nand ( n228456 , n228447 , n228455 );
xor ( n228457 , n228444 , n228456 );
not ( n228458 , n227260 );
not ( n228459 , n227929 );
or ( n228460 , n228458 , n228459 );
and ( n228461 , n225556 , n218736 );
not ( n228462 , n225556 );
and ( n228463 , n228462 , n226655 );
or ( n228464 , n228461 , n228463 );
nand ( n228465 , n228464 , n223949 );
nand ( n228466 , n228460 , n228465 );
xor ( n228467 , n228457 , n228466 );
xor ( n228468 , n228434 , n228467 );
xor ( n228469 , n227688 , n228433 );
and ( n228470 , n228469 , n228467 );
and ( n228471 , n227688 , n228433 );
or ( n228472 , n228470 , n228471 );
not ( n228473 , n214086 );
not ( n228474 , n227902 );
or ( n228475 , n228473 , n228474 );
and ( n228476 , n39812 , n219390 );
not ( n228477 , n39812 );
and ( n228478 , n228477 , n217573 );
or ( n228479 , n228476 , n228478 );
nand ( n228480 , n228479 , n215383 );
nand ( n228481 , n228475 , n228480 );
xor ( n228482 , n228481 , n227624 );
xor ( n228483 , n228482 , n227662 );
xor ( n228484 , n228202 , n228483 );
xor ( n228485 , n228484 , n228175 );
xor ( n228486 , n228202 , n228483 );
and ( n228487 , n228486 , n228175 );
and ( n228488 , n228202 , n228483 );
or ( n228489 , n228487 , n228488 );
xor ( n228490 , n227807 , n227706 );
xor ( n228491 , n228490 , n228285 );
xor ( n228492 , n227807 , n227706 );
and ( n228493 , n228492 , n228285 );
and ( n228494 , n227807 , n227706 );
or ( n228495 , n228493 , n228494 );
xor ( n228496 , n227846 , n228365 );
xor ( n228497 , n228496 , n227910 );
xor ( n228498 , n227846 , n228365 );
and ( n228499 , n228498 , n227910 );
and ( n228500 , n227846 , n228365 );
or ( n228501 , n228499 , n228500 );
xor ( n228502 , n228337 , n228351 );
and ( n228503 , n228502 , n228362 );
and ( n228504 , n228337 , n228351 );
or ( n228505 , n228503 , n228504 );
xor ( n228506 , n227952 , n228371 );
xor ( n228507 , n228506 , n227997 );
xor ( n228508 , n227952 , n228371 );
and ( n228509 , n228508 , n227997 );
and ( n228510 , n227952 , n228371 );
or ( n228511 , n228509 , n228510 );
xor ( n228512 , n228398 , n227989 );
xor ( n228513 , n228512 , n228468 );
xor ( n228514 , n228398 , n227989 );
and ( n228515 , n228514 , n228468 );
and ( n228516 , n228398 , n227989 );
or ( n228517 , n228515 , n228516 );
xor ( n228518 , n228003 , n228491 );
xor ( n228519 , n228518 , n228485 );
xor ( n228520 , n228003 , n228491 );
and ( n228521 , n228520 , n228485 );
and ( n228522 , n228003 , n228491 );
or ( n228523 , n228521 , n228522 );
xor ( n228524 , n228497 , n228009 );
xor ( n228525 , n228524 , n228507 );
xor ( n228526 , n228497 , n228009 );
and ( n228527 , n228526 , n228507 );
and ( n228528 , n228497 , n228009 );
or ( n228529 , n228527 , n228528 );
xor ( n228530 , n228019 , n228025 );
xor ( n228531 , n228530 , n228513 );
xor ( n228532 , n228019 , n228025 );
and ( n228533 , n228532 , n228513 );
and ( n228534 , n228019 , n228025 );
or ( n228535 , n228533 , n228534 );
xor ( n228536 , n228519 , n228031 );
xor ( n228537 , n228536 , n228525 );
xor ( n228538 , n228519 , n228031 );
and ( n228539 , n228538 , n228525 );
and ( n228540 , n228519 , n228031 );
or ( n228541 , n228539 , n228540 );
xor ( n228542 , n228037 , n228531 );
xor ( n228543 , n228542 , n228043 );
xor ( n228544 , n228037 , n228531 );
and ( n228545 , n228544 , n228043 );
and ( n228546 , n228037 , n228531 );
or ( n228547 , n228545 , n228546 );
xor ( n228548 , n228537 , n228543 );
xor ( n228549 , n228548 , n228049 );
xor ( n228550 , n228537 , n228543 );
and ( n228551 , n228550 , n228049 );
and ( n228552 , n228537 , n228543 );
or ( n228553 , n228551 , n228552 );
xor ( n228554 , n228299 , n228310 );
and ( n228555 , n228554 , n228321 );
and ( n228556 , n228299 , n228310 );
or ( n228557 , n228555 , n228556 );
xor ( n228558 , n228257 , n228268 );
and ( n228559 , n228558 , n228283 );
and ( n228560 , n228257 , n228268 );
or ( n228561 , n228559 , n228560 );
xor ( n228562 , n228232 , n228233 );
and ( n228563 , n228562 , n228244 );
and ( n228564 , n228232 , n228233 );
or ( n228565 , n228563 , n228564 );
xor ( n228566 , n228412 , n228421 );
and ( n228567 , n228566 , n228432 );
and ( n228568 , n228412 , n228421 );
or ( n228569 , n228567 , n228568 );
xor ( n228570 , n228444 , n228456 );
and ( n228571 , n228570 , n228466 );
and ( n228572 , n228444 , n228456 );
or ( n228573 , n228571 , n228572 );
xor ( n228574 , n228118 , n228385 );
and ( n228575 , n228574 , n228395 );
and ( n228576 , n228118 , n228385 );
or ( n228577 , n228575 , n228576 );
xor ( n228578 , n228481 , n227624 );
and ( n228579 , n228578 , n227662 );
and ( n228580 , n228481 , n227624 );
or ( n228581 , n228579 , n228580 );
not ( n228582 , n217388 );
not ( n228583 , n216929 );
not ( n228584 , n220077 );
or ( n228585 , n228583 , n228584 );
nand ( n228586 , n41164 , n217076 );
nand ( n228587 , n228585 , n228586 );
not ( n228588 , n228587 );
or ( n228589 , n228582 , n228588 );
nand ( n228590 , n228090 , n222270 );
nand ( n228591 , n228589 , n228590 );
not ( n228592 , n228132 );
not ( n228593 , n218221 );
or ( n228594 , n228592 , n228593 );
not ( n228595 , n224881 );
not ( n228596 , n218226 );
or ( n228597 , n228595 , n228596 );
nand ( n228598 , n218771 , n41249 );
nand ( n228599 , n228597 , n228598 );
nand ( n228600 , n228599 , n218231 );
nand ( n228601 , n228594 , n228600 );
xor ( n228602 , n228591 , n228601 );
not ( n228603 , n228143 );
not ( n228604 , n218835 );
or ( n228605 , n228603 , n228604 );
not ( n228606 , n41396 );
not ( n228607 , n218814 );
or ( n228608 , n228606 , n228607 );
nand ( n228609 , n227631 , n219581 );
nand ( n228610 , n228608 , n228609 );
nand ( n228611 , n218455 , n228610 );
nand ( n228612 , n228605 , n228611 );
xor ( n228613 , n228602 , n228612 );
xor ( n228614 , n228591 , n228601 );
and ( n228615 , n228614 , n228612 );
and ( n228616 , n228591 , n228601 );
or ( n228617 , n228615 , n228616 );
not ( n228618 , n228154 );
not ( n228619 , n221575 );
or ( n228620 , n228618 , n228619 );
and ( n228621 , n41565 , n221227 );
not ( n228622 , n41565 );
and ( n228623 , n228622 , n219423 );
nor ( n228624 , n228621 , n228623 );
nand ( n228625 , n219075 , n228624 );
nand ( n228626 , n228620 , n228625 );
not ( n228627 , n228335 );
not ( n228628 , n220163 );
or ( n228629 , n228627 , n228628 );
not ( n228630 , n225768 );
not ( n228631 , n222412 );
or ( n228632 , n228630 , n228631 );
not ( n228633 , n224562 );
nand ( n228634 , n228633 , n225763 );
nand ( n228635 , n228632 , n228634 );
nand ( n228636 , n219779 , n228635 );
nand ( n228637 , n228629 , n228636 );
xor ( n228638 , n228626 , n228637 );
not ( n228639 , n221265 );
not ( n228640 , n228349 );
or ( n228641 , n228639 , n228640 );
not ( n228642 , n214837 );
not ( n228643 , n224112 );
or ( n228644 , n228642 , n228643 );
nand ( n228645 , n226377 , n218670 );
nand ( n228646 , n228644 , n228645 );
not ( n228647 , n228646 );
not ( n228648 , n220636 );
or ( n228649 , n228647 , n228648 );
nand ( n228650 , n228641 , n228649 );
xor ( n228651 , n228638 , n228650 );
xor ( n228652 , n228626 , n228637 );
and ( n228653 , n228652 , n228650 );
and ( n228654 , n228626 , n228637 );
or ( n228655 , n228653 , n228654 );
not ( n228656 , n217142 );
not ( n228657 , n38531 );
and ( n228658 , n216262 , n228657 );
not ( n228659 , n216262 );
and ( n228660 , n228659 , n38531 );
nor ( n228661 , n228658 , n228660 );
not ( n228662 , n228661 );
not ( n228663 , n228662 );
or ( n228664 , n228656 , n228663 );
nand ( n228665 , n228188 , n213152 );
nand ( n228666 , n228664 , n228665 );
xor ( n228667 , n228666 , n228561 );
not ( n228668 , n218855 );
not ( n228669 , n39926 );
or ( n228670 , n228668 , n228669 );
nand ( n228671 , n225097 , n217944 );
nand ( n228672 , n228670 , n228671 );
not ( n228673 , n228672 );
not ( n228674 , n220985 );
or ( n228675 , n228673 , n228674 );
not ( n228676 , n214717 );
or ( n228677 , n228199 , n228676 );
nand ( n228678 , n228675 , n228677 );
xor ( n228679 , n228667 , n228678 );
xor ( n228680 , n228666 , n228561 );
and ( n228681 , n228680 , n228678 );
and ( n228682 , n228666 , n228561 );
or ( n228683 , n228681 , n228682 );
not ( n228684 , n213577 );
not ( n228685 , n228220 );
or ( n228686 , n228684 , n228685 );
and ( n228687 , n39606 , n213732 );
not ( n228688 , n39606 );
and ( n228689 , n228688 , n213735 );
or ( n228690 , n228687 , n228689 );
nand ( n228691 , n228690 , n216336 );
nand ( n228692 , n228686 , n228691 );
not ( n228693 , n217969 );
not ( n228694 , n228169 );
or ( n228695 , n228693 , n228694 );
or ( n228696 , n213381 , n39286 );
nand ( n228697 , n213381 , n39286 );
nand ( n228698 , n228696 , n228697 );
nand ( n228699 , n228698 , n214319 );
nand ( n228700 , n228695 , n228699 );
xor ( n228701 , n228692 , n228700 );
xor ( n228702 , n228701 , n228565 );
xor ( n228703 , n228692 , n228700 );
and ( n228704 , n228703 , n228565 );
and ( n228705 , n228692 , n228700 );
or ( n228706 , n228704 , n228705 );
nand ( n228707 , n227732 , n227728 );
or ( n228708 , n228281 , n228707 );
and ( n228709 , n228278 , n213583 );
and ( n228710 , n227595 , n214134 );
nor ( n228711 , n228709 , n228710 );
or ( n228712 , n228711 , n227164 );
nand ( n228713 , n228708 , n228712 );
not ( n228714 , n228111 );
and ( n228715 , n228714 , n215999 );
not ( n228716 , n37618 );
not ( n228717 , n37488 );
nor ( n228718 , n36730 , n37687 );
nand ( n228719 , n228718 , n219064 );
nand ( n228720 , n228717 , n228719 , n37689 );
not ( n228721 , n228720 );
not ( n228722 , n228721 );
or ( n228723 , n228716 , n228722 );
nand ( n228724 , n228720 , n37619 );
nand ( n228725 , n228723 , n228724 );
buf ( n228726 , n228725 );
not ( n228727 , n228726 );
nor ( n228728 , n228715 , n228727 );
or ( n228729 , n228714 , n215999 );
nand ( n228730 , n228729 , n228274 );
nand ( n228731 , n228728 , n228730 );
not ( n228732 , n228731 );
not ( n228733 , n228732 );
not ( n228734 , n217230 );
not ( n228735 , n217614 );
not ( n228736 , n227747 );
or ( n228737 , n228735 , n228736 );
nand ( n228738 , n208259 , n217473 );
nand ( n228739 , n228737 , n228738 );
not ( n228740 , n228739 );
or ( n228741 , n228734 , n228740 );
not ( n228742 , n217629 );
nand ( n228743 , n228742 , n228100 );
nand ( n228744 , n228741 , n228743 );
not ( n228745 , n228744 );
not ( n228746 , n228745 );
or ( n228747 , n228733 , n228746 );
or ( n228748 , n228745 , n228732 );
nand ( n228749 , n228747 , n228748 );
xor ( n228750 , n228713 , n228749 );
not ( n228751 , n227241 );
and ( n228752 , n217044 , n226888 );
not ( n228753 , n217044 );
and ( n228754 , n228753 , n227245 );
or ( n228755 , n228752 , n228754 );
not ( n228756 , n228755 );
or ( n228757 , n228751 , n228756 );
or ( n228758 , n227848 , n228229 );
nand ( n228759 , n228757 , n228758 );
xor ( n228760 , n228750 , n228759 );
xor ( n228761 , n228613 , n228760 );
not ( n228762 , n228319 );
not ( n228763 , n226742 );
or ( n228764 , n228762 , n228763 );
not ( n228765 , n215075 );
not ( n228766 , n224844 );
or ( n228767 , n228765 , n228766 );
nand ( n228768 , n224929 , n215899 );
nand ( n228769 , n228767 , n228768 );
nand ( n228770 , n224449 , n228769 );
nand ( n228771 , n228764 , n228770 );
not ( n228772 , n228255 );
not ( n228773 , n226755 );
or ( n228774 , n228772 , n228773 );
not ( n228775 , n225316 );
not ( n228776 , n216964 );
not ( n228777 , n225743 );
or ( n228778 , n228776 , n228777 );
nand ( n228779 , n225952 , n214678 );
nand ( n228780 , n228778 , n228779 );
nand ( n228781 , n228775 , n228780 );
nand ( n228782 , n228774 , n228781 );
xor ( n228783 , n228771 , n228782 );
not ( n228784 , n228265 );
not ( n228785 , n228784 );
not ( n228786 , n223197 );
or ( n228787 , n228785 , n228786 );
not ( n228788 , n219343 );
not ( n228789 , n223156 );
or ( n228790 , n228788 , n228789 );
nand ( n228791 , n223182 , n219348 );
nand ( n228792 , n228790 , n228791 );
nand ( n228793 , n227294 , n228792 );
nand ( n228794 , n228787 , n228793 );
xor ( n228795 , n228783 , n228794 );
xor ( n228796 , n228761 , n228795 );
xor ( n228797 , n228613 , n228760 );
and ( n228798 , n228797 , n228795 );
and ( n228799 , n228613 , n228760 );
or ( n228800 , n228798 , n228799 );
not ( n228801 , n228360 );
not ( n228802 , n224120 );
or ( n228803 , n228801 , n228802 );
not ( n228804 , n224037 );
not ( n228805 , n221632 );
or ( n228806 , n228804 , n228805 );
nand ( n228807 , n221607 , n214821 );
nand ( n228808 , n228806 , n228807 );
nand ( n228809 , n228808 , n223587 );
nand ( n228810 , n228803 , n228809 );
not ( n228811 , n228297 );
not ( n228812 , n222453 );
or ( n228813 , n228811 , n228812 );
not ( n228814 , n215533 );
not ( n228815 , n225418 );
or ( n228816 , n228814 , n228815 );
not ( n228817 , n228295 );
nand ( n228818 , n228817 , n220022 );
nand ( n228819 , n228816 , n228818 );
nand ( n228820 , n228819 , n222465 );
nand ( n228821 , n228813 , n228820 );
xor ( n228822 , n228810 , n228821 );
not ( n228823 , n228308 );
not ( n228824 , n224086 );
or ( n228825 , n228823 , n228824 );
and ( n228826 , n216934 , n224069 );
not ( n228827 , n216934 );
not ( n228828 , n224975 );
and ( n228829 , n228827 , n228828 );
or ( n228830 , n228826 , n228829 );
nand ( n228831 , n227782 , n228830 );
nand ( n228832 , n228825 , n228831 );
xor ( n228833 , n228822 , n228832 );
xor ( n228834 , n228833 , n228651 );
xor ( n228835 , n228834 , n228573 );
xor ( n228836 , n228833 , n228651 );
and ( n228837 , n228836 , n228573 );
and ( n228838 , n228833 , n228651 );
or ( n228839 , n228837 , n228838 );
xor ( n228840 , n228569 , n228577 );
not ( n228841 , n213750 );
not ( n228842 , n37618 );
not ( n228843 , n228721 );
or ( n228844 , n228842 , n228843 );
nand ( n228845 , n228844 , n228724 );
not ( n228846 , n228845 );
buf ( n228847 , n228846 );
not ( n228848 , n228847 );
or ( n228849 , n228841 , n228848 );
not ( n228850 , n228847 );
nand ( n228851 , n228850 , n213751 );
nand ( n228852 , n228849 , n228851 );
not ( n228853 , n228852 );
and ( n228854 , n228111 , n228846 );
and ( n228855 , n228110 , n228845 );
nor ( n228856 , n228854 , n228855 );
nand ( n228857 , n228115 , n228856 );
not ( n228858 , n228857 );
not ( n228859 , n228858 );
not ( n228860 , n228859 );
not ( n228861 , n228860 );
or ( n228862 , n228853 , n228861 );
and ( n228863 , n228846 , n218224 );
and ( n228864 , n228726 , n216076 );
nor ( n228865 , n228863 , n228864 );
not ( n228866 , n228865 );
not ( n228867 , n228116 );
buf ( n228868 , n228867 );
nand ( n228869 , n228866 , n228868 );
nand ( n228870 , n228862 , n228869 );
xor ( n228871 , n228870 , n228122 );
not ( n228872 , n217552 );
not ( n228873 , n228410 );
or ( n228874 , n228872 , n228873 );
and ( n228875 , n40413 , n219358 );
not ( n228876 , n40413 );
and ( n228877 , n228876 , n215955 );
or ( n228878 , n228875 , n228877 );
nand ( n228879 , n228878 , n220272 );
nand ( n228880 , n228874 , n228879 );
xor ( n228881 , n228871 , n228880 );
xor ( n228882 , n228840 , n228881 );
xor ( n228883 , n228569 , n228577 );
and ( n228884 , n228883 , n228881 );
and ( n228885 , n228569 , n228577 );
or ( n228886 , n228884 , n228885 );
not ( n228887 , n227260 );
not ( n228888 , n228464 );
or ( n228889 , n228887 , n228888 );
and ( n228890 , n208078 , n218736 );
not ( n228891 , n208078 );
and ( n228892 , n228891 , n226655 );
or ( n228893 , n228890 , n228892 );
nand ( n228894 , n228893 , n223949 );
nand ( n228895 , n228889 , n228894 );
not ( n228896 , n219501 );
not ( n228897 , n216422 );
not ( n228898 , n218883 );
or ( n228899 , n228897 , n228898 );
nand ( n228900 , n218882 , n227599 );
nand ( n228901 , n228899 , n228900 );
not ( n228902 , n228901 );
or ( n228903 , n228896 , n228902 );
nand ( n228904 , n228242 , n225478 );
nand ( n228905 , n228903 , n228904 );
xor ( n228906 , n228895 , n228905 );
not ( n228907 , n217571 );
and ( n228908 , n39713 , n219390 );
not ( n228909 , n39713 );
and ( n228910 , n228909 , n213960 );
or ( n228911 , n228908 , n228910 );
not ( n228912 , n228911 );
or ( n228913 , n228907 , n228912 );
nand ( n228914 , n228479 , n218467 );
nand ( n228915 , n228913 , n228914 );
xor ( n228916 , n228906 , n228915 );
xor ( n228917 , n228916 , n228581 );
xor ( n228918 , n228917 , n228179 );
xor ( n228919 , n228916 , n228581 );
and ( n228920 , n228919 , n228179 );
and ( n228921 , n228916 , n228581 );
or ( n228922 , n228920 , n228921 );
not ( n228923 , n219731 );
not ( n228924 , n228419 );
or ( n228925 , n228923 , n228924 );
and ( n228926 , n40180 , n226002 );
not ( n228927 , n40180 );
and ( n228928 , n228927 , n219033 );
or ( n228929 , n228926 , n228928 );
nand ( n228930 , n228929 , n214458 );
nand ( n228931 , n228925 , n228930 );
not ( n228932 , n217023 );
not ( n228933 , n228393 );
or ( n228934 , n228932 , n228933 );
not ( n228935 , n217017 );
not ( n228936 , n224285 );
or ( n228937 , n228935 , n228936 );
nand ( n228938 , n40545 , n218661 );
nand ( n228939 , n228937 , n228938 );
nand ( n228940 , n228939 , n219175 );
nand ( n228941 , n228934 , n228940 );
xor ( n228942 , n228931 , n228941 );
not ( n228943 , n219314 );
not ( n228944 , n219687 );
not ( n228945 , n40258 );
or ( n228946 , n228944 , n228945 );
nand ( n228947 , n223383 , n221283 );
nand ( n228948 , n228946 , n228947 );
not ( n228949 , n228948 );
or ( n228950 , n228943 , n228949 );
nand ( n228951 , n228430 , n224624 );
nand ( n228952 , n228950 , n228951 );
xor ( n228953 , n228942 , n228952 );
xor ( n228954 , n228953 , n228206 );
not ( n228955 , n215183 );
not ( n228956 , n228442 );
or ( n228957 , n228955 , n228956 );
not ( n228958 , n221935 );
not ( n228959 , n222500 );
or ( n228960 , n228958 , n228959 );
nand ( n228961 , n40668 , n218994 );
nand ( n228962 , n228960 , n228961 );
nand ( n228963 , n228962 , n221933 );
nand ( n228964 , n228957 , n228963 );
not ( n228965 , n216299 );
not ( n228966 , n228383 );
or ( n228967 , n228965 , n228966 );
not ( n228968 , n215290 );
not ( n228969 , n39996 );
or ( n228970 , n228968 , n228969 );
nand ( n228971 , n39995 , n215289 );
nand ( n228972 , n228970 , n228971 );
nand ( n228973 , n228972 , n214694 );
nand ( n228974 , n228967 , n228973 );
xor ( n228975 , n228964 , n228974 );
not ( n228976 , n228454 );
or ( n228977 , n228976 , n226942 );
not ( n228978 , n227912 );
not ( n228979 , n221040 );
or ( n228980 , n228978 , n228979 );
nand ( n228981 , n221690 , n220038 );
nand ( n228982 , n228980 , n228981 );
not ( n228983 , n228982 );
or ( n228984 , n228983 , n226940 );
nand ( n228985 , n228977 , n228984 );
xor ( n228986 , n228975 , n228985 );
xor ( n228987 , n228954 , n228986 );
xor ( n228988 , n228953 , n228206 );
and ( n228989 , n228988 , n228986 );
and ( n228990 , n228953 , n228206 );
or ( n228991 , n228989 , n228990 );
xor ( n228992 , n228369 , n228702 );
xor ( n228993 , n228161 , n228505 );
xor ( n228994 , n228993 , n228557 );
xor ( n228995 , n228992 , n228994 );
xor ( n228996 , n228369 , n228702 );
and ( n228997 , n228996 , n228994 );
and ( n228998 , n228369 , n228702 );
or ( n228999 , n228997 , n228998 );
xor ( n229000 , n228679 , n228289 );
xor ( n229001 , n229000 , n228375 );
xor ( n229002 , n228679 , n228289 );
and ( n229003 , n229002 , n228375 );
and ( n229004 , n228679 , n228289 );
or ( n229005 , n229003 , n229004 );
xor ( n229006 , n228796 , n228835 );
xor ( n229007 , n229006 , n228472 );
xor ( n229008 , n228796 , n228835 );
and ( n229009 , n229008 , n228472 );
and ( n229010 , n228796 , n228835 );
or ( n229011 , n229009 , n229010 );
xor ( n229012 , n228810 , n228821 );
and ( n229013 , n229012 , n228832 );
and ( n229014 , n228810 , n228821 );
or ( n229015 , n229013 , n229014 );
xor ( n229016 , n228882 , n228402 );
xor ( n229017 , n229016 , n228918 );
xor ( n229018 , n228882 , n228402 );
and ( n229019 , n229018 , n228918 );
and ( n229020 , n228882 , n228402 );
or ( n229021 , n229019 , n229020 );
xor ( n229022 , n228987 , n228489 );
xor ( n229023 , n229022 , n228495 );
xor ( n229024 , n228987 , n228489 );
and ( n229025 , n229024 , n228495 );
and ( n229026 , n228987 , n228489 );
or ( n229027 , n229025 , n229026 );
xor ( n229028 , n228995 , n229001 );
xor ( n229029 , n229028 , n228501 );
xor ( n229030 , n228995 , n229001 );
and ( n229031 , n229030 , n228501 );
and ( n229032 , n228995 , n229001 );
or ( n229033 , n229031 , n229032 );
xor ( n229034 , n229007 , n228517 );
xor ( n229035 , n229034 , n229017 );
xor ( n229036 , n229007 , n228517 );
and ( n229037 , n229036 , n229017 );
and ( n229038 , n229007 , n228517 );
or ( n229039 , n229037 , n229038 );
xor ( n229040 , n228511 , n228523 );
xor ( n229041 , n229040 , n229023 );
xor ( n229042 , n228511 , n228523 );
and ( n229043 , n229042 , n229023 );
and ( n229044 , n228511 , n228523 );
or ( n229045 , n229043 , n229044 );
xor ( n229046 , n229029 , n228529 );
xor ( n229047 , n229046 , n228535 );
xor ( n229048 , n229029 , n228529 );
and ( n229049 , n229048 , n228535 );
and ( n229050 , n229029 , n228529 );
or ( n229051 , n229049 , n229050 );
xor ( n229052 , n229035 , n229041 );
xor ( n229053 , n229052 , n228541 );
xor ( n229054 , n229035 , n229041 );
and ( n229055 , n229054 , n228541 );
and ( n229056 , n229035 , n229041 );
or ( n229057 , n229055 , n229056 );
xor ( n229058 , n229047 , n229053 );
xor ( n229059 , n229058 , n228547 );
xor ( n229060 , n229047 , n229053 );
and ( n229061 , n229060 , n228547 );
and ( n229062 , n229047 , n229053 );
or ( n229063 , n229061 , n229062 );
xor ( n229064 , n228771 , n228782 );
and ( n229065 , n229064 , n228794 );
and ( n229066 , n228771 , n228782 );
or ( n229067 , n229065 , n229066 );
xor ( n229068 , n228713 , n228749 );
and ( n229069 , n229068 , n228759 );
and ( n229070 , n228713 , n228749 );
or ( n229071 , n229069 , n229070 );
xor ( n229072 , n228870 , n228122 );
and ( n229073 , n229072 , n228880 );
and ( n229074 , n228870 , n228122 );
or ( n229075 , n229073 , n229074 );
xor ( n229076 , n228931 , n228941 );
and ( n229077 , n229076 , n228952 );
and ( n229078 , n228931 , n228941 );
or ( n229079 , n229077 , n229078 );
xor ( n229080 , n228964 , n228974 );
and ( n229081 , n229080 , n228985 );
and ( n229082 , n228964 , n228974 );
or ( n229083 , n229081 , n229082 );
xor ( n229084 , n228895 , n228905 );
and ( n229085 , n229084 , n228915 );
and ( n229086 , n228895 , n228905 );
or ( n229087 , n229085 , n229086 );
xor ( n229088 , n228161 , n228505 );
and ( n229089 , n229088 , n228557 );
and ( n229090 , n228161 , n228505 );
or ( n229091 , n229089 , n229090 );
not ( n229092 , n220067 );
not ( n229093 , n217614 );
not ( n229094 , n218420 );
or ( n229095 , n229093 , n229094 );
nand ( n229096 , n41069 , n221924 );
nand ( n229097 , n229095 , n229096 );
not ( n229098 , n229097 );
or ( n229099 , n229092 , n229098 );
nand ( n229100 , n228739 , n220059 );
nand ( n229101 , n229099 , n229100 );
not ( n229102 , n228726 );
buf ( n229103 , n219064 );
not ( n229104 , n37556 );
not ( n229105 , n229104 );
nor ( n229106 , n229105 , n37575 );
nand ( n229107 , n229103 , n229106 );
nand ( n229108 , n229107 , n37693 , n37678 );
nand ( n229109 , n37529 , n37523 );
not ( n229110 , n229109 );
and ( n229111 , n229108 , n229110 );
not ( n229112 , n229108 );
and ( n229113 , n229112 , n229109 );
nor ( n229114 , n229111 , n229113 );
not ( n229115 , n229114 );
not ( n229116 , n229115 );
or ( n229117 , n229102 , n229116 );
and ( n229118 , n229108 , n229110 );
not ( n229119 , n229108 );
and ( n229120 , n229119 , n229109 );
nor ( n229121 , n229118 , n229120 );
nand ( n229122 , n228846 , n229121 );
nand ( n229123 , n229117 , n229122 );
and ( n229124 , n229123 , n215999 );
xor ( n229125 , n229101 , n229124 );
not ( n229126 , n228599 );
not ( n229127 , n218525 );
or ( n229128 , n229126 , n229127 );
not ( n229129 , n223549 );
not ( n229130 , n218772 );
or ( n229131 , n229129 , n229130 );
nand ( n229132 , n218771 , n217314 );
nand ( n229133 , n229131 , n229132 );
nand ( n229134 , n229133 , n218231 );
nand ( n229135 , n229128 , n229134 );
xor ( n229136 , n229125 , n229135 );
xor ( n229137 , n229101 , n229124 );
and ( n229138 , n229137 , n229135 );
and ( n229139 , n229101 , n229124 );
or ( n229140 , n229138 , n229139 );
not ( n229141 , n228610 );
not ( n229142 , n228136 );
or ( n229143 , n229141 , n229142 );
and ( n229144 , n216306 , n218814 );
not ( n229145 , n216306 );
and ( n229146 , n229145 , n220859 );
or ( n229147 , n229144 , n229146 );
nand ( n229148 , n229147 , n218454 );
nand ( n229149 , n229143 , n229148 );
and ( n229150 , n228744 , n228732 );
xor ( n229151 , n229149 , n229150 );
not ( n229152 , n228624 );
not ( n229153 , n219435 );
or ( n229154 , n229152 , n229153 );
not ( n229155 , n208717 );
not ( n229156 , n219419 );
or ( n229157 , n229155 , n229156 );
nand ( n229158 , n216261 , n220180 );
nand ( n229159 , n229157 , n229158 );
nand ( n229160 , n229159 , n219076 );
nand ( n229161 , n229154 , n229160 );
xor ( n229162 , n229151 , n229161 );
xor ( n229163 , n229149 , n229150 );
and ( n229164 , n229163 , n229161 );
and ( n229165 , n229149 , n229150 );
or ( n229166 , n229164 , n229165 );
not ( n229167 , n217142 );
and ( n229168 , n39364 , n216262 );
not ( n229169 , n39364 );
and ( n229170 , n229169 , n214824 );
or ( n229171 , n229168 , n229170 );
not ( n229172 , n229171 );
or ( n229173 , n229167 , n229172 );
not ( n229174 , n228661 );
nand ( n229175 , n229174 , n213874 );
nand ( n229176 , n229173 , n229175 );
xor ( n229177 , n229136 , n229176 );
xor ( n229178 , n229177 , n229067 );
xor ( n229179 , n229136 , n229176 );
and ( n229180 , n229179 , n229067 );
and ( n229181 , n229136 , n229176 );
or ( n229182 , n229180 , n229181 );
not ( n229183 , n214717 );
not ( n229184 , n228672 );
or ( n229185 , n229183 , n229184 );
not ( n229186 , n215113 );
not ( n229187 , n225357 );
or ( n229188 , n229186 , n229187 );
nand ( n229189 , n39812 , n217944 );
nand ( n229190 , n229188 , n229189 );
nand ( n229191 , n229190 , n220985 );
nand ( n229192 , n229185 , n229191 );
xor ( n229193 , n229071 , n229192 );
not ( n229194 , n214694 );
not ( n229195 , n215290 );
not ( n229196 , n39877 );
or ( n229197 , n229195 , n229196 );
not ( n229198 , n39876 );
nand ( n229199 , n229198 , n215289 );
nand ( n229200 , n229197 , n229199 );
not ( n229201 , n229200 );
or ( n229202 , n229194 , n229201 );
nand ( n229203 , n228972 , n216562 );
nand ( n229204 , n229202 , n229203 );
xor ( n229205 , n229193 , n229204 );
xor ( n229206 , n229071 , n229192 );
and ( n229207 , n229206 , n229204 );
and ( n229208 , n229071 , n229192 );
or ( n229209 , n229207 , n229208 );
not ( n229210 , n213784 );
not ( n229211 , n228698 );
or ( n229212 , n229210 , n229211 );
nand ( n229213 , n209768 , n209761 );
not ( n229214 , n229213 );
and ( n229215 , n217715 , n229214 );
not ( n229216 , n217715 );
not ( n229217 , n229214 );
and ( n229218 , n229216 , n229217 );
nor ( n229219 , n229215 , n229218 );
nand ( n229220 , n229219 , n214319 );
nand ( n229221 , n229212 , n229220 );
not ( n229222 , n213577 );
not ( n229223 , n228690 );
or ( n229224 , n229222 , n229223 );
not ( n229225 , n213735 );
not ( n229226 , n228184 );
or ( n229227 , n229225 , n229226 );
nand ( n229228 , n213732 , n39088 );
nand ( n229229 , n229227 , n229228 );
nand ( n229230 , n229229 , n216336 );
nand ( n229231 , n229224 , n229230 );
xor ( n229232 , n229221 , n229231 );
xor ( n229233 , n229232 , n229162 );
xor ( n229234 , n229221 , n229231 );
and ( n229235 , n229234 , n229162 );
and ( n229236 , n229221 , n229231 );
or ( n229237 , n229235 , n229236 );
not ( n229238 , n228755 );
not ( n229239 , n226880 );
or ( n229240 , n229238 , n229239 );
not ( n229241 , n214537 );
not ( n229242 , n226888 );
or ( n229243 , n229241 , n229242 );
nand ( n229244 , n227245 , n214899 );
nand ( n229245 , n229243 , n229244 );
nand ( n229246 , n229245 , n226218 );
nand ( n229247 , n229240 , n229246 );
or ( n229248 , n228857 , n228865 );
not ( n229249 , n228726 );
and ( n229250 , n229249 , n213347 );
and ( n229251 , n228726 , n222031 );
nor ( n229252 , n229250 , n229251 );
or ( n229253 , n229252 , n228116 );
nand ( n229254 , n229248 , n229253 );
xor ( n229255 , n229247 , n229254 );
not ( n229256 , n217388 );
buf ( n229257 , n217076 );
not ( n229258 , n229257 );
not ( n229259 , n40724 );
or ( n229260 , n229258 , n229259 );
buf ( n229261 , n216928 );
not ( n229262 , n229261 );
or ( n229263 , n40724 , n229262 );
nand ( n229264 , n229260 , n229263 );
not ( n229265 , n229264 );
or ( n229266 , n229256 , n229265 );
nand ( n229267 , n228587 , n220046 );
nand ( n229268 , n229266 , n229267 );
xor ( n229269 , n229255 , n229268 );
not ( n229270 , n228780 );
not ( n229271 , n226271 );
not ( n229272 , n229271 );
or ( n229273 , n229270 , n229272 );
not ( n229274 , n216208 );
not ( n229275 , n225743 );
or ( n229276 , n229274 , n229275 );
nand ( n229277 , n225952 , n216207 );
nand ( n229278 , n229276 , n229277 );
nand ( n229279 , n229278 , n225948 );
nand ( n229280 , n229273 , n229279 );
not ( n229281 , n228792 );
not ( n229282 , n223197 );
or ( n229283 , n229281 , n229282 );
not ( n229284 , n221921 );
not ( n229285 , n226806 );
or ( n229286 , n229284 , n229285 );
nand ( n229287 , n223202 , n218980 );
nand ( n229288 , n229286 , n229287 );
nand ( n229289 , n229288 , n222769 );
nand ( n229290 , n229283 , n229289 );
xor ( n229291 , n229280 , n229290 );
or ( n229292 , n228270 , n228711 );
and ( n229293 , n227595 , n214960 );
not ( n229294 , n227595 );
and ( n229295 , n229294 , n214956 );
or ( n229296 , n229293 , n229295 );
not ( n229297 , n229296 );
or ( n229298 , n229297 , n228273 );
nand ( n229299 , n229292 , n229298 );
xor ( n229300 , n229291 , n229299 );
xor ( n229301 , n229269 , n229300 );
not ( n229302 , n228819 );
not ( n229303 , n222453 );
or ( n229304 , n229302 , n229303 );
and ( n229305 , n216293 , n225418 );
not ( n229306 , n216293 );
and ( n229307 , n229306 , n228817 );
or ( n229308 , n229305 , n229307 );
nand ( n229309 , n229308 , n223243 );
nand ( n229310 , n229304 , n229309 );
not ( n229311 , n228830 );
not ( n229312 , n224086 );
or ( n229313 , n229311 , n229312 );
not ( n229314 , n219102 );
not ( n229315 , n224095 );
or ( n229316 , n229314 , n229315 );
nand ( n229317 , n228828 , n220436 );
nand ( n229318 , n229316 , n229317 );
nand ( n229319 , n224090 , n229318 );
nand ( n229320 , n229313 , n229319 );
xor ( n229321 , n229310 , n229320 );
not ( n229322 , n228769 );
not ( n229323 , n226742 );
or ( n229324 , n229322 , n229323 );
not ( n229325 , n218514 );
not ( n229326 , n224844 );
or ( n229327 , n229325 , n229326 );
nand ( n229328 , n224929 , n216170 );
nand ( n229329 , n229327 , n229328 );
nand ( n229330 , n229329 , n224941 );
nand ( n229331 , n229324 , n229330 );
xor ( n229332 , n229321 , n229331 );
xor ( n229333 , n229301 , n229332 );
xor ( n229334 , n229269 , n229300 );
and ( n229335 , n229334 , n229332 );
and ( n229336 , n229269 , n229300 );
or ( n229337 , n229335 , n229336 );
not ( n229338 , n228635 );
not ( n229339 , n220162 );
or ( n229340 , n229338 , n229339 );
not ( n229341 , n41701 );
not ( n229342 , n221256 );
or ( n229343 , n229341 , n229342 );
nand ( n229344 , n225454 , n215428 );
nand ( n229345 , n229343 , n229344 );
nand ( n229346 , n229345 , n219778 );
nand ( n229347 , n229340 , n229346 );
not ( n229348 , n228646 );
not ( n229349 , n223223 );
or ( n229350 , n229348 , n229349 );
not ( n229351 , n225490 );
not ( n229352 , n223227 );
or ( n229353 , n229351 , n229352 );
nand ( n229354 , n220900 , n208726 );
nand ( n229355 , n229353 , n229354 );
nand ( n229356 , n229355 , n220929 );
nand ( n229357 , n229350 , n229356 );
xor ( n229358 , n229347 , n229357 );
not ( n229359 , n228808 );
not ( n229360 , n221625 );
or ( n229361 , n229359 , n229360 );
not ( n229362 , n224492 );
not ( n229363 , n221777 );
or ( n229364 , n229362 , n229363 );
nand ( n229365 , n221608 , n214642 );
nand ( n229366 , n229364 , n229365 );
nand ( n229367 , n229366 , n221387 );
nand ( n229368 , n229361 , n229367 );
xor ( n229369 , n229358 , n229368 );
xor ( n229370 , n229369 , n229075 );
xor ( n229371 , n229370 , n229079 );
xor ( n229372 , n229369 , n229075 );
and ( n229373 , n229372 , n229079 );
and ( n229374 , n229369 , n229075 );
or ( n229375 , n229373 , n229374 );
xor ( n229376 , n229083 , n228683 );
not ( n229377 , n226943 );
not ( n229378 , n228982 );
or ( n229379 , n229377 , n229378 );
and ( n229380 , n207936 , n220038 );
not ( n229381 , n207936 );
and ( n229382 , n229381 , n227912 );
or ( n229383 , n229380 , n229382 );
nand ( n229384 , n229383 , n220033 );
nand ( n229385 , n229379 , n229384 );
not ( n229386 , n228237 );
not ( n229387 , n227599 );
not ( n229388 , n229387 );
not ( n229389 , n220569 );
or ( n229390 , n229388 , n229389 );
nand ( n229391 , n224642 , n227599 );
nand ( n229392 , n229390 , n229391 );
not ( n229393 , n229392 );
or ( n229394 , n229386 , n229393 );
buf ( n229395 , n225478 );
nand ( n229396 , n228901 , n229395 );
nand ( n229397 , n229394 , n229396 );
xor ( n229398 , n229385 , n229397 );
not ( n229399 , n218467 );
not ( n229400 , n228911 );
or ( n229401 , n229399 , n229400 );
not ( n229402 , n217573 );
not ( n229403 , n226243 );
or ( n229404 , n229402 , n229403 );
nand ( n229405 , n228215 , n219390 );
nand ( n229406 , n229404 , n229405 );
nand ( n229407 , n229406 , n215137 );
nand ( n229408 , n229401 , n229407 );
xor ( n229409 , n229398 , n229408 );
xor ( n229410 , n229376 , n229409 );
xor ( n229411 , n229083 , n228683 );
and ( n229412 , n229411 , n229409 );
and ( n229413 , n229083 , n228683 );
or ( n229414 , n229412 , n229413 );
xor ( n229415 , n229087 , n229091 );
not ( n229416 , n215183 );
not ( n229417 , n228962 );
or ( n229418 , n229416 , n229417 );
and ( n229419 , n40409 , n218994 );
not ( n229420 , n40409 );
and ( n229421 , n229420 , n218990 );
or ( n229422 , n229419 , n229421 );
nand ( n229423 , n229422 , n221933 );
nand ( n229424 , n229418 , n229423 );
not ( n229425 , n219175 );
not ( n229426 , n217017 );
not ( n229427 , n223761 );
or ( n229428 , n229426 , n229427 );
nand ( n229429 , n40045 , n219583 );
nand ( n229430 , n229428 , n229429 );
not ( n229431 , n229430 );
or ( n229432 , n229425 , n229431 );
nand ( n229433 , n228939 , n217023 );
nand ( n229434 , n229432 , n229433 );
xor ( n229435 , n229424 , n229434 );
not ( n229436 , n223949 );
not ( n229437 , n226655 );
not ( n229438 , n228449 );
or ( n229439 , n229437 , n229438 );
nand ( n229440 , n219222 , n227927 );
nand ( n229441 , n229439 , n229440 );
not ( n229442 , n229441 );
or ( n229443 , n229436 , n229442 );
nand ( n229444 , n228893 , n227260 );
nand ( n229445 , n229443 , n229444 );
xor ( n229446 , n229435 , n229445 );
xor ( n229447 , n229415 , n229446 );
xor ( n229448 , n229087 , n229091 );
and ( n229449 , n229448 , n229446 );
and ( n229450 , n229087 , n229091 );
or ( n229451 , n229449 , n229450 );
not ( n229452 , n220280 );
not ( n229453 , n228878 );
or ( n229454 , n229452 , n229453 );
not ( n229455 , n215955 );
not ( n229456 , n226444 );
or ( n229457 , n229455 , n229456 );
nand ( n229458 , n40484 , n219358 );
nand ( n229459 , n229457 , n229458 );
nand ( n229460 , n229459 , n219353 );
nand ( n229461 , n229454 , n229460 );
not ( n229462 , n219731 );
not ( n229463 , n228929 );
or ( n229464 , n229462 , n229463 );
and ( n229465 , n40421 , n220538 );
not ( n229466 , n40421 );
and ( n229467 , n229466 , n219033 );
or ( n229468 , n229465 , n229467 );
nand ( n229469 , n229468 , n214458 );
nand ( n229470 , n229464 , n229469 );
xor ( n229471 , n229461 , n229470 );
not ( n229472 , n224624 );
not ( n229473 , n228948 );
or ( n229474 , n229472 , n229473 );
not ( n229475 , n219687 );
not ( n229476 , n222120 );
or ( n229477 , n229475 , n229476 );
nand ( n229478 , n40396 , n221283 );
nand ( n229479 , n229477 , n229478 );
nand ( n229480 , n229479 , n219314 );
nand ( n229481 , n229474 , n229480 );
xor ( n229482 , n229471 , n229481 );
xor ( n229483 , n229482 , n229233 );
xor ( n229484 , n228617 , n228655 );
xor ( n229485 , n229484 , n229015 );
xor ( n229486 , n229483 , n229485 );
xor ( n229487 , n229482 , n229233 );
and ( n229488 , n229487 , n229485 );
and ( n229489 , n229482 , n229233 );
or ( n229490 , n229488 , n229489 );
xor ( n229491 , n229178 , n229205 );
xor ( n229492 , n229491 , n228706 );
xor ( n229493 , n229178 , n229205 );
and ( n229494 , n229493 , n228706 );
and ( n229495 , n229178 , n229205 );
or ( n229496 , n229494 , n229495 );
xor ( n229497 , n228800 , n229333 );
xor ( n229498 , n229497 , n228886 );
xor ( n229499 , n228800 , n229333 );
and ( n229500 , n229499 , n228886 );
and ( n229501 , n228800 , n229333 );
or ( n229502 , n229500 , n229501 );
xor ( n229503 , n229347 , n229357 );
and ( n229504 , n229503 , n229368 );
and ( n229505 , n229347 , n229357 );
or ( n229506 , n229504 , n229505 );
xor ( n229507 , n228839 , n228991 );
xor ( n229508 , n229507 , n228922 );
xor ( n229509 , n228839 , n228991 );
and ( n229510 , n229509 , n228922 );
and ( n229511 , n228839 , n228991 );
or ( n229512 , n229510 , n229511 );
xor ( n229513 , n229371 , n228999 );
xor ( n229514 , n229513 , n229410 );
xor ( n229515 , n229371 , n228999 );
and ( n229516 , n229515 , n229410 );
and ( n229517 , n229371 , n228999 );
or ( n229518 , n229516 , n229517 );
xor ( n229519 , n229447 , n229005 );
xor ( n229520 , n229519 , n229492 );
xor ( n229521 , n229447 , n229005 );
and ( n229522 , n229521 , n229492 );
and ( n229523 , n229447 , n229005 );
or ( n229524 , n229522 , n229523 );
xor ( n229525 , n229486 , n229498 );
xor ( n229526 , n229525 , n229011 );
xor ( n229527 , n229486 , n229498 );
and ( n229528 , n229527 , n229011 );
and ( n229529 , n229486 , n229498 );
or ( n229530 , n229528 , n229529 );
xor ( n229531 , n229508 , n229021 );
xor ( n229532 , n229531 , n229514 );
xor ( n229533 , n229508 , n229021 );
and ( n229534 , n229533 , n229514 );
and ( n229535 , n229508 , n229021 );
or ( n229536 , n229534 , n229535 );
xor ( n229537 , n229027 , n229033 );
xor ( n229538 , n229537 , n229520 );
xor ( n229539 , n229027 , n229033 );
and ( n229540 , n229539 , n229520 );
and ( n229541 , n229027 , n229033 );
or ( n229542 , n229540 , n229541 );
xor ( n229543 , n229039 , n229526 );
xor ( n229544 , n229543 , n229532 );
xor ( n229545 , n229039 , n229526 );
and ( n229546 , n229545 , n229532 );
and ( n229547 , n229039 , n229526 );
or ( n229548 , n229546 , n229547 );
xor ( n229549 , n229045 , n229538 );
xor ( n229550 , n229549 , n229051 );
xor ( n229551 , n229045 , n229538 );
and ( n229552 , n229551 , n229051 );
and ( n229553 , n229045 , n229538 );
or ( n229554 , n229552 , n229553 );
xor ( n229555 , n229544 , n229057 );
xor ( n229556 , n229555 , n229550 );
xor ( n229557 , n229544 , n229057 );
and ( n229558 , n229557 , n229550 );
and ( n229559 , n229544 , n229057 );
or ( n229560 , n229558 , n229559 );
xor ( n229561 , n229310 , n229320 );
and ( n229562 , n229561 , n229331 );
and ( n229563 , n229310 , n229320 );
or ( n229564 , n229562 , n229563 );
xor ( n229565 , n229280 , n229290 );
and ( n229566 , n229565 , n229299 );
and ( n229567 , n229280 , n229290 );
or ( n229568 , n229566 , n229567 );
xor ( n229569 , n229247 , n229254 );
and ( n229570 , n229569 , n229268 );
and ( n229571 , n229247 , n229254 );
or ( n229572 , n229570 , n229571 );
xor ( n229573 , n229461 , n229470 );
and ( n229574 , n229573 , n229481 );
and ( n229575 , n229461 , n229470 );
or ( n229576 , n229574 , n229575 );
xor ( n229577 , n229424 , n229434 );
and ( n229578 , n229577 , n229445 );
and ( n229579 , n229424 , n229434 );
or ( n229580 , n229578 , n229579 );
xor ( n229581 , n229385 , n229397 );
and ( n229582 , n229581 , n229408 );
and ( n229583 , n229385 , n229397 );
or ( n229584 , n229582 , n229583 );
xor ( n229585 , n228617 , n228655 );
and ( n229586 , n229585 , n229015 );
and ( n229587 , n228617 , n228655 );
or ( n229588 , n229586 , n229587 );
not ( n229589 , n229133 );
not ( n229590 , n218221 );
or ( n229591 , n229589 , n229590 );
not ( n229592 , n218137 );
not ( n229593 , n218226 );
or ( n229594 , n229592 , n229593 );
nand ( n229595 , n218775 , n217116 );
nand ( n229596 , n229594 , n229595 );
nand ( n229597 , n229596 , n218533 );
nand ( n229598 , n229591 , n229597 );
not ( n229599 , n229147 );
not ( n229600 , n220480 );
or ( n229601 , n229599 , n229600 );
not ( n229602 , n218876 );
not ( n229603 , n221016 );
or ( n229604 , n229602 , n229603 );
nand ( n229605 , n220859 , n41249 );
nand ( n229606 , n229604 , n229605 );
nand ( n229607 , n229606 , n222376 );
nand ( n229608 , n229601 , n229607 );
xor ( n229609 , n229598 , n229608 );
not ( n229610 , n229159 );
or ( n229611 , n219791 , n229610 );
not ( n229612 , n219076 );
not ( n229613 , n218786 );
not ( n229614 , n219440 );
or ( n229615 , n229613 , n229614 );
nand ( n229616 , n221227 , n215989 );
nand ( n229617 , n229615 , n229616 );
not ( n229618 , n229617 );
or ( n229619 , n229612 , n229618 );
nand ( n229620 , n229611 , n229619 );
xor ( n229621 , n229609 , n229620 );
xor ( n229622 , n229598 , n229608 );
and ( n229623 , n229622 , n229620 );
and ( n229624 , n229598 , n229608 );
or ( n229625 , n229623 , n229624 );
not ( n229626 , n229345 );
not ( n229627 , n220163 );
or ( n229628 , n229626 , n229627 );
not ( n229629 , n216543 );
not ( n229630 , n229629 );
not ( n229631 , n220147 );
or ( n229632 , n229630 , n229631 );
nand ( n229633 , n220150 , n216543 );
nand ( n229634 , n229632 , n229633 );
nand ( n229635 , n220881 , n229634 );
nand ( n229636 , n229628 , n229635 );
not ( n229637 , n229355 );
not ( n229638 , n220919 );
or ( n229639 , n229637 , n229638 );
not ( n229640 , n225768 );
not ( n229641 , n220901 );
or ( n229642 , n229640 , n229641 );
nand ( n229643 , n222399 , n225769 );
nand ( n229644 , n229642 , n229643 );
nand ( n229645 , n229644 , n220636 );
nand ( n229646 , n229639 , n229645 );
xor ( n229647 , n229636 , n229646 );
not ( n229648 , n224120 );
not ( n229649 , n229366 );
or ( n229650 , n229648 , n229649 );
not ( n229651 , n214837 );
not ( n229652 , n221777 );
or ( n229653 , n229651 , n229652 );
nand ( n229654 , n221607 , n226698 );
nand ( n229655 , n229653 , n229654 );
not ( n229656 , n229655 );
or ( n229657 , n223176 , n229656 );
nand ( n229658 , n229650 , n229657 );
xor ( n229659 , n229647 , n229658 );
xor ( n229660 , n229636 , n229646 );
and ( n229661 , n229660 , n229658 );
and ( n229662 , n229636 , n229646 );
or ( n229663 , n229661 , n229662 );
xor ( n229664 , n229564 , n229568 );
not ( n229665 , n220985 );
not ( n229666 , n215113 );
not ( n229667 , n225795 );
not ( n229668 , n229667 );
or ( n229669 , n229666 , n229668 );
nand ( n229670 , n39713 , n217944 );
nand ( n229671 , n229669 , n229670 );
not ( n229672 , n229671 );
or ( n229673 , n229665 , n229672 );
nand ( n229674 , n229190 , n214717 );
nand ( n229675 , n229673 , n229674 );
xor ( n229676 , n229664 , n229675 );
xor ( n229677 , n229564 , n229568 );
and ( n229678 , n229677 , n229675 );
and ( n229679 , n229564 , n229568 );
or ( n229680 , n229678 , n229679 );
not ( n229681 , n216299 );
not ( n229682 , n229200 );
or ( n229683 , n229681 , n229682 );
or ( n229684 , n216810 , n39926 );
nand ( n229685 , n39926 , n216810 );
nand ( n229686 , n229684 , n229685 );
nand ( n229687 , n229686 , n220820 );
nand ( n229688 , n229683 , n229687 );
not ( n229689 , n213912 );
not ( n229690 , n213382 );
not ( n229691 , n209707 );
not ( n229692 , n229691 );
or ( n229693 , n229690 , n229692 );
not ( n229694 , n209708 );
nand ( n229695 , n229694 , n217715 );
nand ( n229696 , n229693 , n229695 );
not ( n229697 , n229696 );
or ( n229698 , n229689 , n229697 );
nand ( n229699 , n229219 , n217969 );
nand ( n229700 , n229698 , n229699 );
xor ( n229701 , n229688 , n229700 );
not ( n229702 , n216336 );
not ( n229703 , n213735 );
buf ( n229704 , n228657 );
not ( n229705 , n229704 );
or ( n229706 , n229703 , n229705 );
or ( n229707 , n227667 , n213735 );
nand ( n229708 , n229706 , n229707 );
not ( n229709 , n229708 );
or ( n229710 , n229702 , n229709 );
nand ( n229711 , n229229 , n213577 );
nand ( n229712 , n229710 , n229711 );
xor ( n229713 , n229701 , n229712 );
xor ( n229714 , n229688 , n229700 );
and ( n229715 , n229714 , n229712 );
and ( n229716 , n229688 , n229700 );
or ( n229717 , n229715 , n229716 );
xor ( n229718 , n229572 , n229621 );
not ( n229719 , n229296 );
not ( n229720 , n227734 );
or ( n229721 , n229719 , n229720 );
not ( n229722 , n217044 );
not ( n229723 , n228278 );
or ( n229724 , n229722 , n229723 );
nand ( n229725 , n227595 , n215131 );
nand ( n229726 , n229724 , n229725 );
nand ( n229727 , n227737 , n229726 );
nand ( n229728 , n229721 , n229727 );
not ( n229729 , n229252 );
not ( n229730 , n229729 );
not ( n229731 , n228858 );
or ( n229732 , n229730 , n229731 );
not ( n229733 , n213583 );
not ( n229734 , n229249 );
or ( n229735 , n229733 , n229734 );
nand ( n229736 , n228726 , n214134 );
nand ( n229737 , n229735 , n229736 );
not ( n229738 , n228116 );
nand ( n229739 , n229737 , n229738 );
nand ( n229740 , n229732 , n229739 );
xor ( n229741 , n229728 , n229740 );
not ( n229742 , n37672 );
not ( n229743 , n37577 );
nand ( n229744 , n229743 , n37100 );
nor ( n229745 , n36730 , n37577 );
nand ( n229746 , n229745 , n36320 );
not ( n229747 , n36580 );
not ( n229748 , n37576 );
or ( n229749 , n229747 , n229748 );
nand ( n229750 , n229749 , n37534 );
not ( n229751 , n229750 );
nand ( n229752 , n229744 , n229746 , n229751 );
not ( n229753 , n229752 );
or ( n229754 , n229742 , n229753 );
not ( n229755 , n37672 );
nand ( n229756 , n229744 , n229751 , n229746 , n229755 );
nand ( n229757 , n229754 , n229756 );
buf ( n229758 , n229757 );
buf ( n229759 , n229758 );
or ( n229760 , n229759 , n213751 );
buf ( n229761 , n229758 );
not ( n229762 , n229761 );
or ( n229763 , n229762 , n215999 );
nand ( n229764 , n229760 , n229763 );
not ( n229765 , n229764 );
not ( n229766 , n229757 );
not ( n229767 , n229766 );
not ( n229768 , n229115 );
or ( n229769 , n229767 , n229768 );
nand ( n229770 , n229758 , n229121 );
nand ( n229771 , n229769 , n229770 );
nor ( n229772 , n229123 , n229771 );
buf ( n229773 , n229772 );
not ( n229774 , n229773 );
or ( n229775 , n229765 , n229774 );
not ( n229776 , n229123 );
not ( n229777 , n229776 );
not ( n229778 , n218224 );
not ( n229779 , n229762 );
or ( n229780 , n229778 , n229779 );
nand ( n229781 , n229761 , n216076 );
nand ( n229782 , n229780 , n229781 );
nand ( n229783 , n229777 , n229782 );
nand ( n229784 , n229775 , n229783 );
xor ( n229785 , n229741 , n229784 );
xor ( n229786 , n229718 , n229785 );
xor ( n229787 , n229572 , n229621 );
and ( n229788 , n229787 , n229785 );
and ( n229789 , n229572 , n229621 );
or ( n229790 , n229788 , n229789 );
not ( n229791 , n229329 );
not ( n229792 , n226742 );
or ( n229793 , n229791 , n229792 );
not ( n229794 , n216934 );
not ( n229795 , n224929 );
not ( n229796 , n229795 );
or ( n229797 , n229794 , n229796 );
nand ( n229798 , n224929 , n216940 );
nand ( n229799 , n229797 , n229798 );
nand ( n229800 , n229799 , n226745 );
nand ( n229801 , n229793 , n229800 );
not ( n229802 , n229278 );
not ( n229803 , n229271 );
or ( n229804 , n229802 , n229803 );
not ( n229805 , n215075 );
not ( n229806 , n225940 );
not ( n229807 , n229806 );
not ( n229808 , n229807 );
or ( n229809 , n229805 , n229808 );
nand ( n229810 , n225952 , n215899 );
nand ( n229811 , n229809 , n229810 );
nand ( n229812 , n228775 , n229811 );
nand ( n229813 , n229804 , n229812 );
xor ( n229814 , n229801 , n229813 );
not ( n229815 , n229245 );
not ( n229816 , n227848 );
not ( n229817 , n229816 );
or ( n229818 , n229815 , n229817 );
not ( n229819 , n216964 );
not ( n229820 , n226648 );
not ( n229821 , n229820 );
or ( n229822 , n229819 , n229821 );
buf ( n229823 , n226647 );
nand ( n229824 , n229823 , n214678 );
nand ( n229825 , n229822 , n229824 );
nand ( n229826 , n226885 , n229825 );
nand ( n229827 , n229818 , n229826 );
xor ( n229828 , n229814 , n229827 );
xor ( n229829 , n229828 , n229659 );
not ( n229830 , n229308 );
not ( n229831 , n222453 );
or ( n229832 , n229830 , n229831 );
not ( n229833 , n224037 );
not ( n229834 , n222458 );
or ( n229835 , n229833 , n229834 );
not ( n229836 , n225418 );
nand ( n229837 , n229836 , n214821 );
nand ( n229838 , n229835 , n229837 );
nand ( n229839 , n229838 , n222158 );
nand ( n229840 , n229832 , n229839 );
not ( n229841 , n229288 );
not ( n229842 , n223591 );
or ( n229843 , n229841 , n229842 );
not ( n229844 , n214468 );
not ( n229845 , n225914 );
or ( n229846 , n229844 , n229845 );
nand ( n229847 , n223182 , n221494 );
nand ( n229848 , n229846 , n229847 );
nand ( n229849 , n229848 , n222769 );
nand ( n229850 , n229843 , n229849 );
xor ( n229851 , n229840 , n229850 );
not ( n229852 , n229318 );
not ( n229853 , n224087 );
or ( n229854 , n229852 , n229853 );
not ( n229855 , n219343 );
not ( n229856 , n224975 );
or ( n229857 , n229855 , n229856 );
nand ( n229858 , n224974 , n219348 );
nand ( n229859 , n229857 , n229858 );
nand ( n229860 , n227782 , n229859 );
nand ( n229861 , n229854 , n229860 );
xor ( n229862 , n229851 , n229861 );
xor ( n229863 , n229829 , n229862 );
xor ( n229864 , n229828 , n229659 );
and ( n229865 , n229864 , n229862 );
and ( n229866 , n229828 , n229659 );
or ( n229867 , n229865 , n229866 );
xor ( n229868 , n229576 , n229580 );
xor ( n229869 , n229868 , n229182 );
xor ( n229870 , n229576 , n229580 );
and ( n229871 , n229870 , n229182 );
and ( n229872 , n229576 , n229580 );
or ( n229873 , n229871 , n229872 );
not ( n229874 , n221933 );
and ( n229875 , n221742 , n218994 );
not ( n229876 , n221742 );
and ( n229877 , n229876 , n218990 );
or ( n229878 , n229875 , n229877 );
not ( n229879 , n229878 );
or ( n229880 , n229874 , n229879 );
nand ( n229881 , n219332 , n229422 );
nand ( n229882 , n229880 , n229881 );
not ( n229883 , n220033 );
not ( n229884 , n226292 );
not ( n229885 , n222500 );
or ( n229886 , n229884 , n229885 );
not ( n229887 , n226292 );
nand ( n229888 , n40668 , n229887 );
nand ( n229889 , n229886 , n229888 );
not ( n229890 , n229889 );
or ( n229891 , n229883 , n229890 );
nand ( n229892 , n229383 , n226943 );
nand ( n229893 , n229891 , n229892 );
xor ( n229894 , n229882 , n229893 );
not ( n229895 , n223949 );
not ( n229896 , n226655 );
not ( n229897 , n221687 );
or ( n229898 , n229896 , n229897 );
nand ( n229899 , n219522 , n227927 );
nand ( n229900 , n229898 , n229899 );
not ( n229901 , n229900 );
or ( n229902 , n229895 , n229901 );
nand ( n229903 , n229441 , n227260 );
nand ( n229904 , n229902 , n229903 );
xor ( n229905 , n229894 , n229904 );
xor ( n229906 , n229905 , n229584 );
xor ( n229907 , n229906 , n229588 );
xor ( n229908 , n229905 , n229584 );
and ( n229909 , n229908 , n229588 );
and ( n229910 , n229905 , n229584 );
or ( n229911 , n229909 , n229910 );
not ( n229912 , n222185 );
not ( n229913 , n219033 );
not ( n229914 , n223368 );
or ( n229915 , n229913 , n229914 );
nand ( n229916 , n222513 , n219034 );
nand ( n229917 , n229915 , n229916 );
not ( n229918 , n229917 );
or ( n229919 , n229912 , n229918 );
nand ( n229920 , n229468 , n219731 );
nand ( n229921 , n229919 , n229920 );
not ( n229922 , n217023 );
not ( n229923 , n229430 );
or ( n229924 , n229922 , n229923 );
not ( n229925 , n217017 );
not ( n229926 , n226961 );
or ( n229927 , n229925 , n229926 );
not ( n229928 , n226961 );
nand ( n229929 , n229928 , n218661 );
nand ( n229930 , n229927 , n229929 );
nand ( n229931 , n229930 , n219175 );
nand ( n229932 , n229924 , n229931 );
xor ( n229933 , n229921 , n229932 );
not ( n229934 , n219314 );
not ( n229935 , n219687 );
buf ( n229936 , n40181 );
not ( n229937 , n229936 );
or ( n229938 , n229935 , n229937 );
nand ( n229939 , n40182 , n221283 );
nand ( n229940 , n229938 , n229939 );
not ( n229941 , n229940 );
or ( n229942 , n229934 , n229941 );
nand ( n229943 , n229479 , n216204 );
nand ( n229944 , n229942 , n229943 );
xor ( n229945 , n229933 , n229944 );
xor ( n229946 , n229209 , n229945 );
nand ( n229947 , n229121 , n213750 );
not ( n229948 , n213751 );
not ( n229949 , n229115 );
or ( n229950 , n229948 , n229949 );
nand ( n229951 , n229950 , n228726 );
and ( n229952 , n229947 , n229761 , n229951 );
not ( n229953 , n220067 );
not ( n229954 , n217616 );
not ( n229955 , n220823 );
or ( n229956 , n229954 , n229955 );
nand ( n229957 , n217714 , n218253 );
nand ( n229958 , n229956 , n229957 );
not ( n229959 , n229958 );
or ( n229960 , n229953 , n229959 );
nand ( n229961 , n229097 , n217631 );
nand ( n229962 , n229960 , n229961 );
xor ( n229963 , n229952 , n229962 );
buf ( n229964 , n217388 );
not ( n229965 , n229964 );
not ( n229966 , n229261 );
not ( n229967 , n218268 );
or ( n229968 , n229966 , n229967 );
nand ( n229969 , n219594 , n229262 );
nand ( n229970 , n229968 , n229969 );
not ( n229971 , n229970 );
or ( n229972 , n229965 , n229971 );
not ( n229973 , n219368 );
not ( n229974 , n229973 );
nand ( n229975 , n229264 , n229974 );
nand ( n229976 , n229972 , n229975 );
xor ( n229977 , n229963 , n229976 );
not ( n229978 , n220272 );
not ( n229979 , n217542 );
not ( n229980 , n223330 );
or ( n229981 , n229979 , n229980 );
nand ( n229982 , n223333 , n216989 );
nand ( n229983 , n229981 , n229982 );
not ( n229984 , n229983 );
or ( n229985 , n229978 , n229984 );
nand ( n229986 , n229459 , n220280 );
nand ( n229987 , n229985 , n229986 );
xor ( n229988 , n229977 , n229987 );
xor ( n229989 , n229946 , n229988 );
xor ( n229990 , n229209 , n229945 );
and ( n229991 , n229990 , n229988 );
and ( n229992 , n229209 , n229945 );
or ( n229993 , n229991 , n229992 );
not ( n229994 , n225478 );
not ( n229995 , n229392 );
or ( n229996 , n229994 , n229995 );
not ( n229997 , n216422 );
not ( n229998 , n220204 );
or ( n229999 , n229997 , n229998 );
nand ( n230000 , n218911 , n227602 );
nand ( n230001 , n229999 , n230000 );
nand ( n230002 , n230001 , n219501 );
nand ( n230003 , n229996 , n230002 );
not ( n230004 , n215137 );
not ( n230005 , n217573 );
not ( n230006 , n226712 );
or ( n230007 , n230005 , n230006 );
nand ( n230008 , n39607 , n215388 );
nand ( n230009 , n230007 , n230008 );
not ( n230010 , n230009 );
or ( n230011 , n230004 , n230010 );
nand ( n230012 , n229406 , n218467 );
nand ( n230013 , n230011 , n230012 );
xor ( n230014 , n230003 , n230013 );
xor ( n230015 , n230014 , n229140 );
xor ( n230016 , n230015 , n229713 );
xor ( n230017 , n230016 , n229676 );
xor ( n230018 , n230015 , n229713 );
and ( n230019 , n230018 , n229676 );
and ( n230020 , n230015 , n229713 );
or ( n230021 , n230019 , n230020 );
xor ( n230022 , n229166 , n229506 );
not ( n230023 , n217142 );
not ( n230024 , n214818 );
not ( n230025 , n39286 );
not ( n230026 , n230025 );
or ( n230027 , n230024 , n230026 );
nand ( n230028 , n39286 , n214824 );
nand ( n230029 , n230027 , n230028 );
not ( n230030 , n230029 );
or ( n230031 , n230023 , n230030 );
nand ( n230032 , n229171 , n213874 );
nand ( n230033 , n230031 , n230032 );
xor ( n230034 , n230022 , n230033 );
xor ( n230035 , n230034 , n229337 );
xor ( n230036 , n230035 , n229237 );
xor ( n230037 , n230034 , n229337 );
and ( n230038 , n230037 , n229237 );
and ( n230039 , n230034 , n229337 );
or ( n230040 , n230038 , n230039 );
xor ( n230041 , n229863 , n229786 );
xor ( n230042 , n230041 , n229375 );
xor ( n230043 , n229863 , n229786 );
and ( n230044 , n230043 , n229375 );
and ( n230045 , n229863 , n229786 );
or ( n230046 , n230044 , n230045 );
xor ( n230047 , n229840 , n229850 );
and ( n230048 , n230047 , n229861 );
and ( n230049 , n229840 , n229850 );
or ( n230050 , n230048 , n230049 );
xor ( n230051 , n229451 , n229414 );
xor ( n230052 , n230051 , n229869 );
xor ( n230053 , n229451 , n229414 );
and ( n230054 , n230053 , n229869 );
and ( n230055 , n229451 , n229414 );
or ( n230056 , n230054 , n230055 );
xor ( n230057 , n229490 , n229907 );
xor ( n230058 , n230057 , n229496 );
xor ( n230059 , n229490 , n229907 );
and ( n230060 , n230059 , n229496 );
and ( n230061 , n229490 , n229907 );
or ( n230062 , n230060 , n230061 );
xor ( n230063 , n229989 , n230036 );
xor ( n230064 , n230063 , n230017 );
xor ( n230065 , n229989 , n230036 );
and ( n230066 , n230065 , n230017 );
and ( n230067 , n229989 , n230036 );
or ( n230068 , n230066 , n230067 );
xor ( n230069 , n229502 , n229512 );
xor ( n230070 , n230069 , n230042 );
xor ( n230071 , n229502 , n229512 );
and ( n230072 , n230071 , n230042 );
and ( n230073 , n229502 , n229512 );
or ( n230074 , n230072 , n230073 );
xor ( n230075 , n230052 , n229518 );
xor ( n230076 , n230075 , n230058 );
xor ( n230077 , n230052 , n229518 );
and ( n230078 , n230077 , n230058 );
and ( n230079 , n230052 , n229518 );
or ( n230080 , n230078 , n230079 );
xor ( n230081 , n229524 , n229530 );
xor ( n230082 , n230081 , n230064 );
xor ( n230083 , n229524 , n229530 );
and ( n230084 , n230083 , n230064 );
and ( n230085 , n229524 , n229530 );
or ( n230086 , n230084 , n230085 );
xor ( n230087 , n230070 , n229536 );
xor ( n230088 , n230087 , n230076 );
xor ( n230089 , n230070 , n229536 );
and ( n230090 , n230089 , n230076 );
and ( n230091 , n230070 , n229536 );
or ( n230092 , n230090 , n230091 );
xor ( n230093 , n229542 , n230082 );
xor ( n230094 , n230093 , n229548 );
xor ( n230095 , n229542 , n230082 );
and ( n230096 , n230095 , n229548 );
and ( n230097 , n229542 , n230082 );
or ( n230098 , n230096 , n230097 );
xor ( n230099 , n230088 , n230094 );
xor ( n230100 , n230099 , n229554 );
xor ( n230101 , n230088 , n230094 );
and ( n230102 , n230101 , n229554 );
and ( n230103 , n230088 , n230094 );
or ( n230104 , n230102 , n230103 );
xor ( n230105 , n229801 , n229813 );
and ( n230106 , n230105 , n229827 );
and ( n230107 , n229801 , n229813 );
or ( n230108 , n230106 , n230107 );
xor ( n230109 , n229728 , n229740 );
and ( n230110 , n230109 , n229784 );
and ( n230111 , n229728 , n229740 );
or ( n230112 , n230110 , n230111 );
xor ( n230113 , n229963 , n229976 );
and ( n230114 , n230113 , n229987 );
and ( n230115 , n229963 , n229976 );
or ( n230116 , n230114 , n230115 );
xor ( n230117 , n229921 , n229932 );
and ( n230118 , n230117 , n229944 );
and ( n230119 , n229921 , n229932 );
or ( n230120 , n230118 , n230119 );
xor ( n230121 , n229882 , n229893 );
and ( n230122 , n230121 , n229904 );
and ( n230123 , n229882 , n229893 );
or ( n230124 , n230122 , n230123 );
xor ( n230125 , n230003 , n230013 );
and ( n230126 , n230125 , n229140 );
and ( n230127 , n230003 , n230013 );
or ( n230128 , n230126 , n230127 );
xor ( n230129 , n229166 , n229506 );
and ( n230130 , n230129 , n230033 );
and ( n230131 , n229166 , n229506 );
or ( n230132 , n230130 , n230131 );
not ( n230133 , n37574 );
nand ( n230134 , n37100 , n230133 );
nor ( n230135 , n229105 , n37574 );
nand ( n230136 , n229103 , n230135 );
and ( n230137 , n37573 , n36580 );
nor ( n230138 , n230137 , n37528 );
nand ( n230139 , n230134 , n230136 , n230138 );
not ( n230140 , n37540 );
nand ( n230141 , n230140 , n37412 );
not ( n230142 , n230141 );
and ( n230143 , n230139 , n230142 );
not ( n230144 , n230139 );
and ( n230145 , n230144 , n230141 );
nor ( n230146 , n230143 , n230145 );
not ( n230147 , n230146 );
or ( n230148 , n229766 , n230147 );
not ( n230149 , n230146 );
not ( n230150 , n229757 );
nand ( n230151 , n230149 , n230150 );
nand ( n230152 , n230148 , n230151 );
not ( n230153 , n230152 );
and ( n230154 , n230153 , n215999 );
not ( n230155 , n229596 );
not ( n230156 , n219836 );
or ( n230157 , n230155 , n230156 );
and ( n230158 , n41069 , n224497 );
not ( n230159 , n41069 );
and ( n230160 , n230159 , n218256 );
nor ( n230161 , n230158 , n230160 );
nand ( n230162 , n230161 , n218533 );
nand ( n230163 , n230157 , n230162 );
xor ( n230164 , n230154 , n230163 );
not ( n230165 , n229606 );
or ( n230166 , n225499 , n230165 );
not ( n230167 , n216859 );
not ( n230168 , n223671 );
not ( n230169 , n230168 );
or ( n230170 , n230167 , n230169 );
not ( n230171 , n219050 );
nand ( n230172 , n230171 , n220126 );
nand ( n230173 , n230170 , n230172 );
not ( n230174 , n230173 );
or ( n230175 , n218456 , n230174 );
nand ( n230176 , n230166 , n230175 );
xor ( n230177 , n230164 , n230176 );
xor ( n230178 , n230154 , n230163 );
and ( n230179 , n230178 , n230176 );
and ( n230180 , n230154 , n230163 );
or ( n230181 , n230179 , n230180 );
not ( n230182 , n229617 );
not ( n230183 , n219435 );
or ( n230184 , n230182 , n230183 );
not ( n230185 , n219902 );
not ( n230186 , n219419 );
or ( n230187 , n230185 , n230186 );
nand ( n230188 , n220180 , n219899 );
nand ( n230189 , n230187 , n230188 );
nand ( n230190 , n219076 , n230189 );
nand ( n230191 , n230184 , n230190 );
not ( n230192 , n229634 );
not ( n230193 , n220163 );
or ( n230194 , n230192 , n230193 );
not ( n230195 , n208717 );
not ( n230196 , n222412 );
or ( n230197 , n230195 , n230196 );
nand ( n230198 , n220145 , n215793 );
nand ( n230199 , n230197 , n230198 );
nand ( n230200 , n219779 , n230199 );
nand ( n230201 , n230194 , n230200 );
xor ( n230202 , n230191 , n230201 );
not ( n230203 , n229644 );
or ( n230204 , n228639 , n230203 );
not ( n230205 , n41701 );
not ( n230206 , n220904 );
or ( n230207 , n230205 , n230206 );
nand ( n230208 , n220899 , n216339 );
nand ( n230209 , n230207 , n230208 );
not ( n230210 , n230209 );
or ( n230211 , n220928 , n230210 );
nand ( n230212 , n230204 , n230211 );
xor ( n230213 , n230202 , n230212 );
xor ( n230214 , n230191 , n230201 );
and ( n230215 , n230214 , n230212 );
and ( n230216 , n230191 , n230201 );
or ( n230217 , n230215 , n230216 );
not ( n230218 , n214818 );
not ( n230219 , n229217 );
not ( n230220 , n230219 );
or ( n230221 , n230218 , n230220 );
not ( n230222 , n229214 );
buf ( n230223 , n230222 );
nand ( n230224 , n230223 , n220300 );
nand ( n230225 , n230221 , n230224 );
not ( n230226 , n230225 );
not ( n230227 , n217142 );
or ( n230228 , n230226 , n230227 );
nand ( n230229 , n230029 , n213874 );
nand ( n230230 , n230228 , n230229 );
xor ( n230231 , n230230 , n230050 );
xor ( n230232 , n230231 , n230108 );
xor ( n230233 , n230230 , n230050 );
and ( n230234 , n230233 , n230108 );
and ( n230235 , n230230 , n230050 );
or ( n230236 , n230234 , n230235 );
not ( n230237 , n214717 );
not ( n230238 , n229671 );
or ( n230239 , n230237 , n230238 );
not ( n230240 , n218855 );
not ( n230241 , n39747 );
not ( n230242 , n230241 );
or ( n230243 , n230240 , n230242 );
nand ( n230244 , n228215 , n216037 );
nand ( n230245 , n230243 , n230244 );
nand ( n230246 , n230245 , n220985 );
nand ( n230247 , n230239 , n230246 );
xor ( n230248 , n230112 , n230247 );
not ( n230249 , n229686 );
not ( n230250 , n216299 );
or ( n230251 , n230249 , n230250 );
not ( n230252 , n216810 );
not ( n230253 , n227224 );
or ( n230254 , n230252 , n230253 );
nand ( n230255 , n227223 , n221307 );
nand ( n230256 , n230254 , n230255 );
not ( n230257 , n230256 );
or ( n230258 , n230257 , n220819 );
nand ( n230259 , n230251 , n230258 );
xor ( n230260 , n230248 , n230259 );
xor ( n230261 , n230112 , n230247 );
and ( n230262 , n230261 , n230259 );
and ( n230263 , n230112 , n230247 );
or ( n230264 , n230262 , n230263 );
not ( n230265 , n213577 );
not ( n230266 , n229708 );
or ( n230267 , n230265 , n230266 );
not ( n230268 , n213735 );
not ( n230269 , n228164 );
buf ( n230270 , n230269 );
not ( n230271 , n230270 );
or ( n230272 , n230268 , n230271 );
not ( n230273 , n230269 );
nand ( n230274 , n230273 , n213732 );
nand ( n230275 , n230272 , n230274 );
nand ( n230276 , n230275 , n216336 );
nand ( n230277 , n230267 , n230276 );
not ( n230278 , n219175 );
not ( n230279 , n219577 );
not ( n230280 , n225344 );
not ( n230281 , n230280 );
or ( n230282 , n230279 , n230281 );
nand ( n230283 , n228195 , n218661 );
nand ( n230284 , n230282 , n230283 );
not ( n230285 , n230284 );
or ( n230286 , n230278 , n230285 );
nand ( n230287 , n229930 , n217023 );
nand ( n230288 , n230286 , n230287 );
xor ( n230289 , n230277 , n230288 );
xor ( n230290 , n230289 , n230213 );
xor ( n230291 , n230277 , n230288 );
and ( n230292 , n230291 , n230213 );
and ( n230293 , n230277 , n230288 );
or ( n230294 , n230292 , n230293 );
not ( n230295 , n229655 );
not ( n230296 , n223579 );
or ( n230297 , n230295 , n230296 );
not ( n230298 , n225490 );
not ( n230299 , n221777 );
or ( n230300 , n230298 , n230299 );
nand ( n230301 , n219690 , n223584 );
nand ( n230302 , n230300 , n230301 );
nand ( n230303 , n223587 , n230302 );
nand ( n230304 , n230297 , n230303 );
not ( n230305 , n229838 );
not ( n230306 , n222453 );
or ( n230307 , n230305 , n230306 );
not ( n230308 , n222428 );
not ( n230309 , n221894 );
or ( n230310 , n230308 , n230309 );
or ( n230311 , n228817 , n224496 );
nand ( n230312 , n230310 , n230311 );
nand ( n230313 , n222158 , n230312 );
nand ( n230314 , n230307 , n230313 );
xor ( n230315 , n230304 , n230314 );
not ( n230316 , n229848 );
not ( n230317 , n223591 );
or ( n230318 , n230316 , n230317 );
not ( n230319 , n216293 );
not ( n230320 , n223595 );
or ( n230321 , n230319 , n230320 );
nand ( n230322 , n223201 , n216290 );
nand ( n230323 , n230321 , n230322 );
nand ( n230324 , n222769 , n230323 );
nand ( n230325 , n230318 , n230324 );
xor ( n230326 , n230315 , n230325 );
xor ( n230327 , n230177 , n230326 );
not ( n230328 , n229825 );
not ( n230329 , n227849 );
or ( n230330 , n230328 , n230329 );
not ( n230331 , n216208 );
not ( n230332 , n229820 );
or ( n230333 , n230331 , n230332 );
nand ( n230334 , n229823 , n216207 );
nand ( n230335 , n230333 , n230334 );
nand ( n230336 , n230335 , n227241 );
nand ( n230337 , n230330 , n230336 );
not ( n230338 , n229726 );
not ( n230339 , n228270 );
not ( n230340 , n230339 );
or ( n230341 , n230338 , n230340 );
not ( n230342 , n214537 );
not ( n230343 , n228278 );
or ( n230344 , n230342 , n230343 );
nand ( n230345 , n228274 , n214899 );
nand ( n230346 , n230344 , n230345 );
nand ( n230347 , n227737 , n230346 );
nand ( n230348 , n230341 , n230347 );
xor ( n230349 , n230337 , n230348 );
not ( n230350 , n229737 );
not ( n230351 , n228860 );
or ( n230352 , n230350 , n230351 );
not ( n230353 , n214956 );
not ( n230354 , n228847 );
or ( n230355 , n230353 , n230354 );
nand ( n230356 , n228726 , n214960 );
nand ( n230357 , n230355 , n230356 );
nand ( n230358 , n229738 , n230357 );
nand ( n230359 , n230352 , n230358 );
xor ( n230360 , n230349 , n230359 );
xor ( n230361 , n230327 , n230360 );
xor ( n230362 , n230177 , n230326 );
and ( n230363 , n230362 , n230360 );
and ( n230364 , n230177 , n230326 );
or ( n230365 , n230363 , n230364 );
not ( n230366 , n229859 );
not ( n230367 , n224086 );
or ( n230368 , n230366 , n230367 );
not ( n230369 , n223989 );
not ( n230370 , n230369 );
not ( n230371 , n221921 );
or ( n230372 , n230370 , n230371 );
nand ( n230373 , n224974 , n218980 );
nand ( n230374 , n230372 , n230373 );
nand ( n230375 , n224090 , n230374 );
nand ( n230376 , n230368 , n230375 );
not ( n230377 , n229799 );
not ( n230378 , n226742 );
or ( n230379 , n230377 , n230378 );
not ( n230380 , n219102 );
not ( n230381 , n226747 );
or ( n230382 , n230380 , n230381 );
nand ( n230383 , n224929 , n220436 );
nand ( n230384 , n230382 , n230383 );
nand ( n230385 , n230384 , n226745 );
nand ( n230386 , n230379 , n230385 );
xor ( n230387 , n230376 , n230386 );
not ( n230388 , n229811 );
not ( n230389 , n226272 );
not ( n230390 , n230389 );
not ( n230391 , n230390 );
or ( n230392 , n230388 , n230391 );
not ( n230393 , n218514 );
not ( n230394 , n226276 );
or ( n230395 , n230393 , n230394 );
nand ( n230396 , n229806 , n216170 );
nand ( n230397 , n230395 , n230396 );
nand ( n230398 , n228775 , n230397 );
nand ( n230399 , n230392 , n230398 );
xor ( n230400 , n230387 , n230399 );
xor ( n230401 , n230400 , n230116 );
xor ( n230402 , n230401 , n230120 );
xor ( n230403 , n230400 , n230116 );
and ( n230404 , n230403 , n230120 );
and ( n230405 , n230400 , n230116 );
or ( n230406 , n230404 , n230405 );
not ( n230407 , n229782 );
not ( n230408 , n229773 );
or ( n230409 , n230407 , n230408 );
and ( n230410 , n213347 , n229766 );
not ( n230411 , n213347 );
and ( n230412 , n230411 , n229758 );
nor ( n230413 , n230410 , n230412 );
not ( n230414 , n230413 );
nand ( n230415 , n230414 , n229777 );
nand ( n230416 , n230409 , n230415 );
and ( n230417 , n229952 , n229962 );
xor ( n230418 , n230416 , n230417 );
not ( n230419 , n220067 );
not ( n230420 , n217614 );
not ( n230421 , n217964 );
or ( n230422 , n230420 , n230421 );
nand ( n230423 , n208002 , n218253 );
nand ( n230424 , n230422 , n230423 );
not ( n230425 , n230424 );
or ( n230426 , n230419 , n230425 );
nand ( n230427 , n229958 , n220059 );
nand ( n230428 , n230426 , n230427 );
xor ( n230429 , n230418 , n230428 );
xor ( n230430 , n230124 , n230429 );
xor ( n230431 , n230430 , n229717 );
xor ( n230432 , n230124 , n230429 );
and ( n230433 , n230432 , n229717 );
and ( n230434 , n230124 , n230429 );
or ( n230435 , n230433 , n230434 );
not ( n230436 , n228237 );
not ( n230437 , n229387 );
not ( n230438 , n219880 );
or ( n230439 , n230437 , n230438 );
not ( n230440 , n222081 );
nand ( n230441 , n230440 , n227599 );
nand ( n230442 , n230439 , n230441 );
not ( n230443 , n230442 );
or ( n230444 , n230436 , n230443 );
nand ( n230445 , n230001 , n229395 );
nand ( n230446 , n230444 , n230445 );
not ( n230447 , n229964 );
not ( n230448 , n229261 );
not ( n230449 , n219238 );
or ( n230450 , n230448 , n230449 );
nand ( n230451 , n220568 , n229257 );
nand ( n230452 , n230450 , n230451 );
not ( n230453 , n230452 );
or ( n230454 , n230447 , n230453 );
nand ( n230455 , n229970 , n219368 );
nand ( n230456 , n230454 , n230455 );
xor ( n230457 , n230446 , n230456 );
not ( n230458 , n215383 );
not ( n230459 , n217573 );
not ( n230460 , n227201 );
or ( n230461 , n230459 , n230460 );
not ( n230462 , n228184 );
nand ( n230463 , n230462 , n217397 );
nand ( n230464 , n230461 , n230463 );
not ( n230465 , n230464 );
or ( n230466 , n230458 , n230465 );
nand ( n230467 , n230009 , n218467 );
nand ( n230468 , n230466 , n230467 );
xor ( n230469 , n230457 , n230468 );
xor ( n230470 , n230132 , n230469 );
xor ( n230471 , n230470 , n230128 );
xor ( n230472 , n230132 , n230469 );
and ( n230473 , n230472 , n230128 );
and ( n230474 , n230132 , n230469 );
or ( n230475 , n230473 , n230474 );
not ( n230476 , n222185 );
not ( n230477 , n219033 );
not ( n230478 , n223721 );
or ( n230479 , n230477 , n230478 );
nand ( n230480 , n223722 , n226002 );
nand ( n230481 , n230479 , n230480 );
not ( n230482 , n230481 );
or ( n230483 , n230476 , n230482 );
nand ( n230484 , n229917 , n219731 );
nand ( n230485 , n230483 , n230484 );
not ( n230486 , n217552 );
not ( n230487 , n229983 );
or ( n230488 , n230486 , n230487 );
not ( n230489 , n215955 );
not ( n230490 , n223765 );
not ( n230491 , n230490 );
or ( n230492 , n230489 , n230491 );
nand ( n230493 , n223765 , n219358 );
nand ( n230494 , n230492 , n230493 );
nand ( n230495 , n230494 , n220272 );
nand ( n230496 , n230488 , n230495 );
xor ( n230497 , n230485 , n230496 );
not ( n230498 , n219314 );
and ( n230499 , n223748 , n219687 );
not ( n230500 , n223748 );
and ( n230501 , n230500 , n221283 );
or ( n230502 , n230499 , n230501 );
not ( n230503 , n230502 );
or ( n230504 , n230498 , n230503 );
nand ( n230505 , n229940 , n224624 );
nand ( n230506 , n230504 , n230505 );
xor ( n230507 , n230497 , n230506 );
xor ( n230508 , n229680 , n230507 );
not ( n230509 , n221933 );
not ( n230510 , n226484 );
not ( n230511 , n40397 );
not ( n230512 , n230511 );
or ( n230513 , n230510 , n230512 );
not ( n230514 , n222121 );
nand ( n230515 , n230514 , n221938 );
nand ( n230516 , n230513 , n230515 );
not ( n230517 , n230516 );
or ( n230518 , n230509 , n230517 );
nand ( n230519 , n229878 , n215183 );
nand ( n230520 , n230518 , n230519 );
not ( n230521 , n226943 );
not ( n230522 , n229889 );
or ( n230523 , n230521 , n230522 );
not ( n230524 , n226292 );
not ( n230525 , n220599 );
or ( n230526 , n230524 , n230525 );
not ( n230527 , n221330 );
nand ( n230528 , n230527 , n229887 );
nand ( n230529 , n230526 , n230528 );
nand ( n230530 , n230529 , n226287 );
nand ( n230531 , n230523 , n230530 );
xor ( n230532 , n230520 , n230531 );
not ( n230533 , n223949 );
not ( n230534 , n226655 );
not ( n230535 , n220581 );
or ( n230536 , n230534 , n230535 );
nand ( n230537 , n207938 , n227927 );
nand ( n230538 , n230536 , n230537 );
not ( n230539 , n230538 );
or ( n230540 , n230533 , n230539 );
nand ( n230541 , n229900 , n227260 );
nand ( n230542 , n230540 , n230541 );
xor ( n230543 , n230532 , n230542 );
xor ( n230544 , n230508 , n230543 );
xor ( n230545 , n229680 , n230507 );
and ( n230546 , n230545 , n230543 );
and ( n230547 , n229680 , n230507 );
or ( n230548 , n230546 , n230547 );
not ( n230549 , n217969 );
not ( n230550 , n229696 );
or ( n230551 , n230549 , n230550 );
not ( n230552 , n213382 );
and ( n230553 , n831 , n39013 );
not ( n230554 , n831 );
and ( n230555 , n230554 , n209861 );
nor ( n230556 , n230553 , n230555 );
not ( n230557 , n230556 );
or ( n230558 , n230552 , n230557 );
nand ( n230559 , n209864 , n217715 );
nand ( n230560 , n230558 , n230559 );
nand ( n230561 , n230560 , n213912 );
nand ( n230562 , n230551 , n230561 );
xor ( n230563 , n230562 , n229625 );
xor ( n230564 , n230563 , n229663 );
xor ( n230565 , n230564 , n230232 );
xor ( n230566 , n230565 , n230290 );
xor ( n230567 , n230564 , n230232 );
and ( n230568 , n230567 , n230290 );
and ( n230569 , n230564 , n230232 );
or ( n230570 , n230568 , n230569 );
xor ( n230571 , n230260 , n229790 );
xor ( n230572 , n230571 , n229867 );
xor ( n230573 , n230260 , n229790 );
and ( n230574 , n230573 , n229867 );
and ( n230575 , n230260 , n229790 );
or ( n230576 , n230574 , n230575 );
xor ( n230577 , n230304 , n230314 );
and ( n230578 , n230577 , n230325 );
and ( n230579 , n230304 , n230314 );
or ( n230580 , n230578 , n230579 );
xor ( n230581 , n230361 , n230402 );
xor ( n230582 , n230581 , n229993 );
xor ( n230583 , n230361 , n230402 );
and ( n230584 , n230583 , n229993 );
and ( n230585 , n230361 , n230402 );
or ( n230586 , n230584 , n230585 );
xor ( n230587 , n230431 , n229873 );
xor ( n230588 , n230587 , n229911 );
xor ( n230589 , n230431 , n229873 );
and ( n230590 , n230589 , n229911 );
and ( n230591 , n230431 , n229873 );
or ( n230592 , n230590 , n230591 );
xor ( n230593 , n230040 , n230021 );
xor ( n230594 , n230593 , n230544 );
xor ( n230595 , n230040 , n230021 );
and ( n230596 , n230595 , n230544 );
and ( n230597 , n230040 , n230021 );
or ( n230598 , n230596 , n230597 );
xor ( n230599 , n230471 , n230046 );
xor ( n230600 , n230599 , n230572 );
xor ( n230601 , n230471 , n230046 );
and ( n230602 , n230601 , n230572 );
and ( n230603 , n230471 , n230046 );
or ( n230604 , n230602 , n230603 );
xor ( n230605 , n230566 , n230056 );
xor ( n230606 , n230605 , n230588 );
xor ( n230607 , n230566 , n230056 );
and ( n230608 , n230607 , n230588 );
and ( n230609 , n230566 , n230056 );
or ( n230610 , n230608 , n230609 );
xor ( n230611 , n230062 , n230582 );
xor ( n230612 , n230611 , n230594 );
xor ( n230613 , n230062 , n230582 );
and ( n230614 , n230613 , n230594 );
and ( n230615 , n230062 , n230582 );
or ( n230616 , n230614 , n230615 );
xor ( n230617 , n230068 , n230600 );
xor ( n230618 , n230617 , n230074 );
xor ( n230619 , n230068 , n230600 );
and ( n230620 , n230619 , n230074 );
and ( n230621 , n230068 , n230600 );
or ( n230622 , n230620 , n230621 );
xor ( n230623 , n230606 , n230612 );
xor ( n230624 , n230623 , n230080 );
xor ( n230625 , n230606 , n230612 );
and ( n230626 , n230625 , n230080 );
and ( n230627 , n230606 , n230612 );
or ( n230628 , n230626 , n230627 );
xor ( n230629 , n230086 , n230618 );
xor ( n230630 , n230629 , n230092 );
xor ( n230631 , n230086 , n230618 );
and ( n230632 , n230631 , n230092 );
and ( n230633 , n230086 , n230618 );
or ( n230634 , n230632 , n230633 );
xor ( n230635 , n230624 , n230630 );
xor ( n230636 , n230635 , n230098 );
xor ( n230637 , n230624 , n230630 );
and ( n230638 , n230637 , n230098 );
and ( n230639 , n230624 , n230630 );
or ( n230640 , n230638 , n230639 );
xor ( n230641 , n230376 , n230386 );
and ( n230642 , n230641 , n230399 );
and ( n230643 , n230376 , n230386 );
or ( n230644 , n230642 , n230643 );
xor ( n230645 , n230337 , n230348 );
and ( n230646 , n230645 , n230359 );
and ( n230647 , n230337 , n230348 );
or ( n230648 , n230646 , n230647 );
xor ( n230649 , n230416 , n230417 );
and ( n230650 , n230649 , n230428 );
and ( n230651 , n230416 , n230417 );
or ( n230652 , n230650 , n230651 );
xor ( n230653 , n230485 , n230496 );
and ( n230654 , n230653 , n230506 );
and ( n230655 , n230485 , n230496 );
or ( n230656 , n230654 , n230655 );
xor ( n230657 , n230520 , n230531 );
and ( n230658 , n230657 , n230542 );
and ( n230659 , n230520 , n230531 );
or ( n230660 , n230658 , n230659 );
xor ( n230661 , n230446 , n230456 );
and ( n230662 , n230661 , n230468 );
and ( n230663 , n230446 , n230456 );
or ( n230664 , n230662 , n230663 );
xor ( n230665 , n230562 , n229625 );
and ( n230666 , n230665 , n229663 );
and ( n230667 , n230562 , n229625 );
or ( n230668 , n230666 , n230667 );
not ( n230669 , n230173 );
not ( n230670 , n220479 );
or ( n230671 , n230669 , n230670 );
not ( n230672 , n218137 );
not ( n230673 , n230168 );
or ( n230674 , n230672 , n230673 );
nand ( n230675 , n217119 , n218815 );
nand ( n230676 , n230674 , n230675 );
nand ( n230677 , n230676 , n218455 );
nand ( n230678 , n230671 , n230677 );
not ( n230679 , n230189 );
not ( n230680 , n223620 );
or ( n230681 , n230679 , n230680 );
not ( n230682 , n217148 );
not ( n230683 , n219440 );
or ( n230684 , n230682 , n230683 );
nand ( n230685 , n219418 , n217147 );
nand ( n230686 , n230684 , n230685 );
nand ( n230687 , n219076 , n230686 );
nand ( n230688 , n230681 , n230687 );
xor ( n230689 , n230678 , n230688 );
not ( n230690 , n213126 );
not ( n230691 , n37670 );
not ( n230692 , n37556 );
nand ( n230693 , n230692 , n36320 , n37415 );
nand ( n230694 , n37416 , n37680 , n230693 );
not ( n230695 , n230694 );
or ( n230696 , n230691 , n230695 );
not ( n230697 , n37670 );
nand ( n230698 , n37416 , n37680 , n230693 , n230697 );
nand ( n230699 , n230696 , n230698 );
not ( n230700 , n230699 );
not ( n230701 , n230700 );
or ( n230702 , n230690 , n230701 );
not ( n230703 , n230699 );
not ( n230704 , n230703 );
nand ( n230705 , n230704 , n216076 );
nand ( n230706 , n230702 , n230705 );
not ( n230707 , n230706 );
buf ( n230708 , n230153 );
not ( n230709 , n230708 );
or ( n230710 , n230707 , n230709 );
not ( n230711 , n230703 );
not ( n230712 , n230147 );
not ( n230713 , n230712 );
or ( n230714 , n230711 , n230713 );
not ( n230715 , n230699 );
not ( n230716 , n230147 );
or ( n230717 , n230715 , n230716 );
nand ( n230718 , n230714 , n230717 );
nand ( n230719 , n230152 , n230718 );
not ( n230720 , n230719 );
not ( n230721 , n230720 );
buf ( n230722 , n230715 );
and ( n230723 , n213750 , n230722 );
not ( n230724 , n213750 );
buf ( n230725 , n230700 );
not ( n230726 , n230725 );
and ( n230727 , n230724 , n230726 );
nor ( n230728 , n230723 , n230727 );
or ( n230729 , n230721 , n230728 );
nand ( n230730 , n230710 , n230729 );
xor ( n230731 , n230689 , n230730 );
xor ( n230732 , n230678 , n230688 );
and ( n230733 , n230732 , n230730 );
and ( n230734 , n230678 , n230688 );
or ( n230735 , n230733 , n230734 );
not ( n230736 , n230199 );
not ( n230737 , n228326 );
or ( n230738 , n230736 , n230737 );
not ( n230739 , n224562 );
not ( n230740 , n41396 );
or ( n230741 , n230739 , n230740 );
not ( n230742 , n41396 );
nand ( n230743 , n230742 , n220146 );
nand ( n230744 , n230741 , n230743 );
nand ( n230745 , n230744 , n219777 );
nand ( n230746 , n230738 , n230745 );
not ( n230747 , n230209 );
not ( n230748 , n228342 );
or ( n230749 , n230747 , n230748 );
not ( n230750 , n225866 );
not ( n230751 , n230750 );
not ( n230752 , n220904 );
or ( n230753 , n230751 , n230752 );
nand ( n230754 , n220899 , n41563 );
nand ( n230755 , n230753 , n230754 );
nand ( n230756 , n230755 , n220635 );
nand ( n230757 , n230749 , n230756 );
xor ( n230758 , n230746 , n230757 );
not ( n230759 , n230302 );
not ( n230760 , n221623 );
or ( n230761 , n230759 , n230760 );
not ( n230762 , n227639 );
not ( n230763 , n221611 );
or ( n230764 , n230762 , n230763 );
nand ( n230765 , n223584 , n225769 );
nand ( n230766 , n230764 , n230765 );
nand ( n230767 , n230766 , n221387 );
nand ( n230768 , n230761 , n230767 );
xor ( n230769 , n230758 , n230768 );
xor ( n230770 , n230746 , n230757 );
and ( n230771 , n230770 , n230768 );
and ( n230772 , n230746 , n230757 );
or ( n230773 , n230771 , n230772 );
xor ( n230774 , n230580 , n230644 );
xor ( n230775 , n230774 , n230648 );
xor ( n230776 , n230580 , n230644 );
and ( n230777 , n230776 , n230648 );
and ( n230778 , n230580 , n230644 );
or ( n230779 , n230777 , n230778 );
not ( n230780 , n214717 );
not ( n230781 , n230245 );
or ( n230782 , n230780 , n230781 );
not ( n230783 , n218855 );
not ( n230784 , n226712 );
or ( n230785 , n230783 , n230784 );
nand ( n230786 , n39607 , n217944 );
nand ( n230787 , n230785 , n230786 );
nand ( n230788 , n230787 , n220985 );
nand ( n230789 , n230782 , n230788 );
not ( n230790 , n216562 );
not ( n230791 , n230256 );
or ( n230792 , n230790 , n230791 );
not ( n230793 , n215290 );
not ( n230794 , n39712 );
or ( n230795 , n230793 , n230794 );
or ( n230796 , n39712 , n215290 );
nand ( n230797 , n230795 , n230796 );
nand ( n230798 , n230797 , n220820 );
nand ( n230799 , n230792 , n230798 );
xor ( n230800 , n230789 , n230799 );
not ( n230801 , n213577 );
not ( n230802 , n230275 );
or ( n230803 , n230801 , n230802 );
not ( n230804 , n213735 );
not ( n230805 , n230025 );
or ( n230806 , n230804 , n230805 );
nand ( n230807 , n39286 , n213732 );
nand ( n230808 , n230806 , n230807 );
nand ( n230809 , n230808 , n216336 );
nand ( n230810 , n230803 , n230809 );
xor ( n230811 , n230800 , n230810 );
xor ( n230812 , n230789 , n230799 );
and ( n230813 , n230812 , n230810 );
and ( n230814 , n230789 , n230799 );
or ( n230815 , n230813 , n230814 );
not ( n230816 , n217023 );
not ( n230817 , n230284 );
or ( n230818 , n230816 , n230817 );
not ( n230819 , n225097 );
not ( n230820 , n230819 );
and ( n230821 , n218661 , n230820 );
not ( n230822 , n218661 );
and ( n230823 , n230822 , n39927 );
nor ( n230824 , n230821 , n230823 );
not ( n230825 , n230824 );
nand ( n230826 , n230825 , n219175 );
nand ( n230827 , n230818 , n230826 );
xor ( n230828 , n230827 , n230652 );
xor ( n230829 , n230828 , n230731 );
xor ( n230830 , n230827 , n230652 );
and ( n230831 , n230830 , n230731 );
and ( n230832 , n230827 , n230652 );
or ( n230833 , n230831 , n230832 );
not ( n230834 , n230346 );
not ( n230835 , n228707 );
not ( n230836 , n230835 );
or ( n230837 , n230834 , n230836 );
not ( n230838 , n216964 );
not ( n230839 , n228278 );
or ( n230840 , n230838 , n230839 );
nand ( n230841 , n227595 , n214678 );
nand ( n230842 , n230840 , n230841 );
nand ( n230843 , n227165 , n230842 );
nand ( n230844 , n230837 , n230843 );
not ( n230845 , n230357 );
not ( n230846 , n228858 );
or ( n230847 , n230845 , n230846 );
not ( n230848 , n214357 );
not ( n230849 , n228847 );
or ( n230850 , n230848 , n230849 );
not ( n230851 , n228846 );
nand ( n230852 , n230851 , n215131 );
nand ( n230853 , n230850 , n230852 );
nand ( n230854 , n228867 , n230853 );
nand ( n230855 , n230847 , n230854 );
xor ( n230856 , n230844 , n230855 );
not ( n230857 , n229771 );
and ( n230858 , n228726 , n229115 );
not ( n230859 , n228726 );
and ( n230860 , n230859 , n229114 );
nor ( n230861 , n230858 , n230860 );
nand ( n230862 , n230857 , n230861 );
or ( n230863 , n230862 , n230413 );
and ( n230864 , n229758 , n214134 );
not ( n230865 , n229758 );
and ( n230866 , n230865 , n213583 );
nor ( n230867 , n230864 , n230866 );
or ( n230868 , n230867 , n230861 );
nand ( n230869 , n230863 , n230868 );
xor ( n230870 , n230856 , n230869 );
xor ( n230871 , n230870 , n230769 );
not ( n230872 , n230384 );
not ( n230873 , n225851 );
or ( n230874 , n230872 , n230873 );
not ( n230875 , n219343 );
not ( n230876 , n224844 );
or ( n230877 , n230875 , n230876 );
nand ( n230878 , n224944 , n223269 );
nand ( n230879 , n230877 , n230878 );
nand ( n230880 , n230879 , n224449 );
nand ( n230881 , n230874 , n230880 );
not ( n230882 , n230397 );
not ( n230883 , n226272 );
or ( n230884 , n230882 , n230883 );
not ( n230885 , n225940 );
not ( n230886 , n216934 );
or ( n230887 , n230885 , n230886 );
nand ( n230888 , n225936 , n216940 );
nand ( n230889 , n230887 , n230888 );
nand ( n230890 , n230889 , n227710 );
nand ( n230891 , n230884 , n230890 );
xor ( n230892 , n230881 , n230891 );
not ( n230893 , n230335 );
not ( n230894 , n227849 );
or ( n230895 , n230893 , n230894 );
not ( n230896 , n215075 );
buf ( n230897 , n226888 );
not ( n230898 , n230897 );
or ( n230899 , n230896 , n230898 );
nand ( n230900 , n229823 , n215899 );
nand ( n230901 , n230899 , n230900 );
nand ( n230902 , n230901 , n227241 );
nand ( n230903 , n230895 , n230902 );
xor ( n230904 , n230892 , n230903 );
xor ( n230905 , n230871 , n230904 );
xor ( n230906 , n230870 , n230769 );
and ( n230907 , n230906 , n230904 );
and ( n230908 , n230870 , n230769 );
or ( n230909 , n230907 , n230908 );
not ( n230910 , n230312 );
not ( n230911 , n225902 );
or ( n230912 , n230910 , n230911 );
not ( n230913 , n214837 );
not ( n230914 , n228295 );
or ( n230915 , n230913 , n230914 );
nand ( n230916 , n222428 , n218670 );
nand ( n230917 , n230915 , n230916 );
nand ( n230918 , n230917 , n222157 );
nand ( n230919 , n230912 , n230918 );
not ( n230920 , n230323 );
not ( n230921 , n225380 );
or ( n230922 , n230920 , n230921 );
not ( n230923 , n215228 );
not ( n230924 , n224986 );
or ( n230925 , n230923 , n230924 );
nand ( n230926 , n223155 , n216555 );
nand ( n230927 , n230925 , n230926 );
nand ( n230928 , n222768 , n230927 );
nand ( n230929 , n230922 , n230928 );
xor ( n230930 , n230919 , n230929 );
not ( n230931 , n230374 );
not ( n230932 , n224086 );
or ( n230933 , n230931 , n230932 );
not ( n230934 , n221495 );
not ( n230935 , n224975 );
or ( n230936 , n230934 , n230935 );
nand ( n230937 , n223989 , n220022 );
nand ( n230938 , n230936 , n230937 );
nand ( n230939 , n224090 , n230938 );
nand ( n230940 , n230933 , n230939 );
xor ( n230941 , n230930 , n230940 );
xor ( n230942 , n230941 , n230656 );
xor ( n230943 , n230942 , n230660 );
xor ( n230944 , n230941 , n230656 );
and ( n230945 , n230944 , n230660 );
and ( n230946 , n230941 , n230656 );
or ( n230947 , n230945 , n230946 );
xor ( n230948 , n230264 , n230668 );
xor ( n230949 , n230948 , n230664 );
xor ( n230950 , n230264 , n230668 );
and ( n230951 , n230950 , n230664 );
and ( n230952 , n230264 , n230668 );
or ( n230953 , n230951 , n230952 );
not ( n230954 , n226287 );
not ( n230955 , n226292 );
not ( n230956 , n40258 );
or ( n230957 , n230955 , n230956 );
nand ( n230958 , n223383 , n229887 );
nand ( n230959 , n230957 , n230958 );
not ( n230960 , n230959 );
or ( n230961 , n230954 , n230960 );
nand ( n230962 , n230529 , n220414 );
nand ( n230963 , n230961 , n230962 );
not ( n230964 , n223949 );
not ( n230965 , n226655 );
buf ( n230966 , n220216 );
not ( n230967 , n230966 );
or ( n230968 , n230965 , n230967 );
nand ( n230969 , n226922 , n227927 );
nand ( n230970 , n230968 , n230969 );
not ( n230971 , n230970 );
or ( n230972 , n230964 , n230971 );
nand ( n230973 , n230538 , n227260 );
nand ( n230974 , n230972 , n230973 );
xor ( n230975 , n230963 , n230974 );
not ( n230976 , n229395 );
not ( n230977 , n230442 );
or ( n230978 , n230976 , n230977 );
not ( n230979 , n229387 );
not ( n230980 , n221687 );
or ( n230981 , n230979 , n230980 );
nand ( n230982 , n219522 , n227599 );
nand ( n230983 , n230981 , n230982 );
nand ( n230984 , n230983 , n228237 );
nand ( n230985 , n230978 , n230984 );
xor ( n230986 , n230975 , n230985 );
xor ( n230987 , n230236 , n230986 );
not ( n230988 , n230147 );
or ( n230989 , n230988 , n213750 );
nand ( n230990 , n230989 , n229761 );
not ( n230991 , n230722 );
nand ( n230992 , n230988 , n215999 );
and ( n230993 , n230990 , n230991 , n230992 );
not ( n230994 , n230993 );
not ( n230995 , n230161 );
not ( n230996 , n218525 );
or ( n230997 , n230995 , n230996 );
not ( n230998 , n218771 );
not ( n230999 , n220077 );
or ( n231000 , n230998 , n230999 );
nand ( n231001 , n218772 , n221559 );
nand ( n231002 , n231000 , n231001 );
nand ( n231003 , n231002 , n218231 );
nand ( n231004 , n230997 , n231003 );
not ( n231005 , n231004 );
not ( n231006 , n231005 );
or ( n231007 , n230994 , n231006 );
or ( n231008 , n231005 , n230993 );
nand ( n231009 , n231007 , n231008 );
not ( n231010 , n217614 );
not ( n231011 , n218268 );
or ( n231012 , n231010 , n231011 );
nand ( n231013 , n219594 , n218253 );
nand ( n231014 , n231012 , n231013 );
not ( n231015 , n231014 );
not ( n231016 , n220067 );
or ( n231017 , n231015 , n231016 );
not ( n231018 , n227130 );
nand ( n231019 , n230424 , n231018 );
nand ( n231020 , n231017 , n231019 );
xor ( n231021 , n231009 , n231020 );
not ( n231022 , n230494 );
or ( n231023 , n231022 , n217551 );
not ( n231024 , n225120 );
not ( n231025 , n39996 );
or ( n231026 , n231024 , n231025 );
nand ( n231027 , n225111 , n216989 );
nand ( n231028 , n231026 , n231027 );
not ( n231029 , n231028 );
or ( n231030 , n231029 , n217549 );
nand ( n231031 , n231023 , n231030 );
xor ( n231032 , n231021 , n231031 );
xor ( n231033 , n230987 , n231032 );
xor ( n231034 , n230236 , n230986 );
and ( n231035 , n231034 , n231032 );
and ( n231036 , n230236 , n230986 );
or ( n231037 , n231035 , n231036 );
not ( n231038 , n222185 );
not ( n231039 , n216166 );
not ( n231040 , n223330 );
or ( n231041 , n231039 , n231040 );
not ( n231042 , n40546 );
nand ( n231043 , n231042 , n226002 );
nand ( n231044 , n231041 , n231043 );
not ( n231045 , n231044 );
or ( n231046 , n231038 , n231045 );
nand ( n231047 , n230481 , n219731 );
nand ( n231048 , n231046 , n231047 );
not ( n231049 , n219314 );
not ( n231050 , n219687 );
not ( n231051 , n222509 );
or ( n231052 , n231050 , n231051 );
nand ( n231053 , n222513 , n221283 );
nand ( n231054 , n231052 , n231053 );
not ( n231055 , n231054 );
or ( n231056 , n231049 , n231055 );
nand ( n231057 , n230502 , n216204 );
nand ( n231058 , n231056 , n231057 );
xor ( n231059 , n231048 , n231058 );
not ( n231060 , n215183 );
not ( n231061 , n230516 );
or ( n231062 , n231060 , n231061 );
not ( n231063 , n226484 );
not ( n231064 , n221715 );
or ( n231065 , n231063 , n231064 );
nand ( n231066 , n221716 , n221938 );
nand ( n231067 , n231065 , n231066 );
nand ( n231068 , n231067 , n221933 );
nand ( n231069 , n231062 , n231068 );
xor ( n231070 , n231059 , n231069 );
xor ( n231071 , n231070 , n230294 );
not ( n231072 , n219368 );
not ( n231073 , n230452 );
or ( n231074 , n231072 , n231073 );
not ( n231075 , n229261 );
not ( n231076 , n219532 );
or ( n231077 , n231075 , n231076 );
nand ( n231078 , n220203 , n229262 );
nand ( n231079 , n231077 , n231078 );
nand ( n231080 , n231079 , n217388 );
nand ( n231081 , n231074 , n231080 );
not ( n231082 , n214086 );
not ( n231083 , n230464 );
or ( n231084 , n231082 , n231083 );
not ( n231085 , n217573 );
not ( n231086 , n227667 );
or ( n231087 , n231085 , n231086 );
not ( n231088 , n228657 );
nand ( n231089 , n231088 , n215388 );
nand ( n231090 , n231087 , n231089 );
nand ( n231091 , n231090 , n217571 );
nand ( n231092 , n231084 , n231091 );
xor ( n231093 , n231081 , n231092 );
not ( n231094 , n217969 );
not ( n231095 , n230560 );
or ( n231096 , n231094 , n231095 );
not ( n231097 , n209962 );
and ( n231098 , n213382 , n231097 );
not ( n231099 , n213382 );
not ( n231100 , n831 );
not ( n231101 , n39465 );
or ( n231102 , n231100 , n231101 );
nand ( n231103 , n231102 , n209960 );
buf ( n231104 , n231103 );
and ( n231105 , n231099 , n231104 );
nor ( n231106 , n231098 , n231105 );
or ( n231107 , n231106 , n213171 );
nand ( n231108 , n231096 , n231107 );
xor ( n231109 , n231093 , n231108 );
xor ( n231110 , n231071 , n231109 );
xor ( n231111 , n231070 , n230294 );
and ( n231112 , n231111 , n231109 );
and ( n231113 , n231070 , n230294 );
or ( n231114 , n231112 , n231113 );
xor ( n231115 , n230181 , n230217 );
not ( n231116 , n213874 );
not ( n231117 , n230225 );
or ( n231118 , n231116 , n231117 );
not ( n231119 , n216262 );
not ( n231120 , n209708 );
or ( n231121 , n231119 , n231120 );
nand ( n231122 , n209707 , n220300 );
nand ( n231123 , n231121 , n231122 );
nand ( n231124 , n231123 , n217142 );
nand ( n231125 , n231118 , n231124 );
xor ( n231126 , n231115 , n231125 );
xor ( n231127 , n231126 , n230811 );
xor ( n231128 , n231127 , n230775 );
xor ( n231129 , n231126 , n230811 );
and ( n231130 , n231129 , n230775 );
and ( n231131 , n231126 , n230811 );
or ( n231132 , n231130 , n231131 );
xor ( n231133 , n230365 , n230905 );
xor ( n231134 , n231133 , n230829 );
xor ( n231135 , n230365 , n230905 );
and ( n231136 , n231135 , n230829 );
and ( n231137 , n230365 , n230905 );
or ( n231138 , n231136 , n231137 );
xor ( n231139 , n230919 , n230929 );
and ( n231140 , n231139 , n230940 );
and ( n231141 , n230919 , n230929 );
or ( n231142 , n231140 , n231141 );
xor ( n231143 , n230406 , n230943 );
xor ( n231144 , n231143 , n230548 );
xor ( n231145 , n230406 , n230943 );
and ( n231146 , n231145 , n230548 );
and ( n231147 , n230406 , n230943 );
or ( n231148 , n231146 , n231147 );
xor ( n231149 , n230475 , n230435 );
xor ( n231150 , n231149 , n231033 );
xor ( n231151 , n230475 , n230435 );
and ( n231152 , n231151 , n231033 );
and ( n231153 , n230475 , n230435 );
or ( n231154 , n231152 , n231153 );
xor ( n231155 , n230949 , n230570 );
xor ( n231156 , n231155 , n230576 );
xor ( n231157 , n230949 , n230570 );
and ( n231158 , n231157 , n230576 );
and ( n231159 , n230949 , n230570 );
or ( n231160 , n231158 , n231159 );
xor ( n231161 , n231128 , n231110 );
xor ( n231162 , n231161 , n230586 );
xor ( n231163 , n231128 , n231110 );
and ( n231164 , n231163 , n230586 );
and ( n231165 , n231128 , n231110 );
or ( n231166 , n231164 , n231165 );
xor ( n231167 , n231134 , n230592 );
xor ( n231168 , n231167 , n231150 );
xor ( n231169 , n231134 , n230592 );
and ( n231170 , n231169 , n231150 );
and ( n231171 , n231134 , n230592 );
or ( n231172 , n231170 , n231171 );
xor ( n231173 , n230598 , n231144 );
xor ( n231174 , n231173 , n231156 );
xor ( n231175 , n230598 , n231144 );
and ( n231176 , n231175 , n231156 );
and ( n231177 , n230598 , n231144 );
or ( n231178 , n231176 , n231177 );
xor ( n231179 , n230604 , n231162 );
xor ( n231180 , n231179 , n230610 );
xor ( n231181 , n230604 , n231162 );
and ( n231182 , n231181 , n230610 );
and ( n231183 , n230604 , n231162 );
or ( n231184 , n231182 , n231183 );
xor ( n231185 , n231168 , n230616 );
xor ( n231186 , n231185 , n231174 );
xor ( n231187 , n231168 , n230616 );
and ( n231188 , n231187 , n231174 );
and ( n231189 , n231168 , n230616 );
or ( n231190 , n231188 , n231189 );
xor ( n231191 , n230622 , n231180 );
xor ( n231192 , n231191 , n230628 );
xor ( n231193 , n230622 , n231180 );
and ( n231194 , n231193 , n230628 );
and ( n231195 , n230622 , n231180 );
or ( n231196 , n231194 , n231195 );
xor ( n231197 , n231186 , n231192 );
xor ( n231198 , n231197 , n230634 );
xor ( n231199 , n231186 , n231192 );
and ( n231200 , n231199 , n230634 );
and ( n231201 , n231186 , n231192 );
or ( n231202 , n231200 , n231201 );
xor ( n231203 , n230881 , n230891 );
and ( n231204 , n231203 , n230903 );
and ( n231205 , n230881 , n230891 );
or ( n231206 , n231204 , n231205 );
xor ( n231207 , n230844 , n230855 );
and ( n231208 , n231207 , n230869 );
and ( n231209 , n230844 , n230855 );
or ( n231210 , n231208 , n231209 );
xor ( n231211 , n231009 , n231020 );
and ( n231212 , n231211 , n231031 );
and ( n231213 , n231009 , n231020 );
or ( n231214 , n231212 , n231213 );
xor ( n231215 , n231048 , n231058 );
and ( n231216 , n231215 , n231069 );
and ( n231217 , n231048 , n231058 );
or ( n231218 , n231216 , n231217 );
xor ( n231219 , n230963 , n230974 );
and ( n231220 , n231219 , n230985 );
and ( n231221 , n230963 , n230974 );
or ( n231222 , n231220 , n231221 );
xor ( n231223 , n231081 , n231092 );
and ( n231224 , n231223 , n231108 );
and ( n231225 , n231081 , n231092 );
or ( n231226 , n231224 , n231225 );
xor ( n231227 , n230181 , n230217 );
and ( n231228 , n231227 , n231125 );
and ( n231229 , n230181 , n230217 );
or ( n231230 , n231228 , n231229 );
buf ( n231231 , n230699 );
buf ( n231232 , n231231 );
and ( n231233 , n231232 , n215999 );
not ( n231234 , n230676 );
not ( n231235 , n220480 );
or ( n231236 , n231234 , n231235 );
not ( n231237 , n41071 );
not ( n231238 , n218814 );
or ( n231239 , n231237 , n231238 );
not ( n231240 , n219201 );
nand ( n231241 , n231240 , n220859 );
nand ( n231242 , n231239 , n231241 );
nand ( n231243 , n218843 , n231242 );
nand ( n231244 , n231236 , n231243 );
xor ( n231245 , n231233 , n231244 );
not ( n231246 , n230686 );
not ( n231247 , n219792 );
or ( n231248 , n231246 , n231247 );
not ( n231249 , n223549 );
not ( n231250 , n219423 );
or ( n231251 , n231249 , n231250 );
nand ( n231252 , n220180 , n230171 );
nand ( n231253 , n231251 , n231252 );
not ( n231254 , n231253 );
or ( n231255 , n231254 , n229612 );
nand ( n231256 , n231248 , n231255 );
xor ( n231257 , n231245 , n231256 );
xor ( n231258 , n231233 , n231244 );
and ( n231259 , n231258 , n231256 );
and ( n231260 , n231233 , n231244 );
or ( n231261 , n231259 , n231260 );
not ( n231262 , n230706 );
not ( n231263 , n230719 );
not ( n231264 , n231263 );
or ( n231265 , n231262 , n231264 );
not ( n231266 , n230700 );
not ( n231267 , n213347 );
or ( n231268 , n231266 , n231267 );
not ( n231269 , n230703 );
nand ( n231270 , n231269 , n222031 );
nand ( n231271 , n231268 , n231270 );
nand ( n231272 , n231271 , n230153 );
nand ( n231273 , n231265 , n231272 );
not ( n231274 , n230744 );
not ( n231275 , n220163 );
or ( n231276 , n231274 , n231275 );
and ( n231277 , n216311 , n224563 );
not ( n231278 , n216311 );
and ( n231279 , n231278 , n222413 );
or ( n231280 , n231277 , n231279 );
nand ( n231281 , n231280 , n219779 );
nand ( n231282 , n231276 , n231281 );
xor ( n231283 , n231273 , n231282 );
not ( n231284 , n230755 );
or ( n231285 , n228639 , n231284 );
and ( n231286 , n220901 , n215796 );
and ( n231287 , n220900 , n216261 );
nor ( n231288 , n231286 , n231287 );
or ( n231289 , n231288 , n220928 );
nand ( n231290 , n231285 , n231289 );
xor ( n231291 , n231283 , n231290 );
xor ( n231292 , n231273 , n231282 );
and ( n231293 , n231292 , n231290 );
and ( n231294 , n231273 , n231282 );
or ( n231295 , n231293 , n231294 );
xor ( n231296 , n230773 , n231142 );
xor ( n231297 , n231296 , n231206 );
xor ( n231298 , n230773 , n231142 );
and ( n231299 , n231298 , n231206 );
and ( n231300 , n230773 , n231142 );
or ( n231301 , n231299 , n231300 );
not ( n231302 , n220985 );
not ( n231303 , n215113 );
not ( n231304 , n228184 );
or ( n231305 , n231303 , n231304 );
nand ( n231306 , n39089 , n217944 );
nand ( n231307 , n231305 , n231306 );
not ( n231308 , n231307 );
or ( n231309 , n231302 , n231308 );
nand ( n231310 , n230787 , n214717 );
nand ( n231311 , n231309 , n231310 );
xor ( n231312 , n231210 , n231311 );
not ( n231313 , n217969 );
not ( n231314 , n231106 );
not ( n231315 , n231314 );
or ( n231316 , n231313 , n231315 );
nand ( n231317 , n213382 , n211314 );
nand ( n231318 , n231316 , n231317 );
xor ( n231319 , n231312 , n231318 );
xor ( n231320 , n231210 , n231311 );
and ( n231321 , n231320 , n231318 );
and ( n231322 , n231210 , n231311 );
or ( n231323 , n231321 , n231322 );
not ( n231324 , n216562 );
not ( n231325 , n230797 );
or ( n231326 , n231324 , n231325 );
not ( n231327 , n216810 );
not ( n231328 , n228216 );
or ( n231329 , n231327 , n231328 );
nand ( n231330 , n39746 , n215289 );
nand ( n231331 , n231329 , n231330 );
nand ( n231332 , n231331 , n214694 );
nand ( n231333 , n231326 , n231332 );
not ( n231334 , n213577 );
not ( n231335 , n230808 );
or ( n231336 , n231334 , n231335 );
not ( n231337 , n213735 );
not ( n231338 , n229214 );
or ( n231339 , n231337 , n231338 );
nand ( n231340 , n230222 , n213732 );
nand ( n231341 , n231339 , n231340 );
nand ( n231342 , n231341 , n216336 );
nand ( n231343 , n231336 , n231342 );
xor ( n231344 , n231333 , n231343 );
not ( n231345 , n219577 );
not ( n231346 , n225357 );
or ( n231347 , n231345 , n231346 );
nand ( n231348 , n39812 , n215971 );
nand ( n231349 , n231347 , n231348 );
not ( n231350 , n231349 );
not ( n231351 , n219175 );
or ( n231352 , n231350 , n231351 );
or ( n231353 , n217367 , n230824 );
nand ( n231354 , n231352 , n231353 );
xor ( n231355 , n231344 , n231354 );
xor ( n231356 , n231333 , n231343 );
and ( n231357 , n231356 , n231354 );
and ( n231358 , n231333 , n231343 );
or ( n231359 , n231357 , n231358 );
xor ( n231360 , n231291 , n231257 );
not ( n231361 , n230766 );
not ( n231362 , n221625 );
or ( n231363 , n231361 , n231362 );
not ( n231364 , n221608 );
not ( n231365 , n226224 );
and ( n231366 , n231364 , n231365 );
not ( n231367 , n41701 );
and ( n231368 , n223584 , n231367 );
nor ( n231369 , n231366 , n231368 );
not ( n231370 , n231369 );
nand ( n231371 , n231370 , n223587 );
nand ( n231372 , n231363 , n231371 );
not ( n231373 , n222453 );
not ( n231374 , n230917 );
or ( n231375 , n231373 , n231374 );
not ( n231376 , n219689 );
not ( n231377 , n222458 );
or ( n231378 , n231376 , n231377 );
nand ( n231379 , n222892 , n225489 );
nand ( n231380 , n231378 , n231379 );
nand ( n231381 , n231380 , n222158 );
nand ( n231382 , n231375 , n231381 );
xor ( n231383 , n231372 , n231382 );
not ( n231384 , n223197 );
not ( n231385 , n230927 );
or ( n231386 , n231384 , n231385 );
not ( n231387 , n224496 );
not ( n231388 , n223202 );
or ( n231389 , n231387 , n231388 );
or ( n231390 , n223182 , n224496 );
nand ( n231391 , n231389 , n231390 );
nand ( n231392 , n231391 , n222769 );
nand ( n231393 , n231386 , n231392 );
xor ( n231394 , n231383 , n231393 );
xor ( n231395 , n231360 , n231394 );
xor ( n231396 , n231291 , n231257 );
and ( n231397 , n231396 , n231394 );
and ( n231398 , n231291 , n231257 );
or ( n231399 , n231397 , n231398 );
not ( n231400 , n230901 );
not ( n231401 , n227849 );
or ( n231402 , n231400 , n231401 );
not ( n231403 , n218514 );
not ( n231404 , n229820 );
or ( n231405 , n231403 , n231404 );
nand ( n231406 , n227245 , n216170 );
nand ( n231407 , n231405 , n231406 );
nand ( n231408 , n226218 , n231407 );
nand ( n231409 , n231402 , n231408 );
not ( n231410 , n230842 );
or ( n231411 , n228270 , n231410 );
not ( n231412 , n227595 );
and ( n231413 , n216208 , n231412 );
not ( n231414 , n216208 );
and ( n231415 , n231414 , n227595 );
nor ( n231416 , n231413 , n231415 );
or ( n231417 , n228273 , n231416 );
nand ( n231418 , n231411 , n231417 );
xor ( n231419 , n231409 , n231418 );
not ( n231420 , n230853 );
buf ( n231421 , n228858 );
not ( n231422 , n231421 );
or ( n231423 , n231420 , n231422 );
nand ( n231424 , n228847 , n214537 );
not ( n231425 , n231424 );
nand ( n231426 , n228726 , n214899 );
not ( n231427 , n231426 );
or ( n231428 , n231425 , n231427 );
nand ( n231429 , n231428 , n229738 );
nand ( n231430 , n231423 , n231429 );
xor ( n231431 , n231419 , n231430 );
not ( n231432 , n230938 );
not ( n231433 , n224086 );
or ( n231434 , n231432 , n231433 );
not ( n231435 , n216293 );
not ( n231436 , n225844 );
or ( n231437 , n231435 , n231436 );
nand ( n231438 , n224974 , n223658 );
nand ( n231439 , n231437 , n231438 );
nand ( n231440 , n224090 , n231439 );
nand ( n231441 , n231434 , n231440 );
not ( n231442 , n224938 );
not ( n231443 , n230879 );
or ( n231444 , n231442 , n231443 );
not ( n231445 , n222821 );
not ( n231446 , n229795 );
or ( n231447 , n231445 , n231446 );
nand ( n231448 , n224929 , n218980 );
nand ( n231449 , n231447 , n231448 );
nand ( n231450 , n226745 , n231449 );
nand ( n231451 , n231444 , n231450 );
xor ( n231452 , n231441 , n231451 );
not ( n231453 , n230390 );
not ( n231454 , n230889 );
or ( n231455 , n231453 , n231454 );
not ( n231456 , n228775 );
not ( n231457 , n219102 );
not ( n231458 , n229807 );
or ( n231459 , n231457 , n231458 );
nand ( n231460 , n225952 , n216139 );
nand ( n231461 , n231459 , n231460 );
not ( n231462 , n231461 );
or ( n231463 , n231456 , n231462 );
nand ( n231464 , n231455 , n231463 );
xor ( n231465 , n231452 , n231464 );
xor ( n231466 , n231431 , n231465 );
xor ( n231467 , n231466 , n231214 );
xor ( n231468 , n231431 , n231465 );
and ( n231469 , n231468 , n231214 );
and ( n231470 , n231431 , n231465 );
or ( n231471 , n231469 , n231470 );
xor ( n231472 , n231218 , n231222 );
not ( n231473 , n230862 );
not ( n231474 , n231473 );
or ( n231475 , n231474 , n230867 );
buf ( n231476 , n230861 );
not ( n231477 , n229761 );
and ( n231478 , n214956 , n231477 );
not ( n231479 , n214956 );
buf ( n231480 , n229761 );
and ( n231481 , n231479 , n231480 );
nor ( n231482 , n231478 , n231481 );
or ( n231483 , n231476 , n231482 );
nand ( n231484 , n231475 , n231483 );
not ( n231485 , n218533 );
not ( n231486 , n40724 );
not ( n231487 , n218256 );
or ( n231488 , n231486 , n231487 );
or ( n231489 , n218256 , n40724 );
nand ( n231490 , n231488 , n231489 );
not ( n231491 , n231490 );
or ( n231492 , n231485 , n231491 );
nand ( n231493 , n219836 , n231002 );
nand ( n231494 , n231492 , n231493 );
xor ( n231495 , n231484 , n231494 );
not ( n231496 , n220067 );
not ( n231497 , n217616 );
not ( n231498 , n226486 );
or ( n231499 , n231497 , n231498 );
buf ( n231500 , n217616 );
not ( n231501 , n231500 );
nand ( n231502 , n224642 , n231501 );
nand ( n231503 , n231499 , n231502 );
not ( n231504 , n231503 );
or ( n231505 , n231496 , n231504 );
nand ( n231506 , n231014 , n231018 );
nand ( n231507 , n231505 , n231506 );
xor ( n231508 , n231495 , n231507 );
xor ( n231509 , n231472 , n231508 );
xor ( n231510 , n231218 , n231222 );
and ( n231511 , n231510 , n231508 );
and ( n231512 , n231218 , n231222 );
or ( n231513 , n231511 , n231512 );
not ( n231514 , n228237 );
not ( n231515 , n216422 );
not ( n231516 , n221356 );
or ( n231517 , n231515 , n231516 );
nand ( n231518 , n207936 , n227599 );
nand ( n231519 , n231517 , n231518 );
not ( n231520 , n231519 );
or ( n231521 , n231514 , n231520 );
nand ( n231522 , n230983 , n229395 );
nand ( n231523 , n231521 , n231522 );
not ( n231524 , n219368 );
not ( n231525 , n231079 );
or ( n231526 , n231524 , n231525 );
not ( n231527 , n229261 );
not ( n231528 , n40560 );
or ( n231529 , n231527 , n231528 );
nand ( n231530 , n219226 , n229262 );
nand ( n231531 , n231529 , n231530 );
nand ( n231532 , n231531 , n229964 );
nand ( n231533 , n231526 , n231532 );
xor ( n231534 , n231523 , n231533 );
not ( n231535 , n219353 );
not ( n231536 , n215955 );
not ( n231537 , n39877 );
or ( n231538 , n231536 , n231537 );
nand ( n231539 , n225344 , n216989 );
nand ( n231540 , n231538 , n231539 );
not ( n231541 , n231540 );
or ( n231542 , n231535 , n231541 );
nand ( n231543 , n231028 , n217552 );
nand ( n231544 , n231542 , n231543 );
xor ( n231545 , n231534 , n231544 );
xor ( n231546 , n231226 , n231545 );
xor ( n231547 , n231546 , n230815 );
xor ( n231548 , n231226 , n231545 );
and ( n231549 , n231548 , n230815 );
and ( n231550 , n231226 , n231545 );
or ( n231551 , n231549 , n231550 );
xor ( n231552 , n230779 , n231230 );
not ( n231553 , n215183 );
not ( n231554 , n231067 );
or ( n231555 , n231553 , n231554 );
not ( n231556 , n218994 );
not ( n231557 , n223751 );
or ( n231558 , n231556 , n231557 );
nand ( n231559 , n222100 , n226484 );
nand ( n231560 , n231558 , n231559 );
nand ( n231561 , n231560 , n221933 );
nand ( n231562 , n231555 , n231561 );
not ( n231563 , n226943 );
not ( n231564 , n230959 );
or ( n231565 , n231563 , n231564 );
and ( n231566 , n221194 , n227912 );
not ( n231567 , n221194 );
and ( n231568 , n231567 , n229887 );
or ( n231569 , n231566 , n231568 );
nand ( n231570 , n231569 , n226287 );
nand ( n231571 , n231565 , n231570 );
xor ( n231572 , n231562 , n231571 );
not ( n231573 , n227260 );
not ( n231574 , n230970 );
or ( n231575 , n231573 , n231574 );
not ( n231576 , n226655 );
not ( n231577 , n223786 );
or ( n231578 , n231576 , n231577 );
nand ( n231579 , n40410 , n227927 );
nand ( n231580 , n231578 , n231579 );
nand ( n231581 , n231580 , n223949 );
nand ( n231582 , n231575 , n231581 );
xor ( n231583 , n231572 , n231582 );
xor ( n231584 , n231552 , n231583 );
xor ( n231585 , n230779 , n231230 );
and ( n231586 , n231585 , n231583 );
and ( n231587 , n230779 , n231230 );
or ( n231588 , n231586 , n231587 );
and ( n231589 , n231004 , n230993 );
not ( n231590 , n219731 );
not ( n231591 , n231044 );
or ( n231592 , n231590 , n231591 );
not ( n231593 , n219033 );
not ( n231594 , n223761 );
or ( n231595 , n231593 , n231594 );
nand ( n231596 , n40045 , n220538 );
nand ( n231597 , n231595 , n231596 );
nand ( n231598 , n231597 , n222185 );
nand ( n231599 , n231592 , n231598 );
xor ( n231600 , n231589 , n231599 );
not ( n231601 , n224624 );
not ( n231602 , n231054 );
or ( n231603 , n231601 , n231602 );
not ( n231604 , n219687 );
not ( n231605 , n223721 );
or ( n231606 , n231604 , n231605 );
nand ( n231607 , n40485 , n221283 );
nand ( n231608 , n231606 , n231607 );
nand ( n231609 , n231608 , n219314 );
nand ( n231610 , n231603 , n231609 );
xor ( n231611 , n231600 , n231610 );
xor ( n231612 , n231611 , n230833 );
xor ( n231613 , n231612 , n231355 );
xor ( n231614 , n231611 , n230833 );
and ( n231615 , n231614 , n231355 );
and ( n231616 , n231611 , n230833 );
or ( n231617 , n231615 , n231616 );
not ( n231618 , n213874 );
not ( n231619 , n231123 );
or ( n231620 , n231618 , n231619 );
and ( n231621 , n220300 , n209863 );
not ( n231622 , n220300 );
not ( n231623 , n230556 );
and ( n231624 , n231622 , n231623 );
nor ( n231625 , n231621 , n231624 );
nand ( n231626 , n231625 , n217142 );
nand ( n231627 , n231620 , n231626 );
xor ( n231628 , n231627 , n230735 );
not ( n231629 , n215137 );
and ( n231630 , n39364 , n213960 );
not ( n231631 , n39364 );
and ( n231632 , n231631 , n217397 );
or ( n231633 , n231630 , n231632 );
not ( n231634 , n231633 );
or ( n231635 , n231629 , n231634 );
nand ( n231636 , n231090 , n218467 );
nand ( n231637 , n231635 , n231636 );
xor ( n231638 , n231628 , n231637 );
xor ( n231639 , n231297 , n231638 );
xor ( n231640 , n231639 , n230909 );
xor ( n231641 , n231297 , n231638 );
and ( n231642 , n231641 , n230909 );
and ( n231643 , n231297 , n231638 );
or ( n231644 , n231642 , n231643 );
xor ( n231645 , n231372 , n231382 );
and ( n231646 , n231645 , n231393 );
and ( n231647 , n231372 , n231382 );
or ( n231648 , n231646 , n231647 );
xor ( n231649 , n231319 , n231467 );
xor ( n231650 , n231649 , n231395 );
xor ( n231651 , n231319 , n231467 );
and ( n231652 , n231651 , n231395 );
and ( n231653 , n231319 , n231467 );
or ( n231654 , n231652 , n231653 );
xor ( n231655 , n230947 , n231509 );
xor ( n231656 , n231655 , n231037 );
xor ( n231657 , n230947 , n231509 );
and ( n231658 , n231657 , n231037 );
and ( n231659 , n230947 , n231509 );
or ( n231660 , n231658 , n231659 );
xor ( n231661 , n230953 , n231547 );
xor ( n231662 , n231661 , n231114 );
xor ( n231663 , n230953 , n231547 );
and ( n231664 , n231663 , n231114 );
and ( n231665 , n230953 , n231547 );
or ( n231666 , n231664 , n231665 );
xor ( n231667 , n231132 , n231584 );
xor ( n231668 , n231667 , n231138 );
xor ( n231669 , n231132 , n231584 );
and ( n231670 , n231669 , n231138 );
and ( n231671 , n231132 , n231584 );
or ( n231672 , n231670 , n231671 );
xor ( n231673 , n231613 , n231640 );
xor ( n231674 , n231673 , n231650 );
xor ( n231675 , n231613 , n231640 );
and ( n231676 , n231675 , n231650 );
and ( n231677 , n231613 , n231640 );
or ( n231678 , n231676 , n231677 );
xor ( n231679 , n231148 , n231154 );
xor ( n231680 , n231679 , n231160 );
xor ( n231681 , n231148 , n231154 );
and ( n231682 , n231681 , n231160 );
and ( n231683 , n231148 , n231154 );
or ( n231684 , n231682 , n231683 );
xor ( n231685 , n231656 , n231668 );
xor ( n231686 , n231685 , n231662 );
xor ( n231687 , n231656 , n231668 );
and ( n231688 , n231687 , n231662 );
and ( n231689 , n231656 , n231668 );
or ( n231690 , n231688 , n231689 );
xor ( n231691 , n231166 , n231674 );
xor ( n231692 , n231691 , n231172 );
xor ( n231693 , n231166 , n231674 );
and ( n231694 , n231693 , n231172 );
and ( n231695 , n231166 , n231674 );
or ( n231696 , n231694 , n231695 );
xor ( n231697 , n231680 , n231178 );
xor ( n231698 , n231697 , n231686 );
xor ( n231699 , n231680 , n231178 );
and ( n231700 , n231699 , n231686 );
and ( n231701 , n231680 , n231178 );
or ( n231702 , n231700 , n231701 );
xor ( n231703 , n231692 , n231184 );
xor ( n231704 , n231703 , n231190 );
xor ( n231705 , n231692 , n231184 );
and ( n231706 , n231705 , n231190 );
and ( n231707 , n231692 , n231184 );
or ( n231708 , n231706 , n231707 );
xor ( n231709 , n231441 , n231451 );
and ( n231710 , n231709 , n231464 );
and ( n231711 , n231441 , n231451 );
or ( n231712 , n231710 , n231711 );
xor ( n231713 , n231698 , n231704 );
xor ( n231714 , n231713 , n231196 );
xor ( n231715 , n231698 , n231704 );
and ( n231716 , n231715 , n231196 );
and ( n231717 , n231698 , n231704 );
or ( n231718 , n231716 , n231717 );
xor ( n231719 , n231409 , n231418 );
and ( n231720 , n231719 , n231430 );
and ( n231721 , n231409 , n231418 );
or ( n231722 , n231720 , n231721 );
xor ( n231723 , n231484 , n231494 );
and ( n231724 , n231723 , n231507 );
and ( n231725 , n231484 , n231494 );
or ( n231726 , n231724 , n231725 );
xor ( n231727 , n231589 , n231599 );
and ( n231728 , n231727 , n231610 );
and ( n231729 , n231589 , n231599 );
or ( n231730 , n231728 , n231729 );
xor ( n231731 , n231562 , n231571 );
and ( n231732 , n231731 , n231582 );
and ( n231733 , n231562 , n231571 );
or ( n231734 , n231732 , n231733 );
xor ( n231735 , n231523 , n231533 );
and ( n231736 , n231735 , n231544 );
and ( n231737 , n231523 , n231533 );
or ( n231738 , n231736 , n231737 );
xor ( n231739 , n231627 , n230735 );
and ( n231740 , n231739 , n231637 );
and ( n231741 , n231627 , n230735 );
or ( n231742 , n231740 , n231741 );
not ( n231743 , n231242 );
not ( n231744 , n220853 );
or ( n231745 , n231743 , n231744 );
not ( n231746 , n220859 );
not ( n231747 , n220823 );
or ( n231748 , n231746 , n231747 );
nand ( n231749 , n41165 , n218876 );
nand ( n231750 , n231748 , n231749 );
nand ( n231751 , n231750 , n218455 );
nand ( n231752 , n231745 , n231751 );
buf ( n231753 , n230725 );
not ( n231754 , n231753 );
and ( n231755 , n231754 , n218224 );
xor ( n231756 , n231752 , n231755 );
not ( n231757 , n231253 );
not ( n231758 , n221576 );
or ( n231759 , n231757 , n231758 );
not ( n231760 , n219440 );
buf ( n231761 , n217119 );
not ( n231762 , n231761 );
not ( n231763 , n231762 );
or ( n231764 , n231760 , n231763 );
nand ( n231765 , n231761 , n219796 );
nand ( n231766 , n231764 , n231765 );
nand ( n231767 , n219076 , n231766 );
nand ( n231768 , n231759 , n231767 );
xor ( n231769 , n231756 , n231768 );
xor ( n231770 , n231752 , n231755 );
and ( n231771 , n231770 , n231768 );
and ( n231772 , n231752 , n231755 );
or ( n231773 , n231771 , n231772 );
not ( n231774 , n217142 );
not ( n231775 , n214818 );
not ( n231776 , n209961 );
not ( n231777 , n231776 );
or ( n231778 , n231775 , n231777 );
not ( n231779 , n209961 );
or ( n231780 , n231779 , n214818 );
nand ( n231781 , n231778 , n231780 );
not ( n231782 , n231781 );
or ( n231783 , n231774 , n231782 );
nand ( n231784 , n213874 , n231625 );
nand ( n231785 , n231783 , n231784 );
not ( n231786 , n218467 );
not ( n231787 , n231633 );
or ( n231788 , n231786 , n231787 );
not ( n231789 , n213261 );
not ( n231790 , n230025 );
or ( n231791 , n231789 , n231790 );
nand ( n231792 , n39286 , n217397 );
nand ( n231793 , n231791 , n231792 );
nand ( n231794 , n231793 , n213204 );
nand ( n231795 , n231788 , n231794 );
xor ( n231796 , n231785 , n231795 );
xor ( n231797 , n231796 , n231261 );
xor ( n231798 , n231785 , n231795 );
and ( n231799 , n231798 , n231261 );
and ( n231800 , n231785 , n231795 );
or ( n231801 , n231799 , n231800 );
xor ( n231802 , n231295 , n231648 );
xor ( n231803 , n231802 , n231712 );
xor ( n231804 , n231295 , n231648 );
and ( n231805 , n231804 , n231712 );
and ( n231806 , n231295 , n231648 );
or ( n231807 , n231805 , n231806 );
not ( n231808 , n228676 );
not ( n231809 , n231808 );
not ( n231810 , n231307 );
or ( n231811 , n231809 , n231810 );
not ( n231812 , n215113 );
not ( n231813 , n38530 );
or ( n231814 , n231812 , n231813 );
not ( n231815 , n215113 );
nand ( n231816 , n231815 , n38531 );
nand ( n231817 , n231814 , n231816 );
nand ( n231818 , n231817 , n220985 );
nand ( n231819 , n231811 , n231818 );
xor ( n231820 , n231819 , n231722 );
not ( n231821 , n220820 );
not ( n231822 , n216810 );
not ( n231823 , n226712 );
or ( n231824 , n231822 , n231823 );
nand ( n231825 , n39607 , n221307 );
nand ( n231826 , n231824 , n231825 );
not ( n231827 , n231826 );
or ( n231828 , n231821 , n231827 );
buf ( n231829 , n231331 );
nand ( n231830 , n231829 , n216299 );
nand ( n231831 , n231828 , n231830 );
xor ( n231832 , n231820 , n231831 );
xor ( n231833 , n231819 , n231722 );
and ( n231834 , n231833 , n231831 );
and ( n231835 , n231819 , n231722 );
or ( n231836 , n231834 , n231835 );
not ( n231837 , n216336 );
not ( n231838 , n213735 );
not ( n231839 , n229691 );
or ( n231840 , n231838 , n231839 );
nand ( n231841 , n229694 , n213732 );
nand ( n231842 , n231840 , n231841 );
not ( n231843 , n231842 );
or ( n231844 , n231837 , n231843 );
nand ( n231845 , n231341 , n213577 );
nand ( n231846 , n231844 , n231845 );
not ( n231847 , n219175 );
not ( n231848 , n219577 );
not ( n231849 , n225792 );
or ( n231850 , n231848 , n231849 );
nand ( n231851 , n225795 , n218661 );
nand ( n231852 , n231850 , n231851 );
not ( n231853 , n231852 );
or ( n231854 , n231847 , n231853 );
nand ( n231855 , n231349 , n217023 );
nand ( n231856 , n231854 , n231855 );
xor ( n231857 , n231846 , n231856 );
not ( n231858 , n231271 );
not ( n231859 , n231263 );
or ( n231860 , n231858 , n231859 );
and ( n231861 , n213583 , n230700 );
not ( n231862 , n213583 );
and ( n231863 , n231862 , n231231 );
or ( n231864 , n231861 , n231863 );
nand ( n231865 , n231864 , n230153 );
nand ( n231866 , n231860 , n231865 );
and ( n231867 , n224881 , n221256 );
not ( n231868 , n224881 );
and ( n231869 , n231868 , n220150 );
or ( n231870 , n231867 , n231869 );
not ( n231871 , n231870 );
not ( n231872 , n220881 );
or ( n231873 , n231871 , n231872 );
nand ( n231874 , n231280 , n220163 );
nand ( n231875 , n231873 , n231874 );
xor ( n231876 , n231866 , n231875 );
or ( n231877 , n228639 , n231288 );
and ( n231878 , n223228 , n219582 );
and ( n231879 , n220900 , n216500 );
nor ( n231880 , n231878 , n231879 );
or ( n231881 , n231880 , n220928 );
nand ( n231882 , n231877 , n231881 );
xor ( n231883 , n231876 , n231882 );
xor ( n231884 , n231857 , n231883 );
xor ( n231885 , n231846 , n231856 );
and ( n231886 , n231885 , n231883 );
and ( n231887 , n231846 , n231856 );
or ( n231888 , n231886 , n231887 );
or ( n231889 , n221624 , n231369 );
and ( n231890 , n230750 , n221632 );
not ( n231891 , n230750 );
and ( n231892 , n231891 , n221608 );
nor ( n231893 , n231890 , n231892 );
or ( n231894 , n231893 , n223176 );
nand ( n231895 , n231889 , n231894 );
not ( n231896 , n222453 );
not ( n231897 , n231380 );
or ( n231898 , n231896 , n231897 );
not ( n231899 , n225768 );
not ( n231900 , n222458 );
or ( n231901 , n231899 , n231900 );
nand ( n231902 , n222462 , n225769 );
nand ( n231903 , n231901 , n231902 );
nand ( n231904 , n231903 , n222465 );
nand ( n231905 , n231898 , n231904 );
xor ( n231906 , n231895 , n231905 );
not ( n231907 , n223197 );
not ( n231908 , n231391 );
or ( n231909 , n231907 , n231908 );
not ( n231910 , n214837 );
not ( n231911 , n223186 );
or ( n231912 , n231910 , n231911 );
not ( n231913 , n214837 );
nand ( n231914 , n223202 , n231913 );
nand ( n231915 , n231912 , n231914 );
nand ( n231916 , n231915 , n222768 );
nand ( n231917 , n231909 , n231916 );
xor ( n231918 , n231906 , n231917 );
xor ( n231919 , n231769 , n231918 );
not ( n231920 , n216934 );
not ( n231921 , n229820 );
or ( n231922 , n231920 , n231921 );
nand ( n231923 , n227245 , n216940 );
nand ( n231924 , n231922 , n231923 );
not ( n231925 , n231924 );
not ( n231926 , n226218 );
or ( n231927 , n231925 , n231926 );
nand ( n231928 , n231407 , n226880 );
nand ( n231929 , n231927 , n231928 );
or ( n231930 , n228270 , n231416 );
xnor ( n231931 , n215075 , n227595 );
or ( n231932 , n228273 , n231931 );
nand ( n231933 , n231930 , n231932 );
xor ( n231934 , n231929 , n231933 );
not ( n231935 , n228858 );
nand ( n231936 , n231424 , n231426 );
not ( n231937 , n231936 );
or ( n231938 , n231935 , n231937 );
not ( n231939 , n219475 );
not ( n231940 , n228726 );
not ( n231941 , n231940 );
or ( n231942 , n231939 , n231941 );
not ( n231943 , n228847 );
nand ( n231944 , n231943 , n214678 );
nand ( n231945 , n231942 , n231944 );
nand ( n231946 , n231945 , n228867 );
nand ( n231947 , n231938 , n231946 );
xor ( n231948 , n231934 , n231947 );
xor ( n231949 , n231919 , n231948 );
xor ( n231950 , n231769 , n231918 );
and ( n231951 , n231950 , n231948 );
and ( n231952 , n231769 , n231918 );
or ( n231953 , n231951 , n231952 );
not ( n231954 , n231439 );
not ( n231955 , n224085 );
or ( n231956 , n231954 , n231955 );
not ( n231957 , n223811 );
not ( n231958 , n215228 );
not ( n231959 , n225844 );
or ( n231960 , n231958 , n231959 );
nand ( n231961 , n224068 , n216555 );
nand ( n231962 , n231960 , n231961 );
nand ( n231963 , n231957 , n231962 );
nand ( n231964 , n231956 , n231963 );
not ( n231965 , n231449 );
not ( n231966 , n224938 );
or ( n231967 , n231965 , n231966 );
not ( n231968 , n224448 );
not ( n231969 , n221495 );
not ( n231970 , n224943 );
or ( n231971 , n231969 , n231970 );
nand ( n231972 , n224929 , n220022 );
nand ( n231973 , n231971 , n231972 );
nand ( n231974 , n231968 , n231973 );
nand ( n231975 , n231967 , n231974 );
xor ( n231976 , n231964 , n231975 );
not ( n231977 , n231461 );
not ( n231978 , n226755 );
or ( n231979 , n231977 , n231978 );
not ( n231980 , n219343 );
not ( n231981 , n226276 );
or ( n231982 , n231980 , n231981 );
nand ( n231983 , n225952 , n219348 );
nand ( n231984 , n231982 , n231983 );
nand ( n231985 , n228775 , n231984 );
nand ( n231986 , n231979 , n231985 );
xor ( n231987 , n231976 , n231986 );
xor ( n231988 , n231987 , n231734 );
xor ( n231989 , n231988 , n231726 );
xor ( n231990 , n231987 , n231734 );
and ( n231991 , n231990 , n231726 );
and ( n231992 , n231987 , n231734 );
or ( n231993 , n231991 , n231992 );
buf ( n231994 , n230862 );
or ( n231995 , n231994 , n231482 );
not ( n231996 , n217044 );
buf ( n231997 , n229766 );
not ( n231998 , n231997 );
or ( n231999 , n231996 , n231998 );
nand ( n232000 , n229759 , n215131 );
nand ( n232001 , n231999 , n232000 );
not ( n232002 , n232001 );
or ( n232003 , n231476 , n232002 );
nand ( n232004 , n231995 , n232003 );
not ( n232005 , n213171 );
not ( n232006 , n213784 );
not ( n232007 , n232006 );
or ( n232008 , n232005 , n232007 );
nand ( n232009 , n232008 , n213382 );
not ( n232010 , n232009 );
xor ( n232011 , n232004 , n232010 );
not ( n232012 , n218232 );
not ( n232013 , n218208 );
not ( n232014 , n218268 );
or ( n232015 , n232013 , n232014 );
nand ( n232016 , n40710 , n221214 );
nand ( n232017 , n232015 , n232016 );
not ( n232018 , n232017 );
or ( n232019 , n232012 , n232018 );
nand ( n232020 , n231490 , n218221 );
nand ( n232021 , n232019 , n232020 );
xor ( n232022 , n232011 , n232021 );
xor ( n232023 , n231730 , n232022 );
xor ( n232024 , n232023 , n231323 );
xor ( n232025 , n231730 , n232022 );
and ( n232026 , n232025 , n231323 );
and ( n232027 , n231730 , n232022 );
or ( n232028 , n232026 , n232027 );
not ( n232029 , n225478 );
not ( n232030 , n231519 );
or ( n232031 , n232029 , n232030 );
not ( n232032 , n216422 );
not ( n232033 , n221031 );
or ( n232034 , n232032 , n232033 );
nand ( n232035 , n40668 , n227599 );
nand ( n232036 , n232034 , n232035 );
nand ( n232037 , n232036 , n219501 );
nand ( n232038 , n232031 , n232037 );
not ( n232039 , n229964 );
not ( n232040 , n229261 );
not ( n232041 , n221040 );
or ( n232042 , n232040 , n232041 );
nand ( n232043 , n40624 , n229262 );
nand ( n232044 , n232042 , n232043 );
not ( n232045 , n232044 );
or ( n232046 , n232039 , n232045 );
not ( n232047 , n229973 );
nand ( n232048 , n232047 , n231531 );
nand ( n232049 , n232046 , n232048 );
xor ( n232050 , n232038 , n232049 );
not ( n232051 , n217552 );
not ( n232052 , n231540 );
or ( n232053 , n232051 , n232052 );
not ( n232054 , n217542 );
not ( n232055 , n230819 );
or ( n232056 , n232054 , n232055 );
not ( n232057 , n39926 );
nand ( n232058 , n232057 , n216989 );
nand ( n232059 , n232056 , n232058 );
nand ( n232060 , n232059 , n220272 );
nand ( n232061 , n232053 , n232060 );
xor ( n232062 , n232050 , n232061 );
xor ( n232063 , n231742 , n232062 );
xor ( n232064 , n232063 , n231738 );
xor ( n232065 , n231742 , n232062 );
and ( n232066 , n232065 , n231738 );
and ( n232067 , n231742 , n232062 );
or ( n232068 , n232066 , n232067 );
xor ( n232069 , n231301 , n231359 );
not ( n232070 , n219731 );
not ( n232071 , n231597 );
or ( n232072 , n232070 , n232071 );
not ( n232073 , n216166 );
not ( n232074 , n224272 );
or ( n232075 , n232073 , n232074 );
nand ( n232076 , n39995 , n220538 );
nand ( n232077 , n232075 , n232076 );
nand ( n232078 , n232077 , n222185 );
nand ( n232079 , n232072 , n232078 );
not ( n232080 , n231018 );
not ( n232081 , n231503 );
or ( n232082 , n232080 , n232081 );
not ( n232083 , n217614 );
not ( n232084 , n219532 );
or ( n232085 , n232083 , n232084 );
nand ( n232086 , n219533 , n218253 );
nand ( n232087 , n232085 , n232086 );
nand ( n232088 , n232087 , n220067 );
nand ( n232089 , n232082 , n232088 );
xor ( n232090 , n232079 , n232089 );
not ( n232091 , n224624 );
not ( n232092 , n231608 );
or ( n232093 , n232091 , n232092 );
not ( n232094 , n219687 );
not ( n232095 , n224285 );
or ( n232096 , n232094 , n232095 );
nand ( n232097 , n40545 , n221283 );
nand ( n232098 , n232096 , n232097 );
nand ( n232099 , n232098 , n219314 );
nand ( n232100 , n232093 , n232099 );
xor ( n232101 , n232090 , n232100 );
xor ( n232102 , n232069 , n232101 );
xor ( n232103 , n231301 , n231359 );
and ( n232104 , n232103 , n232101 );
and ( n232105 , n231301 , n231359 );
or ( n232106 , n232104 , n232105 );
not ( n232107 , n221933 );
not ( n232108 , n226484 );
not ( n232109 , n222509 );
or ( n232110 , n232108 , n232109 );
nand ( n232111 , n40414 , n222333 );
nand ( n232112 , n232110 , n232111 );
not ( n232113 , n232112 );
or ( n232114 , n232107 , n232113 );
nand ( n232115 , n231560 , n215183 );
nand ( n232116 , n232114 , n232115 );
not ( n232117 , n220414 );
not ( n232118 , n231569 );
or ( n232119 , n232117 , n232118 );
not ( n232120 , n227912 );
not ( n232121 , n40181 );
or ( n232122 , n232120 , n232121 );
nand ( n232123 , n221716 , n220038 );
nand ( n232124 , n232122 , n232123 );
nand ( n232125 , n232124 , n220033 );
nand ( n232126 , n232119 , n232125 );
xor ( n232127 , n232116 , n232126 );
not ( n232128 , n223949 );
not ( n232129 , n226655 );
not ( n232130 , n40258 );
or ( n232131 , n232129 , n232130 );
nand ( n232132 , n221742 , n227927 );
nand ( n232133 , n232131 , n232132 );
not ( n232134 , n232133 );
or ( n232135 , n232128 , n232134 );
nand ( n232136 , n231580 , n227260 );
nand ( n232137 , n232135 , n232136 );
xor ( n232138 , n232127 , n232137 );
xor ( n232139 , n232138 , n231797 );
xor ( n232140 , n232139 , n231803 );
xor ( n232141 , n232138 , n231797 );
and ( n232142 , n232141 , n231803 );
and ( n232143 , n232138 , n231797 );
or ( n232144 , n232142 , n232143 );
xor ( n232145 , n231866 , n231875 );
and ( n232146 , n232145 , n231882 );
and ( n232147 , n231866 , n231875 );
or ( n232148 , n232146 , n232147 );
xor ( n232149 , n231832 , n231884 );
xor ( n232150 , n232149 , n231399 );
xor ( n232151 , n231832 , n231884 );
and ( n232152 , n232151 , n231399 );
and ( n232153 , n231832 , n231884 );
or ( n232154 , n232152 , n232153 );
xor ( n232155 , n231471 , n231949 );
xor ( n232156 , n232155 , n231513 );
xor ( n232157 , n231471 , n231949 );
and ( n232158 , n232157 , n231513 );
and ( n232159 , n231471 , n231949 );
or ( n232160 , n232158 , n232159 );
xor ( n232161 , n232024 , n231989 );
xor ( n232162 , n232161 , n231588 );
xor ( n232163 , n232024 , n231989 );
and ( n232164 , n232163 , n231588 );
and ( n232165 , n232024 , n231989 );
or ( n232166 , n232164 , n232165 );
xor ( n232167 , n231551 , n232102 );
xor ( n232168 , n232167 , n231617 );
xor ( n232169 , n231551 , n232102 );
and ( n232170 , n232169 , n231617 );
and ( n232171 , n231551 , n232102 );
or ( n232172 , n232170 , n232171 );
xor ( n232173 , n232064 , n231644 );
xor ( n232174 , n232173 , n231654 );
xor ( n232175 , n232064 , n231644 );
and ( n232176 , n232175 , n231654 );
and ( n232177 , n232064 , n231644 );
or ( n232178 , n232176 , n232177 );
xor ( n232179 , n232150 , n232140 );
xor ( n232180 , n232179 , n231660 );
xor ( n232181 , n232150 , n232140 );
and ( n232182 , n232181 , n231660 );
and ( n232183 , n232150 , n232140 );
or ( n232184 , n232182 , n232183 );
xor ( n232185 , n232156 , n231666 );
xor ( n232186 , n232185 , n232162 );
xor ( n232187 , n232156 , n231666 );
and ( n232188 , n232187 , n232162 );
and ( n232189 , n232156 , n231666 );
or ( n232190 , n232188 , n232189 );
xor ( n232191 , n231672 , n232168 );
xor ( n232192 , n232191 , n232174 );
xor ( n232193 , n231672 , n232168 );
and ( n232194 , n232193 , n232174 );
and ( n232195 , n231672 , n232168 );
or ( n232196 , n232194 , n232195 );
xor ( n232197 , n232180 , n231678 );
xor ( n232198 , n232197 , n231684 );
xor ( n232199 , n232180 , n231678 );
and ( n232200 , n232199 , n231684 );
and ( n232201 , n232180 , n231678 );
or ( n232202 , n232200 , n232201 );
xor ( n232203 , n231690 , n232186 );
xor ( n232204 , n232203 , n232192 );
xor ( n232205 , n231690 , n232186 );
and ( n232206 , n232205 , n232192 );
and ( n232207 , n231690 , n232186 );
or ( n232208 , n232206 , n232207 );
xor ( n232209 , n231895 , n231905 );
and ( n232210 , n232209 , n231917 );
and ( n232211 , n231895 , n231905 );
or ( n232212 , n232210 , n232211 );
xor ( n232213 , n232198 , n231696 );
xor ( n232214 , n232213 , n232204 );
xor ( n232215 , n232198 , n231696 );
and ( n232216 , n232215 , n232204 );
and ( n232217 , n232198 , n231696 );
or ( n232218 , n232216 , n232217 );
xor ( n232219 , n231702 , n231708 );
xor ( n232220 , n232219 , n232214 );
xor ( n232221 , n231702 , n231708 );
and ( n232222 , n232221 , n232214 );
and ( n232223 , n231702 , n231708 );
or ( n232224 , n232222 , n232223 );
xor ( n232225 , n231964 , n231975 );
and ( n232226 , n232225 , n231986 );
and ( n232227 , n231964 , n231975 );
or ( n232228 , n232226 , n232227 );
xor ( n232229 , n231929 , n231933 );
and ( n232230 , n232229 , n231947 );
and ( n232231 , n231929 , n231933 );
or ( n232232 , n232230 , n232231 );
xor ( n232233 , n232004 , n232010 );
and ( n232234 , n232233 , n232021 );
and ( n232235 , n232004 , n232010 );
or ( n232236 , n232234 , n232235 );
xor ( n232237 , n232079 , n232089 );
and ( n232238 , n232237 , n232100 );
and ( n232239 , n232079 , n232089 );
or ( n232240 , n232238 , n232239 );
xor ( n232241 , n232116 , n232126 );
and ( n232242 , n232241 , n232137 );
and ( n232243 , n232116 , n232126 );
or ( n232244 , n232242 , n232243 );
xor ( n232245 , n232038 , n232049 );
and ( n232246 , n232245 , n232061 );
and ( n232247 , n232038 , n232049 );
or ( n232248 , n232246 , n232247 );
not ( n232249 , n231870 );
not ( n232250 , n220163 );
or ( n232251 , n232249 , n232250 );
not ( n232252 , n216855 );
not ( n232253 , n232252 );
not ( n232254 , n220147 );
or ( n232255 , n232253 , n232254 );
nand ( n232256 , n222791 , n217314 );
nand ( n232257 , n232255 , n232256 );
nand ( n232258 , n220881 , n232257 );
nand ( n232259 , n232251 , n232258 );
and ( n232260 , n231232 , n222032 );
xor ( n232261 , n232259 , n232260 );
not ( n232262 , n220919 );
not ( n232263 , n231880 );
not ( n232264 , n232263 );
or ( n232265 , n232262 , n232264 );
not ( n232266 , n216311 );
not ( n232267 , n220901 );
or ( n232268 , n232266 , n232267 );
not ( n232269 , n223227 );
nand ( n232270 , n232269 , n216307 );
nand ( n232271 , n232268 , n232270 );
nand ( n232272 , n232271 , n220636 );
nand ( n232273 , n232265 , n232272 );
xor ( n232274 , n232261 , n232273 );
xor ( n232275 , n232259 , n232260 );
and ( n232276 , n232275 , n232273 );
and ( n232277 , n232259 , n232260 );
or ( n232278 , n232276 , n232277 );
or ( n232279 , n229648 , n231893 );
not ( n232280 , n223584 );
and ( n232281 , n232280 , n215796 );
not ( n232282 , n215796 );
and ( n232283 , n221608 , n232282 );
nor ( n232284 , n232281 , n232283 );
or ( n232285 , n221636 , n232284 );
nand ( n232286 , n232279 , n232285 );
not ( n232287 , n231903 );
not ( n232288 , n222886 );
or ( n232289 , n232287 , n232288 );
not ( n232290 , n226225 );
not ( n232291 , n222458 );
or ( n232292 , n232290 , n232291 );
nand ( n232293 , n222428 , n226224 );
nand ( n232294 , n232292 , n232293 );
nand ( n232295 , n232294 , n222467 );
nand ( n232296 , n232289 , n232295 );
xor ( n232297 , n232286 , n232296 );
not ( n232298 , n223591 );
not ( n232299 , n231915 );
or ( n232300 , n232298 , n232299 );
not ( n232301 , n225490 );
not ( n232302 , n223203 );
or ( n232303 , n232301 , n232302 );
nand ( n232304 , n223202 , n208726 );
nand ( n232305 , n232303 , n232304 );
nand ( n232306 , n232305 , n227294 );
nand ( n232307 , n232300 , n232306 );
xor ( n232308 , n232297 , n232307 );
xor ( n232309 , n232286 , n232296 );
and ( n232310 , n232309 , n232307 );
and ( n232311 , n232286 , n232296 );
or ( n232312 , n232310 , n232311 );
xor ( n232313 , n232228 , n232232 );
not ( n232314 , n220820 );
not ( n232315 , n216810 );
not ( n232316 , n39089 );
not ( n232317 , n232316 );
or ( n232318 , n232315 , n232317 );
nand ( n232319 , n39089 , n215289 );
nand ( n232320 , n232318 , n232319 );
not ( n232321 , n232320 );
or ( n232322 , n232314 , n232321 );
nand ( n232323 , n231826 , n216299 );
nand ( n232324 , n232322 , n232323 );
xor ( n232325 , n232313 , n232324 );
xor ( n232326 , n232228 , n232232 );
and ( n232327 , n232326 , n232324 );
and ( n232328 , n232228 , n232232 );
or ( n232329 , n232327 , n232328 );
not ( n232330 , n222185 );
not ( n232331 , n216166 );
not ( n232332 , n39877 );
or ( n232333 , n232331 , n232332 );
nand ( n232334 , n229198 , n220538 );
nand ( n232335 , n232333 , n232334 );
not ( n232336 , n232335 );
or ( n232337 , n232330 , n232336 );
nand ( n232338 , n232077 , n219731 );
nand ( n232339 , n232337 , n232338 );
not ( n232340 , n213152 );
not ( n232341 , n231781 );
or ( n232342 , n232340 , n232341 );
nand ( n232343 , n214818 , n217142 );
nand ( n232344 , n232342 , n232343 );
xor ( n232345 , n232339 , n232344 );
not ( n232346 , n219175 );
not ( n232347 , n219577 );
not ( n232348 , n228216 );
or ( n232349 , n232347 , n232348 );
nand ( n232350 , n39747 , n218661 );
nand ( n232351 , n232349 , n232350 );
not ( n232352 , n232351 );
or ( n232353 , n232346 , n232352 );
nand ( n232354 , n231852 , n217023 );
nand ( n232355 , n232353 , n232354 );
xor ( n232356 , n232345 , n232355 );
xor ( n232357 , n232339 , n232344 );
and ( n232358 , n232357 , n232355 );
and ( n232359 , n232339 , n232344 );
or ( n232360 , n232358 , n232359 );
not ( n232361 , n215383 );
not ( n232362 , n217573 );
not ( n232363 , n230219 );
or ( n232364 , n232362 , n232363 );
nand ( n232365 , n230223 , n219390 );
nand ( n232366 , n232364 , n232365 );
not ( n232367 , n232366 );
or ( n232368 , n232361 , n232367 );
nand ( n232369 , n231793 , n215605 );
nand ( n232370 , n232368 , n232369 );
not ( n232371 , n217552 );
not ( n232372 , n232059 );
or ( n232373 , n232371 , n232372 );
not ( n232374 , n215955 );
not ( n232375 , n225357 );
or ( n232376 , n232374 , n232375 );
nand ( n232377 , n39812 , n216989 );
nand ( n232378 , n232376 , n232377 );
nand ( n232379 , n220272 , n232378 );
nand ( n232380 , n232373 , n232379 );
xor ( n232381 , n232370 , n232380 );
xor ( n232382 , n232381 , n232274 );
xor ( n232383 , n232370 , n232380 );
and ( n232384 , n232383 , n232274 );
and ( n232385 , n232370 , n232380 );
or ( n232386 , n232384 , n232385 );
not ( n232387 , n232001 );
not ( n232388 , n229773 );
or ( n232389 , n232387 , n232388 );
not ( n232390 , n214537 );
not ( n232391 , n231477 );
or ( n232392 , n232390 , n232391 );
not ( n232393 , n231997 );
nand ( n232394 , n232393 , n214899 );
nand ( n232395 , n232392 , n232394 );
nand ( n232396 , n232395 , n229777 );
nand ( n232397 , n232389 , n232396 );
not ( n232398 , n231864 );
not ( n232399 , n230721 );
not ( n232400 , n232399 );
or ( n232401 , n232398 , n232400 );
buf ( n232402 , n230708 );
not ( n232403 , n214956 );
not ( n232404 , n231232 );
not ( n232405 , n232404 );
or ( n232406 , n232403 , n232405 );
nand ( n232407 , n231232 , n214960 );
nand ( n232408 , n232406 , n232407 );
nand ( n232409 , n232402 , n232408 );
nand ( n232410 , n232401 , n232409 );
xor ( n232411 , n232397 , n232410 );
not ( n232412 , n218843 );
buf ( n232413 , n218815 );
not ( n232414 , n232413 );
not ( n232415 , n217964 );
or ( n232416 , n232414 , n232415 );
nand ( n232417 , n208002 , n221238 );
nand ( n232418 , n232416 , n232417 );
not ( n232419 , n232418 );
or ( n232420 , n232412 , n232419 );
not ( n232421 , n223665 );
not ( n232422 , n232421 );
nand ( n232423 , n232422 , n231750 );
nand ( n232424 , n232420 , n232423 );
xor ( n232425 , n232411 , n232424 );
xor ( n232426 , n232308 , n232425 );
not ( n232427 , n231924 );
not ( n232428 , n227849 );
or ( n232429 , n232427 , n232428 );
not ( n232430 , n219102 );
not ( n232431 , n229823 );
not ( n232432 , n232431 );
or ( n232433 , n232430 , n232432 );
nand ( n232434 , n226651 , n216139 );
nand ( n232435 , n232433 , n232434 );
nand ( n232436 , n226885 , n232435 );
nand ( n232437 , n232429 , n232436 );
not ( n232438 , n231931 );
not ( n232439 , n232438 );
not ( n232440 , n228270 );
not ( n232441 , n232440 );
or ( n232442 , n232439 , n232441 );
and ( n232443 , n218514 , n231412 );
not ( n232444 , n218514 );
and ( n232445 , n232444 , n227595 );
nor ( n232446 , n232443 , n232445 );
not ( n232447 , n232446 );
nand ( n232448 , n232447 , n227737 );
nand ( n232449 , n232442 , n232448 );
xor ( n232450 , n232437 , n232449 );
not ( n232451 , n231421 );
not ( n232452 , n231945 );
or ( n232453 , n232451 , n232452 );
not ( n232454 , n228867 );
not ( n232455 , n216208 );
not ( n232456 , n231940 );
or ( n232457 , n232455 , n232456 );
not ( n232458 , n228727 );
nand ( n232459 , n232458 , n216207 );
nand ( n232460 , n232457 , n232459 );
not ( n232461 , n232460 );
or ( n232462 , n232454 , n232461 );
nand ( n232463 , n232453 , n232462 );
xor ( n232464 , n232450 , n232463 );
xor ( n232465 , n232426 , n232464 );
xor ( n232466 , n232308 , n232425 );
and ( n232467 , n232466 , n232464 );
and ( n232468 , n232308 , n232425 );
or ( n232469 , n232467 , n232468 );
not ( n232470 , n224086 );
not ( n232471 , n231962 );
or ( n232472 , n232470 , n232471 );
and ( n232473 , n224095 , n224492 );
and ( n232474 , n224096 , n224496 );
nor ( n232475 , n232473 , n232474 );
not ( n232476 , n224090 );
or ( n232477 , n232475 , n232476 );
nand ( n232478 , n232472 , n232477 );
not ( n232479 , n224938 );
not ( n232480 , n231973 );
or ( n232481 , n232479 , n232480 );
not ( n232482 , n226745 );
and ( n232483 , n216293 , n224925 );
not ( n232484 , n216293 );
not ( n232485 , n226747 );
and ( n232486 , n232484 , n232485 );
nor ( n232487 , n232483 , n232486 );
or ( n232488 , n232482 , n232487 );
nand ( n232489 , n232481 , n232488 );
xor ( n232490 , n232478 , n232489 );
not ( n232491 , n231984 );
or ( n232492 , n231453 , n232491 );
buf ( n232493 , n225743 );
not ( n232494 , n232493 );
and ( n232495 , n218980 , n232494 );
not ( n232496 , n218980 );
not ( n232497 , n225952 );
and ( n232498 , n232496 , n232497 );
nor ( n232499 , n232495 , n232498 );
or ( n232500 , n231456 , n232499 );
nand ( n232501 , n232492 , n232500 );
xor ( n232502 , n232490 , n232501 );
xor ( n232503 , n232502 , n232236 );
xor ( n232504 , n232503 , n232240 );
xor ( n232505 , n232502 , n232236 );
and ( n232506 , n232505 , n232240 );
and ( n232507 , n232502 , n232236 );
or ( n232508 , n232506 , n232507 );
xor ( n232509 , n232244 , n231807 );
not ( n232510 , n218533 );
not ( n232511 , n218208 );
not ( n232512 , n226486 );
or ( n232513 , n232511 , n232512 );
nand ( n232514 , n208044 , n218204 );
nand ( n232515 , n232513 , n232514 );
not ( n232516 , n232515 );
or ( n232517 , n232510 , n232516 );
nand ( n232518 , n232017 , n219836 );
nand ( n232519 , n232517 , n232518 );
xor ( n232520 , n232009 , n232519 );
not ( n232521 , n231766 );
or ( n232522 , n219791 , n232521 );
not ( n232523 , n41070 );
not ( n232524 , n227309 );
or ( n232525 , n232523 , n232524 );
not ( n232526 , n217977 );
nand ( n232527 , n232526 , n219440 );
nand ( n232528 , n232525 , n232527 );
not ( n232529 , n232528 );
or ( n232530 , n229612 , n232529 );
nand ( n232531 , n232522 , n232530 );
not ( n232532 , n232531 );
xor ( n232533 , n232520 , n232532 );
xor ( n232534 , n232509 , n232533 );
xor ( n232535 , n232244 , n231807 );
and ( n232536 , n232535 , n232533 );
and ( n232537 , n232244 , n231807 );
or ( n232538 , n232536 , n232537 );
xor ( n232539 , n232248 , n231801 );
xor ( n232540 , n232539 , n231836 );
xor ( n232541 , n232248 , n231801 );
and ( n232542 , n232541 , n231836 );
and ( n232543 , n232248 , n231801 );
or ( n232544 , n232542 , n232543 );
not ( n232545 , n224624 );
not ( n232546 , n232098 );
or ( n232547 , n232545 , n232546 );
not ( n232548 , n219687 );
not ( n232549 , n223764 );
or ( n232550 , n232548 , n232549 );
nand ( n232551 , n40045 , n222323 );
nand ( n232552 , n232550 , n232551 );
nand ( n232553 , n232552 , n219314 );
nand ( n232554 , n232547 , n232553 );
not ( n232555 , n221933 );
not ( n232556 , n218990 );
not ( n232557 , n223721 );
or ( n232558 , n232556 , n232557 );
nand ( n232559 , n223722 , n218994 );
nand ( n232560 , n232558 , n232559 );
not ( n232561 , n232560 );
or ( n232562 , n232555 , n232561 );
nand ( n232563 , n232112 , n215183 );
nand ( n232564 , n232562 , n232563 );
xor ( n232565 , n232554 , n232564 );
not ( n232566 , n226287 );
not ( n232567 , n226292 );
not ( n232568 , n222951 );
or ( n232569 , n232567 , n232568 );
nand ( n232570 , n40422 , n220038 );
nand ( n232571 , n232569 , n232570 );
not ( n232572 , n232571 );
or ( n232573 , n232566 , n232572 );
nand ( n232574 , n232124 , n220414 );
nand ( n232575 , n232573 , n232574 );
xor ( n232576 , n232565 , n232575 );
not ( n232577 , n227260 );
not ( n232578 , n232133 );
or ( n232579 , n232577 , n232578 );
or ( n232580 , n226655 , n40396 );
nand ( n232581 , n226655 , n40396 );
nand ( n232582 , n232580 , n232581 , n223949 );
nand ( n232583 , n232579 , n232582 );
not ( n232584 , n232036 );
not ( n232585 , n225478 );
or ( n232586 , n232584 , n232585 );
not ( n232587 , n216422 );
not ( n232588 , n221330 );
or ( n232589 , n232587 , n232588 );
nand ( n232590 , n40410 , n227599 );
nand ( n232591 , n232589 , n232590 );
nand ( n232592 , n232591 , n219501 );
nand ( n232593 , n232586 , n232592 );
xor ( n232594 , n232583 , n232593 );
not ( n232595 , n229964 );
not ( n232596 , n229261 );
not ( n232597 , n221356 );
or ( n232598 , n232596 , n232597 );
nand ( n232599 , n207936 , n229257 );
nand ( n232600 , n232598 , n232599 );
not ( n232601 , n232600 );
or ( n232602 , n232595 , n232601 );
nand ( n232603 , n232044 , n229974 );
nand ( n232604 , n232602 , n232603 );
xor ( n232605 , n232594 , n232604 );
xor ( n232606 , n232576 , n232605 );
xor ( n232607 , n232606 , n231888 );
xor ( n232608 , n232576 , n232605 );
and ( n232609 , n232608 , n231888 );
and ( n232610 , n232576 , n232605 );
or ( n232611 , n232609 , n232610 );
not ( n232612 , n231018 );
not ( n232613 , n232087 );
or ( n232614 , n232612 , n232613 );
not ( n232615 , n231500 );
not ( n232616 , n228452 );
or ( n232617 , n232615 , n232616 );
nand ( n232618 , n219226 , n218253 );
nand ( n232619 , n232617 , n232618 );
nand ( n232620 , n232619 , n220067 );
nand ( n232621 , n232614 , n232620 );
not ( n232622 , n213577 );
not ( n232623 , n231842 );
or ( n232624 , n232622 , n232623 );
not ( n232625 , n213735 );
not ( n232626 , n230556 );
or ( n232627 , n232625 , n232626 );
not ( n232628 , n213735 );
nand ( n232629 , n232628 , n209864 );
nand ( n232630 , n232627 , n232629 );
nand ( n232631 , n232630 , n216336 );
nand ( n232632 , n232624 , n232631 );
xor ( n232633 , n232621 , n232632 );
xor ( n232634 , n232633 , n231773 );
xor ( n232635 , n232634 , n231953 );
xor ( n232636 , n232635 , n232356 );
xor ( n232637 , n232634 , n231953 );
and ( n232638 , n232637 , n232356 );
and ( n232639 , n232634 , n231953 );
or ( n232640 , n232638 , n232639 );
xor ( n232641 , n232325 , n232382 );
not ( n232642 , n214717 );
not ( n232643 , n231817 );
or ( n232644 , n232642 , n232643 );
and ( n232645 , n39363 , n216037 );
not ( n232646 , n39363 );
and ( n232647 , n232646 , n221338 );
or ( n232648 , n232645 , n232647 );
nand ( n232649 , n232648 , n220985 );
nand ( n232650 , n232644 , n232649 );
xor ( n232651 , n232650 , n232148 );
xor ( n232652 , n232651 , n232212 );
xor ( n232653 , n232641 , n232652 );
xor ( n232654 , n232325 , n232382 );
and ( n232655 , n232654 , n232652 );
and ( n232656 , n232325 , n232382 );
or ( n232657 , n232655 , n232656 );
xor ( n232658 , n232478 , n232489 );
and ( n232659 , n232658 , n232501 );
and ( n232660 , n232478 , n232489 );
or ( n232661 , n232659 , n232660 );
xor ( n232662 , n231993 , n232465 );
xor ( n232663 , n232662 , n232068 );
xor ( n232664 , n231993 , n232465 );
and ( n232665 , n232664 , n232068 );
and ( n232666 , n231993 , n232465 );
or ( n232667 , n232665 , n232666 );
xor ( n232668 , n232106 , n232504 );
xor ( n232669 , n232668 , n232028 );
xor ( n232670 , n232106 , n232504 );
and ( n232671 , n232670 , n232028 );
and ( n232672 , n232106 , n232504 );
or ( n232673 , n232671 , n232672 );
xor ( n232674 , n232534 , n232540 );
xor ( n232675 , n232674 , n232154 );
xor ( n232676 , n232534 , n232540 );
and ( n232677 , n232676 , n232154 );
and ( n232678 , n232534 , n232540 );
or ( n232679 , n232677 , n232678 );
xor ( n232680 , n232607 , n232144 );
xor ( n232681 , n232680 , n232653 );
xor ( n232682 , n232607 , n232144 );
and ( n232683 , n232682 , n232653 );
and ( n232684 , n232607 , n232144 );
or ( n232685 , n232683 , n232684 );
xor ( n232686 , n232160 , n232636 );
xor ( n232687 , n232686 , n232663 );
xor ( n232688 , n232160 , n232636 );
and ( n232689 , n232688 , n232663 );
and ( n232690 , n232160 , n232636 );
or ( n232691 , n232689 , n232690 );
xor ( n232692 , n232166 , n232172 );
xor ( n232693 , n232692 , n232669 );
xor ( n232694 , n232166 , n232172 );
and ( n232695 , n232694 , n232669 );
and ( n232696 , n232166 , n232172 );
or ( n232697 , n232695 , n232696 );
xor ( n232698 , n232681 , n232178 );
xor ( n232699 , n232698 , n232675 );
xor ( n232700 , n232681 , n232178 );
and ( n232701 , n232700 , n232675 );
and ( n232702 , n232681 , n232178 );
or ( n232703 , n232701 , n232702 );
xor ( n232704 , n232687 , n232184 );
xor ( n232705 , n232704 , n232190 );
xor ( n232706 , n232687 , n232184 );
and ( n232707 , n232706 , n232190 );
and ( n232708 , n232687 , n232184 );
or ( n232709 , n232707 , n232708 );
xor ( n232710 , n232693 , n232196 );
xor ( n232711 , n232710 , n232699 );
xor ( n232712 , n232693 , n232196 );
and ( n232713 , n232712 , n232699 );
and ( n232714 , n232693 , n232196 );
or ( n232715 , n232713 , n232714 );
xor ( n232716 , n232202 , n232705 );
xor ( n232717 , n232716 , n232208 );
xor ( n232718 , n232202 , n232705 );
and ( n232719 , n232718 , n232208 );
and ( n232720 , n232202 , n232705 );
or ( n232721 , n232719 , n232720 );
xor ( n232722 , n232437 , n232449 );
and ( n232723 , n232722 , n232463 );
and ( n232724 , n232437 , n232449 );
or ( n232725 , n232723 , n232724 );
xor ( n232726 , n232711 , n232717 );
xor ( n232727 , n232726 , n232218 );
xor ( n232728 , n232711 , n232717 );
and ( n232729 , n232728 , n232218 );
and ( n232730 , n232711 , n232717 );
or ( n232731 , n232729 , n232730 );
xor ( n232732 , n232397 , n232410 );
and ( n232733 , n232732 , n232424 );
and ( n232734 , n232397 , n232410 );
or ( n232735 , n232733 , n232734 );
xor ( n232736 , n232009 , n232519 );
and ( n232737 , n232736 , n232532 );
and ( n232738 , n232009 , n232519 );
or ( n232739 , n232737 , n232738 );
xor ( n232740 , n232554 , n232564 );
and ( n232741 , n232740 , n232575 );
and ( n232742 , n232554 , n232564 );
or ( n232743 , n232741 , n232742 );
xor ( n232744 , n232583 , n232593 );
and ( n232745 , n232744 , n232604 );
and ( n232746 , n232583 , n232593 );
or ( n232747 , n232745 , n232746 );
xor ( n232748 , n232621 , n232632 );
and ( n232749 , n232748 , n231773 );
and ( n232750 , n232621 , n232632 );
or ( n232751 , n232749 , n232750 );
xor ( n232752 , n232650 , n232148 );
and ( n232753 , n232752 , n232212 );
and ( n232754 , n232650 , n232148 );
or ( n232755 , n232753 , n232754 );
or ( n232756 , n213758 , n213058 );
nand ( n232757 , n232756 , n216262 );
not ( n232758 , n219075 );
not ( n232759 , n217713 );
not ( n232760 , n220180 );
or ( n232761 , n232759 , n232760 );
nand ( n232762 , n219423 , n41164 );
nand ( n232763 , n232761 , n232762 );
not ( n232764 , n232763 );
or ( n232765 , n232758 , n232764 );
nand ( n232766 , n232528 , n223620 );
nand ( n232767 , n232765 , n232766 );
xor ( n232768 , n232757 , n232767 );
not ( n232769 , n232257 );
not ( n232770 , n220162 );
or ( n232771 , n232769 , n232770 );
not ( n232772 , n218137 );
not ( n232773 , n224563 );
or ( n232774 , n232772 , n232773 );
nand ( n232775 , n222791 , n217116 );
nand ( n232776 , n232774 , n232775 );
nand ( n232777 , n220881 , n232776 );
nand ( n232778 , n232771 , n232777 );
xor ( n232779 , n232768 , n232778 );
xor ( n232780 , n232757 , n232767 );
and ( n232781 , n232780 , n232778 );
and ( n232782 , n232757 , n232767 );
or ( n232783 , n232781 , n232782 );
not ( n232784 , n232404 );
and ( n232785 , n232784 , n213583 );
not ( n232786 , n217148 );
not ( n232787 , n224112 );
or ( n232788 , n232786 , n232787 );
nand ( n232789 , n220900 , n216520 );
nand ( n232790 , n232788 , n232789 );
not ( n232791 , n232790 );
not ( n232792 , n220929 );
or ( n232793 , n232791 , n232792 );
not ( n232794 , n228639 );
nand ( n232795 , n232794 , n232271 );
nand ( n232796 , n232793 , n232795 );
xor ( n232797 , n232785 , n232796 );
not ( n232798 , n221625 );
or ( n232799 , n232798 , n232284 );
not ( n232800 , n222586 );
not ( n232801 , n217133 );
or ( n232802 , n232800 , n232801 );
not ( n232803 , n219582 );
nand ( n232804 , n232803 , n221608 );
nand ( n232805 , n232802 , n232804 );
not ( n232806 , n232805 );
or ( n232807 , n232806 , n223176 );
nand ( n232808 , n232799 , n232807 );
xor ( n232809 , n232797 , n232808 );
xor ( n232810 , n232785 , n232796 );
and ( n232811 , n232810 , n232808 );
and ( n232812 , n232785 , n232796 );
or ( n232813 , n232811 , n232812 );
not ( n232814 , n220985 );
not ( n232815 , n215113 );
not ( n232816 , n230025 );
or ( n232817 , n232815 , n232816 );
nand ( n232818 , n39286 , n216037 );
nand ( n232819 , n232817 , n232818 );
not ( n232820 , n232819 );
or ( n232821 , n232814 , n232820 );
nand ( n232822 , n232648 , n214717 );
nand ( n232823 , n232821 , n232822 );
xor ( n232824 , n232823 , n232661 );
xor ( n232825 , n232824 , n232725 );
xor ( n232826 , n232823 , n232661 );
and ( n232827 , n232826 , n232725 );
and ( n232828 , n232823 , n232661 );
or ( n232829 , n232827 , n232828 );
not ( n232830 , n220820 );
not ( n232831 , n216810 );
not ( n232832 , n229704 );
or ( n232833 , n232831 , n232832 );
nand ( n232834 , n38532 , n221307 );
nand ( n232835 , n232833 , n232834 );
not ( n232836 , n232835 );
or ( n232837 , n232830 , n232836 );
nand ( n232838 , n232320 , n216562 );
nand ( n232839 , n232837 , n232838 );
not ( n232840 , n219175 );
not ( n232841 , n217017 );
not ( n232842 , n39607 );
not ( n232843 , n232842 );
or ( n232844 , n232841 , n232843 );
nand ( n232845 , n39607 , n218661 );
nand ( n232846 , n232844 , n232845 );
not ( n232847 , n232846 );
or ( n232848 , n232840 , n232847 );
nand ( n232849 , n232351 , n217023 );
nand ( n232850 , n232848 , n232849 );
xor ( n232851 , n232839 , n232850 );
not ( n232852 , n232366 );
or ( n232853 , n232852 , n214085 );
and ( n232854 , n217573 , n209709 );
not ( n232855 , n217573 );
not ( n232856 , n209709 );
and ( n232857 , n232855 , n232856 );
or ( n232858 , n232854 , n232857 );
not ( n232859 , n232858 );
or ( n232860 , n232859 , n223390 );
nand ( n232861 , n232853 , n232860 );
xor ( n232862 , n232851 , n232861 );
xor ( n232863 , n232839 , n232850 );
and ( n232864 , n232863 , n232861 );
and ( n232865 , n232839 , n232850 );
or ( n232866 , n232864 , n232865 );
not ( n232867 , n220272 );
not ( n232868 , n215955 );
not ( n232869 , n225792 );
or ( n232870 , n232868 , n232869 );
nand ( n232871 , n39713 , n219358 );
nand ( n232872 , n232870 , n232871 );
not ( n232873 , n232872 );
or ( n232874 , n232867 , n232873 );
nand ( n232875 , n232378 , n220280 );
nand ( n232876 , n232874 , n232875 );
xor ( n232877 , n232876 , n232809 );
xor ( n232878 , n232877 , n232735 );
xor ( n232879 , n232876 , n232809 );
and ( n232880 , n232879 , n232735 );
and ( n232881 , n232876 , n232809 );
or ( n232882 , n232880 , n232881 );
not ( n232883 , n232294 );
not ( n232884 , n222453 );
or ( n232885 , n232883 , n232884 );
not ( n232886 , n41565 );
not ( n232887 , n222461 );
or ( n232888 , n232886 , n232887 );
nand ( n232889 , n222428 , n216543 );
nand ( n232890 , n232888 , n232889 );
nand ( n232891 , n232890 , n223243 );
nand ( n232892 , n232885 , n232891 );
not ( n232893 , n232305 );
not ( n232894 , n223591 );
or ( n232895 , n232893 , n232894 );
not ( n232896 , n225764 );
not ( n232897 , n223186 );
or ( n232898 , n232896 , n232897 );
nand ( n232899 , n226809 , n225769 );
nand ( n232900 , n232898 , n232899 );
nand ( n232901 , n232900 , n222768 );
nand ( n232902 , n232895 , n232901 );
xor ( n232903 , n232892 , n232902 );
not ( n232904 , n224086 );
or ( n232905 , n232904 , n232475 );
and ( n232906 , n224975 , n214837 );
and ( n232907 , n226355 , n226698 );
nor ( n232908 , n232906 , n232907 );
or ( n232909 , n232476 , n232908 );
nand ( n232910 , n232905 , n232909 );
xor ( n232911 , n232903 , n232910 );
xor ( n232912 , n232779 , n232911 );
or ( n232913 , n232446 , n227733 );
and ( n232914 , n231412 , n216934 );
and ( n232915 , n228279 , n216940 );
nor ( n232916 , n232914 , n232915 );
not ( n232917 , n227165 );
or ( n232918 , n232916 , n232917 );
nand ( n232919 , n232913 , n232918 );
not ( n232920 , n232460 );
not ( n232921 , n228858 );
or ( n232922 , n232920 , n232921 );
not ( n232923 , n215075 );
not ( n232924 , n228847 );
or ( n232925 , n232923 , n232924 );
nand ( n232926 , n228726 , n215899 );
nand ( n232927 , n232925 , n232926 );
nand ( n232928 , n232927 , n229738 );
nand ( n232929 , n232922 , n232928 );
xor ( n232930 , n232919 , n232929 );
not ( n232931 , n232395 );
not ( n232932 , n229773 );
or ( n232933 , n232931 , n232932 );
not ( n232934 , n216964 );
not ( n232935 , n229762 );
or ( n232936 , n232934 , n232935 );
nand ( n232937 , n229761 , n214678 );
nand ( n232938 , n232936 , n232937 );
nand ( n232939 , n232938 , n229777 );
nand ( n232940 , n232933 , n232939 );
xor ( n232941 , n232930 , n232940 );
xor ( n232942 , n232912 , n232941 );
xor ( n232943 , n232779 , n232911 );
and ( n232944 , n232943 , n232941 );
and ( n232945 , n232779 , n232911 );
or ( n232946 , n232944 , n232945 );
or ( n232947 , n232479 , n232487 );
not ( n232948 , n224941 );
and ( n232949 , n224925 , n224037 );
and ( n232950 , n224929 , n224041 );
nor ( n232951 , n232949 , n232950 );
or ( n232952 , n232948 , n232951 );
nand ( n232953 , n232947 , n232952 );
not ( n232954 , n232499 );
not ( n232955 , n232954 );
not ( n232956 , n230389 );
not ( n232957 , n232956 );
or ( n232958 , n232955 , n232957 );
not ( n232959 , n221495 );
not ( n232960 , n232493 );
or ( n232961 , n232959 , n232960 );
not ( n232962 , n225743 );
nand ( n232963 , n232962 , n220022 );
nand ( n232964 , n232961 , n232963 );
nand ( n232965 , n228775 , n232964 );
nand ( n232966 , n232958 , n232965 );
xor ( n232967 , n232953 , n232966 );
not ( n232968 , n232435 );
not ( n232969 , n229816 );
or ( n232970 , n232968 , n232969 );
not ( n232971 , n219343 );
not ( n232972 , n226650 );
or ( n232973 , n232971 , n232972 );
not ( n232974 , n230897 );
nand ( n232975 , n232974 , n219348 );
nand ( n232976 , n232973 , n232975 );
nand ( n232977 , n226885 , n232976 );
nand ( n232978 , n232970 , n232977 );
xor ( n232979 , n232967 , n232978 );
xor ( n232980 , n232979 , n232739 );
xor ( n232981 , n232980 , n232743 );
xor ( n232982 , n232979 , n232739 );
and ( n232983 , n232982 , n232743 );
and ( n232984 , n232979 , n232739 );
or ( n232985 , n232983 , n232984 );
xor ( n232986 , n232747 , n232360 );
xor ( n232987 , n232986 , n232751 );
xor ( n232988 , n232747 , n232360 );
and ( n232989 , n232988 , n232751 );
and ( n232990 , n232747 , n232360 );
or ( n232991 , n232989 , n232990 );
xor ( n232992 , n232755 , n232329 );
not ( n232993 , n229974 );
not ( n232994 , n232600 );
or ( n232995 , n232993 , n232994 );
not ( n232996 , n229261 );
not ( n232997 , n220216 );
or ( n232998 , n232996 , n232997 );
nand ( n232999 , n220217 , n229257 );
nand ( n233000 , n232998 , n232999 );
nand ( n233001 , n233000 , n229964 );
nand ( n233002 , n232995 , n233001 );
not ( n233003 , n220067 );
not ( n233004 , n221040 );
not ( n233005 , n231500 );
or ( n233006 , n233004 , n233005 );
nand ( n233007 , n219522 , n218253 );
nand ( n233008 , n233006 , n233007 );
not ( n233009 , n233008 );
or ( n233010 , n233003 , n233009 );
nand ( n233011 , n232619 , n231018 );
nand ( n233012 , n233010 , n233011 );
xor ( n233013 , n233002 , n233012 );
not ( n233014 , n222185 );
not ( n233015 , n219033 );
not ( n233016 , n39927 );
or ( n233017 , n233015 , n233016 );
not ( n233018 , n39926 );
nand ( n233019 , n233018 , n220538 );
nand ( n233020 , n233017 , n233019 );
not ( n233021 , n233020 );
or ( n233022 , n233014 , n233021 );
nand ( n233023 , n232335 , n219731 );
nand ( n233024 , n233022 , n233023 );
xor ( n233025 , n233013 , n233024 );
xor ( n233026 , n232992 , n233025 );
xor ( n233027 , n232755 , n232329 );
and ( n233028 , n233027 , n233025 );
and ( n233029 , n232755 , n232329 );
or ( n233030 , n233028 , n233029 );
not ( n233031 , n220414 );
not ( n233032 , n232571 );
or ( n233033 , n233031 , n233032 );
not ( n233034 , n227912 );
not ( n233035 , n40414 );
not ( n233036 , n233035 );
or ( n233037 , n233034 , n233036 );
not ( n233038 , n226292 );
nand ( n233039 , n233038 , n222513 );
nand ( n233040 , n233037 , n233039 );
nand ( n233041 , n233040 , n220033 );
nand ( n233042 , n233033 , n233041 );
not ( n233043 , n223949 );
not ( n233044 , n226655 );
not ( n233045 , n40181 );
or ( n233046 , n233044 , n233045 );
nand ( n233047 , n223320 , n227927 );
nand ( n233048 , n233046 , n233047 );
not ( n233049 , n233048 );
or ( n233050 , n233043 , n233049 );
and ( n233051 , n40396 , n226655 );
not ( n233052 , n40396 );
not ( n233053 , n226655 );
and ( n233054 , n233052 , n233053 );
nor ( n233055 , n233051 , n233054 );
nand ( n233056 , n233055 , n227260 );
nand ( n233057 , n233050 , n233056 );
xor ( n233058 , n233042 , n233057 );
not ( n233059 , n228237 );
not ( n233060 , n216422 );
not ( n233061 , n40258 );
or ( n233062 , n233060 , n233061 );
nand ( n233063 , n226911 , n227602 );
nand ( n233064 , n233062 , n233063 );
not ( n233065 , n233064 );
or ( n233066 , n233059 , n233065 );
nand ( n233067 , n232591 , n225478 );
nand ( n233068 , n233066 , n233067 );
xor ( n233069 , n233058 , n233068 );
not ( n233070 , n216204 );
not ( n233071 , n232552 );
or ( n233072 , n233070 , n233071 );
not ( n233073 , n219687 );
not ( n233074 , n225108 );
or ( n233075 , n233073 , n233074 );
nand ( n233076 , n225111 , n221283 );
nand ( n233077 , n233075 , n233076 );
nand ( n233078 , n219314 , n233077 );
nand ( n233079 , n233072 , n233078 );
not ( n233080 , n219461 );
not ( n233081 , n232515 );
or ( n233082 , n233080 , n233081 );
not ( n233083 , n218226 );
not ( n233084 , n233083 );
not ( n233085 , n219532 );
or ( n233086 , n233084 , n233085 );
nand ( n233087 , n219533 , n220091 );
nand ( n233088 , n233086 , n233087 );
nand ( n233089 , n233088 , n218533 );
nand ( n233090 , n233082 , n233089 );
xor ( n233091 , n233079 , n233090 );
not ( n233092 , n221933 );
not ( n233093 , n218990 );
not ( n233094 , n223330 );
or ( n233095 , n233093 , n233094 );
nand ( n233096 , n224286 , n218994 );
nand ( n233097 , n233095 , n233096 );
not ( n233098 , n233097 );
or ( n233099 , n233092 , n233098 );
nand ( n233100 , n232560 , n219332 );
nand ( n233101 , n233099 , n233100 );
xor ( n233102 , n233091 , n233101 );
xor ( n233103 , n233069 , n233102 );
not ( n233104 , n232408 );
not ( n233105 , n230721 );
not ( n233106 , n233105 );
or ( n233107 , n233104 , n233106 );
and ( n233108 , n214357 , n230722 );
not ( n233109 , n214357 );
and ( n233110 , n233109 , n230726 );
or ( n233111 , n233108 , n233110 );
nand ( n233112 , n232402 , n233111 );
nand ( n233113 , n233107 , n233112 );
not ( n233114 , n232418 );
not ( n233115 , n223665 );
or ( n233116 , n233114 , n233115 );
not ( n233117 , n221237 );
not ( n233118 , n232413 );
not ( n233119 , n219595 );
or ( n233120 , n233118 , n233119 );
nand ( n233121 , n40710 , n221238 );
nand ( n233122 , n233120 , n233121 );
nand ( n233123 , n233117 , n233122 );
nand ( n233124 , n233116 , n233123 );
xor ( n233125 , n233113 , n233124 );
xor ( n233126 , n233125 , n232531 );
xor ( n233127 , n233103 , n233126 );
xor ( n233128 , n233069 , n233102 );
and ( n233129 , n233128 , n233126 );
and ( n233130 , n233069 , n233102 );
or ( n233131 , n233129 , n233130 );
not ( n233132 , n216336 );
not ( n233133 , n213735 );
not ( n233134 , n231103 );
not ( n233135 , n233134 );
or ( n233136 , n233133 , n233135 );
nand ( n233137 , n213732 , n209961 );
nand ( n233138 , n233136 , n233137 );
not ( n233139 , n233138 );
or ( n233140 , n233132 , n233139 );
nand ( n233141 , n232630 , n213577 );
nand ( n233142 , n233140 , n233141 );
xor ( n233143 , n233142 , n232278 );
xor ( n233144 , n233143 , n232312 );
xor ( n233145 , n233144 , n232469 );
xor ( n233146 , n233145 , n232862 );
xor ( n233147 , n233144 , n232469 );
and ( n233148 , n233147 , n232862 );
and ( n233149 , n233144 , n232469 );
or ( n233150 , n233148 , n233149 );
xor ( n233151 , n232386 , n232825 );
xor ( n233152 , n233151 , n232878 );
xor ( n233153 , n232386 , n232825 );
and ( n233154 , n233153 , n232878 );
and ( n233155 , n232386 , n232825 );
or ( n233156 , n233154 , n233155 );
xor ( n233157 , n232892 , n232902 );
and ( n233158 , n233157 , n232910 );
and ( n233159 , n232892 , n232902 );
or ( n233160 , n233158 , n233159 );
xor ( n233161 , n232942 , n232508 );
xor ( n233162 , n233161 , n232981 );
xor ( n233163 , n232942 , n232508 );
and ( n233164 , n233163 , n232981 );
and ( n233165 , n232942 , n232508 );
or ( n233166 , n233164 , n233165 );
xor ( n233167 , n232544 , n232538 );
xor ( n233168 , n233167 , n232640 );
xor ( n233169 , n232544 , n232538 );
and ( n233170 , n233169 , n232640 );
and ( n233171 , n232544 , n232538 );
or ( n233172 , n233170 , n233171 );
xor ( n233173 , n232987 , n233026 );
xor ( n233174 , n233173 , n232657 );
xor ( n233175 , n232987 , n233026 );
and ( n233176 , n233175 , n232657 );
and ( n233177 , n232987 , n233026 );
or ( n233178 , n233176 , n233177 );
xor ( n233179 , n233127 , n232611 );
xor ( n233180 , n233179 , n233146 );
xor ( n233181 , n233127 , n232611 );
and ( n233182 , n233181 , n233146 );
and ( n233183 , n233127 , n232611 );
or ( n233184 , n233182 , n233183 );
xor ( n233185 , n233152 , n232673 );
xor ( n233186 , n233185 , n232667 );
xor ( n233187 , n233152 , n232673 );
and ( n233188 , n233187 , n232667 );
and ( n233189 , n233152 , n232673 );
or ( n233190 , n233188 , n233189 );
xor ( n233191 , n233162 , n232679 );
xor ( n233192 , n233191 , n233168 );
xor ( n233193 , n233162 , n232679 );
and ( n233194 , n233193 , n233168 );
and ( n233195 , n233162 , n232679 );
or ( n233196 , n233194 , n233195 );
xor ( n233197 , n232685 , n233174 );
xor ( n233198 , n233197 , n233180 );
xor ( n233199 , n232685 , n233174 );
and ( n233200 , n233199 , n233180 );
and ( n233201 , n232685 , n233174 );
or ( n233202 , n233200 , n233201 );
xor ( n233203 , n232691 , n232697 );
xor ( n233204 , n233203 , n233186 );
xor ( n233205 , n232691 , n232697 );
and ( n233206 , n233205 , n233186 );
and ( n233207 , n232691 , n232697 );
or ( n233208 , n233206 , n233207 );
xor ( n233209 , n232703 , n233192 );
xor ( n233210 , n233209 , n233198 );
xor ( n233211 , n232703 , n233192 );
and ( n233212 , n233211 , n233198 );
and ( n233213 , n232703 , n233192 );
or ( n233214 , n233212 , n233213 );
xor ( n233215 , n232709 , n233204 );
xor ( n233216 , n233215 , n233210 );
xor ( n233217 , n232709 , n233204 );
and ( n233218 , n233217 , n233210 );
and ( n233219 , n232709 , n233204 );
or ( n233220 , n233218 , n233219 );
xor ( n233221 , n232953 , n232966 );
and ( n233222 , n233221 , n232978 );
and ( n233223 , n232953 , n232966 );
or ( n233224 , n233222 , n233223 );
xor ( n233225 , n232715 , n233216 );
xor ( n233226 , n233225 , n232721 );
xor ( n233227 , n232715 , n233216 );
and ( n233228 , n233227 , n232721 );
and ( n233229 , n232715 , n233216 );
or ( n233230 , n233228 , n233229 );
xor ( n233231 , n232919 , n232929 );
and ( n233232 , n233231 , n232940 );
and ( n233233 , n232919 , n232929 );
or ( n233234 , n233232 , n233233 );
xor ( n233235 , n233113 , n233124 );
and ( n233236 , n233235 , n232531 );
and ( n233237 , n233113 , n233124 );
or ( n233238 , n233236 , n233237 );
xor ( n233239 , n233079 , n233090 );
and ( n233240 , n233239 , n233101 );
and ( n233241 , n233079 , n233090 );
or ( n233242 , n233240 , n233241 );
xor ( n233243 , n233042 , n233057 );
and ( n233244 , n233243 , n233068 );
and ( n233245 , n233042 , n233057 );
or ( n233246 , n233244 , n233245 );
xor ( n233247 , n233002 , n233012 );
and ( n233248 , n233247 , n233024 );
and ( n233249 , n233002 , n233012 );
or ( n233250 , n233248 , n233249 );
xor ( n233251 , n233142 , n232278 );
and ( n233252 , n233251 , n232312 );
and ( n233253 , n233142 , n232278 );
or ( n233254 , n233252 , n233253 );
not ( n233255 , n232790 );
not ( n233256 , n220919 );
or ( n233257 , n233255 , n233256 );
not ( n233258 , n232252 );
not ( n233259 , n223227 );
or ( n233260 , n233258 , n233259 );
nand ( n233261 , n220900 , n217314 );
nand ( n233262 , n233260 , n233261 );
nand ( n233263 , n233262 , n220636 );
nand ( n233264 , n233257 , n233263 );
not ( n233265 , n232805 );
not ( n233266 , n221625 );
or ( n233267 , n233265 , n233266 );
not ( n233268 , n216311 );
not ( n233269 , n232280 );
or ( n233270 , n233268 , n233269 );
nand ( n233271 , n223584 , n216307 );
nand ( n233272 , n233270 , n233271 );
nand ( n233273 , n223177 , n233272 );
nand ( n233274 , n233267 , n233273 );
xor ( n233275 , n233264 , n233274 );
not ( n233276 , n232890 );
not ( n233277 , n222886 );
or ( n233278 , n233276 , n233277 );
not ( n233279 , n217941 );
not ( n233280 , n233279 );
not ( n233281 , n222458 );
or ( n233282 , n233280 , n233281 );
nand ( n233283 , n222462 , n217394 );
nand ( n233284 , n233282 , n233283 );
nand ( n233285 , n233284 , n222158 );
nand ( n233286 , n233278 , n233285 );
xor ( n233287 , n233275 , n233286 );
xor ( n233288 , n233264 , n233274 );
and ( n233289 , n233288 , n233286 );
and ( n233290 , n233264 , n233274 );
or ( n233291 , n233289 , n233290 );
not ( n233292 , n226225 );
not ( n233293 , n223203 );
or ( n233294 , n233292 , n233293 );
nand ( n233295 , n223202 , n226224 );
nand ( n233296 , n233294 , n233295 );
not ( n233297 , n233296 );
not ( n233298 , n222769 );
or ( n233299 , n233297 , n233298 );
nand ( n233300 , n232900 , n223591 );
nand ( n233301 , n233299 , n233300 );
not ( n233302 , n232908 );
not ( n233303 , n233302 );
not ( n233304 , n224086 );
or ( n233305 , n233303 , n233304 );
not ( n233306 , n226304 );
not ( n233307 , n224069 );
or ( n233308 , n233306 , n233307 );
buf ( n233309 , n224974 );
nand ( n233310 , n233309 , n225489 );
nand ( n233311 , n233308 , n233310 );
nand ( n233312 , n224090 , n233311 );
nand ( n233313 , n233305 , n233312 );
xor ( n233314 , n233301 , n233313 );
buf ( n233315 , n226742 );
not ( n233316 , n233315 );
or ( n233317 , n233316 , n232951 );
and ( n233318 , n224925 , n224492 );
and ( n233319 , n224929 , n214642 );
nor ( n233320 , n233318 , n233319 );
or ( n233321 , n232948 , n233320 );
nand ( n233322 , n233317 , n233321 );
xor ( n233323 , n233314 , n233322 );
xor ( n233324 , n233301 , n233313 );
and ( n233325 , n233324 , n233322 );
and ( n233326 , n233301 , n233313 );
or ( n233327 , n233325 , n233326 );
not ( n233328 , n219175 );
not ( n233329 , n217017 );
not ( n233330 , n227201 );
or ( n233331 , n233329 , n233330 );
nand ( n233332 , n230462 , n219583 );
nand ( n233333 , n233331 , n233332 );
not ( n233334 , n233333 );
or ( n233335 , n233328 , n233334 );
nand ( n233336 , n232846 , n217023 );
nand ( n233337 , n233335 , n233336 );
xor ( n233338 , n233234 , n233337 );
not ( n233339 , n233138 );
not ( n233340 , n213577 );
or ( n233341 , n233339 , n233340 );
nand ( n233342 , n216336 , n213735 );
nand ( n233343 , n233341 , n233342 );
xor ( n233344 , n233338 , n233343 );
xor ( n233345 , n233234 , n233337 );
and ( n233346 , n233345 , n233343 );
and ( n233347 , n233234 , n233337 );
or ( n233348 , n233346 , n233347 );
not ( n233349 , n220280 );
not ( n233350 , n232872 );
or ( n233351 , n233349 , n233350 );
and ( n233352 , n228216 , n215955 );
not ( n233353 , n228216 );
and ( n233354 , n233353 , n219358 );
or ( n233355 , n233352 , n233354 );
nand ( n233356 , n233355 , n220272 );
nand ( n233357 , n233351 , n233356 );
not ( n233358 , n220985 );
not ( n233359 , n221338 );
not ( n233360 , n230219 );
or ( n233361 , n233359 , n233360 );
not ( n233362 , n230222 );
not ( n233363 , n233362 );
nand ( n233364 , n233363 , n217944 );
nand ( n233365 , n233361 , n233364 );
not ( n233366 , n233365 );
or ( n233367 , n233358 , n233366 );
nand ( n233368 , n232819 , n214717 );
nand ( n233369 , n233367 , n233368 );
xor ( n233370 , n233357 , n233369 );
not ( n233371 , n219731 );
not ( n233372 , n233020 );
or ( n233373 , n233371 , n233372 );
not ( n233374 , n219033 );
not ( n233375 , n227224 );
or ( n233376 , n233374 , n233375 );
nand ( n233377 , n227223 , n219034 );
nand ( n233378 , n233376 , n233377 );
nand ( n233379 , n233378 , n218077 );
nand ( n233380 , n233373 , n233379 );
xor ( n233381 , n233370 , n233380 );
xor ( n233382 , n233357 , n233369 );
and ( n233383 , n233382 , n233380 );
and ( n233384 , n233357 , n233369 );
or ( n233385 , n233383 , n233384 );
xor ( n233386 , n233287 , n233323 );
not ( n233387 , n232927 );
not ( n233388 , n228858 );
or ( n233389 , n233387 , n233388 );
not ( n233390 , n218514 );
not ( n233391 , n228847 );
or ( n233392 , n233390 , n233391 );
nand ( n233393 , n230851 , n216170 );
nand ( n233394 , n233392 , n233393 );
nand ( n233395 , n233394 , n228867 );
nand ( n233396 , n233389 , n233395 );
not ( n233397 , n232938 );
or ( n233398 , n231994 , n233397 );
not ( n233399 , n229759 );
and ( n233400 , n216208 , n233399 );
not ( n233401 , n216208 );
and ( n233402 , n233401 , n229761 );
nor ( n233403 , n233400 , n233402 );
or ( n233404 , n231476 , n233403 );
nand ( n233405 , n233398 , n233404 );
xor ( n233406 , n233396 , n233405 );
not ( n233407 , n233111 );
not ( n233408 , n232399 );
or ( n233409 , n233407 , n233408 );
not ( n233410 , n214537 );
not ( n233411 , n231753 );
or ( n233412 , n233410 , n233411 );
nand ( n233413 , n230726 , n214899 );
nand ( n233414 , n233412 , n233413 );
nand ( n233415 , n232402 , n233414 );
nand ( n233416 , n233409 , n233415 );
xor ( n233417 , n233406 , n233416 );
xor ( n233418 , n233386 , n233417 );
xor ( n233419 , n233287 , n233323 );
and ( n233420 , n233419 , n233417 );
and ( n233421 , n233287 , n233323 );
or ( n233422 , n233420 , n233421 );
not ( n233423 , n232964 );
not ( n233424 , n229271 );
or ( n233425 , n233423 , n233424 );
not ( n233426 , n216293 );
not ( n233427 , n232493 );
or ( n233428 , n233426 , n233427 );
nand ( n233429 , n232962 , n223658 );
nand ( n233430 , n233428 , n233429 );
nand ( n233431 , n228775 , n233430 );
nand ( n233432 , n233425 , n233431 );
not ( n233433 , n232976 );
not ( n233434 , n226881 );
or ( n233435 , n233433 , n233434 );
not ( n233436 , n222821 );
not ( n233437 , n226650 );
or ( n233438 , n233436 , n233437 );
nand ( n233439 , n227245 , n218980 );
nand ( n233440 , n233438 , n233439 );
nand ( n233441 , n226885 , n233440 );
nand ( n233442 , n233435 , n233441 );
xor ( n233443 , n233432 , n233442 );
not ( n233444 , n232916 );
not ( n233445 , n233444 );
not ( n233446 , n228270 );
not ( n233447 , n233446 );
or ( n233448 , n233445 , n233447 );
not ( n233449 , n219102 );
buf ( n233450 , n227595 );
not ( n233451 , n233450 );
not ( n233452 , n233451 );
or ( n233453 , n233449 , n233452 );
nand ( n233454 , n233450 , n216139 );
nand ( n233455 , n233453 , n233454 );
nand ( n233456 , n227737 , n233455 );
nand ( n233457 , n233448 , n233456 );
xor ( n233458 , n233443 , n233457 );
xor ( n233459 , n233458 , n233238 );
xor ( n233460 , n233459 , n233242 );
xor ( n233461 , n233458 , n233238 );
and ( n233462 , n233461 , n233242 );
and ( n233463 , n233458 , n233238 );
or ( n233464 , n233462 , n233463 );
not ( n233465 , n230725 );
and ( n233466 , n233465 , n214956 );
not ( n233467 , n219076 );
and ( n233468 , n40724 , n219420 );
not ( n233469 , n40724 );
and ( n233470 , n233469 , n221228 );
or ( n233471 , n233468 , n233470 );
not ( n233472 , n233471 );
or ( n233473 , n233467 , n233472 );
nand ( n233474 , n219792 , n232763 );
nand ( n233475 , n233473 , n233474 );
xor ( n233476 , n233466 , n233475 );
not ( n233477 , n218843 );
not ( n233478 , n232413 );
not ( n233479 , n219238 );
or ( n233480 , n233478 , n233479 );
nand ( n233481 , n218590 , n218818 );
nand ( n233482 , n233480 , n233481 );
not ( n233483 , n233482 );
or ( n233484 , n233477 , n233483 );
nand ( n233485 , n233122 , n223665 );
nand ( n233486 , n233484 , n233485 );
xor ( n233487 , n233476 , n233486 );
xor ( n233488 , n233246 , n233487 );
xor ( n233489 , n233488 , n232829 );
xor ( n233490 , n233246 , n233487 );
and ( n233491 , n233490 , n232829 );
and ( n233492 , n233246 , n233487 );
or ( n233493 , n233491 , n233492 );
xor ( n233494 , n233250 , n233254 );
xor ( n233495 , n233494 , n232866 );
xor ( n233496 , n233250 , n233254 );
and ( n233497 , n233496 , n232866 );
and ( n233498 , n233250 , n233254 );
or ( n233499 , n233497 , n233498 );
not ( n233500 , n220067 );
not ( n233501 , n217616 );
not ( n233502 , n40660 );
or ( n233503 , n233501 , n233502 );
nand ( n233504 , n218253 , n207936 );
nand ( n233505 , n233503 , n233504 );
not ( n233506 , n233505 );
or ( n233507 , n233500 , n233506 );
nand ( n233508 , n233008 , n231018 );
nand ( n233509 , n233507 , n233508 );
not ( n233510 , n219836 );
not ( n233511 , n233088 );
or ( n233512 , n233510 , n233511 );
not ( n233513 , n218205 );
not ( n233514 , n219880 );
or ( n233515 , n233513 , n233514 );
nand ( n233516 , n40559 , n218772 );
nand ( n233517 , n233515 , n233516 );
nand ( n233518 , n233517 , n218533 );
nand ( n233519 , n233512 , n233518 );
xor ( n233520 , n233509 , n233519 );
not ( n233521 , n219314 );
not ( n233522 , n219687 );
not ( n233523 , n39879 );
or ( n233524 , n233522 , n233523 );
not ( n233525 , n39877 );
nand ( n233526 , n233525 , n222323 );
nand ( n233527 , n233524 , n233526 );
not ( n233528 , n233527 );
or ( n233529 , n233521 , n233528 );
nand ( n233530 , n233077 , n216204 );
nand ( n233531 , n233529 , n233530 );
xor ( n233532 , n233520 , n233531 );
not ( n233533 , n224171 );
and ( n233534 , n221593 , n217330 );
not ( n233535 , n221593 );
not ( n233536 , n217330 );
and ( n233537 , n233535 , n233536 );
nor ( n233538 , n233534 , n233537 );
not ( n233539 , n233538 );
and ( n233540 , n233533 , n233539 );
not ( n233541 , n232776 );
nor ( n233542 , n233541 , n224163 );
nor ( n233543 , n233540 , n233542 );
buf ( n233544 , n216422 );
not ( n233545 , n233544 );
buf ( n233546 , n226504 );
not ( n233547 , n233546 );
or ( n233548 , n233545 , n233547 );
nand ( n233549 , n226505 , n227602 );
nand ( n233550 , n233548 , n233549 );
not ( n233551 , n233550 );
not ( n233552 , n219501 );
or ( n233553 , n233551 , n233552 );
nand ( n233554 , n233064 , n225478 );
nand ( n233555 , n233553 , n233554 );
xor ( n233556 , n233543 , n233555 );
not ( n233557 , n229974 );
not ( n233558 , n233000 );
or ( n233559 , n233557 , n233558 );
not ( n233560 , n229261 );
not ( n233561 , n223786 );
or ( n233562 , n233560 , n233561 );
nand ( n233563 , n220600 , n229262 );
nand ( n233564 , n233562 , n233563 );
nand ( n233565 , n233564 , n229964 );
nand ( n233566 , n233559 , n233565 );
xor ( n233567 , n233556 , n233566 );
xor ( n233568 , n233532 , n233567 );
not ( n233569 , n215183 );
not ( n233570 , n233097 );
or ( n233571 , n233569 , n233570 );
not ( n233572 , n218990 );
not ( n233573 , n223761 );
or ( n233574 , n233572 , n233573 );
nand ( n233575 , n218994 , n40045 );
nand ( n233576 , n233574 , n233575 );
nand ( n233577 , n233576 , n221933 );
nand ( n233578 , n233571 , n233577 );
not ( n233579 , n220033 );
not ( n233580 , n227912 );
not ( n233581 , n223721 );
or ( n233582 , n233580 , n233581 );
nand ( n233583 , n40485 , n229887 );
nand ( n233584 , n233582 , n233583 );
not ( n233585 , n233584 );
or ( n233586 , n233579 , n233585 );
nand ( n233587 , n233040 , n226943 );
nand ( n233588 , n233586 , n233587 );
xor ( n233589 , n233578 , n233588 );
not ( n233590 , n223949 );
not ( n233591 , n226655 );
not ( n233592 , n222951 );
or ( n233593 , n233591 , n233592 );
nand ( n233594 , n222955 , n227927 );
nand ( n233595 , n233593 , n233594 );
not ( n233596 , n233595 );
or ( n233597 , n233590 , n233596 );
nand ( n233598 , n233048 , n227260 );
nand ( n233599 , n233597 , n233598 );
xor ( n233600 , n233589 , n233599 );
xor ( n233601 , n233568 , n233600 );
xor ( n233602 , n233532 , n233567 );
and ( n233603 , n233602 , n233600 );
and ( n233604 , n233532 , n233567 );
or ( n233605 , n233603 , n233604 );
xor ( n233606 , n232946 , n232882 );
not ( n233607 , n218467 );
not ( n233608 , n232858 );
or ( n233609 , n233607 , n233608 );
not ( n233610 , n217573 );
not ( n233611 , n209864 );
not ( n233612 , n233611 );
or ( n233613 , n233610 , n233612 );
not ( n233614 , n230556 );
nand ( n233615 , n233614 , n219390 );
nand ( n233616 , n233613 , n233615 );
nand ( n233617 , n233616 , n215383 );
nand ( n233618 , n233609 , n233617 );
xor ( n233619 , n232783 , n233618 );
xor ( n233620 , n233619 , n232813 );
xor ( n233621 , n233606 , n233620 );
xor ( n233622 , n232946 , n232882 );
and ( n233623 , n233622 , n233620 );
and ( n233624 , n232946 , n232882 );
or ( n233625 , n233623 , n233624 );
not ( n233626 , n216299 );
not ( n233627 , n232835 );
or ( n233628 , n233626 , n233627 );
not ( n233629 , n216810 );
not ( n233630 , n228165 );
or ( n233631 , n233629 , n233630 );
nand ( n233632 , n230273 , n215289 );
nand ( n233633 , n233631 , n233632 );
nand ( n233634 , n233633 , n220820 );
nand ( n233635 , n233628 , n233634 );
xor ( n233636 , n233160 , n233635 );
xor ( n233637 , n233636 , n233224 );
xor ( n233638 , n233637 , n233381 );
xor ( n233639 , n233638 , n233344 );
xor ( n233640 , n233637 , n233381 );
and ( n233641 , n233640 , n233344 );
and ( n233642 , n233637 , n233381 );
or ( n233643 , n233641 , n233642 );
xor ( n233644 , n232985 , n233418 );
xor ( n233645 , n233644 , n233489 );
xor ( n233646 , n232985 , n233418 );
and ( n233647 , n233646 , n233489 );
and ( n233648 , n232985 , n233418 );
or ( n233649 , n233647 , n233648 );
xor ( n233650 , n233432 , n233442 );
and ( n233651 , n233650 , n233457 );
and ( n233652 , n233432 , n233442 );
or ( n233653 , n233651 , n233652 );
xor ( n233654 , n233131 , n233460 );
xor ( n233655 , n233654 , n232991 );
xor ( n233656 , n233131 , n233460 );
and ( n233657 , n233656 , n232991 );
and ( n233658 , n233131 , n233460 );
or ( n233659 , n233657 , n233658 );
xor ( n233660 , n233030 , n233150 );
xor ( n233661 , n233660 , n233495 );
xor ( n233662 , n233030 , n233150 );
and ( n233663 , n233662 , n233495 );
and ( n233664 , n233030 , n233150 );
or ( n233665 , n233663 , n233664 );
xor ( n233666 , n233601 , n233156 );
xor ( n233667 , n233666 , n233639 );
xor ( n233668 , n233601 , n233156 );
and ( n233669 , n233668 , n233639 );
and ( n233670 , n233601 , n233156 );
or ( n233671 , n233669 , n233670 );
xor ( n233672 , n233621 , n233166 );
xor ( n233673 , n233672 , n233645 );
xor ( n233674 , n233621 , n233166 );
and ( n233675 , n233674 , n233645 );
and ( n233676 , n233621 , n233166 );
or ( n233677 , n233675 , n233676 );
xor ( n233678 , n233178 , n233172 );
xor ( n233679 , n233678 , n233655 );
xor ( n233680 , n233178 , n233172 );
and ( n233681 , n233680 , n233655 );
and ( n233682 , n233178 , n233172 );
or ( n233683 , n233681 , n233682 );
xor ( n233684 , n233661 , n233184 );
xor ( n233685 , n233684 , n233667 );
xor ( n233686 , n233661 , n233184 );
and ( n233687 , n233686 , n233667 );
and ( n233688 , n233661 , n233184 );
or ( n233689 , n233687 , n233688 );
xor ( n233690 , n233190 , n233673 );
xor ( n233691 , n233690 , n233196 );
xor ( n233692 , n233190 , n233673 );
and ( n233693 , n233692 , n233196 );
and ( n233694 , n233190 , n233673 );
or ( n233695 , n233693 , n233694 );
xor ( n233696 , n233679 , n233202 );
xor ( n233697 , n233696 , n233685 );
xor ( n233698 , n233679 , n233202 );
and ( n233699 , n233698 , n233685 );
and ( n233700 , n233679 , n233202 );
or ( n233701 , n233699 , n233700 );
xor ( n233702 , n233208 , n233691 );
xor ( n233703 , n233702 , n233214 );
xor ( n233704 , n233208 , n233691 );
and ( n233705 , n233704 , n233214 );
and ( n233706 , n233208 , n233691 );
or ( n233707 , n233705 , n233706 );
xor ( n233708 , n233697 , n233703 );
xor ( n233709 , n233708 , n233220 );
xor ( n233710 , n233697 , n233703 );
and ( n233711 , n233710 , n233220 );
and ( n233712 , n233697 , n233703 );
or ( n233713 , n233711 , n233712 );
xor ( n233714 , n233396 , n233405 );
and ( n233715 , n233714 , n233416 );
and ( n233716 , n233396 , n233405 );
or ( n233717 , n233715 , n233716 );
xor ( n233718 , n233466 , n233475 );
and ( n233719 , n233718 , n233486 );
and ( n233720 , n233466 , n233475 );
or ( n233721 , n233719 , n233720 );
xor ( n233722 , n233578 , n233588 );
and ( n233723 , n233722 , n233599 );
and ( n233724 , n233578 , n233588 );
or ( n233725 , n233723 , n233724 );
xor ( n233726 , n233543 , n233555 );
and ( n233727 , n233726 , n233566 );
and ( n233728 , n233543 , n233555 );
or ( n233729 , n233727 , n233728 );
xor ( n233730 , n233509 , n233519 );
and ( n233731 , n233730 , n233531 );
and ( n233732 , n233509 , n233519 );
or ( n233733 , n233731 , n233732 );
xor ( n233734 , n232783 , n233618 );
and ( n233735 , n233734 , n232813 );
and ( n233736 , n232783 , n233618 );
or ( n233737 , n233735 , n233736 );
xor ( n233738 , n233160 , n233635 );
and ( n233739 , n233738 , n233224 );
and ( n233740 , n233160 , n233635 );
or ( n233741 , n233739 , n233740 );
or ( n233742 , n213577 , n213498 );
nand ( n233743 , n233742 , n213735 );
not ( n233744 , n233538 );
not ( n233745 , n233744 );
not ( n233746 , n220164 );
or ( n233747 , n233745 , n233746 );
not ( n233748 , n220151 );
not ( n233749 , n220823 );
or ( n233750 , n233748 , n233749 );
nand ( n233751 , n222414 , n219389 );
nand ( n233752 , n233750 , n233751 );
nand ( n233753 , n233752 , n219779 );
nand ( n233754 , n233747 , n233753 );
xor ( n233755 , n233743 , n233754 );
not ( n233756 , n233262 );
not ( n233757 , n221266 );
or ( n233758 , n233756 , n233757 );
not ( n233759 , n231761 );
not ( n233760 , n220925 );
or ( n233761 , n233759 , n233760 );
nand ( n233762 , n231762 , n220905 );
nand ( n233763 , n233761 , n233762 );
nand ( n233764 , n233763 , n221674 );
nand ( n233765 , n233758 , n233764 );
xor ( n233766 , n233755 , n233765 );
xor ( n233767 , n233743 , n233754 );
and ( n233768 , n233767 , n233765 );
and ( n233769 , n233743 , n233754 );
or ( n233770 , n233768 , n233769 );
not ( n233771 , n221387 );
not ( n233772 , n216519 );
not ( n233773 , n221777 );
or ( n233774 , n233772 , n233773 );
nand ( n233775 , n221608 , n217147 );
nand ( n233776 , n233774 , n233775 );
not ( n233777 , n233776 );
or ( n233778 , n233771 , n233777 );
nand ( n233779 , n233272 , n224120 );
nand ( n233780 , n233778 , n233779 );
not ( n233781 , n223244 );
not ( n233782 , n219582 );
not ( n233783 , n222435 );
or ( n233784 , n233782 , n233783 );
nand ( n233785 , n222462 , n217130 );
nand ( n233786 , n233784 , n233785 );
not ( n233787 , n233786 );
or ( n233788 , n233781 , n233787 );
nand ( n233789 , n222886 , n233284 );
nand ( n233790 , n233788 , n233789 );
xor ( n233791 , n233780 , n233790 );
not ( n233792 , n233296 );
not ( n233793 , n223197 );
or ( n233794 , n233792 , n233793 );
and ( n233795 , n41565 , n223156 );
not ( n233796 , n41565 );
and ( n233797 , n233796 , n223182 );
or ( n233798 , n233795 , n233797 );
nand ( n233799 , n233798 , n222768 );
nand ( n233800 , n233794 , n233799 );
xor ( n233801 , n233791 , n233800 );
xor ( n233802 , n233780 , n233790 );
and ( n233803 , n233802 , n233800 );
and ( n233804 , n233780 , n233790 );
or ( n233805 , n233803 , n233804 );
not ( n233806 , n216299 );
not ( n233807 , n233633 );
or ( n233808 , n233806 , n233807 );
not ( n233809 , n216810 );
not ( n233810 , n39286 );
not ( n233811 , n233810 );
or ( n233812 , n233809 , n233811 );
nand ( n233813 , n39286 , n215289 );
nand ( n233814 , n233812 , n233813 );
nand ( n233815 , n233814 , n214694 );
nand ( n233816 , n233808 , n233815 );
xor ( n233817 , n233816 , n233717 );
not ( n233818 , n217023 );
not ( n233819 , n233333 );
or ( n233820 , n233818 , n233819 );
not ( n233821 , n219577 );
not ( n233822 , n229704 );
or ( n233823 , n233821 , n233822 );
nand ( n233824 , n38532 , n218661 );
nand ( n233825 , n233823 , n233824 );
nand ( n233826 , n233825 , n219175 );
nand ( n233827 , n233820 , n233826 );
xor ( n233828 , n233817 , n233827 );
xor ( n233829 , n233816 , n233717 );
and ( n233830 , n233829 , n233827 );
and ( n233831 , n233816 , n233717 );
or ( n233832 , n233830 , n233831 );
not ( n233833 , n220272 );
and ( n233834 , n215955 , n226712 );
not ( n233835 , n215955 );
and ( n233836 , n233835 , n39607 );
or ( n233837 , n233834 , n233836 );
not ( n233838 , n233837 );
or ( n233839 , n233833 , n233838 );
nand ( n233840 , n233355 , n220280 );
nand ( n233841 , n233839 , n233840 );
not ( n233842 , n220985 );
not ( n233843 , n221338 );
not ( n233844 , n209709 );
or ( n233845 , n233843 , n233844 );
not ( n233846 , n209709 );
nand ( n233847 , n233846 , n217944 );
nand ( n233848 , n233845 , n233847 );
not ( n233849 , n233848 );
or ( n233850 , n233842 , n233849 );
nand ( n233851 , n233365 , n231808 );
nand ( n233852 , n233850 , n233851 );
xor ( n233853 , n233841 , n233852 );
not ( n233854 , n222185 );
not ( n233855 , n219033 );
buf ( n233856 , n39713 );
not ( n233857 , n233856 );
not ( n233858 , n233857 );
or ( n233859 , n233855 , n233858 );
nand ( n233860 , n225795 , n219034 );
nand ( n233861 , n233859 , n233860 );
not ( n233862 , n233861 );
or ( n233863 , n233854 , n233862 );
nand ( n233864 , n233378 , n219731 );
nand ( n233865 , n233863 , n233864 );
xor ( n233866 , n233853 , n233865 );
xor ( n233867 , n233841 , n233852 );
and ( n233868 , n233867 , n233865 );
and ( n233869 , n233841 , n233852 );
or ( n233870 , n233868 , n233869 );
or ( n233871 , n231474 , n233403 );
and ( n233872 , n215075 , n229762 );
not ( n233873 , n215075 );
and ( n233874 , n233873 , n231480 );
nor ( n233875 , n233872 , n233874 );
or ( n233876 , n231476 , n233875 );
nand ( n233877 , n233871 , n233876 );
not ( n233878 , n233414 );
buf ( n233879 , n230720 );
not ( n233880 , n233879 );
or ( n233881 , n233878 , n233880 );
not ( n233882 , n216964 );
not ( n233883 , n232404 );
or ( n233884 , n233882 , n233883 );
not ( n233885 , n230722 );
nand ( n233886 , n233885 , n214678 );
nand ( n233887 , n233884 , n233886 );
nand ( n233888 , n233887 , n232402 );
nand ( n233889 , n233881 , n233888 );
xor ( n233890 , n233877 , n233889 );
buf ( n233891 , n233885 );
and ( n233892 , n233891 , n214357 );
xor ( n233893 , n233890 , n233892 );
xor ( n233894 , n233766 , n233893 );
xor ( n233895 , n233894 , n233801 );
xor ( n233896 , n233766 , n233893 );
and ( n233897 , n233896 , n233801 );
and ( n233898 , n233766 , n233893 );
or ( n233899 , n233897 , n233898 );
not ( n233900 , n233440 );
not ( n233901 , n226881 );
or ( n233902 , n233900 , n233901 );
and ( n233903 , n220022 , n226888 );
not ( n233904 , n220022 );
and ( n233905 , n233904 , n226648 );
nor ( n233906 , n233903 , n233905 );
nand ( n233907 , n233906 , n227241 );
nand ( n233908 , n233902 , n233907 );
not ( n233909 , n233455 );
not ( n233910 , n232440 );
or ( n233911 , n233909 , n233910 );
not ( n233912 , n228273 );
not ( n233913 , n219343 );
not ( n233914 , n233451 );
or ( n233915 , n233913 , n233914 );
nand ( n233916 , n233450 , n219348 );
nand ( n233917 , n233915 , n233916 );
nand ( n233918 , n233912 , n233917 );
nand ( n233919 , n233911 , n233918 );
xor ( n233920 , n233908 , n233919 );
not ( n233921 , n233394 );
not ( n233922 , n228860 );
or ( n233923 , n233921 , n233922 );
not ( n233924 , n216934 );
buf ( n233925 , n231943 );
not ( n233926 , n233925 );
not ( n233927 , n233926 );
or ( n233928 , n233924 , n233927 );
not ( n233929 , n228847 );
nand ( n233930 , n233929 , n216940 );
nand ( n233931 , n233928 , n233930 );
nand ( n233932 , n228868 , n233931 );
nand ( n233933 , n233923 , n233932 );
xor ( n233934 , n233920 , n233933 );
not ( n233935 , n233311 );
not ( n233936 , n224086 );
or ( n233937 , n233935 , n233936 );
not ( n233938 , n225768 );
not ( n233939 , n224095 );
or ( n233940 , n233938 , n233939 );
nand ( n233941 , n224096 , n225769 );
nand ( n233942 , n233940 , n233941 );
nand ( n233943 , n224090 , n233942 );
nand ( n233944 , n233937 , n233943 );
not ( n233945 , n233320 );
not ( n233946 , n233945 );
not ( n233947 , n233315 );
or ( n233948 , n233946 , n233947 );
not ( n233949 , n214837 );
not ( n233950 , n226747 );
or ( n233951 , n233949 , n233950 );
buf ( n233952 , n224944 );
nand ( n233953 , n233952 , n231913 );
nand ( n233954 , n233951 , n233953 );
nand ( n233955 , n226745 , n233954 );
nand ( n233956 , n233948 , n233955 );
xor ( n233957 , n233944 , n233956 );
not ( n233958 , n233430 );
not ( n233959 , n230390 );
or ( n233960 , n233958 , n233959 );
not ( n233961 , n224037 );
buf ( n233962 , n226276 );
not ( n233963 , n233962 );
or ( n233964 , n233961 , n233963 );
not ( n233965 , n229807 );
nand ( n233966 , n233965 , n224041 );
nand ( n233967 , n233964 , n233966 );
nand ( n233968 , n228775 , n233967 );
nand ( n233969 , n233960 , n233968 );
xor ( n233970 , n233957 , n233969 );
xor ( n233971 , n233934 , n233970 );
xor ( n233972 , n233971 , n233721 );
xor ( n233973 , n233934 , n233970 );
and ( n233974 , n233973 , n233721 );
and ( n233975 , n233934 , n233970 );
or ( n233976 , n233974 , n233975 );
xor ( n233977 , n233725 , n233729 );
xor ( n233978 , n233977 , n233348 );
xor ( n233979 , n233725 , n233729 );
and ( n233980 , n233979 , n233348 );
and ( n233981 , n233725 , n233729 );
or ( n233982 , n233980 , n233981 );
xor ( n233983 , n233733 , n233737 );
xor ( n233984 , n233983 , n233741 );
xor ( n233985 , n233733 , n233737 );
and ( n233986 , n233985 , n233741 );
and ( n233987 , n233733 , n233737 );
or ( n233988 , n233986 , n233987 );
not ( n233989 , n225478 );
not ( n233990 , n233550 );
or ( n233991 , n233989 , n233990 );
not ( n233992 , n229387 );
not ( n233993 , n40181 );
or ( n233994 , n233992 , n233993 );
nand ( n233995 , n221716 , n227602 );
nand ( n233996 , n233994 , n233995 );
nand ( n233997 , n233996 , n228237 );
nand ( n233998 , n233991 , n233997 );
not ( n233999 , n229964 );
buf ( n234000 , n220050 );
or ( n234001 , n234000 , n226911 );
nand ( n234002 , n220970 , n234000 );
nand ( n234003 , n234001 , n234002 );
not ( n234004 , n234003 );
or ( n234005 , n233999 , n234004 );
buf ( n234006 , n219368 );
nand ( n234007 , n233564 , n234006 );
nand ( n234008 , n234005 , n234007 );
xor ( n234009 , n233998 , n234008 );
not ( n234010 , n220067 );
not ( n234011 , n217616 );
not ( n234012 , n226921 );
or ( n234013 , n234011 , n234012 );
not ( n234014 , n230966 );
not ( n234015 , n217616 );
nand ( n234016 , n234014 , n234015 );
nand ( n234017 , n234013 , n234016 );
not ( n234018 , n234017 );
or ( n234019 , n234010 , n234018 );
nand ( n234020 , n233505 , n231018 );
nand ( n234021 , n234019 , n234020 );
xor ( n234022 , n234009 , n234021 );
xor ( n234023 , n233385 , n234022 );
not ( n234024 , n219076 );
not ( n234025 , n221228 );
not ( n234026 , n218268 );
or ( n234027 , n234025 , n234026 );
nand ( n234028 , n40710 , n219423 );
nand ( n234029 , n234027 , n234028 );
not ( n234030 , n234029 );
or ( n234031 , n234024 , n234030 );
nand ( n234032 , n233471 , n219792 );
nand ( n234033 , n234031 , n234032 );
not ( n234034 , n233543 );
xor ( n234035 , n234033 , n234034 );
not ( n234036 , n221933 );
not ( n234037 , n226484 );
not ( n234038 , n39996 );
or ( n234039 , n234037 , n234038 );
nand ( n234040 , n225111 , n221938 );
nand ( n234041 , n234039 , n234040 );
not ( n234042 , n234041 );
or ( n234043 , n234036 , n234042 );
not ( n234044 , n233576 );
not ( n234045 , n215183 );
or ( n234046 , n234044 , n234045 );
nand ( n234047 , n234043 , n234046 );
xor ( n234048 , n234035 , n234047 );
xor ( n234049 , n234023 , n234048 );
xor ( n234050 , n233385 , n234022 );
and ( n234051 , n234050 , n234048 );
and ( n234052 , n233385 , n234022 );
or ( n234053 , n234051 , n234052 );
not ( n234054 , n218843 );
and ( n234055 , n219532 , n232413 );
not ( n234056 , n219532 );
and ( n234057 , n234056 , n218818 );
or ( n234058 , n234055 , n234057 );
not ( n234059 , n234058 );
or ( n234060 , n234054 , n234059 );
nand ( n234061 , n219449 , n233482 );
nand ( n234062 , n234060 , n234061 );
not ( n234063 , n220414 );
not ( n234064 , n233584 );
or ( n234065 , n234063 , n234064 );
not ( n234066 , n227912 );
not ( n234067 , n40546 );
or ( n234068 , n234066 , n234067 );
nand ( n234069 , n40547 , n229887 );
nand ( n234070 , n234068 , n234069 );
nand ( n234071 , n234070 , n226287 );
nand ( n234072 , n234065 , n234071 );
xor ( n234073 , n234062 , n234072 );
not ( n234074 , n223949 );
not ( n234075 , n226655 );
not ( n234076 , n227004 );
or ( n234077 , n234075 , n234076 );
not ( n234078 , n223368 );
nand ( n234079 , n234078 , n227927 );
nand ( n234080 , n234077 , n234079 );
not ( n234081 , n234080 );
or ( n234082 , n234074 , n234081 );
nand ( n234083 , n233595 , n227260 );
nand ( n234084 , n234082 , n234083 );
xor ( n234085 , n234073 , n234084 );
xor ( n234086 , n234085 , n233422 );
xor ( n234087 , n234086 , n233866 );
xor ( n234088 , n234085 , n233422 );
and ( n234089 , n234088 , n233866 );
and ( n234090 , n234085 , n233422 );
or ( n234091 , n234089 , n234090 );
not ( n234092 , n220941 );
not ( n234093 , n217573 );
not ( n234094 , n209962 );
not ( n234095 , n234094 );
or ( n234096 , n234093 , n234095 );
nand ( n234097 , n231104 , n219390 );
nand ( n234098 , n234096 , n234097 );
not ( n234099 , n234098 );
or ( n234100 , n234092 , n234099 );
nand ( n234101 , n233616 , n218467 );
nand ( n234102 , n234100 , n234101 );
xor ( n234103 , n234102 , n233327 );
xor ( n234104 , n234103 , n233653 );
xor ( n234105 , n233828 , n234104 );
not ( n234106 , n218533 );
not ( n234107 , n218205 );
buf ( n234108 , n221687 );
not ( n234109 , n234108 );
or ( n234110 , n234107 , n234109 );
nand ( n234111 , n40625 , n220091 );
nand ( n234112 , n234110 , n234111 );
not ( n234113 , n234112 );
or ( n234114 , n234106 , n234113 );
nand ( n234115 , n233517 , n219461 );
nand ( n234116 , n234114 , n234115 );
not ( n234117 , n224624 );
not ( n234118 , n233527 );
or ( n234119 , n234117 , n234118 );
not ( n234120 , n219687 );
not ( n234121 , n39927 );
or ( n234122 , n234120 , n234121 );
nand ( n234123 , n233018 , n222323 );
nand ( n234124 , n234122 , n234123 );
nand ( n234125 , n234124 , n219314 );
nand ( n234126 , n234119 , n234125 );
xor ( n234127 , n234116 , n234126 );
xor ( n234128 , n234127 , n233291 );
xor ( n234129 , n234105 , n234128 );
xor ( n234130 , n233828 , n234104 );
and ( n234131 , n234130 , n234128 );
and ( n234132 , n233828 , n234104 );
or ( n234133 , n234131 , n234132 );
xor ( n234134 , n233972 , n233464 );
xor ( n234135 , n234134 , n233895 );
xor ( n234136 , n233972 , n233464 );
and ( n234137 , n234136 , n233895 );
and ( n234138 , n233972 , n233464 );
or ( n234139 , n234137 , n234138 );
xor ( n234140 , n233944 , n233956 );
and ( n234141 , n234140 , n233969 );
and ( n234142 , n233944 , n233956 );
or ( n234143 , n234141 , n234142 );
xor ( n234144 , n233978 , n233605 );
xor ( n234145 , n234144 , n233493 );
xor ( n234146 , n233978 , n233605 );
and ( n234147 , n234146 , n233493 );
and ( n234148 , n233978 , n233605 );
or ( n234149 , n234147 , n234148 );
xor ( n234150 , n233499 , n233984 );
xor ( n234151 , n234150 , n233643 );
xor ( n234152 , n233499 , n233984 );
and ( n234153 , n234152 , n233643 );
and ( n234154 , n233499 , n233984 );
or ( n234155 , n234153 , n234154 );
xor ( n234156 , n233625 , n234049 );
xor ( n234157 , n234156 , n234129 );
xor ( n234158 , n233625 , n234049 );
and ( n234159 , n234158 , n234129 );
and ( n234160 , n233625 , n234049 );
or ( n234161 , n234159 , n234160 );
xor ( n234162 , n234087 , n233649 );
xor ( n234163 , n234162 , n233659 );
xor ( n234164 , n234087 , n233649 );
and ( n234165 , n234164 , n233659 );
and ( n234166 , n234087 , n233649 );
or ( n234167 , n234165 , n234166 );
xor ( n234168 , n234135 , n233665 );
xor ( n234169 , n234168 , n234145 );
xor ( n234170 , n234135 , n233665 );
and ( n234171 , n234170 , n234145 );
and ( n234172 , n234135 , n233665 );
or ( n234173 , n234171 , n234172 );
xor ( n234174 , n234157 , n233671 );
xor ( n234175 , n234174 , n234151 );
xor ( n234176 , n234157 , n233671 );
and ( n234177 , n234176 , n234151 );
and ( n234178 , n234157 , n233671 );
or ( n234179 , n234177 , n234178 );
xor ( n234180 , n233677 , n233683 );
xor ( n234181 , n234180 , n234163 );
xor ( n234182 , n233677 , n233683 );
and ( n234183 , n234182 , n234163 );
and ( n234184 , n233677 , n233683 );
or ( n234185 , n234183 , n234184 );
xor ( n234186 , n234169 , n233689 );
xor ( n234187 , n234186 , n234175 );
xor ( n234188 , n234169 , n233689 );
and ( n234189 , n234188 , n234175 );
and ( n234190 , n234169 , n233689 );
or ( n234191 , n234189 , n234190 );
xor ( n234192 , n233695 , n234181 );
xor ( n234193 , n234192 , n233701 );
xor ( n234194 , n233695 , n234181 );
and ( n234195 , n234194 , n233701 );
and ( n234196 , n233695 , n234181 );
or ( n234197 , n234195 , n234196 );
xor ( n234198 , n234187 , n234193 );
xor ( n234199 , n234198 , n233707 );
xor ( n234200 , n234187 , n234193 );
and ( n234201 , n234200 , n233707 );
and ( n234202 , n234187 , n234193 );
or ( n234203 , n234201 , n234202 );
xor ( n234204 , n233908 , n233919 );
and ( n234205 , n234204 , n233933 );
and ( n234206 , n233908 , n233919 );
or ( n234207 , n234205 , n234206 );
xor ( n234208 , n233877 , n233889 );
and ( n234209 , n234208 , n233892 );
and ( n234210 , n233877 , n233889 );
or ( n234211 , n234209 , n234210 );
xor ( n234212 , n234033 , n234034 );
and ( n234213 , n234212 , n234047 );
and ( n234214 , n234033 , n234034 );
or ( n234215 , n234213 , n234214 );
xor ( n234216 , n234062 , n234072 );
and ( n234217 , n234216 , n234084 );
and ( n234218 , n234062 , n234072 );
or ( n234219 , n234217 , n234218 );
xor ( n234220 , n233998 , n234008 );
and ( n234221 , n234220 , n234021 );
and ( n234222 , n233998 , n234008 );
or ( n234223 , n234221 , n234222 );
xor ( n234224 , n234116 , n234126 );
and ( n234225 , n234224 , n233291 );
and ( n234226 , n234116 , n234126 );
or ( n234227 , n234225 , n234226 );
xor ( n234228 , n234102 , n233327 );
and ( n234229 , n234228 , n233653 );
and ( n234230 , n234102 , n233327 );
or ( n234231 , n234229 , n234230 );
not ( n234232 , n233786 );
not ( n234233 , n222886 );
or ( n234234 , n234232 , n234233 );
and ( n234235 , n219902 , n222435 );
not ( n234236 , n219902 );
and ( n234237 , n234236 , n222462 );
or ( n234238 , n234235 , n234237 );
nand ( n234239 , n234238 , n222158 );
nand ( n234240 , n234234 , n234239 );
not ( n234241 , n233798 );
not ( n234242 , n223591 );
or ( n234243 , n234241 , n234242 );
not ( n234244 , n215796 );
not ( n234245 , n223595 );
or ( n234246 , n234244 , n234245 );
nand ( n234247 , n223201 , n217394 );
nand ( n234248 , n234246 , n234247 );
nand ( n234249 , n234248 , n227294 );
nand ( n234250 , n234243 , n234249 );
xor ( n234251 , n234240 , n234250 );
not ( n234252 , n233942 );
not ( n234253 , n224087 );
or ( n234254 , n234252 , n234253 );
not ( n234255 , n230369 );
buf ( n234256 , n215428 );
not ( n234257 , n234256 );
not ( n234258 , n234257 );
or ( n234259 , n234255 , n234258 );
nand ( n234260 , n224096 , n234256 );
nand ( n234261 , n234259 , n234260 );
nand ( n234262 , n224090 , n234261 );
nand ( n234263 , n234254 , n234262 );
xor ( n234264 , n234251 , n234263 );
xor ( n234265 , n234240 , n234250 );
and ( n234266 , n234265 , n234263 );
and ( n234267 , n234240 , n234250 );
or ( n234268 , n234266 , n234267 );
not ( n234269 , n233954 );
not ( n234270 , n233315 );
or ( n234271 , n234269 , n234270 );
not ( n234272 , n219689 );
not ( n234273 , n233952 );
not ( n234274 , n234273 );
or ( n234275 , n234272 , n234274 );
nand ( n234276 , n232485 , n208726 );
nand ( n234277 , n234275 , n234276 );
nand ( n234278 , n224941 , n234277 );
nand ( n234279 , n234271 , n234278 );
not ( n234280 , n233763 );
not ( n234281 , n221266 );
or ( n234282 , n234280 , n234281 );
and ( n234283 , n220925 , n217330 );
not ( n234284 , n220925 );
and ( n234285 , n234284 , n233536 );
or ( n234286 , n234283 , n234285 );
nand ( n234287 , n234286 , n220930 );
nand ( n234288 , n234282 , n234287 );
xor ( n234289 , n234279 , n234288 );
not ( n234290 , n226881 );
not ( n234291 , n233906 );
or ( n234292 , n234290 , n234291 );
buf ( n234293 , n232431 );
and ( n234294 , n234293 , n216293 );
not ( n234295 , n234293 );
and ( n234296 , n234295 , n223658 );
nor ( n234297 , n234294 , n234296 );
or ( n234298 , n226884 , n234297 );
nand ( n234299 , n234292 , n234298 );
xor ( n234300 , n234289 , n234299 );
xor ( n234301 , n234279 , n234288 );
and ( n234302 , n234301 , n234299 );
and ( n234303 , n234279 , n234288 );
or ( n234304 , n234302 , n234303 );
not ( n234305 , n219353 );
not ( n234306 , n215955 );
not ( n234307 , n232316 );
or ( n234308 , n234306 , n234307 );
nand ( n234309 , n39089 , n216989 );
nand ( n234310 , n234308 , n234309 );
not ( n234311 , n234310 );
or ( n234312 , n234305 , n234311 );
nand ( n234313 , n233837 , n220280 );
nand ( n234314 , n234312 , n234313 );
not ( n234315 , n214086 );
not ( n234316 , n234098 );
or ( n234317 , n234315 , n234316 );
nand ( n234318 , n215137 , n217573 );
nand ( n234319 , n234317 , n234318 );
xor ( n234320 , n234314 , n234319 );
not ( n234321 , n219731 );
not ( n234322 , n233861 );
or ( n234323 , n234321 , n234322 );
buf ( n234324 , n226243 );
and ( n234325 , n219033 , n234324 );
not ( n234326 , n219033 );
and ( n234327 , n234326 , n228215 );
or ( n234328 , n234325 , n234327 );
nand ( n234329 , n222185 , n234328 );
nand ( n234330 , n234323 , n234329 );
xor ( n234331 , n234320 , n234330 );
xor ( n234332 , n234314 , n234319 );
and ( n234333 , n234332 , n234330 );
and ( n234334 , n234314 , n234319 );
or ( n234335 , n234333 , n234334 );
not ( n234336 , n214694 );
and ( n234337 , n216810 , n233362 );
not ( n234338 , n216810 );
and ( n234339 , n234338 , n233363 );
or ( n234340 , n234337 , n234339 );
not ( n234341 , n234340 );
or ( n234342 , n234336 , n234341 );
nand ( n234343 , n233814 , n216299 );
nand ( n234344 , n234342 , n234343 );
not ( n234345 , n219314 );
not ( n234346 , n219687 );
not ( n234347 , n39812 );
not ( n234348 , n234347 );
or ( n234349 , n234346 , n234348 );
buf ( n234350 , n225357 );
not ( n234351 , n234350 );
nand ( n234352 , n234351 , n222323 );
nand ( n234353 , n234349 , n234352 );
not ( n234354 , n234353 );
or ( n234355 , n234345 , n234354 );
nand ( n234356 , n234124 , n224624 );
nand ( n234357 , n234355 , n234356 );
xor ( n234358 , n234344 , n234357 );
not ( n234359 , n233887 );
not ( n234360 , n232399 );
or ( n234361 , n234359 , n234360 );
not ( n234362 , n216208 );
not ( n234363 , n230722 );
or ( n234364 , n234362 , n234363 );
nand ( n234365 , n231232 , n216207 );
nand ( n234366 , n234364 , n234365 );
nand ( n234367 , n234366 , n232402 );
nand ( n234368 , n234361 , n234367 );
not ( n234369 , n233875 );
not ( n234370 , n234369 );
buf ( n234371 , n229773 );
not ( n234372 , n234371 );
or ( n234373 , n234370 , n234372 );
and ( n234374 , n233399 , n218514 );
and ( n234375 , n229761 , n216170 );
nor ( n234376 , n234374 , n234375 );
not ( n234377 , n234376 );
not ( n234378 , n229776 );
nand ( n234379 , n234377 , n234378 );
nand ( n234380 , n234373 , n234379 );
xor ( n234381 , n234368 , n234380 );
buf ( n234382 , n231232 );
and ( n234383 , n234382 , n214537 );
xor ( n234384 , n234381 , n234383 );
xor ( n234385 , n234358 , n234384 );
xor ( n234386 , n234344 , n234357 );
and ( n234387 , n234386 , n234384 );
and ( n234388 , n234344 , n234357 );
or ( n234389 , n234387 , n234388 );
not ( n234390 , n233917 );
not ( n234391 , n232440 );
or ( n234392 , n234390 , n234391 );
not ( n234393 , n221921 );
not ( n234394 , n233450 );
not ( n234395 , n234394 );
or ( n234396 , n234393 , n234395 );
nand ( n234397 , n233450 , n218980 );
nand ( n234398 , n234396 , n234397 );
nand ( n234399 , n227737 , n234398 );
nand ( n234400 , n234392 , n234399 );
not ( n234401 , n233931 );
not ( n234402 , n231421 );
or ( n234403 , n234401 , n234402 );
not ( n234404 , n232454 );
and ( n234405 , n219102 , n228847 );
not ( n234406 , n219102 );
and ( n234407 , n234406 , n233925 );
or ( n234408 , n234405 , n234407 );
nand ( n234409 , n234404 , n234408 );
nand ( n234410 , n234403 , n234409 );
xor ( n234411 , n234400 , n234410 );
not ( n234412 , n233967 );
not ( n234413 , n232956 );
or ( n234414 , n234412 , n234413 );
not ( n234415 , n224492 );
not ( n234416 , n233962 );
or ( n234417 , n234415 , n234416 );
nand ( n234418 , n232494 , n225505 );
nand ( n234419 , n234417 , n234418 );
nand ( n234420 , n228775 , n234419 );
nand ( n234421 , n234414 , n234420 );
xor ( n234422 , n234411 , n234421 );
xor ( n234423 , n234264 , n234422 );
xor ( n234424 , n234423 , n234300 );
xor ( n234425 , n234264 , n234422 );
and ( n234426 , n234425 , n234300 );
and ( n234427 , n234264 , n234422 );
or ( n234428 , n234426 , n234427 );
xor ( n234429 , n234215 , n234219 );
xor ( n234430 , n234429 , n234223 );
xor ( n234431 , n234215 , n234219 );
and ( n234432 , n234431 , n234223 );
and ( n234433 , n234215 , n234219 );
or ( n234434 , n234432 , n234433 );
xor ( n234435 , n233870 , n234227 );
xor ( n234436 , n234435 , n234231 );
xor ( n234437 , n233870 , n234227 );
and ( n234438 , n234437 , n234231 );
and ( n234439 , n233870 , n234227 );
or ( n234440 , n234438 , n234439 );
not ( n234441 , n229964 );
not ( n234442 , n229261 );
not ( n234443 , n233546 );
or ( n234444 , n234442 , n234443 );
nand ( n234445 , n40397 , n234000 );
nand ( n234446 , n234444 , n234445 );
not ( n234447 , n234446 );
or ( n234448 , n234441 , n234447 );
not ( n234449 , n234000 );
not ( n234450 , n234449 );
not ( n234451 , n40258 );
or ( n234452 , n234450 , n234451 );
nand ( n234453 , n234452 , n234002 );
nand ( n234454 , n234453 , n234006 );
nand ( n234455 , n234448 , n234454 );
not ( n234456 , n231018 );
not ( n234457 , n234017 );
or ( n234458 , n234456 , n234457 );
not ( n234459 , n217616 );
not ( n234460 , n220599 );
or ( n234461 , n234459 , n234460 );
nand ( n234462 , n221956 , n234015 );
nand ( n234463 , n234461 , n234462 );
nand ( n234464 , n234463 , n220067 );
nand ( n234465 , n234458 , n234464 );
xor ( n234466 , n234455 , n234465 );
not ( n234467 , n219461 );
not ( n234468 , n234112 );
or ( n234469 , n234467 , n234468 );
not ( n234470 , n218775 );
not ( n234471 , n220581 );
or ( n234472 , n234470 , n234471 );
nand ( n234473 , n207936 , n218209 );
nand ( n234474 , n234472 , n234473 );
nand ( n234475 , n234474 , n218232 );
nand ( n234476 , n234469 , n234475 );
xor ( n234477 , n234466 , n234476 );
xor ( n234478 , n233832 , n234477 );
not ( n234479 , n219779 );
not ( n234480 , n220290 );
not ( n234481 , n208002 );
or ( n234482 , n234480 , n234481 );
or ( n234483 , n208002 , n220499 );
nand ( n234484 , n234482 , n234483 );
not ( n234485 , n234484 );
or ( n234486 , n234479 , n234485 );
not ( n234487 , n224163 );
nand ( n234488 , n234487 , n233752 );
nand ( n234489 , n234486 , n234488 );
not ( n234490 , n219076 );
not ( n234491 , n221228 );
not ( n234492 , n226486 );
or ( n234493 , n234491 , n234492 );
nand ( n234494 , n226489 , n219420 );
nand ( n234495 , n234493 , n234494 );
not ( n234496 , n234495 );
or ( n234497 , n234490 , n234496 );
nand ( n234498 , n234029 , n220507 );
nand ( n234499 , n234497 , n234498 );
xor ( n234500 , n234489 , n234499 );
not ( n234501 , n226287 );
not ( n234502 , n227912 );
buf ( n234503 , n223764 );
not ( n234504 , n234503 );
or ( n234505 , n234502 , n234504 );
buf ( n234506 , n40045 );
nand ( n234507 , n234506 , n220038 );
nand ( n234508 , n234505 , n234507 );
not ( n234509 , n234508 );
or ( n234510 , n234501 , n234509 );
nand ( n234511 , n234070 , n220414 );
nand ( n234512 , n234510 , n234511 );
xor ( n234513 , n234500 , n234512 );
xor ( n234514 , n234478 , n234513 );
xor ( n234515 , n233832 , n234477 );
and ( n234516 , n234515 , n234513 );
and ( n234517 , n233832 , n234477 );
or ( n234518 , n234516 , n234517 );
not ( n234519 , n223949 );
not ( n234520 , n226655 );
not ( n234521 , n223717 );
or ( n234522 , n234520 , n234521 );
nand ( n234523 , n223722 , n227927 );
nand ( n234524 , n234522 , n234523 );
not ( n234525 , n234524 );
or ( n234526 , n234519 , n234525 );
nand ( n234527 , n234080 , n227260 );
nand ( n234528 , n234526 , n234527 );
not ( n234529 , n228237 );
not ( n234530 , n216422 );
not ( n234531 , n222951 );
or ( n234532 , n234530 , n234531 );
nand ( n234533 , n223751 , n227602 );
nand ( n234534 , n234532 , n234533 );
not ( n234535 , n234534 );
or ( n234536 , n234529 , n234535 );
nand ( n234537 , n233996 , n225478 );
nand ( n234538 , n234536 , n234537 );
xor ( n234539 , n234528 , n234538 );
not ( n234540 , n233776 );
or ( n234541 , n222471 , n234540 );
and ( n234542 , n230171 , n226388 );
not ( n234543 , n230171 );
and ( n234544 , n234543 , n221632 );
nor ( n234545 , n234542 , n234544 );
or ( n234546 , n221636 , n234545 );
nand ( n234547 , n234541 , n234546 );
not ( n234548 , n234547 );
xor ( n234549 , n234539 , n234548 );
not ( n234550 , n222376 );
not ( n234551 , n220126 );
not ( n234552 , n227448 );
or ( n234553 , n234551 , n234552 );
not ( n234554 , n219880 );
nand ( n234555 , n234554 , n221238 );
nand ( n234556 , n234553 , n234555 );
not ( n234557 , n234556 );
or ( n234558 , n234550 , n234557 );
nand ( n234559 , n234058 , n223665 );
nand ( n234560 , n234558 , n234559 );
not ( n234561 , n221933 );
not ( n234562 , n221935 );
not ( n234563 , n227477 );
or ( n234564 , n234562 , n234563 );
not ( n234565 , n230280 );
nand ( n234566 , n234565 , n222333 );
nand ( n234567 , n234564 , n234566 );
not ( n234568 , n234567 );
or ( n234569 , n234561 , n234568 );
nand ( n234570 , n234041 , n219332 );
nand ( n234571 , n234569 , n234570 );
xor ( n234572 , n234560 , n234571 );
xor ( n234573 , n234572 , n233770 );
xor ( n234574 , n234549 , n234573 );
not ( n234575 , n231808 );
not ( n234576 , n233848 );
or ( n234577 , n234575 , n234576 );
not ( n234578 , n221338 );
not ( n234579 , n233614 );
not ( n234580 , n234579 );
or ( n234581 , n234578 , n234580 );
nand ( n234582 , n209865 , n217944 );
nand ( n234583 , n234581 , n234582 );
nand ( n234584 , n234583 , n220985 );
nand ( n234585 , n234577 , n234584 );
xor ( n234586 , n233805 , n234585 );
xor ( n234587 , n234586 , n234143 );
xor ( n234588 , n234574 , n234587 );
xor ( n234589 , n234549 , n234573 );
and ( n234590 , n234589 , n234587 );
and ( n234591 , n234549 , n234573 );
or ( n234592 , n234590 , n234591 );
not ( n234593 , n219175 );
not ( n234594 , n219577 );
not ( n234595 , n39364 );
or ( n234596 , n234594 , n234595 );
nand ( n234597 , n39365 , n218661 );
nand ( n234598 , n234596 , n234597 );
not ( n234599 , n234598 );
or ( n234600 , n234593 , n234599 );
nand ( n234601 , n233825 , n217023 );
nand ( n234602 , n234600 , n234601 );
xor ( n234603 , n234207 , n234602 );
xor ( n234604 , n234603 , n234211 );
xor ( n234605 , n234604 , n233899 );
xor ( n234606 , n234605 , n234331 );
xor ( n234607 , n234604 , n233899 );
and ( n234608 , n234607 , n234331 );
and ( n234609 , n234604 , n233899 );
or ( n234610 , n234608 , n234609 );
xor ( n234611 , n234385 , n233976 );
xor ( n234612 , n234611 , n234424 );
xor ( n234613 , n234385 , n233976 );
and ( n234614 , n234613 , n234424 );
and ( n234615 , n234385 , n233976 );
or ( n234616 , n234614 , n234615 );
xor ( n234617 , n234430 , n233982 );
xor ( n234618 , n234617 , n233988 );
xor ( n234619 , n234430 , n233982 );
and ( n234620 , n234619 , n233988 );
and ( n234621 , n234430 , n233982 );
or ( n234622 , n234620 , n234621 );
xor ( n234623 , n234400 , n234410 );
and ( n234624 , n234623 , n234421 );
and ( n234625 , n234400 , n234410 );
or ( n234626 , n234624 , n234625 );
xor ( n234627 , n234053 , n234514 );
xor ( n234628 , n234627 , n234436 );
xor ( n234629 , n234053 , n234514 );
and ( n234630 , n234629 , n234436 );
and ( n234631 , n234053 , n234514 );
or ( n234632 , n234630 , n234631 );
xor ( n234633 , n234091 , n234133 );
xor ( n234634 , n234633 , n234139 );
xor ( n234635 , n234091 , n234133 );
and ( n234636 , n234635 , n234139 );
and ( n234637 , n234091 , n234133 );
or ( n234638 , n234636 , n234637 );
xor ( n234639 , n234588 , n234606 );
xor ( n234640 , n234639 , n234612 );
xor ( n234641 , n234588 , n234606 );
and ( n234642 , n234641 , n234612 );
and ( n234643 , n234588 , n234606 );
or ( n234644 , n234642 , n234643 );
xor ( n234645 , n234149 , n234155 );
xor ( n234646 , n234645 , n234618 );
xor ( n234647 , n234149 , n234155 );
and ( n234648 , n234647 , n234618 );
and ( n234649 , n234149 , n234155 );
or ( n234650 , n234648 , n234649 );
xor ( n234651 , n234161 , n234628 );
xor ( n234652 , n234651 , n234634 );
xor ( n234653 , n234161 , n234628 );
and ( n234654 , n234653 , n234634 );
and ( n234655 , n234161 , n234628 );
or ( n234656 , n234654 , n234655 );
xor ( n234657 , n234167 , n234640 );
xor ( n234658 , n234657 , n234173 );
xor ( n234659 , n234167 , n234640 );
and ( n234660 , n234659 , n234173 );
and ( n234661 , n234167 , n234640 );
or ( n234662 , n234660 , n234661 );
xor ( n234663 , n234646 , n234179 );
xor ( n234664 , n234663 , n234652 );
xor ( n234665 , n234646 , n234179 );
and ( n234666 , n234665 , n234652 );
and ( n234667 , n234646 , n234179 );
or ( n234668 , n234666 , n234667 );
xor ( n234669 , n234185 , n234658 );
xor ( n234670 , n234669 , n234664 );
xor ( n234671 , n234185 , n234658 );
and ( n234672 , n234671 , n234664 );
and ( n234673 , n234185 , n234658 );
or ( n234674 , n234672 , n234673 );
xor ( n234675 , n234191 , n234670 );
xor ( n234676 , n234675 , n234197 );
xor ( n234677 , n234191 , n234670 );
and ( n234678 , n234677 , n234197 );
and ( n234679 , n234191 , n234670 );
or ( n234680 , n234678 , n234679 );
xor ( n234681 , n234368 , n234380 );
and ( n234682 , n234681 , n234383 );
and ( n234683 , n234368 , n234380 );
or ( n234684 , n234682 , n234683 );
xor ( n234685 , n234489 , n234499 );
and ( n234686 , n234685 , n234512 );
and ( n234687 , n234489 , n234499 );
or ( n234688 , n234686 , n234687 );
xor ( n234689 , n234528 , n234538 );
and ( n234690 , n234689 , n234548 );
and ( n234691 , n234528 , n234538 );
or ( n234692 , n234690 , n234691 );
xor ( n234693 , n234455 , n234465 );
and ( n234694 , n234693 , n234476 );
and ( n234695 , n234455 , n234465 );
or ( n234696 , n234694 , n234695 );
xor ( n234697 , n234560 , n234571 );
and ( n234698 , n234697 , n233770 );
and ( n234699 , n234560 , n234571 );
or ( n234700 , n234698 , n234699 );
xor ( n234701 , n233805 , n234585 );
and ( n234702 , n234701 , n234143 );
and ( n234703 , n233805 , n234585 );
or ( n234704 , n234702 , n234703 );
xor ( n234705 , n234207 , n234602 );
and ( n234706 , n234705 , n234211 );
and ( n234707 , n234207 , n234602 );
or ( n234708 , n234706 , n234707 );
or ( n234709 , n215605 , n220941 );
nand ( n234710 , n234709 , n217573 );
not ( n234711 , n234286 );
not ( n234712 , n221266 );
or ( n234713 , n234711 , n234712 );
not ( n234714 , n220901 );
not ( n234715 , n219389 );
or ( n234716 , n234714 , n234715 );
not ( n234717 , n221559 );
nand ( n234718 , n234717 , n220925 );
nand ( n234719 , n234716 , n234718 );
nand ( n234720 , n234719 , n220929 );
nand ( n234721 , n234713 , n234720 );
xor ( n234722 , n234710 , n234721 );
or ( n234723 , n222471 , n234545 );
not ( n234724 , n231762 );
not ( n234725 , n222586 );
or ( n234726 , n234724 , n234725 );
not ( n234727 , n232280 );
nand ( n234728 , n234727 , n231761 );
nand ( n234729 , n234726 , n234728 );
not ( n234730 , n234729 );
or ( n234731 , n234730 , n221636 );
nand ( n234732 , n234723 , n234731 );
xor ( n234733 , n234722 , n234732 );
xor ( n234734 , n234710 , n234721 );
and ( n234735 , n234734 , n234732 );
and ( n234736 , n234710 , n234721 );
or ( n234737 , n234735 , n234736 );
not ( n234738 , n234238 );
not ( n234739 , n222454 );
or ( n234740 , n234738 , n234739 );
not ( n234741 , n217148 );
not ( n234742 , n222458 );
or ( n234743 , n234741 , n234742 );
nand ( n234744 , n222892 , n220106 );
nand ( n234745 , n234743 , n234744 );
nand ( n234746 , n222467 , n234745 );
nand ( n234747 , n234740 , n234746 );
not ( n234748 , n234248 );
not ( n234749 , n223591 );
or ( n234750 , n234748 , n234749 );
not ( n234751 , n216500 );
nand ( n234752 , n223156 , n234751 );
not ( n234753 , n234752 );
nand ( n234754 , n223202 , n216500 );
not ( n234755 , n234754 );
or ( n234756 , n234753 , n234755 );
nand ( n234757 , n234756 , n222768 );
nand ( n234758 , n234750 , n234757 );
xor ( n234759 , n234747 , n234758 );
not ( n234760 , n234261 );
not ( n234761 , n224087 );
or ( n234762 , n234760 , n234761 );
not ( n234763 , n41565 );
not ( n234764 , n233309 );
not ( n234765 , n234764 );
or ( n234766 , n234763 , n234765 );
nand ( n234767 , n224096 , n211422 );
nand ( n234768 , n234766 , n234767 );
nand ( n234769 , n227782 , n234768 );
nand ( n234770 , n234762 , n234769 );
xor ( n234771 , n234759 , n234770 );
xor ( n234772 , n234747 , n234758 );
and ( n234773 , n234772 , n234770 );
and ( n234774 , n234747 , n234758 );
or ( n234775 , n234773 , n234774 );
not ( n234776 , n217023 );
not ( n234777 , n234598 );
or ( n234778 , n234776 , n234777 );
not ( n234779 , n219577 );
not ( n234780 , n233810 );
or ( n234781 , n234779 , n234780 );
nand ( n234782 , n39286 , n215971 );
nand ( n234783 , n234781 , n234782 );
nand ( n234784 , n234783 , n219175 );
nand ( n234785 , n234778 , n234784 );
not ( n234786 , n220272 );
buf ( n234787 , n216989 );
not ( n234788 , n234787 );
not ( n234789 , n234788 );
not ( n234790 , n229704 );
or ( n234791 , n234789 , n234790 );
not ( n234792 , n229704 );
nand ( n234793 , n234792 , n219358 );
nand ( n234794 , n234791 , n234793 );
not ( n234795 , n234794 );
or ( n234796 , n234786 , n234795 );
nand ( n234797 , n234310 , n220280 );
nand ( n234798 , n234796 , n234797 );
xor ( n234799 , n234785 , n234798 );
not ( n234800 , n219731 );
not ( n234801 , n234328 );
or ( n234802 , n234800 , n234801 );
not ( n234803 , n219033 );
not ( n234804 , n226712 );
or ( n234805 , n234803 , n234804 );
not ( n234806 , n216166 );
nand ( n234807 , n234806 , n226713 );
nand ( n234808 , n234805 , n234807 );
nand ( n234809 , n234808 , n222185 );
nand ( n234810 , n234802 , n234809 );
xor ( n234811 , n234799 , n234810 );
xor ( n234812 , n234785 , n234798 );
and ( n234813 , n234812 , n234810 );
and ( n234814 , n234785 , n234798 );
or ( n234815 , n234813 , n234814 );
not ( n234816 , n214694 );
not ( n234817 , n216810 );
not ( n234818 , n209709 );
or ( n234819 , n234817 , n234818 );
nand ( n234820 , n232856 , n221307 );
nand ( n234821 , n234819 , n234820 );
not ( n234822 , n234821 );
or ( n234823 , n234816 , n234822 );
nand ( n234824 , n234340 , n216299 );
nand ( n234825 , n234823 , n234824 );
not ( n234826 , n219314 );
not ( n234827 , n219687 );
not ( n234828 , n227693 );
or ( n234829 , n234827 , n234828 );
nand ( n234830 , n233856 , n222323 );
nand ( n234831 , n234829 , n234830 );
not ( n234832 , n234831 );
or ( n234833 , n234826 , n234832 );
nand ( n234834 , n234353 , n224624 );
nand ( n234835 , n234833 , n234834 );
xor ( n234836 , n234825 , n234835 );
xor ( n234837 , n234836 , n234733 );
xor ( n234838 , n234825 , n234835 );
and ( n234839 , n234838 , n234733 );
and ( n234840 , n234825 , n234835 );
or ( n234841 , n234839 , n234840 );
not ( n234842 , n234398 );
not ( n234843 , n230339 );
or ( n234844 , n234842 , n234843 );
not ( n234845 , n221495 );
not ( n234846 , n234394 );
or ( n234847 , n234845 , n234846 );
nand ( n234848 , n233450 , n221494 );
nand ( n234849 , n234847 , n234848 );
nand ( n234850 , n233912 , n234849 );
nand ( n234851 , n234844 , n234850 );
not ( n234852 , n234408 );
not ( n234853 , n231421 );
or ( n234854 , n234852 , n234853 );
not ( n234855 , n219343 );
not ( n234856 , n228847 );
or ( n234857 , n234855 , n234856 );
nand ( n234858 , n233929 , n223269 );
nand ( n234859 , n234857 , n234858 );
nand ( n234860 , n228867 , n234859 );
nand ( n234861 , n234854 , n234860 );
xor ( n234862 , n234851 , n234861 );
or ( n234863 , n231474 , n234376 );
and ( n234864 , n233399 , n216934 );
not ( n234865 , n231477 );
and ( n234866 , n234865 , n216940 );
nor ( n234867 , n234864 , n234866 );
or ( n234868 , n231476 , n234867 );
nand ( n234869 , n234863 , n234868 );
xor ( n234870 , n234862 , n234869 );
xor ( n234871 , n234870 , n234771 );
not ( n234872 , n234277 );
not ( n234873 , n227792 );
or ( n234874 , n234872 , n234873 );
not ( n234875 , n225768 );
not ( n234876 , n234273 );
or ( n234877 , n234875 , n234876 );
buf ( n234878 , n233952 );
nand ( n234879 , n234878 , n225769 );
nand ( n234880 , n234877 , n234879 );
nand ( n234881 , n224941 , n234880 );
nand ( n234882 , n234874 , n234881 );
not ( n234883 , n234419 );
not ( n234884 , n230390 );
or ( n234885 , n234883 , n234884 );
not ( n234886 , n214837 );
not ( n234887 , n232497 );
or ( n234888 , n234886 , n234887 );
nand ( n234889 , n225952 , n226698 );
nand ( n234890 , n234888 , n234889 );
nand ( n234891 , n228775 , n234890 );
nand ( n234892 , n234885 , n234891 );
xor ( n234893 , n234882 , n234892 );
not ( n234894 , n229816 );
or ( n234895 , n234894 , n234297 );
not ( n234896 , n227852 );
and ( n234897 , n224041 , n232974 );
not ( n234898 , n224041 );
and ( n234899 , n234898 , n230897 );
nor ( n234900 , n234897 , n234899 );
or ( n234901 , n234896 , n234900 );
nand ( n234902 , n234895 , n234901 );
xor ( n234903 , n234893 , n234902 );
xor ( n234904 , n234871 , n234903 );
xor ( n234905 , n234870 , n234771 );
and ( n234906 , n234905 , n234903 );
and ( n234907 , n234870 , n234771 );
or ( n234908 , n234906 , n234907 );
xor ( n234909 , n234688 , n234692 );
xor ( n234910 , n234909 , n234696 );
xor ( n234911 , n234688 , n234692 );
and ( n234912 , n234911 , n234696 );
and ( n234913 , n234688 , n234692 );
or ( n234914 , n234912 , n234913 );
not ( n234915 , n234366 );
not ( n234916 , n233105 );
or ( n234917 , n234915 , n234916 );
not ( n234918 , n215075 );
not ( n234919 , n230722 );
or ( n234920 , n234918 , n234919 );
nand ( n234921 , n233885 , n215899 );
nand ( n234922 , n234920 , n234921 );
nand ( n234923 , n232402 , n234922 );
nand ( n234924 , n234917 , n234923 );
not ( n234925 , n233891 );
nor ( n234926 , n234925 , n214678 );
xor ( n234927 , n234924 , n234926 );
not ( n234928 , n220881 );
not ( n234929 , n221593 );
not ( n234930 , n218884 );
or ( n234931 , n234929 , n234930 );
nand ( n234932 , n219594 , n220290 );
nand ( n234933 , n234931 , n234932 );
not ( n234934 , n234933 );
or ( n234935 , n234928 , n234934 );
nand ( n234936 , n234484 , n220164 );
nand ( n234937 , n234935 , n234936 );
xor ( n234938 , n234927 , n234937 );
xor ( n234939 , n234938 , n234704 );
xor ( n234940 , n234939 , n234708 );
xor ( n234941 , n234938 , n234704 );
and ( n234942 , n234941 , n234708 );
and ( n234943 , n234938 , n234704 );
or ( n234944 , n234942 , n234943 );
not ( n234945 , n218533 );
not ( n234946 , n218775 );
not ( n234947 , n230966 );
or ( n234948 , n234946 , n234947 );
not ( n234949 , n233083 );
nand ( n234950 , n226922 , n234949 );
nand ( n234951 , n234948 , n234950 );
not ( n234952 , n234951 );
or ( n234953 , n234945 , n234952 );
nand ( n234954 , n234474 , n219461 );
nand ( n234955 , n234953 , n234954 );
not ( n234956 , n222376 );
not ( n234957 , n232413 );
not ( n234958 , n221040 );
or ( n234959 , n234957 , n234958 );
nand ( n234960 , n40625 , n218876 );
nand ( n234961 , n234959 , n234960 );
not ( n234962 , n234961 );
or ( n234963 , n234956 , n234962 );
nand ( n234964 , n234556 , n223665 );
nand ( n234965 , n234963 , n234964 );
xor ( n234966 , n234955 , n234965 );
xor ( n234967 , n234966 , n234547 );
xor ( n234968 , n234335 , n234967 );
not ( n234969 , n228237 );
not ( n234970 , n229387 );
not ( n234971 , n233035 );
or ( n234972 , n234970 , n234971 );
nand ( n234973 , n227007 , n227602 );
nand ( n234974 , n234972 , n234973 );
not ( n234975 , n234974 );
or ( n234976 , n234969 , n234975 );
nand ( n234977 , n229395 , n234534 );
nand ( n234978 , n234976 , n234977 );
not ( n234979 , n219368 );
not ( n234980 , n234446 );
or ( n234981 , n234979 , n234980 );
not ( n234982 , n229261 );
not ( n234983 , n229936 );
or ( n234984 , n234982 , n234983 );
buf ( n234985 , n221716 );
nand ( n234986 , n234985 , n229262 );
nand ( n234987 , n234984 , n234986 );
nand ( n234988 , n234987 , n229964 );
nand ( n234989 , n234981 , n234988 );
xor ( n234990 , n234978 , n234989 );
not ( n234991 , n234463 );
not ( n234992 , n231018 );
or ( n234993 , n234991 , n234992 );
and ( n234994 , n231501 , n221743 );
not ( n234995 , n231501 );
and ( n234996 , n234995 , n223384 );
nor ( n234997 , n234994 , n234996 );
or ( n234998 , n234997 , n227138 );
nand ( n234999 , n234993 , n234998 );
xor ( n235000 , n234990 , n234999 );
xor ( n235001 , n234968 , n235000 );
xor ( n235002 , n234335 , n234967 );
and ( n235003 , n235002 , n235000 );
and ( n235004 , n234335 , n234967 );
or ( n235005 , n235003 , n235004 );
not ( n235006 , n220414 );
not ( n235007 , n234508 );
or ( n235008 , n235006 , n235007 );
not ( n235009 , n226292 );
not ( n235010 , n226961 );
or ( n235011 , n235009 , n235010 );
not ( n235012 , n226961 );
nand ( n235013 , n235012 , n220038 );
nand ( n235014 , n235011 , n235013 );
nand ( n235015 , n235014 , n226287 );
nand ( n235016 , n235008 , n235015 );
not ( n235017 , n219800 );
not ( n235018 , n218912 );
or ( n235019 , n235017 , n235018 );
nand ( n235020 , n218911 , n219420 );
nand ( n235021 , n235019 , n235020 );
not ( n235022 , n235021 );
not ( n235023 , n219076 );
or ( n235024 , n235022 , n235023 );
nand ( n235025 , n234495 , n219792 );
nand ( n235026 , n235024 , n235025 );
xor ( n235027 , n235016 , n235026 );
not ( n235028 , n226655 );
not ( n235029 , n223330 );
or ( n235030 , n235028 , n235029 );
not ( n235031 , n40546 );
nand ( n235032 , n235031 , n233053 );
nand ( n235033 , n235030 , n235032 );
nand ( n235034 , n235033 , n223949 );
nand ( n235035 , n234524 , n227260 );
nand ( n235036 , n235034 , n235035 );
xor ( n235037 , n235027 , n235036 );
xor ( n235038 , n235037 , n234700 );
xor ( n235039 , n235038 , n234389 );
xor ( n235040 , n235037 , n234700 );
and ( n235041 , n235040 , n234389 );
and ( n235042 , n235037 , n234700 );
or ( n235043 , n235041 , n235042 );
not ( n235044 , n219332 );
not ( n235045 , n234567 );
or ( n235046 , n235044 , n235045 );
not ( n235047 , n221935 );
not ( n235048 , n39926 );
or ( n235049 , n235047 , n235048 );
nand ( n235050 , n225097 , n221938 );
nand ( n235051 , n235049 , n235050 );
nand ( n235052 , n235051 , n221933 );
nand ( n235053 , n235046 , n235052 );
xor ( n235054 , n235053 , n234268 );
xor ( n235055 , n235054 , n234304 );
xor ( n235056 , n234428 , n235055 );
not ( n235057 , n231808 );
not ( n235058 , n234583 );
or ( n235059 , n235057 , n235058 );
not ( n235060 , n215113 );
not ( n235061 , n209963 );
or ( n235062 , n235060 , n235061 );
nand ( n235063 , n231104 , n216037 );
nand ( n235064 , n235062 , n235063 );
nand ( n235065 , n235064 , n220985 );
nand ( n235066 , n235059 , n235065 );
xor ( n235067 , n235066 , n234626 );
xor ( n235068 , n235067 , n234684 );
xor ( n235069 , n235056 , n235068 );
xor ( n235070 , n234428 , n235055 );
and ( n235071 , n235070 , n235068 );
and ( n235072 , n234428 , n235055 );
or ( n235073 , n235071 , n235072 );
xor ( n235074 , n234811 , n234837 );
xor ( n235075 , n235074 , n234904 );
xor ( n235076 , n234811 , n234837 );
and ( n235077 , n235076 , n234904 );
and ( n235078 , n234811 , n234837 );
or ( n235079 , n235077 , n235078 );
xor ( n235080 , n234434 , n234910 );
xor ( n235081 , n235080 , n234440 );
xor ( n235082 , n234434 , n234910 );
and ( n235083 , n235082 , n234440 );
and ( n235084 , n234434 , n234910 );
or ( n235085 , n235083 , n235084 );
xor ( n235086 , n234882 , n234892 );
and ( n235087 , n235086 , n234902 );
and ( n235088 , n234882 , n234892 );
or ( n235089 , n235087 , n235088 );
xor ( n235090 , n234518 , n234610 );
xor ( n235091 , n235090 , n235039 );
xor ( n235092 , n234518 , n234610 );
and ( n235093 , n235092 , n235039 );
and ( n235094 , n234518 , n234610 );
or ( n235095 , n235093 , n235094 );
xor ( n235096 , n234940 , n234592 );
xor ( n235097 , n235096 , n235001 );
xor ( n235098 , n234940 , n234592 );
and ( n235099 , n235098 , n235001 );
and ( n235100 , n234940 , n234592 );
or ( n235101 , n235099 , n235100 );
xor ( n235102 , n234616 , n235075 );
xor ( n235103 , n235102 , n235069 );
xor ( n235104 , n234616 , n235075 );
and ( n235105 , n235104 , n235069 );
and ( n235106 , n234616 , n235075 );
or ( n235107 , n235105 , n235106 );
xor ( n235108 , n234622 , n235081 );
xor ( n235109 , n235108 , n234632 );
xor ( n235110 , n234622 , n235081 );
and ( n235111 , n235110 , n234632 );
and ( n235112 , n234622 , n235081 );
or ( n235113 , n235111 , n235112 );
xor ( n235114 , n234638 , n235097 );
xor ( n235115 , n235114 , n235091 );
xor ( n235116 , n234638 , n235097 );
and ( n235117 , n235116 , n235091 );
and ( n235118 , n234638 , n235097 );
or ( n235119 , n235117 , n235118 );
xor ( n235120 , n235103 , n234644 );
xor ( n235121 , n235120 , n234650 );
xor ( n235122 , n235103 , n234644 );
and ( n235123 , n235122 , n234650 );
and ( n235124 , n235103 , n234644 );
or ( n235125 , n235123 , n235124 );
xor ( n235126 , n235109 , n234656 );
xor ( n235127 , n235126 , n235115 );
xor ( n235128 , n235109 , n234656 );
and ( n235129 , n235128 , n235115 );
and ( n235130 , n235109 , n234656 );
or ( n235131 , n235129 , n235130 );
xor ( n235132 , n235121 , n234662 );
xor ( n235133 , n235132 , n234668 );
xor ( n235134 , n235121 , n234662 );
and ( n235135 , n235134 , n234668 );
and ( n235136 , n235121 , n234662 );
or ( n235137 , n235135 , n235136 );
xor ( n235138 , n235127 , n235133 );
xor ( n235139 , n235138 , n234674 );
xor ( n235140 , n235127 , n235133 );
and ( n235141 , n235140 , n234674 );
and ( n235142 , n235127 , n235133 );
or ( n235143 , n235141 , n235142 );
xor ( n235144 , n234851 , n234861 );
and ( n235145 , n235144 , n234869 );
and ( n235146 , n234851 , n234861 );
or ( n235147 , n235145 , n235146 );
xor ( n235148 , n234924 , n234926 );
and ( n235149 , n235148 , n234937 );
and ( n235150 , n234924 , n234926 );
or ( n235151 , n235149 , n235150 );
xor ( n235152 , n235016 , n235026 );
and ( n235153 , n235152 , n235036 );
and ( n235154 , n235016 , n235026 );
or ( n235155 , n235153 , n235154 );
xor ( n235156 , n234978 , n234989 );
and ( n235157 , n235156 , n234999 );
and ( n235158 , n234978 , n234989 );
or ( n235159 , n235157 , n235158 );
xor ( n235160 , n234955 , n234965 );
and ( n235161 , n235160 , n234547 );
and ( n235162 , n234955 , n234965 );
or ( n235163 , n235161 , n235162 );
xor ( n235164 , n235053 , n234268 );
and ( n235165 , n235164 , n234304 );
and ( n235166 , n235053 , n234268 );
or ( n235167 , n235165 , n235166 );
xor ( n235168 , n235066 , n234626 );
and ( n235169 , n235168 , n234684 );
and ( n235170 , n235066 , n234626 );
or ( n235171 , n235169 , n235170 );
buf ( n235172 , n223197 );
not ( n235173 , n235172 );
nand ( n235174 , n234754 , n234752 );
not ( n235175 , n235174 );
or ( n235176 , n235173 , n235175 );
not ( n235177 , n219902 );
not ( n235178 , n225914 );
or ( n235179 , n235177 , n235178 );
nand ( n235180 , n224059 , n208597 );
nand ( n235181 , n235179 , n235180 );
nand ( n235182 , n222768 , n235181 );
nand ( n235183 , n235176 , n235182 );
not ( n235184 , n234768 );
not ( n235185 , n224087 );
or ( n235186 , n235184 , n235185 );
not ( n235187 , n208717 );
not ( n235188 , n234764 );
or ( n235189 , n235187 , n235188 );
nand ( n235190 , n223989 , n232282 );
nand ( n235191 , n235189 , n235190 );
nand ( n235192 , n224090 , n235191 );
nand ( n235193 , n235186 , n235192 );
xor ( n235194 , n235183 , n235193 );
not ( n235195 , n227792 );
not ( n235196 , n234880 );
or ( n235197 , n235195 , n235196 );
and ( n235198 , n234256 , n233952 );
not ( n235199 , n234256 );
buf ( n235200 , n226747 );
and ( n235201 , n235199 , n235200 );
nor ( n235202 , n235198 , n235201 );
or ( n235203 , n232948 , n235202 );
nand ( n235204 , n235197 , n235203 );
xor ( n235205 , n235194 , n235204 );
xor ( n235206 , n235183 , n235193 );
and ( n235207 , n235206 , n235204 );
and ( n235208 , n235183 , n235193 );
or ( n235209 , n235207 , n235208 );
not ( n235210 , n234890 );
not ( n235211 , n226755 );
or ( n235212 , n235210 , n235211 );
not ( n235213 , n226304 );
not ( n235214 , n226276 );
or ( n235215 , n235213 , n235214 );
not ( n235216 , n226304 );
nand ( n235217 , n225952 , n235216 );
nand ( n235218 , n235215 , n235217 );
nand ( n235219 , n228775 , n235218 );
nand ( n235220 , n235212 , n235219 );
not ( n235221 , n234729 );
not ( n235222 , n221626 );
or ( n235223 , n235221 , n235222 );
not ( n235224 , n217330 );
not ( n235225 , n226388 );
or ( n235226 , n235224 , n235225 );
not ( n235227 , n234727 );
nand ( n235228 , n235227 , n219201 );
nand ( n235229 , n235226 , n235228 );
nand ( n235230 , n221387 , n235229 );
nand ( n235231 , n235223 , n235230 );
xor ( n235232 , n235220 , n235231 );
not ( n235233 , n234849 );
not ( n235234 , n233446 );
or ( n235235 , n235233 , n235234 );
not ( n235236 , n216293 );
not ( n235237 , n233451 );
or ( n235238 , n235236 , n235237 );
nand ( n235239 , n233450 , n223658 );
nand ( n235240 , n235238 , n235239 );
nand ( n235241 , n233912 , n235240 );
nand ( n235242 , n235235 , n235241 );
xor ( n235243 , n235232 , n235242 );
xor ( n235244 , n235220 , n235231 );
and ( n235245 , n235244 , n235242 );
and ( n235246 , n235220 , n235231 );
or ( n235247 , n235245 , n235246 );
not ( n235248 , n217023 );
not ( n235249 , n234783 );
or ( n235250 , n235248 , n235249 );
not ( n235251 , n219577 );
not ( n235252 , n233362 );
or ( n235253 , n235251 , n235252 );
nand ( n235254 , n229217 , n218661 );
nand ( n235255 , n235253 , n235254 );
nand ( n235256 , n235255 , n219175 );
nand ( n235257 , n235250 , n235256 );
not ( n235258 , n219332 );
not ( n235259 , n235051 );
or ( n235260 , n235258 , n235259 );
nor ( n235261 , n221938 , n221932 );
nand ( n235262 , n235261 , n234347 );
not ( n235263 , n221932 );
nand ( n235264 , n235263 , n227223 , n221938 );
and ( n235265 , n235262 , n235264 );
nand ( n235266 , n235260 , n235265 );
xor ( n235267 , n235257 , n235266 );
xor ( n235268 , n235267 , n234737 );
xor ( n235269 , n235257 , n235266 );
and ( n235270 , n235269 , n234737 );
and ( n235271 , n235257 , n235266 );
or ( n235272 , n235270 , n235271 );
and ( n235273 , n234382 , n216208 );
not ( n235274 , n234922 );
not ( n235275 , n232399 );
or ( n235276 , n235274 , n235275 );
and ( n235277 , n218514 , n230725 );
not ( n235278 , n218514 );
not ( n235279 , n230722 );
and ( n235280 , n235278 , n235279 );
or ( n235281 , n235277 , n235280 );
nand ( n235282 , n232402 , n235281 );
nand ( n235283 , n235276 , n235282 );
xor ( n235284 , n235273 , n235283 );
not ( n235285 , n221674 );
and ( n235286 , n40724 , n220901 );
not ( n235287 , n40724 );
and ( n235288 , n235287 , n220906 );
or ( n235289 , n235286 , n235288 );
not ( n235290 , n235289 );
or ( n235291 , n235285 , n235290 );
not ( n235292 , n228639 );
nand ( n235293 , n235292 , n234719 );
nand ( n235294 , n235291 , n235293 );
xor ( n235295 , n235284 , n235294 );
not ( n235296 , n234859 );
not ( n235297 , n228858 );
or ( n235298 , n235296 , n235297 );
not ( n235299 , n222821 );
not ( n235300 , n228847 );
or ( n235301 , n235299 , n235300 );
nand ( n235302 , n230851 , n218980 );
nand ( n235303 , n235301 , n235302 );
nand ( n235304 , n229738 , n235303 );
nand ( n235305 , n235298 , n235304 );
or ( n235306 , n231474 , n234867 );
not ( n235307 , n219102 );
not ( n235308 , n229762 );
or ( n235309 , n235307 , n235308 );
nand ( n235310 , n229761 , n216139 );
nand ( n235311 , n235309 , n235310 );
not ( n235312 , n235311 );
or ( n235313 , n231476 , n235312 );
nand ( n235314 , n235306 , n235313 );
xor ( n235315 , n235305 , n235314 );
not ( n235316 , n226885 );
not ( n235317 , n224492 );
not ( n235318 , n230897 );
or ( n235319 , n235317 , n235318 );
nand ( n235320 , n229823 , n214642 );
nand ( n235321 , n235319 , n235320 );
not ( n235322 , n235321 );
or ( n235323 , n235316 , n235322 );
or ( n235324 , n234290 , n234900 );
nand ( n235325 , n235323 , n235324 );
xor ( n235326 , n235315 , n235325 );
xor ( n235327 , n235295 , n235326 );
xor ( n235328 , n235327 , n235205 );
xor ( n235329 , n235295 , n235326 );
and ( n235330 , n235329 , n235205 );
and ( n235331 , n235295 , n235326 );
or ( n235332 , n235330 , n235331 );
xor ( n235333 , n235243 , n235151 );
xor ( n235334 , n235333 , n235155 );
xor ( n235335 , n235243 , n235151 );
and ( n235336 , n235335 , n235155 );
and ( n235337 , n235243 , n235151 );
or ( n235338 , n235336 , n235337 );
xor ( n235339 , n235159 , n235163 );
xor ( n235340 , n235339 , n235171 );
xor ( n235341 , n235159 , n235163 );
and ( n235342 , n235341 , n235171 );
and ( n235343 , n235159 , n235163 );
or ( n235344 , n235342 , n235343 );
not ( n235345 , n219461 );
not ( n235346 , n234951 );
or ( n235347 , n235345 , n235346 );
not ( n235348 , n218208 );
not ( n235349 , n220599 );
or ( n235350 , n235348 , n235349 );
nand ( n235351 , n221956 , n234949 );
nand ( n235352 , n235350 , n235351 );
nand ( n235353 , n235352 , n218533 );
nand ( n235354 , n235347 , n235353 );
not ( n235355 , n218843 );
not ( n235356 , n232413 );
not ( n235357 , n40660 );
or ( n235358 , n235356 , n235357 );
buf ( n235359 , n207936 );
nand ( n235360 , n235359 , n221238 );
nand ( n235361 , n235358 , n235360 );
not ( n235362 , n235361 );
or ( n235363 , n235355 , n235362 );
nand ( n235364 , n234961 , n223665 );
nand ( n235365 , n235363 , n235364 );
xor ( n235366 , n235354 , n235365 );
not ( n235367 , n220507 );
not ( n235368 , n235021 );
or ( n235369 , n235367 , n235368 );
not ( n235370 , n219424 );
not ( n235371 , n227448 );
or ( n235372 , n235370 , n235371 );
nand ( n235373 , n219226 , n219420 );
nand ( n235374 , n235372 , n235373 );
nand ( n235375 , n235374 , n219076 );
nand ( n235376 , n235369 , n235375 );
xor ( n235377 , n235366 , n235376 );
xor ( n235378 , n234815 , n235377 );
not ( n235379 , n234006 );
not ( n235380 , n234987 );
or ( n235381 , n235379 , n235380 );
not ( n235382 , n229261 );
not ( n235383 , n40422 );
not ( n235384 , n235383 );
or ( n235385 , n235382 , n235384 );
nand ( n235386 , n40422 , n229262 );
nand ( n235387 , n235385 , n235386 );
nand ( n235388 , n235387 , n229964 );
nand ( n235389 , n235381 , n235388 );
not ( n235390 , n234745 );
not ( n235391 , n222454 );
or ( n235392 , n235390 , n235391 );
and ( n235393 , n208164 , n222435 );
not ( n235394 , n208164 );
and ( n235395 , n235394 , n222430 );
nor ( n235396 , n235393 , n235395 );
not ( n235397 , n235396 );
nand ( n235398 , n235397 , n222158 );
nand ( n235399 , n235392 , n235398 );
not ( n235400 , n235399 );
xor ( n235401 , n235389 , n235400 );
or ( n235402 , n234997 , n227130 );
not ( n235403 , n217616 );
not ( n235404 , n222121 );
or ( n235405 , n235403 , n235404 );
nand ( n235406 , n40397 , n218253 );
nand ( n235407 , n235405 , n235406 );
not ( n235408 , n235407 );
or ( n235409 , n235408 , n227138 );
nand ( n235410 , n235402 , n235409 );
xor ( n235411 , n235401 , n235410 );
xor ( n235412 , n235378 , n235411 );
xor ( n235413 , n234815 , n235377 );
and ( n235414 , n235413 , n235411 );
and ( n235415 , n234815 , n235377 );
or ( n235416 , n235414 , n235415 );
not ( n235417 , n220164 );
not ( n235418 , n234933 );
or ( n235419 , n235417 , n235418 );
not ( n235420 , n40766 );
not ( n235421 , n220500 );
or ( n235422 , n235420 , n235421 );
nand ( n235423 , n226489 , n221257 );
nand ( n235424 , n235422 , n235423 );
nand ( n235425 , n220881 , n235424 );
nand ( n235426 , n235419 , n235425 );
not ( n235427 , n227260 );
not ( n235428 , n235033 );
or ( n235429 , n235427 , n235428 );
not ( n235430 , n226655 );
not ( n235431 , n234503 );
or ( n235432 , n235430 , n235431 );
nand ( n235433 , n234506 , n233053 );
nand ( n235434 , n235432 , n235433 );
nand ( n235435 , n235434 , n223949 );
nand ( n235436 , n235429 , n235435 );
xor ( n235437 , n235426 , n235436 );
not ( n235438 , n229395 );
not ( n235439 , n234974 );
or ( n235440 , n235438 , n235439 );
not ( n235441 , n229387 );
not ( n235442 , n223721 );
or ( n235443 , n235441 , n235442 );
nand ( n235444 , n40485 , n227599 );
nand ( n235445 , n235443 , n235444 );
nand ( n235446 , n235445 , n228237 );
nand ( n235447 , n235440 , n235446 );
xor ( n235448 , n235437 , n235447 );
xor ( n235449 , n235167 , n235448 );
not ( n235450 , n226287 );
not ( n235451 , n227912 );
not ( n235452 , n225344 );
not ( n235453 , n235452 );
or ( n235454 , n235451 , n235453 );
not ( n235455 , n39877 );
nand ( n235456 , n235455 , n229887 );
nand ( n235457 , n235454 , n235456 );
not ( n235458 , n235457 );
or ( n235459 , n235450 , n235458 );
nand ( n235460 , n235014 , n226943 );
nand ( n235461 , n235459 , n235460 );
xor ( n235462 , n235461 , n234775 );
xor ( n235463 , n235462 , n235089 );
xor ( n235464 , n235449 , n235463 );
xor ( n235465 , n235167 , n235448 );
and ( n235466 , n235465 , n235463 );
and ( n235467 , n235167 , n235448 );
or ( n235468 , n235466 , n235467 );
xor ( n235469 , n234908 , n235268 );
not ( n235470 , n216562 );
not ( n235471 , n234821 );
or ( n235472 , n235470 , n235471 );
and ( n235473 , n216810 , n233611 );
not ( n235474 , n216810 );
and ( n235475 , n235474 , n209865 );
or ( n235476 , n235473 , n235475 );
nand ( n235477 , n235476 , n214694 );
nand ( n235478 , n235472 , n235477 );
xor ( n235479 , n235478 , n235147 );
not ( n235480 , n220272 );
not ( n235481 , n234788 );
not ( n235482 , n228165 );
or ( n235483 , n235481 , n235482 );
or ( n235484 , n228165 , n215955 );
nand ( n235485 , n235483 , n235484 );
not ( n235486 , n235485 );
or ( n235487 , n235480 , n235486 );
nand ( n235488 , n234794 , n220280 );
nand ( n235489 , n235487 , n235488 );
xor ( n235490 , n235479 , n235489 );
xor ( n235491 , n235469 , n235490 );
xor ( n235492 , n234908 , n235268 );
and ( n235493 , n235492 , n235490 );
and ( n235494 , n234908 , n235268 );
or ( n235495 , n235493 , n235494 );
not ( n235496 , n222185 );
not ( n235497 , n219033 );
not ( n235498 , n228184 );
or ( n235499 , n235497 , n235498 );
nand ( n235500 , n39089 , n220538 );
nand ( n235501 , n235499 , n235500 );
not ( n235502 , n235501 );
or ( n235503 , n235496 , n235502 );
nand ( n235504 , n234808 , n219731 );
nand ( n235505 , n235503 , n235504 );
not ( n235506 , n214717 );
not ( n235507 , n235064 );
or ( n235508 , n235506 , n235507 );
nand ( n235509 , n220985 , n221338 );
nand ( n235510 , n235508 , n235509 );
xor ( n235511 , n235505 , n235510 );
not ( n235512 , n216204 );
not ( n235513 , n234831 );
or ( n235514 , n235512 , n235513 );
not ( n235515 , n219687 );
buf ( n235516 , n228216 );
not ( n235517 , n235516 );
or ( n235518 , n235515 , n235517 );
nand ( n235519 , n39747 , n222323 );
nand ( n235520 , n235518 , n235519 );
nand ( n235521 , n235520 , n219314 );
nand ( n235522 , n235514 , n235521 );
xor ( n235523 , n235511 , n235522 );
xor ( n235524 , n234841 , n235523 );
xor ( n235525 , n235524 , n235328 );
xor ( n235526 , n234841 , n235523 );
and ( n235527 , n235526 , n235328 );
and ( n235528 , n234841 , n235523 );
or ( n235529 , n235527 , n235528 );
xor ( n235530 , n234914 , n235005 );
xor ( n235531 , n235530 , n235334 );
xor ( n235532 , n234914 , n235005 );
and ( n235533 , n235532 , n235334 );
and ( n235534 , n234914 , n235005 );
or ( n235535 , n235533 , n235534 );
xor ( n235536 , n234944 , n235340 );
xor ( n235537 , n235536 , n235073 );
xor ( n235538 , n234944 , n235340 );
and ( n235539 , n235538 , n235073 );
and ( n235540 , n234944 , n235340 );
or ( n235541 , n235539 , n235540 );
xor ( n235542 , n235305 , n235314 );
and ( n235543 , n235542 , n235325 );
and ( n235544 , n235305 , n235314 );
or ( n235545 , n235543 , n235544 );
xor ( n235546 , n235043 , n235464 );
xor ( n235547 , n235546 , n235412 );
xor ( n235548 , n235043 , n235464 );
and ( n235549 , n235548 , n235412 );
and ( n235550 , n235043 , n235464 );
or ( n235551 , n235549 , n235550 );
xor ( n235552 , n235079 , n235525 );
xor ( n235553 , n235552 , n235491 );
xor ( n235554 , n235079 , n235525 );
and ( n235555 , n235554 , n235491 );
and ( n235556 , n235079 , n235525 );
or ( n235557 , n235555 , n235556 );
xor ( n235558 , n235085 , n235101 );
xor ( n235559 , n235558 , n235095 );
xor ( n235560 , n235085 , n235101 );
and ( n235561 , n235560 , n235095 );
and ( n235562 , n235085 , n235101 );
or ( n235563 , n235561 , n235562 );
xor ( n235564 , n235531 , n235537 );
xor ( n235565 , n235564 , n235547 );
xor ( n235566 , n235531 , n235537 );
and ( n235567 , n235566 , n235547 );
and ( n235568 , n235531 , n235537 );
or ( n235569 , n235567 , n235568 );
xor ( n235570 , n235107 , n235553 );
xor ( n235571 , n235570 , n235113 );
xor ( n235572 , n235107 , n235553 );
and ( n235573 , n235572 , n235113 );
and ( n235574 , n235107 , n235553 );
or ( n235575 , n235573 , n235574 );
xor ( n235576 , n235119 , n235565 );
xor ( n235577 , n235576 , n235559 );
xor ( n235578 , n235119 , n235565 );
and ( n235579 , n235578 , n235559 );
and ( n235580 , n235119 , n235565 );
or ( n235581 , n235579 , n235580 );
xor ( n235582 , n235571 , n235125 );
xor ( n235583 , n235582 , n235131 );
xor ( n235584 , n235571 , n235125 );
and ( n235585 , n235584 , n235131 );
and ( n235586 , n235571 , n235125 );
or ( n235587 , n235585 , n235586 );
xor ( n235588 , n235577 , n235583 );
xor ( n235589 , n235588 , n235137 );
xor ( n235590 , n235577 , n235583 );
and ( n235591 , n235590 , n235137 );
and ( n235592 , n235577 , n235583 );
or ( n235593 , n235591 , n235592 );
xor ( n235594 , n235273 , n235283 );
and ( n235595 , n235594 , n235294 );
and ( n235596 , n235273 , n235283 );
or ( n235597 , n235595 , n235596 );
xor ( n235598 , n235426 , n235436 );
and ( n235599 , n235598 , n235447 );
and ( n235600 , n235426 , n235436 );
or ( n235601 , n235599 , n235600 );
xor ( n235602 , n235389 , n235400 );
and ( n235603 , n235602 , n235410 );
and ( n235604 , n235389 , n235400 );
or ( n235605 , n235603 , n235604 );
xor ( n235606 , n235354 , n235365 );
and ( n235607 , n235606 , n235376 );
and ( n235608 , n235354 , n235365 );
or ( n235609 , n235607 , n235608 );
xor ( n235610 , n235461 , n234775 );
and ( n235611 , n235610 , n235089 );
and ( n235612 , n235461 , n234775 );
or ( n235613 , n235611 , n235612 );
xor ( n235614 , n235478 , n235147 );
and ( n235615 , n235614 , n235489 );
and ( n235616 , n235478 , n235147 );
or ( n235617 , n235615 , n235616 );
xor ( n235618 , n235505 , n235510 );
and ( n235619 , n235618 , n235522 );
and ( n235620 , n235505 , n235510 );
or ( n235621 , n235619 , n235620 );
or ( n235622 , n214717 , n216239 );
nand ( n235623 , n235622 , n221338 );
not ( n235624 , n235229 );
not ( n235625 , n221626 );
or ( n235626 , n235624 , n235625 );
not ( n235627 , n223584 );
not ( n235628 , n220823 );
or ( n235629 , n235627 , n235628 );
nand ( n235630 , n222586 , n221559 );
nand ( n235631 , n235629 , n235630 );
nand ( n235632 , n235631 , n221387 );
nand ( n235633 , n235626 , n235632 );
xor ( n235634 , n235623 , n235633 );
not ( n235635 , n231762 );
not ( n235636 , n222458 );
or ( n235637 , n235635 , n235636 );
not ( n235638 , n220226 );
nand ( n235639 , n235638 , n222892 );
nand ( n235640 , n235637 , n235639 );
not ( n235641 , n235640 );
not ( n235642 , n222158 );
or ( n235643 , n235641 , n235642 );
not ( n235644 , n222886 );
or ( n235645 , n235644 , n235396 );
nand ( n235646 , n235643 , n235645 );
xor ( n235647 , n235634 , n235646 );
xor ( n235648 , n235623 , n235633 );
and ( n235649 , n235648 , n235646 );
and ( n235650 , n235623 , n235633 );
or ( n235651 , n235649 , n235650 );
not ( n235652 , n235181 );
not ( n235653 , n223591 );
or ( n235654 , n235652 , n235653 );
not ( n235655 , n217148 );
not ( n235656 , n223183 );
or ( n235657 , n235655 , n235656 );
nand ( n235658 , n224059 , n220106 );
nand ( n235659 , n235657 , n235658 );
nand ( n235660 , n235659 , n222768 );
nand ( n235661 , n235654 , n235660 );
not ( n235662 , n235191 );
not ( n235663 , n224087 );
or ( n235664 , n235662 , n235663 );
not ( n235665 , n224095 );
not ( n235666 , n219582 );
or ( n235667 , n235665 , n235666 );
nand ( n235668 , n219581 , n224068 );
nand ( n235669 , n235667 , n235668 );
nand ( n235670 , n224090 , n235669 );
nand ( n235671 , n235664 , n235670 );
xor ( n235672 , n235661 , n235671 );
or ( n235673 , n233316 , n235202 );
not ( n235674 , n41565 );
not ( n235675 , n229795 );
or ( n235676 , n235674 , n235675 );
nand ( n235677 , n224929 , n216543 );
nand ( n235678 , n235676 , n235677 );
not ( n235679 , n235678 );
or ( n235680 , n232948 , n235679 );
nand ( n235681 , n235673 , n235680 );
xor ( n235682 , n235672 , n235681 );
xor ( n235683 , n235661 , n235671 );
and ( n235684 , n235683 , n235681 );
and ( n235685 , n235661 , n235671 );
or ( n235686 , n235684 , n235685 );
not ( n235687 , n219175 );
not ( n235688 , n217017 );
not ( n235689 , n209709 );
or ( n235690 , n235688 , n235689 );
not ( n235691 , n229691 );
nand ( n235692 , n235691 , n215971 );
nand ( n235693 , n235690 , n235692 );
not ( n235694 , n235693 );
or ( n235695 , n235687 , n235694 );
nand ( n235696 , n235255 , n217023 );
nand ( n235697 , n235695 , n235696 );
not ( n235698 , n221935 );
not ( n235699 , n225792 );
or ( n235700 , n235698 , n235699 );
nand ( n235701 , n39713 , n222333 );
nand ( n235702 , n235700 , n235701 );
not ( n235703 , n235702 );
not ( n235704 , n221933 );
or ( n235705 , n235703 , n235704 );
or ( n235706 , n234347 , n221938 );
not ( n235707 , n227223 );
nand ( n235708 , n235707 , n221938 );
nand ( n235709 , n235706 , n235708 , n219332 );
nand ( n235710 , n235705 , n235709 );
xor ( n235711 , n235697 , n235710 );
xor ( n235712 , n235711 , n235209 );
xor ( n235713 , n235697 , n235710 );
and ( n235714 , n235713 , n235209 );
and ( n235715 , n235697 , n235710 );
or ( n235716 , n235714 , n235715 );
xor ( n235717 , n235597 , n235647 );
not ( n235718 , n235303 );
not ( n235719 , n228858 );
or ( n235720 , n235718 , n235719 );
not ( n235721 , n220022 );
not ( n235722 , n231943 );
or ( n235723 , n235721 , n235722 );
not ( n235724 , n230851 );
nand ( n235725 , n235724 , n221495 );
nand ( n235726 , n235723 , n235725 );
nand ( n235727 , n235726 , n228867 );
nand ( n235728 , n235720 , n235727 );
not ( n235729 , n235311 );
not ( n235730 , n229773 );
or ( n235731 , n235729 , n235730 );
not ( n235732 , n219348 );
not ( n235733 , n229759 );
or ( n235734 , n235732 , n235733 );
not ( n235735 , n229761 );
nand ( n235736 , n235735 , n219343 );
nand ( n235737 , n235734 , n235736 );
nand ( n235738 , n229777 , n235737 );
nand ( n235739 , n235731 , n235738 );
xor ( n235740 , n235728 , n235739 );
not ( n235741 , n235281 );
not ( n235742 , n232399 );
or ( n235743 , n235741 , n235742 );
not ( n235744 , n233885 );
nand ( n235745 , n235744 , n216934 );
not ( n235746 , n235745 );
nand ( n235747 , n231232 , n216940 );
not ( n235748 , n235747 );
or ( n235749 , n235746 , n235748 );
nand ( n235750 , n235749 , n232402 );
nand ( n235751 , n235743 , n235750 );
xor ( n235752 , n235740 , n235751 );
xor ( n235753 , n235717 , n235752 );
xor ( n235754 , n235597 , n235647 );
and ( n235755 , n235754 , n235752 );
and ( n235756 , n235597 , n235647 );
or ( n235757 , n235755 , n235756 );
not ( n235758 , n235218 );
not ( n235759 , n229271 );
or ( n235760 , n235758 , n235759 );
not ( n235761 , n225764 );
not ( n235762 , n226276 );
or ( n235763 , n235761 , n235762 );
nand ( n235764 , n225952 , n225769 );
nand ( n235765 , n235763 , n235764 );
nand ( n235766 , n227710 , n235765 );
nand ( n235767 , n235760 , n235766 );
not ( n235768 , n235321 );
not ( n235769 , n227849 );
or ( n235770 , n235768 , n235769 );
not ( n235771 , n214837 );
not ( n235772 , n226888 );
or ( n235773 , n235771 , n235772 );
nand ( n235774 , n229823 , n218670 );
nand ( n235775 , n235773 , n235774 );
nand ( n235776 , n235775 , n227241 );
nand ( n235777 , n235770 , n235776 );
xor ( n235778 , n235767 , n235777 );
not ( n235779 , n235240 );
not ( n235780 , n230339 );
or ( n235781 , n235779 , n235780 );
not ( n235782 , n224037 );
not ( n235783 , n233451 );
or ( n235784 , n235782 , n235783 );
nand ( n235785 , n233450 , n224041 );
nand ( n235786 , n235784 , n235785 );
nand ( n235787 , n233912 , n235786 );
nand ( n235788 , n235781 , n235787 );
xor ( n235789 , n235778 , n235788 );
xor ( n235790 , n235789 , n235682 );
xor ( n235791 , n235790 , n235601 );
xor ( n235792 , n235789 , n235682 );
and ( n235793 , n235792 , n235601 );
and ( n235794 , n235789 , n235682 );
or ( n235795 , n235793 , n235794 );
xor ( n235796 , n235605 , n235609 );
xor ( n235797 , n235796 , n235613 );
xor ( n235798 , n235605 , n235609 );
and ( n235799 , n235798 , n235613 );
and ( n235800 , n235605 , n235609 );
or ( n235801 , n235799 , n235800 );
xor ( n235802 , n235621 , n235272 );
not ( n235803 , n219435 );
not ( n235804 , n235374 );
or ( n235805 , n235803 , n235804 );
not ( n235806 , n219800 );
not ( n235807 , n221040 );
or ( n235808 , n235806 , n235807 );
not ( n235809 , n221228 );
nand ( n235810 , n235809 , n221690 );
nand ( n235811 , n235808 , n235810 );
nand ( n235812 , n235811 , n219076 );
nand ( n235813 , n235805 , n235812 );
xor ( n235814 , n235813 , n235399 );
not ( n235815 , n226287 );
not ( n235816 , n227912 );
not ( n235817 , n226727 );
not ( n235818 , n235817 );
or ( n235819 , n235816 , n235818 );
not ( n235820 , n39927 );
nand ( n235821 , n235820 , n220038 );
nand ( n235822 , n235819 , n235821 );
not ( n235823 , n235822 );
or ( n235824 , n235815 , n235823 );
nand ( n235825 , n235457 , n220414 );
nand ( n235826 , n235824 , n235825 );
xor ( n235827 , n235814 , n235826 );
xor ( n235828 , n235802 , n235827 );
xor ( n235829 , n235621 , n235272 );
and ( n235830 , n235829 , n235827 );
and ( n235831 , n235621 , n235272 );
or ( n235832 , n235830 , n235831 );
not ( n235833 , n220067 );
not ( n235834 , n217614 );
not ( n235835 , n221715 );
or ( n235836 , n235834 , n235835 );
nand ( n235837 , n223320 , n218253 );
nand ( n235838 , n235836 , n235837 );
not ( n235839 , n235838 );
or ( n235840 , n235833 , n235839 );
nand ( n235841 , n235407 , n231018 );
nand ( n235842 , n235840 , n235841 );
not ( n235843 , n218533 );
not ( n235844 , n218775 );
not ( n235845 , n40258 );
or ( n235846 , n235844 , n235845 );
nand ( n235847 , n220970 , n218226 );
nand ( n235848 , n235846 , n235847 );
not ( n235849 , n235848 );
or ( n235850 , n235843 , n235849 );
nand ( n235851 , n235352 , n219461 );
nand ( n235852 , n235850 , n235851 );
xor ( n235853 , n235842 , n235852 );
not ( n235854 , n222376 );
not ( n235855 , n232413 );
not ( n235856 , n226921 );
or ( n235857 , n235855 , n235856 );
nand ( n235858 , n226922 , n221238 );
nand ( n235859 , n235857 , n235858 );
not ( n235860 , n235859 );
or ( n235861 , n235854 , n235860 );
nand ( n235862 , n235361 , n223665 );
nand ( n235863 , n235861 , n235862 );
xor ( n235864 , n235853 , n235863 );
not ( n235865 , n220492 );
not ( n235866 , n235424 );
or ( n235867 , n235865 , n235866 );
not ( n235868 , n220500 );
not ( n235869 , n220204 );
or ( n235870 , n235868 , n235869 );
nand ( n235871 , n218911 , n221257 );
nand ( n235872 , n235870 , n235871 );
nand ( n235873 , n235872 , n219779 );
nand ( n235874 , n235867 , n235873 );
not ( n235875 , n228237 );
not ( n235876 , n233544 );
not ( n235877 , n40546 );
or ( n235878 , n235876 , n235877 );
nand ( n235879 , n223333 , n227599 );
nand ( n235880 , n235878 , n235879 );
not ( n235881 , n235880 );
or ( n235882 , n235875 , n235881 );
nand ( n235883 , n235445 , n225478 );
nand ( n235884 , n235882 , n235883 );
xor ( n235885 , n235874 , n235884 );
not ( n235886 , n229964 );
not ( n235887 , n234449 );
not ( n235888 , n227004 );
or ( n235889 , n235887 , n235888 );
nand ( n235890 , n40415 , n229262 );
nand ( n235891 , n235889 , n235890 );
not ( n235892 , n235891 );
or ( n235893 , n235886 , n235892 );
nand ( n235894 , n235387 , n229974 );
nand ( n235895 , n235893 , n235894 );
xor ( n235896 , n235885 , n235895 );
xor ( n235897 , n235864 , n235896 );
xor ( n235898 , n235897 , n235617 );
xor ( n235899 , n235864 , n235896 );
and ( n235900 , n235899 , n235617 );
and ( n235901 , n235864 , n235896 );
or ( n235902 , n235900 , n235901 );
and ( n235903 , n233465 , n215075 );
not ( n235904 , n221674 );
not ( n235905 , n220906 );
not ( n235906 , n218884 );
or ( n235907 , n235905 , n235906 );
not ( n235908 , n218884 );
nand ( n235909 , n235908 , n220901 );
nand ( n235910 , n235907 , n235909 );
not ( n235911 , n235910 );
or ( n235912 , n235904 , n235911 );
buf ( n235913 , n221266 );
nand ( n235914 , n235289 , n235913 );
nand ( n235915 , n235912 , n235914 );
xor ( n235916 , n235903 , n235915 );
not ( n235917 , n227260 );
not ( n235918 , n235434 );
or ( n235919 , n235917 , n235918 );
not ( n235920 , n226655 );
not ( n235921 , n226964 );
not ( n235922 , n235921 );
or ( n235923 , n235920 , n235922 );
nand ( n235924 , n225111 , n227927 );
nand ( n235925 , n235923 , n235924 );
nand ( n235926 , n235925 , n223949 );
nand ( n235927 , n235919 , n235926 );
xor ( n235928 , n235916 , n235927 );
xor ( n235929 , n235247 , n235545 );
not ( n235930 , n235476 );
or ( n235931 , n235930 , n216298 );
not ( n235932 , n231104 );
not ( n235933 , n215289 );
or ( n235934 , n235932 , n235933 );
nand ( n235935 , n233134 , n216810 );
nand ( n235936 , n235934 , n235935 );
not ( n235937 , n235936 );
or ( n235938 , n235937 , n220819 );
nand ( n235939 , n235931 , n235938 );
xor ( n235940 , n235929 , n235939 );
xor ( n235941 , n235928 , n235940 );
xor ( n235942 , n235941 , n235712 );
xor ( n235943 , n235928 , n235940 );
and ( n235944 , n235943 , n235712 );
and ( n235945 , n235928 , n235940 );
or ( n235946 , n235944 , n235945 );
not ( n235947 , n220280 );
not ( n235948 , n235485 );
or ( n235949 , n235947 , n235948 );
not ( n235950 , n234788 );
not ( n235951 , n39287 );
or ( n235952 , n235950 , n235951 );
buf ( n235953 , n39286 );
nand ( n235954 , n235953 , n219358 );
nand ( n235955 , n235952 , n235954 );
nand ( n235956 , n235955 , n220272 );
nand ( n235957 , n235949 , n235956 );
not ( n235958 , n219731 );
not ( n235959 , n235501 );
or ( n235960 , n235958 , n235959 );
not ( n235961 , n219033 );
not ( n235962 , n38532 );
not ( n235963 , n235962 );
or ( n235964 , n235961 , n235963 );
not ( n235965 , n229704 );
nand ( n235966 , n235965 , n219034 );
nand ( n235967 , n235964 , n235966 );
nand ( n235968 , n235967 , n222185 );
nand ( n235969 , n235960 , n235968 );
xor ( n235970 , n235957 , n235969 );
not ( n235971 , n224624 );
not ( n235972 , n235520 );
or ( n235973 , n235971 , n235972 );
not ( n235974 , n219687 );
not ( n235975 , n226709 );
or ( n235976 , n235974 , n235975 );
not ( n235977 , n232842 );
nand ( n235978 , n235977 , n222323 );
nand ( n235979 , n235976 , n235978 );
nand ( n235980 , n235979 , n219314 );
nand ( n235981 , n235973 , n235980 );
xor ( n235982 , n235970 , n235981 );
xor ( n235983 , n235332 , n235982 );
xor ( n235984 , n235983 , n235791 );
xor ( n235985 , n235332 , n235982 );
and ( n235986 , n235985 , n235791 );
and ( n235987 , n235332 , n235982 );
or ( n235988 , n235986 , n235987 );
xor ( n235989 , n235338 , n235753 );
xor ( n235990 , n235989 , n235797 );
xor ( n235991 , n235338 , n235753 );
and ( n235992 , n235991 , n235797 );
and ( n235993 , n235338 , n235753 );
or ( n235994 , n235992 , n235993 );
xor ( n235995 , n235344 , n235416 );
xor ( n235996 , n235995 , n235495 );
xor ( n235997 , n235344 , n235416 );
and ( n235998 , n235997 , n235495 );
and ( n235999 , n235344 , n235416 );
or ( n236000 , n235998 , n235999 );
xor ( n236001 , n235767 , n235777 );
and ( n236002 , n236001 , n235788 );
and ( n236003 , n235767 , n235777 );
or ( n236004 , n236002 , n236003 );
xor ( n236005 , n235898 , n235468 );
xor ( n236006 , n236005 , n235828 );
xor ( n236007 , n235898 , n235468 );
and ( n236008 , n236007 , n235828 );
and ( n236009 , n235898 , n235468 );
or ( n236010 , n236008 , n236009 );
xor ( n236011 , n235984 , n235529 );
xor ( n236012 , n236011 , n235942 );
xor ( n236013 , n235984 , n235529 );
and ( n236014 , n236013 , n235942 );
and ( n236015 , n235984 , n235529 );
or ( n236016 , n236014 , n236015 );
xor ( n236017 , n235535 , n235990 );
xor ( n236018 , n236017 , n235551 );
xor ( n236019 , n235535 , n235990 );
and ( n236020 , n236019 , n235551 );
and ( n236021 , n235535 , n235990 );
or ( n236022 , n236020 , n236021 );
xor ( n236023 , n235996 , n235541 );
xor ( n236024 , n236023 , n236006 );
xor ( n236025 , n235996 , n235541 );
and ( n236026 , n236025 , n236006 );
and ( n236027 , n235996 , n235541 );
or ( n236028 , n236026 , n236027 );
xor ( n236029 , n235557 , n236012 );
xor ( n236030 , n236029 , n235563 );
xor ( n236031 , n235557 , n236012 );
and ( n236032 , n236031 , n235563 );
and ( n236033 , n235557 , n236012 );
or ( n236034 , n236032 , n236033 );
xor ( n236035 , n236018 , n235569 );
xor ( n236036 , n236035 , n236024 );
xor ( n236037 , n236018 , n235569 );
and ( n236038 , n236037 , n236024 );
and ( n236039 , n236018 , n235569 );
or ( n236040 , n236038 , n236039 );
xor ( n236041 , n236030 , n235575 );
xor ( n236042 , n236041 , n235581 );
xor ( n236043 , n236030 , n235575 );
and ( n236044 , n236043 , n235581 );
and ( n236045 , n236030 , n235575 );
or ( n236046 , n236044 , n236045 );
xor ( n236047 , n236036 , n236042 );
xor ( n236048 , n236047 , n235587 );
xor ( n236049 , n236036 , n236042 );
and ( n236050 , n236049 , n235587 );
and ( n236051 , n236036 , n236042 );
or ( n236052 , n236050 , n236051 );
xor ( n236053 , n235728 , n235739 );
and ( n236054 , n236053 , n235751 );
and ( n236055 , n235728 , n235739 );
or ( n236056 , n236054 , n236055 );
xor ( n236057 , n235903 , n235915 );
and ( n236058 , n236057 , n235927 );
and ( n236059 , n235903 , n235915 );
or ( n236060 , n236058 , n236059 );
xor ( n236061 , n235874 , n235884 );
and ( n236062 , n236061 , n235895 );
and ( n236063 , n235874 , n235884 );
or ( n236064 , n236062 , n236063 );
xor ( n236065 , n235842 , n235852 );
and ( n236066 , n236065 , n235863 );
and ( n236067 , n235842 , n235852 );
or ( n236068 , n236066 , n236067 );
xor ( n236069 , n235813 , n235399 );
and ( n236070 , n236069 , n235826 );
and ( n236071 , n235813 , n235399 );
or ( n236072 , n236070 , n236071 );
xor ( n236073 , n235247 , n235545 );
and ( n236074 , n236073 , n235939 );
and ( n236075 , n235247 , n235545 );
or ( n236076 , n236074 , n236075 );
xor ( n236077 , n235957 , n235969 );
and ( n236078 , n236077 , n235981 );
and ( n236079 , n235957 , n235969 );
or ( n236080 , n236078 , n236079 );
not ( n236081 , n235669 );
not ( n236082 , n224086 );
or ( n236083 , n236081 , n236082 );
not ( n236084 , n216311 );
not ( n236085 , n224095 );
or ( n236086 , n236084 , n236085 );
nand ( n236087 , n219899 , n226355 );
nand ( n236088 , n236086 , n236087 );
nand ( n236089 , n224090 , n236088 );
nand ( n236090 , n236083 , n236089 );
not ( n236091 , n235678 );
not ( n236092 , n233315 );
or ( n236093 , n236091 , n236092 );
not ( n236094 , n233279 );
not ( n236095 , n229795 );
or ( n236096 , n236094 , n236095 );
nand ( n236097 , n224929 , n217394 );
nand ( n236098 , n236096 , n236097 );
nand ( n236099 , n224941 , n236098 );
nand ( n236100 , n236093 , n236099 );
xor ( n236101 , n236090 , n236100 );
not ( n236102 , n235765 );
not ( n236103 , n230390 );
or ( n236104 , n236102 , n236103 );
not ( n236105 , n226225 );
not ( n236106 , n229807 );
or ( n236107 , n236105 , n236106 );
nand ( n236108 , n232962 , n234256 );
nand ( n236109 , n236107 , n236108 );
nand ( n236110 , n228775 , n236109 );
nand ( n236111 , n236104 , n236110 );
xor ( n236112 , n236101 , n236111 );
xor ( n236113 , n236090 , n236100 );
and ( n236114 , n236113 , n236111 );
and ( n236115 , n236090 , n236100 );
or ( n236116 , n236114 , n236115 );
not ( n236117 , n235775 );
not ( n236118 , n227849 );
or ( n236119 , n236117 , n236118 );
not ( n236120 , n226884 );
not ( n236121 , n226304 );
not ( n236122 , n230897 );
or ( n236123 , n236121 , n236122 );
nand ( n236124 , n226648 , n225489 );
nand ( n236125 , n236123 , n236124 );
nand ( n236126 , n236120 , n236125 );
nand ( n236127 , n236119 , n236126 );
not ( n236128 , n235640 );
not ( n236129 , n222454 );
or ( n236130 , n236128 , n236129 );
not ( n236131 , n233536 );
not ( n236132 , n222429 );
or ( n236133 , n236131 , n236132 );
not ( n236134 , n232526 );
nand ( n236135 , n236134 , n222462 );
nand ( n236136 , n236133 , n236135 );
nand ( n236137 , n236136 , n223244 );
nand ( n236138 , n236130 , n236137 );
xor ( n236139 , n236127 , n236138 );
not ( n236140 , n235726 );
not ( n236141 , n231421 );
or ( n236142 , n236140 , n236141 );
not ( n236143 , n216293 );
not ( n236144 , n233926 );
or ( n236145 , n236143 , n236144 );
nand ( n236146 , n233925 , n223658 );
nand ( n236147 , n236145 , n236146 );
nand ( n236148 , n236147 , n228868 );
nand ( n236149 , n236142 , n236148 );
xor ( n236150 , n236139 , n236149 );
xor ( n236151 , n236127 , n236138 );
and ( n236152 , n236151 , n236149 );
and ( n236153 , n236127 , n236138 );
or ( n236154 , n236152 , n236153 );
xor ( n236155 , n235651 , n235686 );
not ( n236156 , n235737 );
not ( n236157 , n229773 );
or ( n236158 , n236156 , n236157 );
not ( n236159 , n229759 );
not ( n236160 , n218980 );
and ( n236161 , n236159 , n236160 );
and ( n236162 , n229761 , n218980 );
nor ( n236163 , n236161 , n236162 );
not ( n236164 , n236163 );
nand ( n236165 , n236164 , n234378 );
nand ( n236166 , n236158 , n236165 );
not ( n236167 , n216934 );
not ( n236168 , n231753 );
or ( n236169 , n236167 , n236168 );
nand ( n236170 , n236169 , n235747 );
not ( n236171 , n236170 );
not ( n236172 , n232399 );
or ( n236173 , n236171 , n236172 );
not ( n236174 , n219102 );
not ( n236175 , n230725 );
or ( n236176 , n236174 , n236175 );
nand ( n236177 , n231232 , n216139 );
nand ( n236178 , n236176 , n236177 );
nand ( n236179 , n236178 , n232402 );
nand ( n236180 , n236173 , n236179 );
xor ( n236181 , n236166 , n236180 );
not ( n236182 , n235786 );
not ( n236183 , n233446 );
or ( n236184 , n236182 , n236183 );
not ( n236185 , n224492 );
not ( n236186 , n234394 );
or ( n236187 , n236185 , n236186 );
not ( n236188 , n227596 );
nand ( n236189 , n236188 , n225505 );
nand ( n236190 , n236187 , n236189 );
nand ( n236191 , n227737 , n236190 );
nand ( n236192 , n236184 , n236191 );
xor ( n236193 , n236181 , n236192 );
xor ( n236194 , n236155 , n236193 );
xor ( n236195 , n235651 , n235686 );
and ( n236196 , n236195 , n236193 );
and ( n236197 , n235651 , n235686 );
or ( n236198 , n236196 , n236197 );
xor ( n236199 , n236150 , n236112 );
xor ( n236200 , n236199 , n236060 );
xor ( n236201 , n236150 , n236112 );
and ( n236202 , n236201 , n236060 );
and ( n236203 , n236150 , n236112 );
or ( n236204 , n236202 , n236203 );
xor ( n236205 , n236064 , n236068 );
and ( n236206 , n233891 , n218514 );
not ( n236207 , n221637 );
and ( n236208 , n40724 , n221632 );
not ( n236209 , n40724 );
and ( n236210 , n236209 , n226388 );
or ( n236211 , n236208 , n236210 );
not ( n236212 , n236211 );
or ( n236213 , n236207 , n236212 );
not ( n236214 , n222471 );
nand ( n236215 , n236214 , n235631 );
nand ( n236216 , n236213 , n236215 );
xor ( n236217 , n236206 , n236216 );
not ( n236218 , n221266 );
not ( n236219 , n235910 );
or ( n236220 , n236218 , n236219 );
not ( n236221 , n220925 );
not ( n236222 , n220569 );
or ( n236223 , n236221 , n236222 );
nand ( n236224 , n221342 , n220901 );
nand ( n236225 , n236223 , n236224 );
nand ( n236226 , n236225 , n220930 );
nand ( n236227 , n236220 , n236226 );
xor ( n236228 , n236217 , n236227 );
xor ( n236229 , n236205 , n236228 );
xor ( n236230 , n236064 , n236068 );
and ( n236231 , n236230 , n236228 );
and ( n236232 , n236064 , n236068 );
or ( n236233 , n236231 , n236232 );
xor ( n236234 , n236072 , n236076 );
xor ( n236235 , n236234 , n236080 );
xor ( n236236 , n236072 , n236076 );
and ( n236237 , n236236 , n236080 );
and ( n236238 , n236072 , n236076 );
or ( n236239 , n236237 , n236238 );
not ( n236240 , n219076 );
not ( n236241 , n219440 );
not ( n236242 , n236241 );
not ( n236243 , n220581 );
or ( n236244 , n236242 , n236243 );
nand ( n236245 , n207936 , n219420 );
nand ( n236246 , n236244 , n236245 );
not ( n236247 , n236246 );
or ( n236248 , n236240 , n236247 );
nand ( n236249 , n235811 , n219792 );
nand ( n236250 , n236248 , n236249 );
not ( n236251 , n220164 );
not ( n236252 , n235872 );
or ( n236253 , n236251 , n236252 );
not ( n236254 , n220151 );
not ( n236255 , n40560 );
or ( n236256 , n236254 , n236255 );
nand ( n236257 , n219222 , n220290 );
nand ( n236258 , n236256 , n236257 );
nand ( n236259 , n236258 , n220881 );
nand ( n236260 , n236253 , n236259 );
xor ( n236261 , n236250 , n236260 );
not ( n236262 , n227260 );
not ( n236263 , n235925 );
or ( n236264 , n236262 , n236263 );
not ( n236265 , n226655 );
not ( n236266 , n39877 );
or ( n236267 , n236265 , n236266 );
nand ( n236268 , n235455 , n227927 );
nand ( n236269 , n236267 , n236268 );
not ( n236270 , n236269 );
not ( n236271 , n223949 );
or ( n236272 , n236270 , n236271 );
nand ( n236273 , n236264 , n236272 );
xor ( n236274 , n236261 , n236273 );
xor ( n236275 , n235716 , n236274 );
not ( n236276 , n225478 );
not ( n236277 , n235880 );
or ( n236278 , n236276 , n236277 );
not ( n236279 , n229387 );
not ( n236280 , n230490 );
or ( n236281 , n236279 , n236280 );
nand ( n236282 , n234506 , n227602 );
nand ( n236283 , n236281 , n236282 );
nand ( n236284 , n236283 , n228237 );
nand ( n236285 , n236278 , n236284 );
not ( n236286 , n229964 );
not ( n236287 , n229261 );
not ( n236288 , n222940 );
or ( n236289 , n236287 , n236288 );
not ( n236290 , n223717 );
nand ( n236291 , n236290 , n229262 );
nand ( n236292 , n236289 , n236291 );
not ( n236293 , n236292 );
or ( n236294 , n236286 , n236293 );
nand ( n236295 , n235891 , n234006 );
nand ( n236296 , n236294 , n236295 );
xor ( n236297 , n236285 , n236296 );
not ( n236298 , n220067 );
not ( n236299 , n231500 );
buf ( n236300 , n222955 );
not ( n236301 , n236300 );
not ( n236302 , n236301 );
or ( n236303 , n236299 , n236302 );
not ( n236304 , n235383 );
nand ( n236305 , n236304 , n234015 );
nand ( n236306 , n236303 , n236305 );
not ( n236307 , n236306 );
or ( n236308 , n236298 , n236307 );
nand ( n236309 , n235838 , n231018 );
nand ( n236310 , n236308 , n236309 );
xor ( n236311 , n236297 , n236310 );
xor ( n236312 , n236275 , n236311 );
xor ( n236313 , n235716 , n236274 );
and ( n236314 , n236313 , n236311 );
and ( n236315 , n235716 , n236274 );
or ( n236316 , n236314 , n236315 );
not ( n236317 , n218232 );
not ( n236318 , n233083 );
not ( n236319 , n233546 );
or ( n236320 , n236318 , n236319 );
nand ( n236321 , n230514 , n220091 );
nand ( n236322 , n236320 , n236321 );
not ( n236323 , n236322 );
or ( n236324 , n236317 , n236323 );
nand ( n236325 , n235848 , n219461 );
nand ( n236326 , n236324 , n236325 );
not ( n236327 , n223665 );
not ( n236328 , n235859 );
or ( n236329 , n236327 , n236328 );
not ( n236330 , n221241 );
not ( n236331 , n223786 );
or ( n236332 , n236330 , n236331 );
nand ( n236333 , n230527 , n221238 );
nand ( n236334 , n236332 , n236333 );
nand ( n236335 , n236334 , n218843 );
nand ( n236336 , n236329 , n236335 );
xor ( n236337 , n236326 , n236336 );
not ( n236338 , n223197 );
not ( n236339 , n235659 );
or ( n236340 , n236338 , n236339 );
not ( n236341 , n40888 );
not ( n236342 , n223182 );
or ( n236343 , n236341 , n236342 );
not ( n236344 , n223202 );
nand ( n236345 , n236344 , n223549 );
nand ( n236346 , n236343 , n236345 );
not ( n236347 , n236346 );
or ( n236348 , n236347 , n225376 );
nand ( n236349 , n236340 , n236348 );
not ( n236350 , n236349 );
xor ( n236351 , n236337 , n236350 );
xor ( n236352 , n236351 , n236194 );
xor ( n236353 , n236352 , n235757 );
xor ( n236354 , n236351 , n236194 );
and ( n236355 , n236354 , n235757 );
and ( n236356 , n236351 , n236194 );
or ( n236357 , n236355 , n236356 );
xor ( n236358 , n236004 , n236056 );
not ( n236359 , n217023 );
not ( n236360 , n235693 );
or ( n236361 , n236359 , n236360 );
not ( n236362 , n219577 );
not ( n236363 , n234579 );
or ( n236364 , n236362 , n236363 );
nand ( n236365 , n209865 , n218661 );
nand ( n236366 , n236364 , n236365 );
nand ( n236367 , n236366 , n219175 );
nand ( n236368 , n236361 , n236367 );
xor ( n236369 , n236358 , n236368 );
not ( n236370 , n222185 );
not ( n236371 , n219033 );
not ( n236372 , n228165 );
or ( n236373 , n236371 , n236372 );
nand ( n236374 , n230273 , n219034 );
nand ( n236375 , n236373 , n236374 );
not ( n236376 , n236375 );
or ( n236377 , n236370 , n236376 );
nand ( n236378 , n235967 , n219731 );
nand ( n236379 , n236377 , n236378 );
not ( n236380 , n219314 );
not ( n236381 , n219687 );
not ( n236382 , n39089 );
not ( n236383 , n236382 );
or ( n236384 , n236381 , n236383 );
nand ( n236385 , n39089 , n222323 );
nand ( n236386 , n236384 , n236385 );
not ( n236387 , n236386 );
or ( n236388 , n236380 , n236387 );
nand ( n236389 , n235979 , n224624 );
nand ( n236390 , n236388 , n236389 );
xor ( n236391 , n236379 , n236390 );
not ( n236392 , n226943 );
not ( n236393 , n235822 );
or ( n236394 , n236392 , n236393 );
not ( n236395 , n226292 );
not ( n236396 , n234350 );
or ( n236397 , n236395 , n236396 );
nand ( n236398 , n227223 , n229887 );
nand ( n236399 , n236397 , n236398 );
nand ( n236400 , n236399 , n226287 );
nand ( n236401 , n236394 , n236400 );
xor ( n236402 , n236391 , n236401 );
xor ( n236403 , n236369 , n236402 );
not ( n236404 , n216299 );
not ( n236405 , n235936 );
or ( n236406 , n236404 , n236405 );
nand ( n236407 , n214694 , n216810 );
nand ( n236408 , n236406 , n236407 );
not ( n236409 , n221933 );
not ( n236410 , n226484 );
not ( n236411 , n228216 );
or ( n236412 , n236410 , n236411 );
nand ( n236413 , n39747 , n221938 );
nand ( n236414 , n236412 , n236413 );
not ( n236415 , n236414 );
or ( n236416 , n236409 , n236415 );
nand ( n236417 , n219332 , n235702 );
nand ( n236418 , n236416 , n236417 );
xor ( n236419 , n236408 , n236418 );
not ( n236420 , n220280 );
not ( n236421 , n235955 );
or ( n236422 , n236420 , n236421 );
not ( n236423 , n234788 );
not ( n236424 , n233362 );
or ( n236425 , n236423 , n236424 );
nand ( n236426 , n229217 , n234787 );
nand ( n236427 , n236425 , n236426 );
nand ( n236428 , n236427 , n220272 );
nand ( n236429 , n236422 , n236428 );
xor ( n236430 , n236419 , n236429 );
xor ( n236431 , n236403 , n236430 );
xor ( n236432 , n236369 , n236402 );
and ( n236433 , n236432 , n236430 );
and ( n236434 , n236369 , n236402 );
or ( n236435 , n236433 , n236434 );
xor ( n236436 , n236200 , n235795 );
xor ( n236437 , n236436 , n235801 );
xor ( n236438 , n236200 , n235795 );
and ( n236439 , n236438 , n235801 );
and ( n236440 , n236200 , n235795 );
or ( n236441 , n236439 , n236440 );
xor ( n236442 , n236229 , n235832 );
xor ( n236443 , n236442 , n235902 );
xor ( n236444 , n236229 , n235832 );
and ( n236445 , n236444 , n235902 );
and ( n236446 , n236229 , n235832 );
or ( n236447 , n236445 , n236446 );
xor ( n236448 , n236235 , n236312 );
xor ( n236449 , n236448 , n235946 );
xor ( n236450 , n236235 , n236312 );
and ( n236451 , n236450 , n235946 );
and ( n236452 , n236235 , n236312 );
or ( n236453 , n236451 , n236452 );
xor ( n236454 , n236166 , n236180 );
and ( n236455 , n236454 , n236192 );
and ( n236456 , n236166 , n236180 );
or ( n236457 , n236455 , n236456 );
xor ( n236458 , n235988 , n236431 );
xor ( n236459 , n236458 , n236353 );
xor ( n236460 , n235988 , n236431 );
and ( n236461 , n236460 , n236353 );
and ( n236462 , n235988 , n236431 );
or ( n236463 , n236461 , n236462 );
xor ( n236464 , n235994 , n236437 );
xor ( n236465 , n236464 , n236000 );
xor ( n236466 , n235994 , n236437 );
and ( n236467 , n236466 , n236000 );
and ( n236468 , n235994 , n236437 );
or ( n236469 , n236467 , n236468 );
xor ( n236470 , n236443 , n236010 );
xor ( n236471 , n236470 , n236449 );
xor ( n236472 , n236443 , n236010 );
and ( n236473 , n236472 , n236449 );
and ( n236474 , n236443 , n236010 );
or ( n236475 , n236473 , n236474 );
xor ( n236476 , n236016 , n236459 );
xor ( n236477 , n236476 , n236022 );
xor ( n236478 , n236016 , n236459 );
and ( n236479 , n236478 , n236022 );
and ( n236480 , n236016 , n236459 );
or ( n236481 , n236479 , n236480 );
xor ( n236482 , n236465 , n236471 );
xor ( n236483 , n236482 , n236028 );
xor ( n236484 , n236465 , n236471 );
and ( n236485 , n236484 , n236028 );
and ( n236486 , n236465 , n236471 );
or ( n236487 , n236485 , n236486 );
xor ( n236488 , n236034 , n236477 );
xor ( n236489 , n236488 , n236040 );
xor ( n236490 , n236034 , n236477 );
and ( n236491 , n236490 , n236040 );
and ( n236492 , n236034 , n236477 );
or ( n236493 , n236491 , n236492 );
xor ( n236494 , n236483 , n236489 );
xor ( n236495 , n236494 , n236046 );
xor ( n236496 , n236483 , n236489 );
and ( n236497 , n236496 , n236046 );
and ( n236498 , n236483 , n236489 );
or ( n236499 , n236497 , n236498 );
xor ( n236500 , n236206 , n236216 );
and ( n236501 , n236500 , n236227 );
and ( n236502 , n236206 , n236216 );
or ( n236503 , n236501 , n236502 );
xor ( n236504 , n236285 , n236296 );
and ( n236505 , n236504 , n236310 );
and ( n236506 , n236285 , n236296 );
or ( n236507 , n236505 , n236506 );
xor ( n236508 , n236326 , n236336 );
and ( n236509 , n236508 , n236350 );
and ( n236510 , n236326 , n236336 );
or ( n236511 , n236509 , n236510 );
xor ( n236512 , n236250 , n236260 );
and ( n236513 , n236512 , n236273 );
and ( n236514 , n236250 , n236260 );
or ( n236515 , n236513 , n236514 );
xor ( n236516 , n236004 , n236056 );
and ( n236517 , n236516 , n236368 );
and ( n236518 , n236004 , n236056 );
or ( n236519 , n236517 , n236518 );
xor ( n236520 , n236379 , n236390 );
and ( n236521 , n236520 , n236401 );
and ( n236522 , n236379 , n236390 );
or ( n236523 , n236521 , n236522 );
xor ( n236524 , n236408 , n236418 );
and ( n236525 , n236524 , n236429 );
and ( n236526 , n236408 , n236418 );
or ( n236527 , n236525 , n236526 );
not ( n236528 , n220819 );
not ( n236529 , n216298 );
or ( n236530 , n236528 , n236529 );
nand ( n236531 , n236530 , n216810 );
not ( n236532 , n236136 );
not ( n236533 , n222886 );
or ( n236534 , n236532 , n236533 );
not ( n236535 , n222892 );
not ( n236536 , n219386 );
or ( n236537 , n236535 , n236536 );
nand ( n236538 , n222435 , n217714 );
nand ( n236539 , n236537 , n236538 );
nand ( n236540 , n236539 , n223244 );
nand ( n236541 , n236534 , n236540 );
xor ( n236542 , n236531 , n236541 );
not ( n236543 , n236346 );
not ( n236544 , n223591 );
or ( n236545 , n236543 , n236544 );
not ( n236546 , n220226 );
not ( n236547 , n223201 );
not ( n236548 , n236547 );
or ( n236549 , n236546 , n236548 );
nand ( n236550 , n223182 , n231761 );
nand ( n236551 , n236549 , n236550 );
nand ( n236552 , n236551 , n227294 );
nand ( n236553 , n236545 , n236552 );
xor ( n236554 , n236542 , n236553 );
xor ( n236555 , n236531 , n236541 );
and ( n236556 , n236555 , n236553 );
and ( n236557 , n236531 , n236541 );
or ( n236558 , n236556 , n236557 );
not ( n236559 , n236088 );
or ( n236560 , n232904 , n236559 );
and ( n236561 , n224975 , n224881 );
and ( n236562 , n217147 , n228828 );
nor ( n236563 , n236561 , n236562 );
or ( n236564 , n232476 , n236563 );
nand ( n236565 , n236560 , n236564 );
not ( n236566 , n236098 );
not ( n236567 , n233315 );
or ( n236568 , n236566 , n236567 );
not ( n236569 , n224929 );
not ( n236570 , n215989 );
and ( n236571 , n236569 , n236570 );
and ( n236572 , n232485 , n215989 );
nor ( n236573 , n236571 , n236572 );
not ( n236574 , n236573 );
nand ( n236575 , n236574 , n224941 );
nand ( n236576 , n236568 , n236575 );
xor ( n236577 , n236565 , n236576 );
not ( n236578 , n236109 );
or ( n236579 , n231453 , n236578 );
not ( n236580 , n41565 );
and ( n236581 , n236580 , n232494 );
not ( n236582 , n236580 );
and ( n236583 , n236582 , n229807 );
nor ( n236584 , n236581 , n236583 );
or ( n236585 , n236584 , n231456 );
nand ( n236586 , n236579 , n236585 );
xor ( n236587 , n236577 , n236586 );
xor ( n236588 , n236565 , n236576 );
and ( n236589 , n236588 , n236586 );
and ( n236590 , n236565 , n236576 );
or ( n236591 , n236589 , n236590 );
xor ( n236592 , n236116 , n236154 );
xor ( n236593 , n236592 , n236554 );
xor ( n236594 , n236116 , n236154 );
and ( n236595 , n236594 , n236554 );
and ( n236596 , n236116 , n236154 );
or ( n236597 , n236595 , n236596 );
or ( n236598 , n231994 , n236163 );
and ( n236599 , n231477 , n221495 );
and ( n236600 , n229761 , n220022 );
nor ( n236601 , n236599 , n236600 );
or ( n236602 , n231476 , n236601 );
nand ( n236603 , n236598 , n236602 );
not ( n236604 , n236178 );
not ( n236605 , n233879 );
or ( n236606 , n236604 , n236605 );
not ( n236607 , n219343 );
not ( n236608 , n230725 );
or ( n236609 , n236607 , n236608 );
nand ( n236610 , n231232 , n223269 );
nand ( n236611 , n236609 , n236610 );
nand ( n236612 , n232402 , n236611 );
nand ( n236613 , n236606 , n236612 );
xor ( n236614 , n236603 , n236613 );
not ( n236615 , n230722 );
and ( n236616 , n236615 , n216934 );
xor ( n236617 , n236614 , n236616 );
not ( n236618 , n236125 );
not ( n236619 , n229816 );
or ( n236620 , n236618 , n236619 );
not ( n236621 , n225768 );
not ( n236622 , n232431 );
or ( n236623 , n236621 , n236622 );
not ( n236624 , n230897 );
nand ( n236625 , n236624 , n225769 );
nand ( n236626 , n236623 , n236625 );
nand ( n236627 , n226885 , n236626 );
nand ( n236628 , n236620 , n236627 );
not ( n236629 , n236190 );
not ( n236630 , n232440 );
or ( n236631 , n236629 , n236630 );
not ( n236632 , n214837 );
not ( n236633 , n233451 );
or ( n236634 , n236632 , n236633 );
nand ( n236635 , n233450 , n231913 );
nand ( n236636 , n236634 , n236635 );
nand ( n236637 , n227737 , n236636 );
nand ( n236638 , n236631 , n236637 );
xor ( n236639 , n236628 , n236638 );
not ( n236640 , n236147 );
not ( n236641 , n231421 );
or ( n236642 , n236640 , n236641 );
not ( n236643 , n233925 );
and ( n236644 , n224037 , n236643 );
not ( n236645 , n224037 );
and ( n236646 , n236645 , n233925 );
or ( n236647 , n236644 , n236646 );
nand ( n236648 , n229738 , n236647 );
nand ( n236649 , n236642 , n236648 );
xor ( n236650 , n236639 , n236649 );
xor ( n236651 , n236617 , n236650 );
xor ( n236652 , n236651 , n236587 );
xor ( n236653 , n236617 , n236650 );
and ( n236654 , n236653 , n236587 );
and ( n236655 , n236617 , n236650 );
or ( n236656 , n236654 , n236655 );
xor ( n236657 , n236503 , n236507 );
xor ( n236658 , n236657 , n236511 );
xor ( n236659 , n236503 , n236507 );
and ( n236660 , n236659 , n236511 );
and ( n236661 , n236503 , n236507 );
or ( n236662 , n236660 , n236661 );
xor ( n236663 , n236515 , n236519 );
xor ( n236664 , n236663 , n236523 );
xor ( n236665 , n236515 , n236519 );
and ( n236666 , n236665 , n236523 );
and ( n236667 , n236515 , n236519 );
or ( n236668 , n236666 , n236667 );
not ( n236669 , n219449 );
not ( n236670 , n236334 );
or ( n236671 , n236669 , n236670 );
not ( n236672 , n218456 );
not ( n236673 , n232413 );
not ( n236674 , n40258 );
or ( n236675 , n236673 , n236674 );
or ( n236676 , n40258 , n232413 );
nand ( n236677 , n236675 , n236676 );
nand ( n236678 , n236672 , n236677 );
nand ( n236679 , n236671 , n236678 );
not ( n236680 , n219076 );
and ( n236681 , n221725 , n219424 );
not ( n236682 , n221725 );
and ( n236683 , n236682 , n219420 );
or ( n236684 , n236681 , n236683 );
not ( n236685 , n236684 );
or ( n236686 , n236680 , n236685 );
nand ( n236687 , n220507 , n236246 );
nand ( n236688 , n236686 , n236687 );
xor ( n236689 , n236679 , n236688 );
xor ( n236690 , n236689 , n236349 );
xor ( n236691 , n236527 , n236690 );
not ( n236692 , n234006 );
not ( n236693 , n236292 );
or ( n236694 , n236692 , n236693 );
not ( n236695 , n229261 );
not ( n236696 , n223330 );
or ( n236697 , n236695 , n236696 );
nand ( n236698 , n223333 , n229262 );
nand ( n236699 , n236697 , n236698 );
nand ( n236700 , n236699 , n229964 );
nand ( n236701 , n236694 , n236700 );
not ( n236702 , n231018 );
not ( n236703 , n236306 );
or ( n236704 , n236702 , n236703 );
not ( n236705 , n217614 );
not ( n236706 , n233035 );
or ( n236707 , n236705 , n236706 );
nand ( n236708 , n222513 , n234015 );
nand ( n236709 , n236707 , n236708 );
nand ( n236710 , n236709 , n220067 );
nand ( n236711 , n236704 , n236710 );
xor ( n236712 , n236701 , n236711 );
not ( n236713 , n219461 );
not ( n236714 , n236322 );
or ( n236715 , n236713 , n236714 );
not ( n236716 , n233083 );
not ( n236717 , n221712 );
or ( n236718 , n236716 , n236717 );
not ( n236719 , n229936 );
nand ( n236720 , n236719 , n234949 );
nand ( n236721 , n236718 , n236720 );
nand ( n236722 , n218232 , n236721 );
nand ( n236723 , n236715 , n236722 );
xor ( n236724 , n236712 , n236723 );
xor ( n236725 , n236691 , n236724 );
xor ( n236726 , n236527 , n236690 );
and ( n236727 , n236726 , n236724 );
and ( n236728 , n236527 , n236690 );
or ( n236729 , n236727 , n236728 );
not ( n236730 , n221637 );
not ( n236731 , n221608 );
not ( n236732 , n219595 );
or ( n236733 , n236731 , n236732 );
nand ( n236734 , n40710 , n221632 );
nand ( n236735 , n236733 , n236734 );
not ( n236736 , n236735 );
or ( n236737 , n236730 , n236736 );
nand ( n236738 , n236211 , n221626 );
nand ( n236739 , n236737 , n236738 );
not ( n236740 , n229395 );
not ( n236741 , n236283 );
or ( n236742 , n236740 , n236741 );
not ( n236743 , n229387 );
not ( n236744 , n225108 );
or ( n236745 , n236743 , n236744 );
nand ( n236746 , n226964 , n227602 );
nand ( n236747 , n236745 , n236746 );
nand ( n236748 , n236747 , n228237 );
nand ( n236749 , n236742 , n236748 );
xor ( n236750 , n236739 , n236749 );
not ( n236751 , n220930 );
buf ( n236752 , n220203 );
not ( n236753 , n236752 );
not ( n236754 , n220906 );
not ( n236755 , n236754 );
or ( n236756 , n236753 , n236755 );
nand ( n236757 , n220925 , n219532 );
nand ( n236758 , n236756 , n236757 );
not ( n236759 , n236758 );
or ( n236760 , n236751 , n236759 );
nand ( n236761 , n236225 , n235913 );
nand ( n236762 , n236760 , n236761 );
xor ( n236763 , n236750 , n236762 );
xor ( n236764 , n236763 , n236593 );
not ( n236765 , n220164 );
not ( n236766 , n236258 );
or ( n236767 , n236765 , n236766 );
not ( n236768 , n222414 );
not ( n236769 , n236768 );
not ( n236770 , n221687 );
or ( n236771 , n236769 , n236770 );
nand ( n236772 , n221690 , n220147 );
nand ( n236773 , n236771 , n236772 );
nand ( n236774 , n236773 , n220881 );
nand ( n236775 , n236767 , n236774 );
not ( n236776 , n227260 );
not ( n236777 , n236269 );
or ( n236778 , n236776 , n236777 );
not ( n236779 , n226655 );
not ( n236780 , n39927 );
or ( n236781 , n236779 , n236780 );
nand ( n236782 , n226723 , n227927 );
nand ( n236783 , n236781 , n236782 );
nand ( n236784 , n236783 , n223949 );
nand ( n236785 , n236778 , n236784 );
xor ( n236786 , n236775 , n236785 );
xor ( n236787 , n236786 , n236457 );
xor ( n236788 , n236764 , n236787 );
xor ( n236789 , n236763 , n236593 );
and ( n236790 , n236789 , n236787 );
and ( n236791 , n236763 , n236593 );
or ( n236792 , n236790 , n236791 );
not ( n236793 , n219332 );
not ( n236794 , n236414 );
or ( n236795 , n236793 , n236794 );
not ( n236796 , n221935 );
not ( n236797 , n226712 );
or ( n236798 , n236796 , n236797 );
nand ( n236799 , n39607 , n222333 );
nand ( n236800 , n236798 , n236799 );
nand ( n236801 , n236800 , n221933 );
nand ( n236802 , n236795 , n236801 );
not ( n236803 , n220280 );
not ( n236804 , n236427 );
or ( n236805 , n236803 , n236804 );
not ( n236806 , n225120 );
not ( n236807 , n209709 );
or ( n236808 , n236806 , n236807 );
nand ( n236809 , n232856 , n234787 );
nand ( n236810 , n236808 , n236809 );
nand ( n236811 , n236810 , n219353 );
nand ( n236812 , n236805 , n236811 );
xor ( n236813 , n236802 , n236812 );
not ( n236814 , n226287 );
not ( n236815 , n227912 );
not ( n236816 , n229667 );
or ( n236817 , n236815 , n236816 );
nand ( n236818 , n233856 , n220038 );
nand ( n236819 , n236817 , n236818 );
not ( n236820 , n236819 );
or ( n236821 , n236814 , n236820 );
nand ( n236822 , n236399 , n220414 );
nand ( n236823 , n236821 , n236822 );
xor ( n236824 , n236813 , n236823 );
xor ( n236825 , n236198 , n236824 );
not ( n236826 , n219175 );
not ( n236827 , n219577 );
not ( n236828 , n233134 );
or ( n236829 , n236827 , n236828 );
not ( n236830 , n231097 );
nand ( n236831 , n236830 , n218661 );
nand ( n236832 , n236829 , n236831 );
not ( n236833 , n236832 );
or ( n236834 , n236826 , n236833 );
nand ( n236835 , n236366 , n217023 );
nand ( n236836 , n236834 , n236835 );
not ( n236837 , n219731 );
not ( n236838 , n236375 );
or ( n236839 , n236837 , n236838 );
buf ( n236840 , n39286 );
not ( n236841 , n236840 );
not ( n236842 , n219034 );
or ( n236843 , n236841 , n236842 );
not ( n236844 , n236840 );
nand ( n236845 , n236844 , n219033 );
nand ( n236846 , n236843 , n236845 );
nand ( n236847 , n236846 , n222185 );
nand ( n236848 , n236839 , n236847 );
xor ( n236849 , n236836 , n236848 );
not ( n236850 , n236386 );
or ( n236851 , n236850 , n223825 );
and ( n236852 , n235962 , n219687 );
not ( n236853 , n235962 );
and ( n236854 , n236853 , n222323 );
or ( n236855 , n236852 , n236854 );
not ( n236856 , n236855 );
or ( n236857 , n236856 , n223833 );
nand ( n236858 , n236851 , n236857 );
xor ( n236859 , n236849 , n236858 );
xor ( n236860 , n236825 , n236859 );
xor ( n236861 , n236198 , n236824 );
and ( n236862 , n236861 , n236859 );
and ( n236863 , n236198 , n236824 );
or ( n236864 , n236862 , n236863 );
xor ( n236865 , n236233 , n236652 );
xor ( n236866 , n236865 , n236204 );
xor ( n236867 , n236233 , n236652 );
and ( n236868 , n236867 , n236204 );
and ( n236869 , n236233 , n236652 );
or ( n236870 , n236868 , n236869 );
xor ( n236871 , n236658 , n236239 );
xor ( n236872 , n236871 , n236316 );
xor ( n236873 , n236658 , n236239 );
and ( n236874 , n236873 , n236316 );
and ( n236875 , n236658 , n236239 );
or ( n236876 , n236874 , n236875 );
xor ( n236877 , n236664 , n236435 );
xor ( n236878 , n236877 , n236357 );
xor ( n236879 , n236664 , n236435 );
and ( n236880 , n236879 , n236357 );
and ( n236881 , n236664 , n236435 );
or ( n236882 , n236880 , n236881 );
xor ( n236883 , n236628 , n236638 );
and ( n236884 , n236883 , n236649 );
and ( n236885 , n236628 , n236638 );
or ( n236886 , n236884 , n236885 );
xor ( n236887 , n236725 , n236860 );
xor ( n236888 , n236887 , n236788 );
xor ( n236889 , n236725 , n236860 );
and ( n236890 , n236889 , n236788 );
and ( n236891 , n236725 , n236860 );
or ( n236892 , n236890 , n236891 );
xor ( n236893 , n236447 , n236866 );
xor ( n236894 , n236893 , n236441 );
xor ( n236895 , n236447 , n236866 );
and ( n236896 , n236895 , n236441 );
and ( n236897 , n236447 , n236866 );
or ( n236898 , n236896 , n236897 );
xor ( n236899 , n236453 , n236872 );
xor ( n236900 , n236899 , n236878 );
xor ( n236901 , n236453 , n236872 );
and ( n236902 , n236901 , n236878 );
and ( n236903 , n236453 , n236872 );
or ( n236904 , n236902 , n236903 );
xor ( n236905 , n236463 , n236888 );
xor ( n236906 , n236905 , n236469 );
xor ( n236907 , n236463 , n236888 );
and ( n236908 , n236907 , n236469 );
and ( n236909 , n236463 , n236888 );
or ( n236910 , n236908 , n236909 );
xor ( n236911 , n236894 , n236475 );
xor ( n236912 , n236911 , n236900 );
xor ( n236913 , n236894 , n236475 );
and ( n236914 , n236913 , n236900 );
and ( n236915 , n236894 , n236475 );
or ( n236916 , n236914 , n236915 );
xor ( n236917 , n236481 , n236906 );
xor ( n236918 , n236917 , n236487 );
xor ( n236919 , n236481 , n236906 );
and ( n236920 , n236919 , n236487 );
and ( n236921 , n236481 , n236906 );
or ( n236922 , n236920 , n236921 );
xor ( n236923 , n236912 , n236918 );
xor ( n236924 , n236923 , n236493 );
xor ( n236925 , n236912 , n236918 );
and ( n236926 , n236925 , n236493 );
and ( n236927 , n236912 , n236918 );
or ( n236928 , n236926 , n236927 );
xor ( n236929 , n236603 , n236613 );
and ( n236930 , n236929 , n236616 );
and ( n236931 , n236603 , n236613 );
or ( n236932 , n236930 , n236931 );
xor ( n236933 , n236739 , n236749 );
and ( n236934 , n236933 , n236762 );
and ( n236935 , n236739 , n236749 );
or ( n236936 , n236934 , n236935 );
xor ( n236937 , n236701 , n236711 );
and ( n236938 , n236937 , n236723 );
and ( n236939 , n236701 , n236711 );
or ( n236940 , n236938 , n236939 );
xor ( n236941 , n236679 , n236688 );
and ( n236942 , n236941 , n236349 );
and ( n236943 , n236679 , n236688 );
or ( n236944 , n236942 , n236943 );
xor ( n236945 , n236775 , n236785 );
and ( n236946 , n236945 , n236457 );
and ( n236947 , n236775 , n236785 );
or ( n236948 , n236946 , n236947 );
xor ( n236949 , n236836 , n236848 );
and ( n236950 , n236949 , n236858 );
and ( n236951 , n236836 , n236848 );
or ( n236952 , n236950 , n236951 );
xor ( n236953 , n236802 , n236812 );
and ( n236954 , n236953 , n236823 );
and ( n236955 , n236802 , n236812 );
or ( n236956 , n236954 , n236955 );
or ( n236957 , n235195 , n236573 );
not ( n236958 , n224941 );
and ( n236959 , n219902 , n229795 );
not ( n236960 , n219902 );
and ( n236961 , n236960 , n232485 );
nor ( n236962 , n236959 , n236961 );
or ( n236963 , n236958 , n236962 );
nand ( n236964 , n236957 , n236963 );
not ( n236965 , n236584 );
not ( n236966 , n236965 );
not ( n236967 , n232956 );
or ( n236968 , n236966 , n236967 );
not ( n236969 , n215796 );
not ( n236970 , n233962 );
or ( n236971 , n236969 , n236970 );
nand ( n236972 , n232494 , n216261 );
nand ( n236973 , n236971 , n236972 );
nand ( n236974 , n228775 , n236973 );
nand ( n236975 , n236968 , n236974 );
xor ( n236976 , n236964 , n236975 );
not ( n236977 , n236626 );
or ( n236978 , n234290 , n236977 );
and ( n236979 , n234257 , n234293 );
not ( n236980 , n234257 );
and ( n236981 , n236980 , n232974 );
nor ( n236982 , n236979 , n236981 );
or ( n236983 , n234896 , n236982 );
nand ( n236984 , n236978 , n236983 );
xor ( n236985 , n236976 , n236984 );
xor ( n236986 , n236964 , n236975 );
and ( n236987 , n236986 , n236984 );
and ( n236988 , n236964 , n236975 );
or ( n236989 , n236987 , n236988 );
not ( n236990 , n236636 );
not ( n236991 , n232440 );
or ( n236992 , n236990 , n236991 );
and ( n236993 , n225490 , n233451 );
not ( n236994 , n225490 );
and ( n236995 , n236994 , n233450 );
nor ( n236996 , n236993 , n236995 );
or ( n236997 , n228273 , n236996 );
nand ( n236998 , n236992 , n236997 );
not ( n236999 , n236551 );
not ( n237000 , n223591 );
or ( n237001 , n236999 , n237000 );
not ( n237002 , n217331 );
not ( n237003 , n223183 );
or ( n237004 , n237002 , n237003 );
not ( n237005 , n223156 );
nand ( n237006 , n217330 , n237005 );
nand ( n237007 , n237004 , n237006 );
nand ( n237008 , n227294 , n237007 );
nand ( n237009 , n237001 , n237008 );
xor ( n237010 , n236998 , n237009 );
or ( n237011 , n231474 , n236601 );
not ( n237012 , n231476 );
not ( n237013 , n237012 );
not ( n237014 , n231480 );
and ( n237015 , n216293 , n237014 );
not ( n237016 , n216293 );
not ( n237017 , n229762 );
and ( n237018 , n237016 , n237017 );
nor ( n237019 , n237015 , n237018 );
or ( n237020 , n237013 , n237019 );
nand ( n237021 , n237011 , n237020 );
xor ( n237022 , n237010 , n237021 );
xor ( n237023 , n236998 , n237009 );
and ( n237024 , n237023 , n237021 );
and ( n237025 , n236998 , n237009 );
or ( n237026 , n237024 , n237025 );
not ( n237027 , n236611 );
not ( n237028 , n232399 );
or ( n237029 , n237027 , n237028 );
and ( n237030 , n221921 , n232404 );
not ( n237031 , n221921 );
and ( n237032 , n237031 , n232784 );
or ( n237033 , n237030 , n237032 );
nand ( n237034 , n237033 , n232402 );
nand ( n237035 , n237029 , n237034 );
and ( n237036 , n234382 , n219102 );
xor ( n237037 , n237035 , n237036 );
buf ( n237038 , n228859 );
not ( n237039 , n236647 );
or ( n237040 , n237038 , n237039 );
not ( n237041 , n228868 );
and ( n237042 , n224492 , n228847 );
not ( n237043 , n224492 );
and ( n237044 , n237043 , n228850 );
or ( n237045 , n237042 , n237044 );
not ( n237046 , n237045 );
or ( n237047 , n237041 , n237046 );
nand ( n237048 , n237040 , n237047 );
xor ( n237049 , n237037 , n237048 );
xor ( n237050 , n236886 , n237049 );
xor ( n237051 , n237050 , n237022 );
xor ( n237052 , n236886 , n237049 );
and ( n237053 , n237052 , n237022 );
and ( n237054 , n236886 , n237049 );
or ( n237055 , n237053 , n237054 );
xor ( n237056 , n236985 , n236936 );
xor ( n237057 , n237056 , n236940 );
xor ( n237058 , n236985 , n236936 );
and ( n237059 , n237058 , n236940 );
and ( n237060 , n236985 , n236936 );
or ( n237061 , n237059 , n237060 );
xor ( n237062 , n236944 , n236948 );
xor ( n237063 , n237062 , n236952 );
xor ( n237064 , n236944 , n236948 );
and ( n237065 , n237064 , n236952 );
and ( n237066 , n236944 , n236948 );
or ( n237067 , n237065 , n237066 );
not ( n237068 , n219449 );
not ( n237069 , n236677 );
or ( n237070 , n237068 , n237069 );
nand ( n237071 , n226505 , n218876 );
not ( n237072 , n237071 );
nand ( n237073 , n233546 , n232413 );
not ( n237074 , n237073 );
or ( n237075 , n237072 , n237074 );
nand ( n237076 , n237075 , n218843 );
nand ( n237077 , n237070 , n237076 );
not ( n237078 , n219435 );
not ( n237079 , n236684 );
or ( n237080 , n237078 , n237079 );
not ( n237081 , n219424 );
not ( n237082 , n220596 );
or ( n237083 , n237081 , n237082 );
not ( n237084 , n221330 );
nand ( n237085 , n237084 , n219420 );
nand ( n237086 , n237083 , n237085 );
nand ( n237087 , n237086 , n219076 );
nand ( n237088 , n237080 , n237087 );
xor ( n237089 , n237077 , n237088 );
not ( n237090 , n220881 );
and ( n237091 , n220581 , n220150 );
not ( n237092 , n220581 );
and ( n237093 , n237092 , n222414 );
or ( n237094 , n237091 , n237093 );
not ( n237095 , n237094 );
or ( n237096 , n237090 , n237095 );
nand ( n237097 , n236773 , n220164 );
nand ( n237098 , n237096 , n237097 );
xor ( n237099 , n237089 , n237098 );
xor ( n237100 , n236956 , n237099 );
not ( n237101 , n220067 );
not ( n237102 , n222940 );
not ( n237103 , n231500 );
or ( n237104 , n237102 , n237103 );
nand ( n237105 , n223722 , n231501 );
nand ( n237106 , n237104 , n237105 );
not ( n237107 , n237106 );
or ( n237108 , n237101 , n237107 );
nand ( n237109 , n236709 , n231018 );
nand ( n237110 , n237108 , n237109 );
not ( n237111 , n219461 );
not ( n237112 , n236721 );
or ( n237113 , n237111 , n237112 );
not ( n237114 , n218771 );
not ( n237115 , n223748 );
or ( n237116 , n237114 , n237115 );
nand ( n237117 , n222101 , n220091 );
nand ( n237118 , n237116 , n237117 );
nand ( n237119 , n237118 , n218232 );
nand ( n237120 , n237113 , n237119 );
xor ( n237121 , n237110 , n237120 );
not ( n237122 , n236563 );
not ( n237123 , n237122 );
not ( n237124 , n224087 );
or ( n237125 , n237123 , n237124 );
not ( n237126 , n219050 );
not ( n237127 , n224095 );
or ( n237128 , n237126 , n237127 );
buf ( n237129 , n224069 );
not ( n237130 , n237129 );
nand ( n237131 , n237130 , n40888 );
nand ( n237132 , n237128 , n237131 );
nand ( n237133 , n224090 , n237132 );
nand ( n237134 , n237125 , n237133 );
not ( n237135 , n237134 );
xor ( n237136 , n237121 , n237135 );
xor ( n237137 , n237100 , n237136 );
xor ( n237138 , n236956 , n237099 );
and ( n237139 , n237138 , n237136 );
and ( n237140 , n236956 , n237099 );
or ( n237141 , n237139 , n237140 );
not ( n237142 , n222158 );
not ( n237143 , n222434 );
not ( n237144 , n217964 );
or ( n237145 , n237143 , n237144 );
nand ( n237146 , n208002 , n222429 );
nand ( n237147 , n237145 , n237146 );
not ( n237148 , n237147 );
or ( n237149 , n237142 , n237148 );
nand ( n237150 , n222886 , n236539 );
nand ( n237151 , n237149 , n237150 );
not ( n237152 , n221637 );
not ( n237153 , n221633 );
not ( n237154 , n40768 );
or ( n237155 , n237153 , n237154 );
not ( n237156 , n226388 );
nand ( n237157 , n237156 , n224642 );
nand ( n237158 , n237155 , n237157 );
not ( n237159 , n237158 );
or ( n237160 , n237152 , n237159 );
nand ( n237161 , n236735 , n221626 );
nand ( n237162 , n237160 , n237161 );
xor ( n237163 , n237151 , n237162 );
not ( n237164 , n234006 );
not ( n237165 , n236699 );
or ( n237166 , n237164 , n237165 );
xor ( n237167 , n229261 , n234506 );
nand ( n237168 , n229964 , n237167 );
nand ( n237169 , n237166 , n237168 );
xor ( n237170 , n237163 , n237169 );
not ( n237171 , n223949 );
not ( n237172 , n226655 );
not ( n237173 , n234347 );
or ( n237174 , n237172 , n237173 );
nand ( n237175 , n227223 , n227927 );
nand ( n237176 , n237174 , n237175 );
not ( n237177 , n237176 );
or ( n237178 , n237171 , n237177 );
nand ( n237179 , n236783 , n227260 );
nand ( n237180 , n237178 , n237179 );
xor ( n237181 , n237180 , n236558 );
xor ( n237182 , n237181 , n236591 );
xor ( n237183 , n237170 , n237182 );
xor ( n237184 , n237183 , n236597 );
xor ( n237185 , n237170 , n237182 );
and ( n237186 , n237185 , n236597 );
and ( n237187 , n237170 , n237182 );
or ( n237188 , n237186 , n237187 );
not ( n237189 , n221266 );
not ( n237190 , n236758 );
or ( n237191 , n237189 , n237190 );
not ( n237192 , n222399 );
not ( n237193 , n40560 );
or ( n237194 , n237192 , n237193 );
nand ( n237195 , n219226 , n236754 );
nand ( n237196 , n237194 , n237195 );
nand ( n237197 , n237196 , n220930 );
nand ( n237198 , n237191 , n237197 );
not ( n237199 , n228237 );
not ( n237200 , n233544 );
not ( n237201 , n230280 );
or ( n237202 , n237200 , n237201 );
not ( n237203 , n233544 );
nand ( n237204 , n39878 , n237203 );
nand ( n237205 , n237202 , n237204 );
not ( n237206 , n237205 );
or ( n237207 , n237199 , n237206 );
nand ( n237208 , n236747 , n225478 );
nand ( n237209 , n237207 , n237208 );
xor ( n237210 , n237198 , n237209 );
xor ( n237211 , n237210 , n236932 );
xor ( n237212 , n237211 , n236656 );
not ( n237213 , n220272 );
not ( n237214 , n234787 );
not ( n237215 , n209865 );
or ( n237216 , n237214 , n237215 );
nand ( n237217 , n225120 , n234579 );
nand ( n237218 , n237216 , n237217 );
not ( n237219 , n237218 );
or ( n237220 , n237213 , n237219 );
nand ( n237221 , n236810 , n220280 );
nand ( n237222 , n237220 , n237221 );
not ( n237223 , n224624 );
not ( n237224 , n236855 );
or ( n237225 , n237223 , n237224 );
not ( n237226 , n219687 );
not ( n237227 , n39366 );
or ( n237228 , n237226 , n237227 );
not ( n237229 , n228165 );
nand ( n237230 , n237229 , n222323 );
nand ( n237231 , n237228 , n237230 );
nand ( n237232 , n237231 , n219314 );
nand ( n237233 , n237225 , n237232 );
xor ( n237234 , n237222 , n237233 );
not ( n237235 , n221933 );
not ( n237236 , n226484 );
not ( n237237 , n228184 );
or ( n237238 , n237236 , n237237 );
nand ( n237239 , n230462 , n221938 );
nand ( n237240 , n237238 , n237239 );
not ( n237241 , n237240 );
or ( n237242 , n237235 , n237241 );
nand ( n237243 , n236800 , n219332 );
nand ( n237244 , n237242 , n237243 );
xor ( n237245 , n237234 , n237244 );
xor ( n237246 , n237212 , n237245 );
xor ( n237247 , n237211 , n236656 );
and ( n237248 , n237247 , n237245 );
and ( n237249 , n237211 , n236656 );
or ( n237250 , n237248 , n237249 );
not ( n237251 , n217023 );
not ( n237252 , n236832 );
or ( n237253 , n237251 , n237252 );
nand ( n237254 , n219175 , n217017 );
nand ( n237255 , n237253 , n237254 );
not ( n237256 , n220414 );
not ( n237257 , n236819 );
or ( n237258 , n237256 , n237257 );
not ( n237259 , n227912 );
not ( n237260 , n230241 );
or ( n237261 , n237259 , n237260 );
nand ( n237262 , n39747 , n229887 );
nand ( n237263 , n237261 , n237262 );
nand ( n237264 , n237263 , n226287 );
nand ( n237265 , n237258 , n237264 );
xor ( n237266 , n237255 , n237265 );
not ( n237267 , n222185 );
not ( n237268 , n219033 );
not ( n237269 , n230219 );
or ( n237270 , n237268 , n237269 );
buf ( n237271 , n230219 );
not ( n237272 , n237271 );
nand ( n237273 , n237272 , n219034 );
nand ( n237274 , n237270 , n237273 );
not ( n237275 , n237274 );
or ( n237276 , n237267 , n237275 );
nand ( n237277 , n219731 , n236846 );
nand ( n237278 , n237276 , n237277 );
xor ( n237279 , n237266 , n237278 );
xor ( n237280 , n237279 , n237051 );
xor ( n237281 , n237280 , n236662 );
xor ( n237282 , n237279 , n237051 );
and ( n237283 , n237282 , n236662 );
and ( n237284 , n237279 , n237051 );
or ( n237285 , n237283 , n237284 );
xor ( n237286 , n236668 , n236729 );
xor ( n237287 , n237286 , n237057 );
xor ( n237288 , n236668 , n236729 );
and ( n237289 , n237288 , n237057 );
and ( n237290 , n236668 , n236729 );
or ( n237291 , n237289 , n237290 );
xor ( n237292 , n236792 , n237063 );
xor ( n237293 , n237292 , n236864 );
xor ( n237294 , n236792 , n237063 );
and ( n237295 , n237294 , n236864 );
and ( n237296 , n236792 , n237063 );
or ( n237297 , n237295 , n237296 );
xor ( n237298 , n237137 , n236870 );
xor ( n237299 , n237298 , n237246 );
xor ( n237300 , n237137 , n236870 );
and ( n237301 , n237300 , n237246 );
and ( n237302 , n237137 , n236870 );
or ( n237303 , n237301 , n237302 );
xor ( n237304 , n237035 , n237036 );
and ( n237305 , n237304 , n237048 );
and ( n237306 , n237035 , n237036 );
or ( n237307 , n237305 , n237306 );
xor ( n237308 , n237184 , n236876 );
xor ( n237309 , n237308 , n237281 );
xor ( n237310 , n237184 , n236876 );
and ( n237311 , n237310 , n237281 );
and ( n237312 , n237184 , n236876 );
or ( n237313 , n237311 , n237312 );
xor ( n237314 , n237287 , n236882 );
xor ( n237315 , n237314 , n237293 );
xor ( n237316 , n237287 , n236882 );
and ( n237317 , n237316 , n237293 );
and ( n237318 , n237287 , n236882 );
or ( n237319 , n237317 , n237318 );
xor ( n237320 , n236892 , n237299 );
xor ( n237321 , n237320 , n236898 );
xor ( n237322 , n236892 , n237299 );
and ( n237323 , n237322 , n236898 );
and ( n237324 , n236892 , n237299 );
or ( n237325 , n237323 , n237324 );
xor ( n237326 , n237309 , n237315 );
xor ( n237327 , n237326 , n236904 );
xor ( n237328 , n237309 , n237315 );
and ( n237329 , n237328 , n236904 );
and ( n237330 , n237309 , n237315 );
or ( n237331 , n237329 , n237330 );
xor ( n237332 , n237321 , n236910 );
xor ( n237333 , n237332 , n236916 );
xor ( n237334 , n237321 , n236910 );
and ( n237335 , n237334 , n236916 );
and ( n237336 , n237321 , n236910 );
or ( n237337 , n237335 , n237336 );
xor ( n237338 , n237327 , n237333 );
xor ( n237339 , n237338 , n236922 );
xor ( n237340 , n237327 , n237333 );
and ( n237341 , n237340 , n236922 );
and ( n237342 , n237327 , n237333 );
or ( n237343 , n237341 , n237342 );
xor ( n237344 , n237151 , n237162 );
and ( n237345 , n237344 , n237169 );
and ( n237346 , n237151 , n237162 );
or ( n237347 , n237345 , n237346 );
xor ( n237348 , n237110 , n237120 );
and ( n237349 , n237348 , n237135 );
and ( n237350 , n237110 , n237120 );
or ( n237351 , n237349 , n237350 );
xor ( n237352 , n237077 , n237088 );
and ( n237353 , n237352 , n237098 );
and ( n237354 , n237077 , n237088 );
or ( n237355 , n237353 , n237354 );
xor ( n237356 , n237198 , n237209 );
and ( n237357 , n237356 , n236932 );
and ( n237358 , n237198 , n237209 );
or ( n237359 , n237357 , n237358 );
xor ( n237360 , n237222 , n237233 );
and ( n237361 , n237360 , n237244 );
and ( n237362 , n237222 , n237233 );
or ( n237363 , n237361 , n237362 );
xor ( n237364 , n237255 , n237265 );
and ( n237365 , n237364 , n237278 );
and ( n237366 , n237255 , n237265 );
or ( n237367 , n237365 , n237366 );
xor ( n237368 , n237180 , n236558 );
and ( n237369 , n237368 , n236591 );
and ( n237370 , n237180 , n236558 );
or ( n237371 , n237369 , n237370 );
not ( n237372 , n227943 );
not ( n237373 , n217367 );
or ( n237374 , n237372 , n237373 );
nand ( n237375 , n237374 , n219577 );
not ( n237376 , n237007 );
not ( n237377 , n223591 );
or ( n237378 , n237376 , n237377 );
not ( n237379 , n223182 );
not ( n237380 , n220823 );
or ( n237381 , n237379 , n237380 );
nand ( n237382 , n219389 , n236547 );
nand ( n237383 , n237381 , n237382 );
nand ( n237384 , n237383 , n222768 );
nand ( n237385 , n237378 , n237384 );
xor ( n237386 , n237375 , n237385 );
not ( n237387 , n237132 );
not ( n237388 , n224087 );
or ( n237389 , n237387 , n237388 );
not ( n237390 , n233309 );
not ( n237391 , n231761 );
or ( n237392 , n237390 , n237391 );
buf ( n237393 , n220226 );
nand ( n237394 , n237129 , n237393 );
nand ( n237395 , n237392 , n237394 );
nand ( n237396 , n224090 , n237395 );
nand ( n237397 , n237389 , n237396 );
xor ( n237398 , n237386 , n237397 );
xor ( n237399 , n237375 , n237385 );
and ( n237400 , n237399 , n237397 );
and ( n237401 , n237375 , n237385 );
or ( n237402 , n237400 , n237401 );
or ( n237403 , n232479 , n236962 );
and ( n237404 , n224925 , n221016 );
not ( n237405 , n224881 );
and ( n237406 , n224929 , n237405 );
nor ( n237407 , n237404 , n237406 );
or ( n237408 , n232948 , n237407 );
nand ( n237409 , n237403 , n237408 );
not ( n237410 , n236973 );
not ( n237411 , n232956 );
or ( n237412 , n237410 , n237411 );
not ( n237413 , n229806 );
not ( n237414 , n217130 );
and ( n237415 , n237413 , n237414 );
and ( n237416 , n219581 , n232962 );
nor ( n237417 , n237415 , n237416 );
not ( n237418 , n237417 );
nand ( n237419 , n237418 , n228775 );
nand ( n237420 , n237412 , n237419 );
xor ( n237421 , n237409 , n237420 );
not ( n237422 , n236982 );
not ( n237423 , n237422 );
not ( n237424 , n229816 );
or ( n237425 , n237423 , n237424 );
not ( n237426 , n41565 );
not ( n237427 , n232431 );
or ( n237428 , n237426 , n237427 );
nand ( n237429 , n232974 , n211422 );
nand ( n237430 , n237428 , n237429 );
nand ( n237431 , n237430 , n226885 );
nand ( n237432 , n237425 , n237431 );
xor ( n237433 , n237421 , n237432 );
xor ( n237434 , n237409 , n237420 );
and ( n237435 , n237434 , n237432 );
and ( n237436 , n237409 , n237420 );
or ( n237437 , n237435 , n237436 );
xor ( n237438 , n237307 , n237398 );
or ( n237439 , n228270 , n236996 );
and ( n237440 , n227596 , n225768 );
and ( n237441 , n233450 , n225769 );
nor ( n237442 , n237440 , n237441 );
or ( n237443 , n228273 , n237442 );
nand ( n237444 , n237439 , n237443 );
not ( n237445 , n237045 );
not ( n237446 , n231421 );
or ( n237447 , n237445 , n237446 );
not ( n237448 , n214837 );
not ( n237449 , n231940 );
or ( n237450 , n237448 , n237449 );
nand ( n237451 , n228850 , n231913 );
nand ( n237452 , n237450 , n237451 );
nand ( n237453 , n228868 , n237452 );
nand ( n237454 , n237447 , n237453 );
xor ( n237455 , n237444 , n237454 );
not ( n237456 , n237019 );
not ( n237457 , n237456 );
not ( n237458 , n234371 );
or ( n237459 , n237457 , n237458 );
not ( n237460 , n229759 );
not ( n237461 , n224041 );
and ( n237462 , n237460 , n237461 );
and ( n237463 , n237017 , n224041 );
nor ( n237464 , n237462 , n237463 );
not ( n237465 , n237464 );
nand ( n237466 , n237465 , n234378 );
nand ( n237467 , n237459 , n237466 );
xor ( n237468 , n237455 , n237467 );
xor ( n237469 , n237438 , n237468 );
xor ( n237470 , n237307 , n237398 );
and ( n237471 , n237470 , n237468 );
and ( n237472 , n237307 , n237398 );
or ( n237473 , n237471 , n237472 );
xor ( n237474 , n237433 , n237347 );
xor ( n237475 , n237474 , n237351 );
xor ( n237476 , n237433 , n237347 );
and ( n237477 , n237476 , n237351 );
and ( n237478 , n237433 , n237347 );
or ( n237479 , n237477 , n237478 );
not ( n237480 , n237033 );
not ( n237481 , n233105 );
or ( n237482 , n237480 , n237481 );
not ( n237483 , n220022 );
not ( n237484 , n237483 );
not ( n237485 , n230722 );
or ( n237486 , n237484 , n237485 );
nand ( n237487 , n236615 , n220022 );
nand ( n237488 , n237486 , n237487 );
nand ( n237489 , n237488 , n232402 );
nand ( n237490 , n237482 , n237489 );
and ( n237491 , n231754 , n219343 );
xor ( n237492 , n237490 , n237491 );
buf ( n237493 , n222158 );
not ( n237494 , n237493 );
not ( n237495 , n222892 );
not ( n237496 , n219599 );
not ( n237497 , n237496 );
or ( n237498 , n237495 , n237497 );
nand ( n237499 , n219599 , n222458 );
nand ( n237500 , n237498 , n237499 );
not ( n237501 , n237500 );
or ( n237502 , n237494 , n237501 );
not ( n237503 , n235644 );
nand ( n237504 , n237147 , n237503 );
nand ( n237505 , n237502 , n237504 );
xor ( n237506 , n237492 , n237505 );
xor ( n237507 , n237355 , n237506 );
xor ( n237508 , n237507 , n237363 );
xor ( n237509 , n237355 , n237506 );
and ( n237510 , n237509 , n237363 );
and ( n237511 , n237355 , n237506 );
or ( n237512 , n237510 , n237511 );
xor ( n237513 , n237367 , n237371 );
not ( n237514 , n218533 );
not ( n237515 , n218771 );
not ( n237516 , n227004 );
or ( n237517 , n237515 , n237516 );
nand ( n237518 , n227007 , n221214 );
nand ( n237519 , n237517 , n237518 );
not ( n237520 , n237519 );
or ( n237521 , n237514 , n237520 );
nand ( n237522 , n237118 , n219836 );
nand ( n237523 , n237521 , n237522 );
not ( n237524 , n218843 );
not ( n237525 , n220126 );
not ( n237526 , n221712 );
or ( n237527 , n237525 , n237526 );
nand ( n237528 , n40182 , n221238 );
nand ( n237529 , n237527 , n237528 );
not ( n237530 , n237529 );
or ( n237531 , n237524 , n237530 );
not ( n237532 , n237073 );
not ( n237533 , n237071 );
or ( n237534 , n237532 , n237533 );
nand ( n237535 , n237534 , n223665 );
nand ( n237536 , n237531 , n237535 );
xor ( n237537 , n237523 , n237536 );
not ( n237538 , n219076 );
not ( n237539 , n219424 );
not ( n237540 , n222552 );
or ( n237541 , n237539 , n237540 );
nand ( n237542 , n220970 , n219420 );
nand ( n237543 , n237541 , n237542 );
not ( n237544 , n237543 );
or ( n237545 , n237538 , n237544 );
nand ( n237546 , n219792 , n237086 );
nand ( n237547 , n237545 , n237546 );
xor ( n237548 , n237537 , n237547 );
xor ( n237549 , n237513 , n237548 );
xor ( n237550 , n237367 , n237371 );
and ( n237551 , n237550 , n237548 );
and ( n237552 , n237367 , n237371 );
or ( n237553 , n237551 , n237552 );
not ( n237554 , n219779 );
not ( n237555 , n220150 );
not ( n237556 , n226921 );
or ( n237557 , n237555 , n237556 );
nand ( n237558 , n226922 , n221257 );
nand ( n237559 , n237557 , n237558 );
not ( n237560 , n237559 );
or ( n237561 , n237554 , n237560 );
nand ( n237562 , n237094 , n220164 );
nand ( n237563 , n237561 , n237562 );
xor ( n237564 , n237563 , n237134 );
not ( n237565 , n237196 );
not ( n237566 , n235913 );
or ( n237567 , n237565 , n237566 );
not ( n237568 , n222399 );
not ( n237569 , n221040 );
or ( n237570 , n237568 , n237569 );
nand ( n237571 , n40625 , n236754 );
nand ( n237572 , n237570 , n237571 );
nand ( n237573 , n221674 , n237572 );
nand ( n237574 , n237567 , n237573 );
xor ( n237575 , n237564 , n237574 );
not ( n237576 , n234006 );
not ( n237577 , n237167 );
or ( n237578 , n237576 , n237577 );
not ( n237579 , n229261 );
not ( n237580 , n226961 );
or ( n237581 , n237579 , n237580 );
nand ( n237582 , n226964 , n229262 );
nand ( n237583 , n237581 , n237582 );
nand ( n237584 , n237583 , n229964 );
nand ( n237585 , n237578 , n237584 );
not ( n237586 , n221637 );
not ( n237587 , n221633 );
not ( n237588 , n236752 );
not ( n237589 , n237588 );
or ( n237590 , n237587 , n237589 );
nand ( n237591 , n236752 , n221778 );
nand ( n237592 , n237590 , n237591 );
not ( n237593 , n237592 );
or ( n237594 , n237586 , n237593 );
nand ( n237595 , n237158 , n221626 );
nand ( n237596 , n237594 , n237595 );
xor ( n237597 , n237585 , n237596 );
not ( n237598 , n220067 );
not ( n237599 , n231500 );
not ( n237600 , n235031 );
not ( n237601 , n237600 );
or ( n237602 , n237599 , n237601 );
nand ( n237603 , n235031 , n234015 );
nand ( n237604 , n237602 , n237603 );
not ( n237605 , n237604 );
or ( n237606 , n237598 , n237605 );
nand ( n237607 , n237106 , n220059 );
nand ( n237608 , n237606 , n237607 );
xor ( n237609 , n237597 , n237608 );
xor ( n237610 , n237575 , n237609 );
xor ( n237611 , n237610 , n237359 );
xor ( n237612 , n237575 , n237609 );
and ( n237613 , n237612 , n237359 );
and ( n237614 , n237575 , n237609 );
or ( n237615 , n237613 , n237614 );
not ( n237616 , n223949 );
not ( n237617 , n226655 );
not ( n237618 , n233857 );
or ( n237619 , n237617 , n237618 );
nand ( n237620 , n233856 , n233053 );
nand ( n237621 , n237619 , n237620 );
not ( n237622 , n237621 );
or ( n237623 , n237616 , n237622 );
nand ( n237624 , n237176 , n227260 );
nand ( n237625 , n237623 , n237624 );
xor ( n237626 , n237625 , n236989 );
xor ( n237627 , n237626 , n237026 );
xor ( n237628 , n237627 , n237055 );
not ( n237629 , n225478 );
not ( n237630 , n237205 );
or ( n237631 , n237629 , n237630 );
not ( n237632 , n229387 );
not ( n237633 , n39928 );
or ( n237634 , n237632 , n237633 );
nand ( n237635 , n235820 , n227599 );
nand ( n237636 , n237634 , n237635 );
nand ( n237637 , n237636 , n219501 );
nand ( n237638 , n237631 , n237637 );
not ( n237639 , n220272 );
not ( n237640 , n234788 );
not ( n237641 , n234094 );
or ( n237642 , n237640 , n237641 );
not ( n237643 , n209963 );
nand ( n237644 , n237643 , n234787 );
nand ( n237645 , n237642 , n237644 );
not ( n237646 , n237645 );
or ( n237647 , n237639 , n237646 );
nand ( n237648 , n237218 , n220280 );
nand ( n237649 , n237647 , n237648 );
xor ( n237650 , n237638 , n237649 );
not ( n237651 , n219314 );
nand ( n237652 , n236840 , n222323 );
nand ( n237653 , n236844 , n219687 );
nand ( n237654 , n237652 , n237653 );
not ( n237655 , n237654 );
or ( n237656 , n237651 , n237655 );
nand ( n237657 , n237231 , n224624 );
nand ( n237658 , n237656 , n237657 );
xor ( n237659 , n237650 , n237658 );
xor ( n237660 , n237628 , n237659 );
xor ( n237661 , n237627 , n237055 );
and ( n237662 , n237661 , n237659 );
and ( n237663 , n237627 , n237055 );
or ( n237664 , n237662 , n237663 );
buf ( n237665 , n215183 );
not ( n237666 , n237665 );
not ( n237667 , n237240 );
or ( n237668 , n237666 , n237667 );
not ( n237669 , n226484 );
not ( n237670 , n229704 );
or ( n237671 , n237669 , n237670 );
nand ( n237672 , n38532 , n222333 );
nand ( n237673 , n237671 , n237672 );
nand ( n237674 , n221933 , n237673 );
nand ( n237675 , n237668 , n237674 );
not ( n237676 , n226287 );
and ( n237677 , n226292 , n39607 );
not ( n237678 , n226292 );
and ( n237679 , n237678 , n226712 );
nor ( n237680 , n237677 , n237679 );
not ( n237681 , n237680 );
or ( n237682 , n237676 , n237681 );
nand ( n237683 , n237263 , n220414 );
nand ( n237684 , n237682 , n237683 );
xor ( n237685 , n237675 , n237684 );
not ( n237686 , n219731 );
not ( n237687 , n237274 );
or ( n237688 , n237686 , n237687 );
not ( n237689 , n219033 );
not ( n237690 , n229691 );
or ( n237691 , n237689 , n237690 );
nand ( n237692 , n233846 , n219034 );
nand ( n237693 , n237691 , n237692 );
nand ( n237694 , n237693 , n222185 );
nand ( n237695 , n237688 , n237694 );
xor ( n237696 , n237685 , n237695 );
xor ( n237697 , n237696 , n237469 );
xor ( n237698 , n237697 , n237061 );
xor ( n237699 , n237696 , n237469 );
and ( n237700 , n237699 , n237061 );
and ( n237701 , n237696 , n237469 );
or ( n237702 , n237700 , n237701 );
xor ( n237703 , n237067 , n237508 );
xor ( n237704 , n237703 , n237141 );
xor ( n237705 , n237067 , n237508 );
and ( n237706 , n237705 , n237141 );
and ( n237707 , n237067 , n237508 );
or ( n237708 , n237706 , n237707 );
xor ( n237709 , n237475 , n237188 );
xor ( n237710 , n237709 , n237250 );
xor ( n237711 , n237475 , n237188 );
and ( n237712 , n237711 , n237250 );
and ( n237713 , n237475 , n237188 );
or ( n237714 , n237712 , n237713 );
xor ( n237715 , n237611 , n237549 );
xor ( n237716 , n237715 , n237285 );
xor ( n237717 , n237611 , n237549 );
and ( n237718 , n237717 , n237285 );
and ( n237719 , n237611 , n237549 );
or ( n237720 , n237718 , n237719 );
xor ( n237721 , n237444 , n237454 );
and ( n237722 , n237721 , n237467 );
and ( n237723 , n237444 , n237454 );
or ( n237724 , n237722 , n237723 );
xor ( n237725 , n237660 , n237291 );
xor ( n237726 , n237725 , n237698 );
xor ( n237727 , n237660 , n237291 );
and ( n237728 , n237727 , n237698 );
and ( n237729 , n237660 , n237291 );
or ( n237730 , n237728 , n237729 );
xor ( n237731 , n237704 , n237297 );
xor ( n237732 , n237731 , n237710 );
xor ( n237733 , n237704 , n237297 );
and ( n237734 , n237733 , n237710 );
and ( n237735 , n237704 , n237297 );
or ( n237736 , n237734 , n237735 );
xor ( n237737 , n237303 , n237716 );
xor ( n237738 , n237737 , n237313 );
xor ( n237739 , n237303 , n237716 );
and ( n237740 , n237739 , n237313 );
and ( n237741 , n237303 , n237716 );
or ( n237742 , n237740 , n237741 );
xor ( n237743 , n237726 , n237319 );
xor ( n237744 , n237743 , n237732 );
xor ( n237745 , n237726 , n237319 );
and ( n237746 , n237745 , n237732 );
and ( n237747 , n237726 , n237319 );
or ( n237748 , n237746 , n237747 );
xor ( n237749 , n237738 , n237325 );
xor ( n237750 , n237749 , n237331 );
xor ( n237751 , n237738 , n237325 );
and ( n237752 , n237751 , n237331 );
and ( n237753 , n237738 , n237325 );
or ( n237754 , n237752 , n237753 );
xor ( n237755 , n237744 , n237750 );
xor ( n237756 , n237755 , n237337 );
xor ( n237757 , n237744 , n237750 );
and ( n237758 , n237757 , n237337 );
and ( n237759 , n237744 , n237750 );
or ( n237760 , n237758 , n237759 );
xor ( n237761 , n237490 , n237491 );
and ( n237762 , n237761 , n237505 );
and ( n237763 , n237490 , n237491 );
or ( n237764 , n237762 , n237763 );
xor ( n237765 , n237585 , n237596 );
and ( n237766 , n237765 , n237608 );
and ( n237767 , n237585 , n237596 );
or ( n237768 , n237766 , n237767 );
xor ( n237769 , n237523 , n237536 );
and ( n237770 , n237769 , n237547 );
and ( n237771 , n237523 , n237536 );
or ( n237772 , n237770 , n237771 );
xor ( n237773 , n237563 , n237134 );
and ( n237774 , n237773 , n237574 );
and ( n237775 , n237563 , n237134 );
or ( n237776 , n237774 , n237775 );
xor ( n237777 , n237638 , n237649 );
and ( n237778 , n237777 , n237658 );
and ( n237779 , n237638 , n237649 );
or ( n237780 , n237778 , n237779 );
xor ( n237781 , n237675 , n237684 );
and ( n237782 , n237781 , n237695 );
and ( n237783 , n237675 , n237684 );
or ( n237784 , n237782 , n237783 );
xor ( n237785 , n237625 , n236989 );
and ( n237786 , n237785 , n237026 );
and ( n237787 , n237625 , n236989 );
or ( n237788 , n237786 , n237787 );
not ( n237789 , n229271 );
or ( n237790 , n237789 , n237417 );
and ( n237791 , n232493 , n41321 );
and ( n237792 , n232962 , n208597 );
nor ( n237793 , n237791 , n237792 );
or ( n237794 , n231456 , n237793 );
nand ( n237795 , n237790 , n237794 );
not ( n237796 , n237430 );
buf ( n237797 , n226881 );
not ( n237798 , n237797 );
or ( n237799 , n237796 , n237798 );
not ( n237800 , n215796 );
not ( n237801 , n234293 );
or ( n237802 , n237800 , n237801 );
nand ( n237803 , n232974 , n216261 );
nand ( n237804 , n237802 , n237803 );
nand ( n237805 , n226885 , n237804 );
nand ( n237806 , n237799 , n237805 );
xor ( n237807 , n237795 , n237806 );
not ( n237808 , n237442 );
not ( n237809 , n237808 );
buf ( n237810 , n232440 );
not ( n237811 , n237810 );
or ( n237812 , n237809 , n237811 );
not ( n237813 , n226225 );
not ( n237814 , n227596 );
or ( n237815 , n237813 , n237814 );
buf ( n237816 , n233450 );
nand ( n237817 , n237816 , n234256 );
nand ( n237818 , n237815 , n237817 );
nand ( n237819 , n227737 , n237818 );
nand ( n237820 , n237812 , n237819 );
xor ( n237821 , n237807 , n237820 );
xor ( n237822 , n237795 , n237806 );
and ( n237823 , n237822 , n237820 );
and ( n237824 , n237795 , n237806 );
or ( n237825 , n237823 , n237824 );
not ( n237826 , n228860 );
not ( n237827 , n237452 );
or ( n237828 , n237826 , n237827 );
not ( n237829 , n219689 );
not ( n237830 , n228847 );
or ( n237831 , n237829 , n237830 );
nand ( n237832 , n233925 , n235216 );
nand ( n237833 , n237831 , n237832 );
nand ( n237834 , n234404 , n237833 );
nand ( n237835 , n237828 , n237834 );
not ( n237836 , n237395 );
not ( n237837 , n224087 );
or ( n237838 , n237836 , n237837 );
not ( n237839 , n217330 );
not ( n237840 , n233309 );
or ( n237841 , n237839 , n237840 );
nand ( n237842 , n237129 , n217331 );
nand ( n237843 , n237841 , n237842 );
nand ( n237844 , n227782 , n237843 );
nand ( n237845 , n237838 , n237844 );
xor ( n237846 , n237835 , n237845 );
or ( n237847 , n231994 , n237464 );
and ( n237848 , n225505 , n237017 );
not ( n237849 , n225505 );
and ( n237850 , n237849 , n233399 );
nor ( n237851 , n237848 , n237850 );
or ( n237852 , n231476 , n237851 );
nand ( n237853 , n237847 , n237852 );
xor ( n237854 , n237846 , n237853 );
xor ( n237855 , n237835 , n237845 );
and ( n237856 , n237855 , n237853 );
and ( n237857 , n237835 , n237845 );
or ( n237858 , n237856 , n237857 );
xor ( n237859 , n237854 , n237821 );
xor ( n237860 , n237859 , n237768 );
xor ( n237861 , n237854 , n237821 );
and ( n237862 , n237861 , n237768 );
and ( n237863 , n237854 , n237821 );
or ( n237864 , n237862 , n237863 );
xor ( n237865 , n237772 , n237776 );
xor ( n237866 , n237865 , n237764 );
xor ( n237867 , n237772 , n237776 );
and ( n237868 , n237867 , n237764 );
and ( n237869 , n237772 , n237776 );
or ( n237870 , n237868 , n237869 );
xor ( n237871 , n237784 , n237788 );
not ( n237872 , n222376 );
not ( n237873 , n232413 );
not ( n237874 , n224700 );
or ( n237875 , n237873 , n237874 );
nand ( n237876 , n236300 , n221238 );
nand ( n237877 , n237875 , n237876 );
not ( n237878 , n237877 );
or ( n237879 , n237872 , n237878 );
nand ( n237880 , n237529 , n223665 );
nand ( n237881 , n237879 , n237880 );
not ( n237882 , n219435 );
not ( n237883 , n237543 );
or ( n237884 , n237882 , n237883 );
not ( n237885 , n219800 );
not ( n237886 , n222121 );
or ( n237887 , n237885 , n237886 );
not ( n237888 , n230511 );
nand ( n237889 , n237888 , n219420 );
nand ( n237890 , n237887 , n237889 );
nand ( n237891 , n237890 , n219076 );
nand ( n237892 , n237884 , n237891 );
xor ( n237893 , n237881 , n237892 );
not ( n237894 , n237559 );
not ( n237895 , n220164 );
or ( n237896 , n237894 , n237895 );
not ( n237897 , n220151 );
not ( n237898 , n221330 );
or ( n237899 , n237897 , n237898 );
nand ( n237900 , n220600 , n220147 );
nand ( n237901 , n237899 , n237900 );
not ( n237902 , n237901 );
or ( n237903 , n237902 , n224171 );
nand ( n237904 , n237896 , n237903 );
xor ( n237905 , n237893 , n237904 );
xor ( n237906 , n237871 , n237905 );
xor ( n237907 , n237784 , n237788 );
and ( n237908 , n237907 , n237905 );
and ( n237909 , n237784 , n237788 );
or ( n237910 , n237908 , n237909 );
not ( n237911 , n235195 );
not ( n237912 , n237407 );
and ( n237913 , n237911 , n237912 );
buf ( n237914 , n224941 );
not ( n237915 , n237914 );
and ( n237916 , n40888 , n234878 );
not ( n237917 , n40888 );
not ( n237918 , n234878 );
and ( n237919 , n237917 , n237918 );
nor ( n237920 , n237916 , n237919 );
nor ( n237921 , n237915 , n237920 );
nor ( n237922 , n237913 , n237921 );
not ( n237923 , n235913 );
not ( n237924 , n237572 );
or ( n237925 , n237923 , n237924 );
not ( n237926 , n222399 );
not ( n237927 , n40660 );
or ( n237928 , n237926 , n237927 );
nand ( n237929 , n207938 , n220901 );
nand ( n237930 , n237928 , n237929 );
nand ( n237931 , n237930 , n220930 );
nand ( n237932 , n237925 , n237931 );
xor ( n237933 , n237922 , n237932 );
not ( n237934 , n221626 );
not ( n237935 , n237592 );
or ( n237936 , n237934 , n237935 );
not ( n237937 , n221778 );
not ( n237938 , n237937 );
not ( n237939 , n227448 );
or ( n237940 , n237938 , n237939 );
nand ( n237941 , n220657 , n222586 );
nand ( n237942 , n237940 , n237941 );
nand ( n237943 , n237942 , n221637 );
nand ( n237944 , n237936 , n237943 );
xor ( n237945 , n237933 , n237944 );
not ( n237946 , n237493 );
not ( n237947 , n222430 );
buf ( n237948 , n40766 );
not ( n237949 , n237948 );
or ( n237950 , n237947 , n237949 );
nand ( n237951 , n224642 , n222458 );
nand ( n237952 , n237950 , n237951 );
not ( n237953 , n237952 );
or ( n237954 , n237946 , n237953 );
nand ( n237955 , n237500 , n222454 );
nand ( n237956 , n237954 , n237955 );
not ( n237957 , n231018 );
not ( n237958 , n237604 );
or ( n237959 , n237957 , n237958 );
not ( n237960 , n231500 );
not ( n237961 , n230490 );
or ( n237962 , n237960 , n237961 );
buf ( n237963 , n234506 );
nand ( n237964 , n237963 , n234015 );
nand ( n237965 , n237962 , n237964 );
nand ( n237966 , n237965 , n220067 );
nand ( n237967 , n237959 , n237966 );
xor ( n237968 , n237956 , n237967 );
not ( n237969 , n218232 );
not ( n237970 , n218205 );
not ( n237971 , n40484 );
not ( n237972 , n237971 );
or ( n237973 , n237970 , n237972 );
nand ( n237974 , n236290 , n234949 );
nand ( n237975 , n237973 , n237974 );
not ( n237976 , n237975 );
or ( n237977 , n237969 , n237976 );
nand ( n237978 , n237519 , n219461 );
nand ( n237979 , n237977 , n237978 );
xor ( n237980 , n237968 , n237979 );
xor ( n237981 , n237945 , n237980 );
xor ( n237982 , n237981 , n237780 );
xor ( n237983 , n237945 , n237980 );
and ( n237984 , n237983 , n237780 );
and ( n237985 , n237945 , n237980 );
or ( n237986 , n237984 , n237985 );
xor ( n237987 , n237437 , n237724 );
not ( n237988 , n237488 );
not ( n237989 , n233105 );
or ( n237990 , n237988 , n237989 );
not ( n237991 , n216293 );
not ( n237992 , n231753 );
or ( n237993 , n237991 , n237992 );
nand ( n237994 , n230726 , n223658 );
nand ( n237995 , n237993 , n237994 );
nand ( n237996 , n237995 , n232402 );
nand ( n237997 , n237990 , n237996 );
and ( n237998 , n234382 , n221921 );
xor ( n237999 , n237997 , n237998 );
not ( n238000 , n227294 );
and ( n238001 , n40724 , n223183 );
not ( n238002 , n40724 );
and ( n238003 , n238002 , n237005 );
or ( n238004 , n238001 , n238003 );
not ( n238005 , n238004 );
or ( n238006 , n238000 , n238005 );
nand ( n238007 , n223197 , n237383 );
nand ( n238008 , n238006 , n238007 );
xor ( n238009 , n237999 , n238008 );
xor ( n238010 , n237987 , n238009 );
xor ( n238011 , n238010 , n237473 );
not ( n238012 , n229964 );
not ( n238013 , n229261 );
not ( n238014 , n39877 );
or ( n238015 , n238013 , n238014 );
nand ( n238016 , n225344 , n229262 );
nand ( n238017 , n238015 , n238016 );
not ( n238018 , n238017 );
or ( n238019 , n238012 , n238018 );
nand ( n238020 , n237583 , n229974 );
nand ( n238021 , n238019 , n238020 );
not ( n238022 , n219731 );
not ( n238023 , n237693 );
or ( n238024 , n238022 , n238023 );
not ( n238025 , n219033 );
not ( n238026 , n233611 );
or ( n238027 , n238025 , n238026 );
nand ( n238028 , n209865 , n219034 );
nand ( n238029 , n238027 , n238028 );
nand ( n238030 , n238029 , n222185 );
nand ( n238031 , n238024 , n238030 );
xor ( n238032 , n238021 , n238031 );
not ( n238033 , n221933 );
not ( n238034 , n226484 );
not ( n238035 , n39366 );
or ( n238036 , n238034 , n238035 );
nand ( n238037 , n39365 , n221938 );
nand ( n238038 , n238036 , n238037 );
not ( n238039 , n238038 );
or ( n238040 , n238033 , n238039 );
nand ( n238041 , n237673 , n219332 );
nand ( n238042 , n238040 , n238041 );
xor ( n238043 , n238032 , n238042 );
xor ( n238044 , n238011 , n238043 );
xor ( n238045 , n238010 , n237473 );
and ( n238046 , n238045 , n238043 );
and ( n238047 , n238010 , n237473 );
or ( n238048 , n238046 , n238047 );
not ( n238049 , n227260 );
not ( n238050 , n237621 );
or ( n238051 , n238049 , n238050 );
not ( n238052 , n226655 );
not ( n238053 , n235516 );
or ( n238054 , n238052 , n238053 );
nand ( n238055 , n39747 , n233053 );
nand ( n238056 , n238054 , n238055 );
nand ( n238057 , n238056 , n223949 );
nand ( n238058 , n238051 , n238057 );
not ( n238059 , n228237 );
not ( n238060 , n233544 );
not ( n238061 , n234350 );
or ( n238062 , n238060 , n238061 );
nand ( n238063 , n227223 , n237203 );
nand ( n238064 , n238062 , n238063 );
not ( n238065 , n238064 );
or ( n238066 , n238059 , n238065 );
nand ( n238067 , n237636 , n229395 );
nand ( n238068 , n238066 , n238067 );
xor ( n238069 , n238058 , n238068 );
xor ( n238070 , n238069 , n237402 );
not ( n238071 , n226287 );
not ( n238072 , n227912 );
not ( n238073 , n228184 );
or ( n238074 , n238072 , n238073 );
nand ( n238075 , n39089 , n229887 );
nand ( n238076 , n238074 , n238075 );
not ( n238077 , n238076 );
or ( n238078 , n238071 , n238077 );
nand ( n238079 , n237680 , n226943 );
nand ( n238080 , n238078 , n238079 );
not ( n238081 , n224624 );
not ( n238082 , n237654 );
or ( n238083 , n238081 , n238082 );
not ( n238084 , n219687 );
not ( n238085 , n233362 );
or ( n238086 , n238084 , n238085 );
nand ( n238087 , n233363 , n222323 );
nand ( n238088 , n238086 , n238087 );
nand ( n238089 , n238088 , n219314 );
nand ( n238090 , n238083 , n238089 );
xor ( n238091 , n238080 , n238090 );
not ( n238092 , n237645 );
or ( n238093 , n238092 , n217551 );
or ( n238094 , n217549 , n234787 );
nand ( n238095 , n238093 , n238094 );
xor ( n238096 , n238091 , n238095 );
xor ( n238097 , n238070 , n238096 );
xor ( n238098 , n238097 , n237479 );
xor ( n238099 , n238070 , n238096 );
and ( n238100 , n238099 , n237479 );
and ( n238101 , n238070 , n238096 );
or ( n238102 , n238100 , n238101 );
xor ( n238103 , n237860 , n237615 );
xor ( n238104 , n238103 , n237553 );
xor ( n238105 , n237860 , n237615 );
and ( n238106 , n238105 , n237553 );
and ( n238107 , n237860 , n237615 );
or ( n238108 , n238106 , n238107 );
xor ( n238109 , n237866 , n237512 );
xor ( n238110 , n238109 , n237664 );
xor ( n238111 , n237866 , n237512 );
and ( n238112 , n238111 , n237664 );
and ( n238113 , n237866 , n237512 );
or ( n238114 , n238112 , n238113 );
xor ( n238115 , n237982 , n237906 );
xor ( n238116 , n238115 , n238098 );
xor ( n238117 , n237982 , n237906 );
and ( n238118 , n238117 , n238098 );
and ( n238119 , n237982 , n237906 );
or ( n238120 , n238118 , n238119 );
xor ( n238121 , n237702 , n238044 );
xor ( n238122 , n238121 , n237708 );
xor ( n238123 , n237702 , n238044 );
and ( n238124 , n238123 , n237708 );
and ( n238125 , n237702 , n238044 );
or ( n238126 , n238124 , n238125 );
xor ( n238127 , n237997 , n237998 );
and ( n238128 , n238127 , n238008 );
and ( n238129 , n237997 , n237998 );
or ( n238130 , n238128 , n238129 );
xor ( n238131 , n237714 , n238104 );
xor ( n238132 , n238131 , n238110 );
xor ( n238133 , n237714 , n238104 );
and ( n238134 , n238133 , n238110 );
and ( n238135 , n237714 , n238104 );
or ( n238136 , n238134 , n238135 );
xor ( n238137 , n238116 , n237720 );
xor ( n238138 , n238137 , n238122 );
xor ( n238139 , n238116 , n237720 );
and ( n238140 , n238139 , n238122 );
and ( n238141 , n238116 , n237720 );
or ( n238142 , n238140 , n238141 );
xor ( n238143 , n237730 , n237736 );
xor ( n238144 , n238143 , n238132 );
xor ( n238145 , n237730 , n237736 );
and ( n238146 , n238145 , n238132 );
and ( n238147 , n237730 , n237736 );
or ( n238148 , n238146 , n238147 );
xor ( n238149 , n238138 , n237742 );
xor ( n238150 , n238149 , n237748 );
xor ( n238151 , n238138 , n237742 );
and ( n238152 , n238151 , n237748 );
and ( n238153 , n238138 , n237742 );
or ( n238154 , n238152 , n238153 );
xor ( n238155 , n238144 , n238150 );
xor ( n238156 , n238155 , n237754 );
xor ( n238157 , n238144 , n238150 );
and ( n238158 , n238157 , n237754 );
and ( n238159 , n238144 , n238150 );
or ( n238160 , n238158 , n238159 );
xor ( n238161 , n237956 , n237967 );
and ( n238162 , n238161 , n237979 );
and ( n238163 , n237956 , n237967 );
or ( n238164 , n238162 , n238163 );
xor ( n238165 , n237881 , n237892 );
and ( n238166 , n238165 , n237904 );
and ( n238167 , n237881 , n237892 );
or ( n238168 , n238166 , n238167 );
xor ( n238169 , n237922 , n237932 );
and ( n238170 , n238169 , n237944 );
and ( n238171 , n237922 , n237932 );
or ( n238172 , n238170 , n238171 );
xor ( n238173 , n238021 , n238031 );
and ( n238174 , n238173 , n238042 );
and ( n238175 , n238021 , n238031 );
or ( n238176 , n238174 , n238175 );
xor ( n238177 , n238080 , n238090 );
and ( n238178 , n238177 , n238095 );
and ( n238179 , n238080 , n238090 );
or ( n238180 , n238178 , n238179 );
xor ( n238181 , n238058 , n238068 );
and ( n238182 , n238181 , n237402 );
and ( n238183 , n238058 , n238068 );
or ( n238184 , n238182 , n238183 );
xor ( n238185 , n237437 , n237724 );
and ( n238186 , n238185 , n238009 );
and ( n238187 , n237437 , n237724 );
or ( n238188 , n238186 , n238187 );
not ( n238189 , n217549 );
not ( n238190 , n217551 );
or ( n238191 , n238189 , n238190 );
nand ( n238192 , n238191 , n215955 );
not ( n238193 , n237843 );
not ( n238194 , n224087 );
or ( n238195 , n238193 , n238194 );
not ( n238196 , n237130 );
not ( n238197 , n219386 );
or ( n238198 , n238196 , n238197 );
not ( n238199 , n219386 );
nand ( n238200 , n238199 , n234764 );
nand ( n238201 , n238198 , n238200 );
nand ( n238202 , n224090 , n238201 );
nand ( n238203 , n238195 , n238202 );
xor ( n238204 , n238192 , n238203 );
or ( n238205 , n237920 , n233316 );
and ( n238206 , n231762 , n234273 );
not ( n238207 , n231762 );
and ( n238208 , n238207 , n234878 );
nor ( n238209 , n238206 , n238208 );
or ( n238210 , n236958 , n238209 );
nand ( n238211 , n238205 , n238210 );
xor ( n238212 , n238204 , n238211 );
xor ( n238213 , n238192 , n238203 );
and ( n238214 , n238213 , n238211 );
and ( n238215 , n238192 , n238203 );
or ( n238216 , n238214 , n238215 );
or ( n238217 , n231453 , n237793 );
not ( n238218 , n41249 );
and ( n238219 , n233962 , n238218 );
and ( n238220 , n225952 , n237405 );
nor ( n238221 , n238219 , n238220 );
or ( n238222 , n231456 , n238221 );
nand ( n238223 , n238217 , n238222 );
not ( n238224 , n237804 );
not ( n238225 , n234290 );
not ( n238226 , n238225 );
or ( n238227 , n238224 , n238226 );
and ( n238228 , n216500 , n234295 );
not ( n238229 , n216500 );
buf ( n238230 , n230897 );
and ( n238231 , n238229 , n238230 );
nor ( n238232 , n238228 , n238231 );
not ( n238233 , n238232 );
nand ( n238234 , n238233 , n227852 );
nand ( n238235 , n238227 , n238234 );
xor ( n238236 , n238223 , n238235 );
not ( n238237 , n237818 );
not ( n238238 , n237810 );
or ( n238239 , n238237 , n238238 );
buf ( n238240 , n233912 );
not ( n238241 , n41565 );
not ( n238242 , n233451 );
or ( n238243 , n238241 , n238242 );
nand ( n238244 , n236188 , n236580 );
nand ( n238245 , n238243 , n238244 );
nand ( n238246 , n238240 , n238245 );
nand ( n238247 , n238239 , n238246 );
xor ( n238248 , n238236 , n238247 );
xor ( n238249 , n238223 , n238235 );
and ( n238250 , n238249 , n238247 );
and ( n238251 , n238223 , n238235 );
or ( n238252 , n238250 , n238251 );
not ( n238253 , n237833 );
not ( n238254 , n228860 );
or ( n238255 , n238253 , n238254 );
not ( n238256 , n225768 );
not ( n238257 , n228847 );
or ( n238258 , n238256 , n238257 );
nand ( n238259 , n233925 , n225769 );
nand ( n238260 , n238258 , n238259 );
nand ( n238261 , n234404 , n238260 );
nand ( n238262 , n238255 , n238261 );
or ( n238263 , n231994 , n237851 );
and ( n238264 , n214837 , n229762 );
not ( n238265 , n214837 );
and ( n238266 , n238265 , n231480 );
nor ( n238267 , n238264 , n238266 );
or ( n238268 , n237013 , n238267 );
nand ( n238269 , n238263 , n238268 );
xor ( n238270 , n238262 , n238269 );
not ( n238271 , n233105 );
not ( n238272 , n237995 );
or ( n238273 , n238271 , n238272 );
buf ( n238274 , n230708 );
not ( n238275 , n238274 );
not ( n238276 , n231232 );
not ( n238277 , n224041 );
and ( n238278 , n238276 , n238277 );
and ( n238279 , n231232 , n224041 );
nor ( n238280 , n238278 , n238279 );
or ( n238281 , n238275 , n238280 );
nand ( n238282 , n238273 , n238281 );
xor ( n238283 , n238270 , n238282 );
xor ( n238284 , n238283 , n238248 );
xor ( n238285 , n238284 , n238130 );
xor ( n238286 , n238283 , n238248 );
and ( n238287 , n238286 , n238130 );
and ( n238288 , n238283 , n238248 );
or ( n238289 , n238287 , n238288 );
xor ( n238290 , n238168 , n238172 );
xor ( n238291 , n238290 , n238164 );
xor ( n238292 , n238168 , n238172 );
and ( n238293 , n238292 , n238164 );
and ( n238294 , n238168 , n238172 );
or ( n238295 , n238293 , n238294 );
xor ( n238296 , n238176 , n238184 );
not ( n238297 , n221674 );
not ( n238298 , n220906 );
not ( n238299 , n230966 );
or ( n238300 , n238298 , n238299 );
not ( n238301 , n220925 );
nand ( n238302 , n226922 , n238301 );
nand ( n238303 , n238300 , n238302 );
not ( n238304 , n238303 );
or ( n238305 , n238297 , n238304 );
nand ( n238306 , n237930 , n235913 );
nand ( n238307 , n238305 , n238306 );
not ( n238308 , n221637 );
not ( n238309 , n221633 );
not ( n238310 , n234108 );
or ( n238311 , n238309 , n238310 );
nand ( n238312 , n40625 , n221778 );
nand ( n238313 , n238311 , n238312 );
not ( n238314 , n238313 );
or ( n238315 , n238308 , n238314 );
nand ( n238316 , n237942 , n221626 );
nand ( n238317 , n238315 , n238316 );
xor ( n238318 , n238307 , n238317 );
not ( n238319 , n229964 );
not ( n238320 , n229261 );
not ( n238321 , n226724 );
or ( n238322 , n238320 , n238321 );
not ( n238323 , n39928 );
nand ( n238324 , n238323 , n234000 );
nand ( n238325 , n238322 , n238324 );
not ( n238326 , n238325 );
or ( n238327 , n238319 , n238326 );
nand ( n238328 , n238017 , n234006 );
nand ( n238329 , n238327 , n238328 );
xor ( n238330 , n238318 , n238329 );
xor ( n238331 , n238296 , n238330 );
xor ( n238332 , n238176 , n238184 );
and ( n238333 , n238332 , n238330 );
and ( n238334 , n238176 , n238184 );
or ( n238335 , n238333 , n238334 );
not ( n238336 , n237493 );
not ( n238337 , n222892 );
not ( n238338 , n237588 );
or ( n238339 , n238337 , n238338 );
nand ( n238340 , n236752 , n222458 );
nand ( n238341 , n238339 , n238340 );
not ( n238342 , n238341 );
or ( n238343 , n238336 , n238342 );
nand ( n238344 , n237952 , n237503 );
nand ( n238345 , n238343 , n238344 );
not ( n238346 , n219461 );
not ( n238347 , n237975 );
or ( n238348 , n238346 , n238347 );
not ( n238349 , n218775 );
not ( n238350 , n237600 );
or ( n238351 , n238349 , n238350 );
not ( n238352 , n218205 );
nand ( n238353 , n235031 , n238352 );
nand ( n238354 , n238351 , n238353 );
nand ( n238355 , n238354 , n218533 );
nand ( n238356 , n238348 , n238355 );
xor ( n238357 , n238345 , n238356 );
not ( n238358 , n218843 );
not ( n238359 , n221241 );
not ( n238360 , n227004 );
or ( n238361 , n238359 , n238360 );
not ( n238362 , n233035 );
not ( n238363 , n221241 );
nand ( n238364 , n238362 , n238363 );
nand ( n238365 , n238361 , n238364 );
not ( n238366 , n238365 );
or ( n238367 , n238358 , n238366 );
nand ( n238368 , n237877 , n223665 );
nand ( n238369 , n238367 , n238368 );
xor ( n238370 , n238357 , n238369 );
not ( n238371 , n220507 );
not ( n238372 , n237890 );
or ( n238373 , n238371 , n238372 );
not ( n238374 , n236241 );
not ( n238375 , n40181 );
or ( n238376 , n238374 , n238375 );
not ( n238377 , n221712 );
nand ( n238378 , n238377 , n219423 );
nand ( n238379 , n238376 , n238378 );
nand ( n238380 , n238379 , n219076 );
nand ( n238381 , n238373 , n238380 );
not ( n238382 , n222414 );
not ( n238383 , n223384 );
not ( n238384 , n238383 );
or ( n238385 , n238382 , n238384 );
not ( n238386 , n226911 );
nand ( n238387 , n238386 , n220150 );
nand ( n238388 , n238385 , n238387 );
not ( n238389 , n238388 );
not ( n238390 , n219779 );
or ( n238391 , n238389 , n238390 );
nand ( n238392 , n220492 , n237901 );
nand ( n238393 , n238391 , n238392 );
xor ( n238394 , n238381 , n238393 );
not ( n238395 , n237922 );
xor ( n238396 , n238394 , n238395 );
xor ( n238397 , n238370 , n238396 );
and ( n238398 , n234382 , n237483 );
not ( n238399 , n227294 );
not ( n238400 , n223182 );
not ( n238401 , n219596 );
or ( n238402 , n238400 , n238401 );
not ( n238403 , n219596 );
not ( n238404 , n223182 );
nand ( n238405 , n238403 , n238404 );
nand ( n238406 , n238402 , n238405 );
not ( n238407 , n238406 );
or ( n238408 , n238399 , n238407 );
not ( n238409 , n236338 );
nand ( n238410 , n238004 , n238409 );
nand ( n238411 , n238408 , n238410 );
xor ( n238412 , n238398 , n238411 );
not ( n238413 , n220059 );
not ( n238414 , n237965 );
or ( n238415 , n238413 , n238414 );
not ( n238416 , n226961 );
not ( n238417 , n217616 );
or ( n238418 , n238416 , n238417 );
nand ( n238419 , n39997 , n234015 );
nand ( n238420 , n238418 , n238419 );
nand ( n238421 , n238420 , n220067 );
nand ( n238422 , n238415 , n238421 );
xor ( n238423 , n238412 , n238422 );
xor ( n238424 , n238397 , n238423 );
xor ( n238425 , n238370 , n238396 );
and ( n238426 , n238425 , n238423 );
and ( n238427 , n238370 , n238396 );
or ( n238428 , n238426 , n238427 );
xor ( n238429 , n237825 , n237858 );
xor ( n238430 , n238429 , n238212 );
xor ( n238431 , n238180 , n238430 );
xor ( n238432 , n238431 , n238188 );
xor ( n238433 , n238180 , n238430 );
and ( n238434 , n238433 , n238188 );
and ( n238435 , n238180 , n238430 );
or ( n238436 , n238434 , n238435 );
not ( n238437 , n223949 );
not ( n238438 , n226655 );
not ( n238439 , n232842 );
or ( n238440 , n238438 , n238439 );
nand ( n238441 , n39607 , n227927 );
nand ( n238442 , n238440 , n238441 );
not ( n238443 , n238442 );
or ( n238444 , n238437 , n238443 );
nand ( n238445 , n238056 , n227260 );
nand ( n238446 , n238444 , n238445 );
not ( n238447 , n219314 );
not ( n238448 , n219687 );
not ( n238449 , n235691 );
not ( n238450 , n238449 );
or ( n238451 , n238448 , n238450 );
nand ( n238452 , n235691 , n222323 );
nand ( n238453 , n238451 , n238452 );
not ( n238454 , n238453 );
or ( n238455 , n238447 , n238454 );
nand ( n238456 , n238088 , n216204 );
nand ( n238457 , n238455 , n238456 );
xor ( n238458 , n238446 , n238457 );
not ( n238459 , n219501 );
not ( n238460 , n229387 );
not ( n238461 , n225792 );
or ( n238462 , n238460 , n238461 );
nand ( n238463 , n227696 , n227599 );
nand ( n238464 , n238462 , n238463 );
not ( n238465 , n238464 );
or ( n238466 , n238459 , n238465 );
nand ( n238467 , n238064 , n225478 );
nand ( n238468 , n238466 , n238467 );
xor ( n238469 , n238458 , n238468 );
not ( n238470 , n222185 );
not ( n238471 , n219033 );
buf ( n238472 , n209961 );
not ( n238473 , n238472 );
not ( n238474 , n238473 );
or ( n238475 , n238471 , n238474 );
nand ( n238476 , n238472 , n219034 );
nand ( n238477 , n238475 , n238476 );
not ( n238478 , n238477 );
or ( n238479 , n238470 , n238478 );
nand ( n238480 , n238029 , n219731 );
nand ( n238481 , n238479 , n238480 );
not ( n238482 , n219332 );
not ( n238483 , n238038 );
or ( n238484 , n238482 , n238483 );
not ( n238485 , n226484 );
not ( n238486 , n236840 );
not ( n238487 , n238486 );
or ( n238488 , n238485 , n238487 );
nand ( n238489 , n236840 , n221938 );
nand ( n238490 , n238488 , n238489 );
nand ( n238491 , n238490 , n221933 );
nand ( n238492 , n238484 , n238491 );
xor ( n238493 , n238481 , n238492 );
not ( n238494 , n226287 );
and ( n238495 , n227912 , n38532 );
not ( n238496 , n227912 );
and ( n238497 , n238496 , n235962 );
nor ( n238498 , n238495 , n238497 );
not ( n238499 , n238498 );
or ( n238500 , n238494 , n238499 );
nand ( n238501 , n238076 , n220414 );
nand ( n238502 , n238500 , n238501 );
xor ( n238503 , n238493 , n238502 );
xor ( n238504 , n238469 , n238503 );
xor ( n238505 , n238504 , n237870 );
xor ( n238506 , n238469 , n238503 );
and ( n238507 , n238506 , n237870 );
and ( n238508 , n238469 , n238503 );
or ( n238509 , n238507 , n238508 );
xor ( n238510 , n237864 , n238285 );
xor ( n238511 , n238510 , n237910 );
xor ( n238512 , n237864 , n238285 );
and ( n238513 , n238512 , n237910 );
and ( n238514 , n237864 , n238285 );
or ( n238515 , n238513 , n238514 );
xor ( n238516 , n237986 , n238291 );
xor ( n238517 , n238516 , n238424 );
xor ( n238518 , n237986 , n238291 );
and ( n238519 , n238518 , n238424 );
and ( n238520 , n237986 , n238291 );
or ( n238521 , n238519 , n238520 );
xor ( n238522 , n238331 , n238048 );
xor ( n238523 , n238522 , n238102 );
xor ( n238524 , n238331 , n238048 );
and ( n238525 , n238524 , n238102 );
and ( n238526 , n238331 , n238048 );
or ( n238527 , n238525 , n238526 );
xor ( n238528 , n238505 , n238432 );
xor ( n238529 , n238528 , n238108 );
xor ( n238530 , n238505 , n238432 );
and ( n238531 , n238530 , n238108 );
and ( n238532 , n238505 , n238432 );
or ( n238533 , n238531 , n238532 );
xor ( n238534 , n238262 , n238269 );
and ( n238535 , n238534 , n238282 );
and ( n238536 , n238262 , n238269 );
or ( n238537 , n238535 , n238536 );
xor ( n238538 , n238511 , n238114 );
xor ( n238539 , n238538 , n238517 );
xor ( n238540 , n238511 , n238114 );
and ( n238541 , n238540 , n238517 );
and ( n238542 , n238511 , n238114 );
or ( n238543 , n238541 , n238542 );
xor ( n238544 , n238120 , n238523 );
xor ( n238545 , n238544 , n238529 );
xor ( n238546 , n238120 , n238523 );
and ( n238547 , n238546 , n238529 );
and ( n238548 , n238120 , n238523 );
or ( n238549 , n238547 , n238548 );
xor ( n238550 , n238126 , n238136 );
xor ( n238551 , n238550 , n238539 );
xor ( n238552 , n238126 , n238136 );
and ( n238553 , n238552 , n238539 );
and ( n238554 , n238126 , n238136 );
or ( n238555 , n238553 , n238554 );
xor ( n238556 , n238545 , n238142 );
xor ( n238557 , n238556 , n238148 );
xor ( n238558 , n238545 , n238142 );
and ( n238559 , n238558 , n238148 );
and ( n238560 , n238545 , n238142 );
or ( n238561 , n238559 , n238560 );
xor ( n238562 , n238551 , n238557 );
xor ( n238563 , n238562 , n238154 );
xor ( n238564 , n238551 , n238557 );
and ( n238565 , n238564 , n238154 );
and ( n238566 , n238551 , n238557 );
or ( n238567 , n238565 , n238566 );
xor ( n238568 , n238398 , n238411 );
and ( n238569 , n238568 , n238422 );
and ( n238570 , n238398 , n238411 );
or ( n238571 , n238569 , n238570 );
xor ( n238572 , n238345 , n238356 );
and ( n238573 , n238572 , n238369 );
and ( n238574 , n238345 , n238356 );
or ( n238575 , n238573 , n238574 );
xor ( n238576 , n238381 , n238393 );
and ( n238577 , n238576 , n238395 );
and ( n238578 , n238381 , n238393 );
or ( n238579 , n238577 , n238578 );
xor ( n238580 , n238307 , n238317 );
and ( n238581 , n238580 , n238329 );
and ( n238582 , n238307 , n238317 );
or ( n238583 , n238581 , n238582 );
xor ( n238584 , n238481 , n238492 );
and ( n238585 , n238584 , n238502 );
and ( n238586 , n238481 , n238492 );
or ( n238587 , n238585 , n238586 );
xor ( n238588 , n238446 , n238457 );
and ( n238589 , n238588 , n238468 );
and ( n238590 , n238446 , n238457 );
or ( n238591 , n238589 , n238590 );
xor ( n238592 , n237825 , n237858 );
and ( n238593 , n238592 , n238212 );
and ( n238594 , n237825 , n237858 );
or ( n238595 , n238593 , n238594 );
or ( n238596 , n234894 , n238232 );
and ( n238597 , n41319 , n230897 );
not ( n238598 , n41319 );
and ( n238599 , n238598 , n229823 );
nor ( n238600 , n238597 , n238599 );
or ( n238601 , n234896 , n238600 );
nand ( n238602 , n238596 , n238601 );
not ( n238603 , n238245 );
not ( n238604 , n237810 );
or ( n238605 , n238603 , n238604 );
not ( n238606 , n215796 );
not ( n238607 , n227596 );
or ( n238608 , n238606 , n238607 );
nand ( n238609 , n237816 , n232282 );
nand ( n238610 , n238608 , n238609 );
nand ( n238611 , n238240 , n238610 );
nand ( n238612 , n238605 , n238611 );
xor ( n238613 , n238602 , n238612 );
not ( n238614 , n231421 );
not ( n238615 , n238260 );
or ( n238616 , n238614 , n238615 );
not ( n238617 , n228850 );
and ( n238618 , n238617 , n226225 );
not ( n238619 , n231940 );
and ( n238620 , n238619 , n226224 );
nor ( n238621 , n238618 , n238620 );
or ( n238622 , n232454 , n238621 );
nand ( n238623 , n238616 , n238622 );
xor ( n238624 , n238613 , n238623 );
xor ( n238625 , n238602 , n238612 );
and ( n238626 , n238625 , n238623 );
and ( n238627 , n238602 , n238612 );
or ( n238628 , n238626 , n238627 );
or ( n238629 , n231474 , n238267 );
and ( n238630 , n226304 , n237014 );
not ( n238631 , n226304 );
and ( n238632 , n238631 , n229759 );
nor ( n238633 , n238630 , n238632 );
or ( n238634 , n231476 , n238633 );
nand ( n238635 , n238629 , n238634 );
not ( n238636 , n238209 );
not ( n238637 , n238636 );
not ( n238638 , n227792 );
or ( n238639 , n238637 , n238638 );
not ( n238640 , n219201 );
not ( n238641 , n238640 );
not ( n238642 , n238641 );
not ( n238643 , n237918 );
or ( n238644 , n238642 , n238643 );
nand ( n238645 , n233952 , n217330 );
nand ( n238646 , n238644 , n238645 );
nand ( n238647 , n237914 , n238646 );
nand ( n238648 , n238639 , n238647 );
xor ( n238649 , n238635 , n238648 );
not ( n238650 , n238280 );
not ( n238651 , n238650 );
not ( n238652 , n232399 );
or ( n238653 , n238651 , n238652 );
not ( n238654 , n224492 );
not ( n238655 , n230722 );
or ( n238656 , n238654 , n238655 );
nand ( n238657 , n234382 , n224496 );
nand ( n238658 , n238656 , n238657 );
nand ( n238659 , n238274 , n238658 );
nand ( n238660 , n238653 , n238659 );
xor ( n238661 , n238649 , n238660 );
xor ( n238662 , n238635 , n238648 );
and ( n238663 , n238662 , n238660 );
and ( n238664 , n238635 , n238648 );
or ( n238665 , n238663 , n238664 );
and ( n238666 , n231754 , n216293 );
not ( n238667 , n227782 );
not ( n238668 , n224096 );
not ( n238669 , n217964 );
or ( n238670 , n238668 , n238669 );
not ( n238671 , n219151 );
buf ( n238672 , n234764 );
nand ( n238673 , n238671 , n238672 );
nand ( n238674 , n238670 , n238673 );
not ( n238675 , n238674 );
or ( n238676 , n238667 , n238675 );
nand ( n238677 , n224087 , n238201 );
nand ( n238678 , n238676 , n238677 );
xor ( n238679 , n238666 , n238678 );
not ( n238680 , n227294 );
not ( n238681 , n223183 );
not ( n238682 , n238681 );
not ( n238683 , n40768 );
or ( n238684 , n238682 , n238683 );
nand ( n238685 , n221342 , n236547 );
nand ( n238686 , n238684 , n238685 );
not ( n238687 , n238686 );
or ( n238688 , n238680 , n238687 );
nand ( n238689 , n238406 , n235172 );
nand ( n238690 , n238688 , n238689 );
xor ( n238691 , n238679 , n238690 );
xor ( n238692 , n238579 , n238691 );
xor ( n238693 , n238692 , n238571 );
xor ( n238694 , n238579 , n238691 );
and ( n238695 , n238694 , n238571 );
and ( n238696 , n238579 , n238691 );
or ( n238697 , n238695 , n238696 );
xor ( n238698 , n238575 , n238583 );
xor ( n238699 , n238698 , n238587 );
xor ( n238700 , n238575 , n238583 );
and ( n238701 , n238700 , n238587 );
and ( n238702 , n238575 , n238583 );
or ( n238703 , n238701 , n238702 );
not ( n238704 , n221637 );
not ( n238705 , n221612 );
not ( n238706 , n238705 );
not ( n238707 , n219742 );
or ( n238708 , n238706 , n238707 );
nand ( n238709 , n235359 , n222586 );
nand ( n238710 , n238708 , n238709 );
not ( n238711 , n238710 );
or ( n238712 , n238704 , n238711 );
nand ( n238713 , n238313 , n221626 );
nand ( n238714 , n238712 , n238713 );
not ( n238715 , n237493 );
not ( n238716 , n222892 );
not ( n238717 , n219880 );
or ( n238718 , n238716 , n238717 );
not ( n238719 , n222430 );
nand ( n238720 , n219226 , n238719 );
nand ( n238721 , n238718 , n238720 );
not ( n238722 , n238721 );
or ( n238723 , n238715 , n238722 );
nand ( n238724 , n238341 , n237503 );
nand ( n238725 , n238723 , n238724 );
xor ( n238726 , n238714 , n238725 );
not ( n238727 , n220067 );
buf ( n238728 , n39877 );
and ( n238729 , n238728 , n231500 );
not ( n238730 , n238728 );
and ( n238731 , n238730 , n234015 );
or ( n238732 , n238729 , n238731 );
not ( n238733 , n238732 );
or ( n238734 , n238727 , n238733 );
nand ( n238735 , n238420 , n220059 );
nand ( n238736 , n238734 , n238735 );
xor ( n238737 , n238726 , n238736 );
not ( n238738 , n219461 );
not ( n238739 , n238354 );
or ( n238740 , n238738 , n238739 );
not ( n238741 , n233083 );
not ( n238742 , n230490 );
or ( n238743 , n238741 , n238742 );
nand ( n238744 , n237963 , n218226 );
nand ( n238745 , n238743 , n238744 );
nand ( n238746 , n238745 , n218232 );
nand ( n238747 , n238740 , n238746 );
not ( n238748 , n223665 );
not ( n238749 , n238365 );
or ( n238750 , n238748 , n238749 );
not ( n238751 , n221241 );
not ( n238752 , n236290 );
not ( n238753 , n238752 );
or ( n238754 , n238751 , n238753 );
not ( n238755 , n232413 );
nand ( n238756 , n236290 , n238755 );
nand ( n238757 , n238754 , n238756 );
nand ( n238758 , n238757 , n218843 );
nand ( n238759 , n238750 , n238758 );
xor ( n238760 , n238747 , n238759 );
not ( n238761 , n219076 );
not ( n238762 , n236241 );
not ( n238763 , n236301 );
or ( n238764 , n238762 , n238763 );
nand ( n238765 , n236304 , n219440 );
nand ( n238766 , n238764 , n238765 );
not ( n238767 , n238766 );
or ( n238768 , n238761 , n238767 );
nand ( n238769 , n238379 , n220507 );
nand ( n238770 , n238768 , n238769 );
xor ( n238771 , n238760 , n238770 );
xor ( n238772 , n238737 , n238771 );
not ( n238773 , n230389 );
not ( n238774 , n238221 );
and ( n238775 , n238773 , n238774 );
buf ( n238776 , n228775 );
not ( n238777 , n238776 );
and ( n238778 , n208164 , n232493 );
not ( n238779 , n208164 );
and ( n238780 , n238779 , n225952 );
nor ( n238781 , n238778 , n238780 );
nor ( n238782 , n238777 , n238781 );
nor ( n238783 , n238775 , n238782 );
not ( n238784 , n219779 );
not ( n238785 , n221593 );
buf ( n238786 , n230511 );
not ( n238787 , n238786 );
or ( n238788 , n238785 , n238787 );
buf ( n238789 , n226505 );
nand ( n238790 , n238789 , n222414 );
nand ( n238791 , n238788 , n238790 );
not ( n238792 , n238791 );
or ( n238793 , n238784 , n238792 );
nand ( n238794 , n238388 , n220164 );
nand ( n238795 , n238793 , n238794 );
xor ( n238796 , n238783 , n238795 );
not ( n238797 , n235913 );
not ( n238798 , n238303 );
or ( n238799 , n238797 , n238798 );
not ( n238800 , n220906 );
not ( n238801 , n221330 );
or ( n238802 , n238800 , n238801 );
nand ( n238803 , n221956 , n238301 );
nand ( n238804 , n238802 , n238803 );
nand ( n238805 , n238804 , n220930 );
nand ( n238806 , n238799 , n238805 );
xor ( n238807 , n238796 , n238806 );
xor ( n238808 , n238772 , n238807 );
xor ( n238809 , n238737 , n238771 );
and ( n238810 , n238809 , n238807 );
and ( n238811 , n238737 , n238771 );
or ( n238812 , n238810 , n238811 );
not ( n238813 , n234006 );
not ( n238814 , n238325 );
or ( n238815 , n238813 , n238814 );
not ( n238816 , n229261 );
not ( n238817 , n234350 );
or ( n238818 , n238816 , n238817 );
not ( n238819 , n234347 );
nand ( n238820 , n238819 , n229262 );
nand ( n238821 , n238818 , n238820 );
nand ( n238822 , n238821 , n229964 );
nand ( n238823 , n238815 , n238822 );
xor ( n238824 , n238216 , n238823 );
xor ( n238825 , n238824 , n238252 );
xor ( n238826 , n238591 , n238825 );
xor ( n238827 , n238826 , n238289 );
xor ( n238828 , n238591 , n238825 );
and ( n238829 , n238828 , n238289 );
and ( n238830 , n238591 , n238825 );
or ( n238831 , n238829 , n238830 );
not ( n238832 , n219314 );
and ( n238833 , n222323 , n234579 );
not ( n238834 , n222323 );
not ( n238835 , n234579 );
and ( n238836 , n238834 , n238835 );
nor ( n238837 , n238833 , n238836 );
not ( n238838 , n238837 );
or ( n238839 , n238832 , n238838 );
nand ( n238840 , n238453 , n216204 );
nand ( n238841 , n238839 , n238840 );
not ( n238842 , n226943 );
not ( n238843 , n238498 );
or ( n238844 , n238842 , n238843 );
not ( n238845 , n227912 );
not ( n238846 , n228165 );
or ( n238847 , n238845 , n238846 );
nand ( n238848 , n39365 , n220038 );
nand ( n238849 , n238847 , n238848 );
nand ( n238850 , n238849 , n226287 );
nand ( n238851 , n238844 , n238850 );
xor ( n238852 , n238841 , n238851 );
not ( n238853 , n223949 );
not ( n238854 , n226655 );
not ( n238855 , n227201 );
or ( n238856 , n238854 , n238855 );
not ( n238857 , n227201 );
nand ( n238858 , n238857 , n233053 );
nand ( n238859 , n238856 , n238858 );
not ( n238860 , n238859 );
or ( n238861 , n238853 , n238860 );
nand ( n238862 , n238442 , n227260 );
nand ( n238863 , n238861 , n238862 );
xor ( n238864 , n238852 , n238863 );
xor ( n238865 , n238595 , n238864 );
not ( n238866 , n219731 );
not ( n238867 , n238477 );
or ( n238868 , n238866 , n238867 );
nand ( n238869 , n222185 , n219033 );
nand ( n238870 , n238868 , n238869 );
not ( n238871 , n229395 );
not ( n238872 , n238464 );
or ( n238873 , n238871 , n238872 );
not ( n238874 , n233544 );
not ( n238875 , n235516 );
or ( n238876 , n238874 , n238875 );
not ( n238877 , n235516 );
nand ( n238878 , n238877 , n237203 );
nand ( n238879 , n238876 , n238878 );
nand ( n238880 , n238879 , n219501 );
nand ( n238881 , n238873 , n238880 );
xor ( n238882 , n238870 , n238881 );
not ( n238883 , n221933 );
not ( n238884 , n226484 );
not ( n238885 , n237271 );
or ( n238886 , n238884 , n238885 );
not ( n238887 , n230219 );
nand ( n238888 , n238887 , n221938 );
nand ( n238889 , n238886 , n238888 );
not ( n238890 , n238889 );
or ( n238891 , n238883 , n238890 );
nand ( n238892 , n238490 , n219332 );
nand ( n238893 , n238891 , n238892 );
xor ( n238894 , n238882 , n238893 );
xor ( n238895 , n238865 , n238894 );
xor ( n238896 , n238595 , n238864 );
and ( n238897 , n238896 , n238894 );
and ( n238898 , n238595 , n238864 );
or ( n238899 , n238897 , n238898 );
xor ( n238900 , n238537 , n238661 );
xor ( n238901 , n238900 , n238624 );
xor ( n238902 , n238295 , n238901 );
xor ( n238903 , n238902 , n238428 );
xor ( n238904 , n238295 , n238901 );
and ( n238905 , n238904 , n238428 );
and ( n238906 , n238295 , n238901 );
or ( n238907 , n238905 , n238906 );
xor ( n238908 , n238335 , n238693 );
xor ( n238909 , n238908 , n238699 );
xor ( n238910 , n238335 , n238693 );
and ( n238911 , n238910 , n238699 );
and ( n238912 , n238335 , n238693 );
or ( n238913 , n238911 , n238912 );
xor ( n238914 , n238436 , n238808 );
xor ( n238915 , n238914 , n238509 );
xor ( n238916 , n238436 , n238808 );
and ( n238917 , n238916 , n238509 );
and ( n238918 , n238436 , n238808 );
or ( n238919 , n238917 , n238918 );
xor ( n238920 , n238895 , n238827 );
xor ( n238921 , n238920 , n238515 );
xor ( n238922 , n238895 , n238827 );
and ( n238923 , n238922 , n238515 );
and ( n238924 , n238895 , n238827 );
or ( n238925 , n238923 , n238924 );
xor ( n238926 , n238903 , n238909 );
xor ( n238927 , n238926 , n238521 );
xor ( n238928 , n238903 , n238909 );
and ( n238929 , n238928 , n238521 );
and ( n238930 , n238903 , n238909 );
or ( n238931 , n238929 , n238930 );
xor ( n238932 , n238666 , n238678 );
and ( n238933 , n238932 , n238690 );
and ( n238934 , n238666 , n238678 );
or ( n238935 , n238933 , n238934 );
xor ( n238936 , n238527 , n238915 );
xor ( n238937 , n238936 , n238533 );
xor ( n238938 , n238527 , n238915 );
and ( n238939 , n238938 , n238533 );
and ( n238940 , n238527 , n238915 );
or ( n238941 , n238939 , n238940 );
xor ( n238942 , n238921 , n238543 );
xor ( n238943 , n238942 , n238927 );
xor ( n238944 , n238921 , n238543 );
and ( n238945 , n238944 , n238927 );
and ( n238946 , n238921 , n238543 );
or ( n238947 , n238945 , n238946 );
xor ( n238948 , n238937 , n238549 );
xor ( n238949 , n238948 , n238555 );
xor ( n238950 , n238937 , n238549 );
and ( n238951 , n238950 , n238555 );
and ( n238952 , n238937 , n238549 );
or ( n238953 , n238951 , n238952 );
xor ( n238954 , n238943 , n238949 );
xor ( n238955 , n238954 , n238561 );
xor ( n238956 , n238943 , n238949 );
and ( n238957 , n238956 , n238561 );
and ( n238958 , n238943 , n238949 );
or ( n238959 , n238957 , n238958 );
xor ( n238960 , n238747 , n238759 );
and ( n238961 , n238960 , n238770 );
and ( n238962 , n238747 , n238759 );
or ( n238963 , n238961 , n238962 );
xor ( n238964 , n238783 , n238795 );
and ( n238965 , n238964 , n238806 );
and ( n238966 , n238783 , n238795 );
or ( n238967 , n238965 , n238966 );
xor ( n238968 , n238714 , n238725 );
and ( n238969 , n238968 , n238736 );
and ( n238970 , n238714 , n238725 );
or ( n238971 , n238969 , n238970 );
xor ( n238972 , n238841 , n238851 );
and ( n238973 , n238972 , n238863 );
and ( n238974 , n238841 , n238851 );
or ( n238975 , n238973 , n238974 );
xor ( n238976 , n238870 , n238881 );
and ( n238977 , n238976 , n238893 );
and ( n238978 , n238870 , n238881 );
or ( n238979 , n238977 , n238978 );
xor ( n238980 , n238216 , n238823 );
and ( n238981 , n238980 , n238252 );
and ( n238982 , n238216 , n238823 );
or ( n238983 , n238981 , n238982 );
xor ( n238984 , n238537 , n238661 );
and ( n238985 , n238984 , n238624 );
and ( n238986 , n238537 , n238661 );
or ( n238987 , n238985 , n238986 );
or ( n238988 , n219731 , n222185 );
nand ( n238989 , n238988 , n219033 );
not ( n238990 , n238646 );
or ( n238991 , n235195 , n238990 );
and ( n238992 , n235200 , n219389 );
not ( n238993 , n235200 );
and ( n238994 , n238993 , n220823 );
nor ( n238995 , n238992 , n238994 );
or ( n238996 , n238995 , n232948 );
nand ( n238997 , n238991 , n238996 );
xor ( n238998 , n238989 , n238997 );
not ( n238999 , n232956 );
or ( n239000 , n238999 , n238781 );
buf ( n239001 , n220226 );
and ( n239002 , n239001 , n232493 );
not ( n239003 , n239001 );
and ( n239004 , n239003 , n229806 );
or ( n239005 , n239002 , n239004 );
not ( n239006 , n239005 );
or ( n239007 , n231456 , n239006 );
nand ( n239008 , n239000 , n239007 );
xor ( n239009 , n238998 , n239008 );
xor ( n239010 , n238989 , n238997 );
and ( n239011 , n239010 , n239008 );
and ( n239012 , n238989 , n238997 );
or ( n239013 , n239011 , n239012 );
not ( n239014 , n238600 );
not ( n239015 , n239014 );
not ( n239016 , n229816 );
or ( n239017 , n239015 , n239016 );
not ( n239018 , n238218 );
not ( n239019 , n234293 );
or ( n239020 , n239018 , n239019 );
not ( n239021 , n226650 );
nand ( n239022 , n239021 , n217697 );
nand ( n239023 , n239020 , n239022 );
nand ( n239024 , n226885 , n239023 );
nand ( n239025 , n239017 , n239024 );
not ( n239026 , n238610 );
not ( n239027 , n237810 );
or ( n239028 , n239026 , n239027 );
not ( n239029 , n234751 );
not ( n239030 , n234394 );
or ( n239031 , n239029 , n239030 );
nand ( n239032 , n237816 , n217130 );
nand ( n239033 , n239031 , n239032 );
nand ( n239034 , n227737 , n239033 );
nand ( n239035 , n239028 , n239034 );
xor ( n239036 , n239025 , n239035 );
or ( n239037 , n237038 , n238621 );
and ( n239038 , n41565 , n229249 );
not ( n239039 , n41565 );
and ( n239040 , n239039 , n238619 );
or ( n239041 , n239038 , n239040 );
not ( n239042 , n239041 );
or ( n239043 , n232454 , n239042 );
nand ( n239044 , n239037 , n239043 );
xor ( n239045 , n239036 , n239044 );
xor ( n239046 , n239025 , n239035 );
and ( n239047 , n239046 , n239044 );
and ( n239048 , n239025 , n239035 );
or ( n239049 , n239047 , n239048 );
xor ( n239050 , n239045 , n238935 );
xor ( n239051 , n239050 , n238963 );
xor ( n239052 , n239045 , n238935 );
and ( n239053 , n239052 , n238963 );
and ( n239054 , n239045 , n238935 );
or ( n239055 , n239053 , n239054 );
xor ( n239056 , n238967 , n238971 );
xor ( n239057 , n239056 , n238975 );
xor ( n239058 , n238967 , n238971 );
and ( n239059 , n239058 , n238975 );
and ( n239060 , n238967 , n238971 );
or ( n239061 , n239059 , n239060 );
not ( n239062 , n220930 );
not ( n239063 , n222399 );
not ( n239064 , n40258 );
or ( n239065 , n239063 , n239064 );
not ( n239066 , n220906 );
nand ( n239067 , n220970 , n239066 );
nand ( n239068 , n239065 , n239067 );
not ( n239069 , n239068 );
or ( n239070 , n239062 , n239069 );
nand ( n239071 , n235913 , n238804 );
nand ( n239072 , n239070 , n239071 );
not ( n239073 , n238783 );
xor ( n239074 , n239072 , n239073 );
not ( n239075 , n221637 );
not ( n239076 , n237937 );
not ( n239077 , n234014 );
not ( n239078 , n239077 );
or ( n239079 , n239076 , n239078 );
not ( n239080 , n226921 );
nand ( n239081 , n239080 , n221612 );
nand ( n239082 , n239079 , n239081 );
not ( n239083 , n239082 );
or ( n239084 , n239075 , n239083 );
nand ( n239085 , n238710 , n221626 );
nand ( n239086 , n239084 , n239085 );
xor ( n239087 , n239074 , n239086 );
xor ( n239088 , n238979 , n239087 );
not ( n239089 , n227782 );
not ( n239090 , n237130 );
not ( n239091 , n237496 );
or ( n239092 , n239090 , n239091 );
nand ( n239093 , n219599 , n224095 );
nand ( n239094 , n239092 , n239093 );
not ( n239095 , n239094 );
or ( n239096 , n239089 , n239095 );
nand ( n239097 , n238674 , n224087 );
nand ( n239098 , n239096 , n239097 );
not ( n239099 , n219461 );
not ( n239100 , n238745 );
or ( n239101 , n239099 , n239100 );
not ( n239102 , n218205 );
not ( n239103 , n235921 );
or ( n239104 , n239102 , n239103 );
nand ( n239105 , n229928 , n218256 );
nand ( n239106 , n239104 , n239105 );
nand ( n239107 , n239106 , n218533 );
nand ( n239108 , n239101 , n239107 );
xor ( n239109 , n239098 , n239108 );
not ( n239110 , n227294 );
and ( n239111 , n238404 , n218912 );
not ( n239112 , n238404 );
and ( n239113 , n239112 , n236752 );
nor ( n239114 , n239111 , n239113 );
not ( n239115 , n239114 );
or ( n239116 , n239110 , n239115 );
nand ( n239117 , n238686 , n235172 );
nand ( n239118 , n239116 , n239117 );
xor ( n239119 , n239109 , n239118 );
xor ( n239120 , n239088 , n239119 );
xor ( n239121 , n238979 , n239087 );
and ( n239122 , n239121 , n239119 );
and ( n239123 , n238979 , n239087 );
or ( n239124 , n239122 , n239123 );
not ( n239125 , n223665 );
not ( n239126 , n238757 );
or ( n239127 , n239125 , n239126 );
not ( n239128 , n221241 );
not ( n239129 , n237600 );
or ( n239130 , n239128 , n239129 );
nand ( n239131 , n235031 , n238755 );
nand ( n239132 , n239130 , n239131 );
nand ( n239133 , n239132 , n218843 );
nand ( n239134 , n239127 , n239133 );
not ( n239135 , n219076 );
not ( n239136 , n236241 );
not ( n239137 , n227004 );
or ( n239138 , n239136 , n239137 );
not ( n239139 , n227004 );
nand ( n239140 , n239139 , n219797 );
nand ( n239141 , n239138 , n239140 );
not ( n239142 , n239141 );
or ( n239143 , n239135 , n239142 );
nand ( n239144 , n238766 , n220507 );
nand ( n239145 , n239143 , n239144 );
xor ( n239146 , n239134 , n239145 );
not ( n239147 , n220164 );
not ( n239148 , n238791 );
or ( n239149 , n239147 , n239148 );
not ( n239150 , n221593 );
not ( n239151 , n229936 );
or ( n239152 , n239150 , n239151 );
nand ( n239153 , n238377 , n222414 );
nand ( n239154 , n239152 , n239153 );
nand ( n239155 , n239154 , n220881 );
nand ( n239156 , n239149 , n239155 );
xor ( n239157 , n239146 , n239156 );
xor ( n239158 , n239157 , n238983 );
not ( n239159 , n237503 );
not ( n239160 , n238721 );
or ( n239161 , n239159 , n239160 );
not ( n239162 , n222430 );
not ( n239163 , n219518 );
or ( n239164 , n239162 , n239163 );
nand ( n239165 , n40625 , n238719 );
nand ( n239166 , n239164 , n239165 );
nand ( n239167 , n239166 , n237493 );
nand ( n239168 , n239161 , n239167 );
not ( n239169 , n220067 );
not ( n239170 , n231500 );
not ( n239171 , n226724 );
or ( n239172 , n239170 , n239171 );
not ( n239173 , n226724 );
nand ( n239174 , n239173 , n231501 );
nand ( n239175 , n239172 , n239174 );
not ( n239176 , n239175 );
or ( n239177 , n239169 , n239176 );
nand ( n239178 , n238732 , n220059 );
nand ( n239179 , n239177 , n239178 );
xor ( n239180 , n239168 , n239179 );
not ( n239181 , n224624 );
not ( n239182 , n238837 );
or ( n239183 , n239181 , n239182 );
not ( n239184 , n222323 );
buf ( n239185 , n231104 );
not ( n239186 , n239185 );
not ( n239187 , n239186 );
or ( n239188 , n239184 , n239187 );
not ( n239189 , n238472 );
or ( n239190 , n239189 , n222323 );
nand ( n239191 , n239188 , n239190 );
not ( n239192 , n239191 );
nand ( n239193 , n239192 , n219314 );
nand ( n239194 , n239183 , n239193 );
xor ( n239195 , n239180 , n239194 );
xor ( n239196 , n239158 , n239195 );
xor ( n239197 , n239157 , n238983 );
and ( n239198 , n239197 , n239195 );
and ( n239199 , n239157 , n238983 );
or ( n239200 , n239198 , n239199 );
not ( n239201 , n219332 );
not ( n239202 , n238889 );
or ( n239203 , n239201 , n239202 );
not ( n239204 , n226484 );
not ( n239205 , n238449 );
or ( n239206 , n239204 , n239205 );
nand ( n239207 , n235691 , n221938 );
nand ( n239208 , n239206 , n239207 );
nand ( n239209 , n239208 , n221933 );
nand ( n239210 , n239203 , n239209 );
xor ( n239211 , n239210 , n238628 );
not ( n239212 , n229964 );
not ( n239213 , n229261 );
not ( n239214 , n227696 );
not ( n239215 , n239214 );
or ( n239216 , n239213 , n239215 );
nand ( n239217 , n39714 , n234000 );
nand ( n239218 , n239216 , n239217 );
not ( n239219 , n239218 );
or ( n239220 , n239212 , n239219 );
nand ( n239221 , n238821 , n234006 );
nand ( n239222 , n239220 , n239221 );
xor ( n239223 , n239211 , n239222 );
xor ( n239224 , n238987 , n239223 );
not ( n239225 , n226943 );
not ( n239226 , n238849 );
or ( n239227 , n239225 , n239226 );
not ( n239228 , n227912 );
not ( n239229 , n39287 );
or ( n239230 , n239228 , n239229 );
nand ( n239231 , n236840 , n220038 );
nand ( n239232 , n239230 , n239231 );
nand ( n239233 , n239232 , n226287 );
nand ( n239234 , n239227 , n239233 );
not ( n239235 , n227260 );
not ( n239236 , n238859 );
or ( n239237 , n239235 , n239236 );
and ( n239238 , n229704 , n226655 );
not ( n239239 , n229704 );
and ( n239240 , n239239 , n233053 );
or ( n239241 , n239238 , n239240 );
nand ( n239242 , n239241 , n223949 );
nand ( n239243 , n239237 , n239242 );
xor ( n239244 , n239234 , n239243 );
not ( n239245 , n219501 );
not ( n239246 , n233544 );
not ( n239247 , n232842 );
or ( n239248 , n239246 , n239247 );
nand ( n239249 , n39608 , n227599 );
nand ( n239250 , n239248 , n239249 );
not ( n239251 , n239250 );
or ( n239252 , n239245 , n239251 );
nand ( n239253 , n238879 , n229395 );
nand ( n239254 , n239252 , n239253 );
xor ( n239255 , n239244 , n239254 );
xor ( n239256 , n239224 , n239255 );
xor ( n239257 , n238987 , n239223 );
and ( n239258 , n239257 , n239255 );
and ( n239259 , n238987 , n239223 );
or ( n239260 , n239258 , n239259 );
or ( n239261 , n231474 , n238633 );
and ( n239262 , n225769 , n231480 );
not ( n239263 , n225769 );
and ( n239264 , n239263 , n233399 );
nor ( n239265 , n239262 , n239264 );
or ( n239266 , n231476 , n239265 );
nand ( n239267 , n239261 , n239266 );
not ( n239268 , n238658 );
not ( n239269 , n233879 );
not ( n239270 , n239269 );
not ( n239271 , n239270 );
or ( n239272 , n239268 , n239271 );
not ( n239273 , n214837 );
not ( n239274 , n230722 );
or ( n239275 , n239273 , n239274 );
nand ( n239276 , n234382 , n226698 );
nand ( n239277 , n239275 , n239276 );
nand ( n239278 , n238274 , n239277 );
nand ( n239279 , n239272 , n239278 );
xor ( n239280 , n239267 , n239279 );
not ( n239281 , n230725 );
and ( n239282 , n239281 , n224037 );
xor ( n239283 , n239280 , n239282 );
xor ( n239284 , n238665 , n239283 );
xor ( n239285 , n239284 , n239009 );
xor ( n239286 , n238697 , n239285 );
xor ( n239287 , n239286 , n239051 );
xor ( n239288 , n238697 , n239285 );
and ( n239289 , n239288 , n239051 );
and ( n239290 , n238697 , n239285 );
or ( n239291 , n239289 , n239290 );
xor ( n239292 , n238703 , n238812 );
xor ( n239293 , n239292 , n238899 );
xor ( n239294 , n238703 , n238812 );
and ( n239295 , n239294 , n238899 );
and ( n239296 , n238703 , n238812 );
or ( n239297 , n239295 , n239296 );
xor ( n239298 , n238831 , n239196 );
xor ( n239299 , n239298 , n239120 );
xor ( n239300 , n238831 , n239196 );
and ( n239301 , n239300 , n239120 );
and ( n239302 , n238831 , n239196 );
or ( n239303 , n239301 , n239302 );
xor ( n239304 , n239057 , n239256 );
xor ( n239305 , n239304 , n239287 );
xor ( n239306 , n239057 , n239256 );
and ( n239307 , n239306 , n239287 );
and ( n239308 , n239057 , n239256 );
or ( n239309 , n239307 , n239308 );
xor ( n239310 , n238907 , n239293 );
xor ( n239311 , n239310 , n238913 );
xor ( n239312 , n238907 , n239293 );
and ( n239313 , n239312 , n238913 );
and ( n239314 , n238907 , n239293 );
or ( n239315 , n239313 , n239314 );
xor ( n239316 , n239267 , n239279 );
and ( n239317 , n239316 , n239282 );
and ( n239318 , n239267 , n239279 );
or ( n239319 , n239317 , n239318 );
xor ( n239320 , n238919 , n239299 );
xor ( n239321 , n239320 , n238925 );
xor ( n239322 , n238919 , n239299 );
and ( n239323 , n239322 , n238925 );
and ( n239324 , n238919 , n239299 );
or ( n239325 , n239323 , n239324 );
xor ( n239326 , n239305 , n238931 );
xor ( n239327 , n239326 , n239311 );
xor ( n239328 , n239305 , n238931 );
and ( n239329 , n239328 , n239311 );
and ( n239330 , n239305 , n238931 );
or ( n239331 , n239329 , n239330 );
xor ( n239332 , n239321 , n238941 );
xor ( n239333 , n239332 , n238947 );
xor ( n239334 , n239321 , n238941 );
and ( n239335 , n239334 , n238947 );
and ( n239336 , n239321 , n238941 );
or ( n239337 , n239335 , n239336 );
xor ( n239338 , n239327 , n239333 );
xor ( n239339 , n239338 , n238953 );
xor ( n239340 , n239327 , n239333 );
and ( n239341 , n239340 , n238953 );
and ( n239342 , n239327 , n239333 );
or ( n239343 , n239341 , n239342 );
xor ( n239344 , n239098 , n239108 );
and ( n239345 , n239344 , n239118 );
and ( n239346 , n239098 , n239108 );
or ( n239347 , n239345 , n239346 );
xor ( n239348 , n239134 , n239145 );
and ( n239349 , n239348 , n239156 );
and ( n239350 , n239134 , n239145 );
or ( n239351 , n239349 , n239350 );
xor ( n239352 , n239072 , n239073 );
and ( n239353 , n239352 , n239086 );
and ( n239354 , n239072 , n239073 );
or ( n239355 , n239353 , n239354 );
xor ( n239356 , n239168 , n239179 );
and ( n239357 , n239356 , n239194 );
and ( n239358 , n239168 , n239179 );
or ( n239359 , n239357 , n239358 );
xor ( n239360 , n239234 , n239243 );
and ( n239361 , n239360 , n239254 );
and ( n239362 , n239234 , n239243 );
or ( n239363 , n239361 , n239362 );
xor ( n239364 , n239210 , n238628 );
and ( n239365 , n239364 , n239222 );
and ( n239366 , n239210 , n238628 );
or ( n239367 , n239365 , n239366 );
xor ( n239368 , n238665 , n239283 );
and ( n239369 , n239368 , n239009 );
and ( n239370 , n238665 , n239283 );
or ( n239371 , n239369 , n239370 );
not ( n239372 , n239033 );
not ( n239373 , n232440 );
or ( n239374 , n239372 , n239373 );
not ( n239375 , n41321 );
not ( n239376 , n233451 );
or ( n239377 , n239375 , n239376 );
nand ( n239378 , n233450 , n216307 );
nand ( n239379 , n239377 , n239378 );
nand ( n239380 , n227737 , n239379 );
nand ( n239381 , n239374 , n239380 );
not ( n239382 , n239041 );
not ( n239383 , n231421 );
or ( n239384 , n239382 , n239383 );
and ( n239385 , n215796 , n236643 );
not ( n239386 , n215796 );
and ( n239387 , n239386 , n238619 );
or ( n239388 , n239385 , n239387 );
nand ( n239389 , n234404 , n239388 );
nand ( n239390 , n239384 , n239389 );
xor ( n239391 , n239381 , n239390 );
or ( n239392 , n231474 , n239265 );
not ( n239393 , n233399 );
and ( n239394 , n234256 , n239393 );
not ( n239395 , n234256 );
and ( n239396 , n239395 , n237014 );
nor ( n239397 , n239394 , n239396 );
or ( n239398 , n237013 , n239397 );
nand ( n239399 , n239392 , n239398 );
xor ( n239400 , n239391 , n239399 );
xor ( n239401 , n239381 , n239390 );
and ( n239402 , n239401 , n239399 );
and ( n239403 , n239381 , n239390 );
or ( n239404 , n239402 , n239403 );
not ( n239405 , n239277 );
not ( n239406 , n233105 );
or ( n239407 , n239405 , n239406 );
not ( n239408 , n209437 );
not ( n239409 , n230725 );
or ( n239410 , n239408 , n239409 );
nand ( n239411 , n232784 , n208726 );
nand ( n239412 , n239410 , n239411 );
nand ( n239413 , n232402 , n239412 );
nand ( n239414 , n239407 , n239413 );
not ( n239415 , n239005 );
buf ( n239416 , n230390 );
not ( n239417 , n239416 );
or ( n239418 , n239415 , n239417 );
not ( n239419 , n217331 );
not ( n239420 , n232497 );
or ( n239421 , n239419 , n239420 );
nand ( n239422 , n225952 , n222984 );
nand ( n239423 , n239421 , n239422 );
nand ( n239424 , n228775 , n239423 );
nand ( n239425 , n239418 , n239424 );
xor ( n239426 , n239414 , n239425 );
and ( n239427 , n233891 , n224492 );
xor ( n239428 , n239426 , n239427 );
xor ( n239429 , n239414 , n239425 );
and ( n239430 , n239429 , n239427 );
and ( n239431 , n239414 , n239425 );
or ( n239432 , n239430 , n239431 );
xor ( n239433 , n239347 , n239351 );
xor ( n239434 , n239433 , n239359 );
xor ( n239435 , n239347 , n239351 );
and ( n239436 , n239435 , n239359 );
and ( n239437 , n239347 , n239351 );
or ( n239438 , n239436 , n239437 );
xor ( n239439 , n239363 , n239367 );
not ( n239440 , n239023 );
buf ( n239441 , n229816 );
not ( n239442 , n239441 );
or ( n239443 , n239440 , n239442 );
not ( n239444 , n238230 );
not ( n239445 , n208166 );
or ( n239446 , n239444 , n239445 );
nand ( n239447 , n226651 , n40888 );
nand ( n239448 , n239446 , n239447 );
nand ( n239449 , n227852 , n239448 );
nand ( n239450 , n239443 , n239449 );
not ( n239451 , n239450 );
not ( n239452 , n222471 );
not ( n239453 , n239452 );
not ( n239454 , n239082 );
or ( n239455 , n239453 , n239454 );
and ( n239456 , n237937 , n223786 );
not ( n239457 , n237937 );
not ( n239458 , n220596 );
and ( n239459 , n239457 , n239458 );
or ( n239460 , n239456 , n239459 );
nand ( n239461 , n239460 , n221637 );
nand ( n239462 , n239455 , n239461 );
xor ( n239463 , n239451 , n239462 );
not ( n239464 , n237503 );
not ( n239465 , n239166 );
or ( n239466 , n239464 , n239465 );
not ( n239467 , n207938 );
not ( n239468 , n238719 );
and ( n239469 , n239467 , n239468 );
not ( n239470 , n220581 );
and ( n239471 , n239470 , n238719 );
nor ( n239472 , n239469 , n239471 );
not ( n239473 , n239472 );
nand ( n239474 , n239473 , n237493 );
nand ( n239475 , n239466 , n239474 );
xor ( n239476 , n239463 , n239475 );
xor ( n239477 , n239439 , n239476 );
xor ( n239478 , n239363 , n239367 );
and ( n239479 , n239478 , n239476 );
and ( n239480 , n239363 , n239367 );
or ( n239481 , n239479 , n239480 );
not ( n239482 , n237914 );
not ( n239483 , n234273 );
not ( n239484 , n40724 );
or ( n239485 , n239483 , n239484 );
not ( n239486 , n238671 );
nand ( n239487 , n239486 , n234878 );
nand ( n239488 , n239485 , n239487 );
not ( n239489 , n239488 );
or ( n239490 , n239482 , n239489 );
not ( n239491 , n238995 );
not ( n239492 , n235195 );
nand ( n239493 , n239491 , n239492 );
nand ( n239494 , n239490 , n239493 );
buf ( n239495 , n227782 );
not ( n239496 , n239495 );
not ( n239497 , n237130 );
not ( n239498 , n237948 );
or ( n239499 , n239497 , n239498 );
nand ( n239500 , n208046 , n224095 );
nand ( n239501 , n239499 , n239500 );
not ( n239502 , n239501 );
or ( n239503 , n239496 , n239502 );
nand ( n239504 , n239094 , n224087 );
nand ( n239505 , n239503 , n239504 );
xor ( n239506 , n239494 , n239505 );
not ( n239507 , n223665 );
not ( n239508 , n239507 );
not ( n239509 , n239508 );
not ( n239510 , n239132 );
or ( n239511 , n239509 , n239510 );
not ( n239512 , n221241 );
not ( n239513 , n234503 );
or ( n239514 , n239512 , n239513 );
not ( n239515 , n230490 );
nand ( n239516 , n239515 , n238363 );
nand ( n239517 , n239514 , n239516 );
nand ( n239518 , n239517 , n218843 );
nand ( n239519 , n239511 , n239518 );
xor ( n239520 , n239506 , n239519 );
not ( n239521 , n219435 );
not ( n239522 , n239141 );
or ( n239523 , n239521 , n239522 );
not ( n239524 , n219424 );
not ( n239525 , n237971 );
or ( n239526 , n239524 , n239525 );
not ( n239527 , n237971 );
nand ( n239528 , n239527 , n219440 );
nand ( n239529 , n239526 , n239528 );
buf ( n239530 , n219076 );
nand ( n239531 , n239529 , n239530 );
nand ( n239532 , n239523 , n239531 );
not ( n239533 , n220164 );
not ( n239534 , n239154 );
or ( n239535 , n239533 , n239534 );
not ( n239536 , n236768 );
not ( n239537 , n224700 );
or ( n239538 , n239536 , n239537 );
nand ( n239539 , n236300 , n222414 );
nand ( n239540 , n239538 , n239539 );
nand ( n239541 , n239540 , n219779 );
nand ( n239542 , n239535 , n239541 );
xor ( n239543 , n239532 , n239542 );
not ( n239544 , n221674 );
not ( n239545 , n222399 );
not ( n239546 , n233546 );
or ( n239547 , n239545 , n239546 );
not ( n239548 , n222399 );
nand ( n239549 , n238789 , n239548 );
nand ( n239550 , n239547 , n239549 );
not ( n239551 , n239550 );
or ( n239552 , n239544 , n239551 );
nand ( n239553 , n239068 , n235913 );
nand ( n239554 , n239552 , n239553 );
xor ( n239555 , n239543 , n239554 );
xor ( n239556 , n239520 , n239555 );
or ( n239557 , n239191 , n223825 );
or ( n239558 , n222323 , n223833 );
nand ( n239559 , n239557 , n239558 );
not ( n239560 , n226287 );
not ( n239561 , n226292 );
buf ( n239562 , n233362 );
not ( n239563 , n239562 );
or ( n239564 , n239561 , n239563 );
not ( n239565 , n227912 );
nand ( n239566 , n239565 , n238887 );
nand ( n239567 , n239564 , n239566 );
not ( n239568 , n239567 );
or ( n239569 , n239560 , n239568 );
nand ( n239570 , n220414 , n239232 );
nand ( n239571 , n239569 , n239570 );
xor ( n239572 , n239559 , n239571 );
xor ( n239573 , n239572 , n239013 );
xor ( n239574 , n239556 , n239573 );
xor ( n239575 , n239520 , n239555 );
and ( n239576 , n239575 , n239573 );
and ( n239577 , n239520 , n239555 );
or ( n239578 , n239576 , n239577 );
not ( n239579 , n231018 );
not ( n239580 , n239175 );
or ( n239581 , n239579 , n239580 );
not ( n239582 , n231500 );
not ( n239583 , n234347 );
or ( n239584 , n239582 , n239583 );
buf ( n239585 , n227223 );
nand ( n239586 , n239585 , n231501 );
nand ( n239587 , n239584 , n239586 );
nand ( n239588 , n239587 , n220067 );
nand ( n239589 , n239581 , n239588 );
xor ( n239590 , n239049 , n239589 );
xor ( n239591 , n239590 , n239319 );
not ( n239592 , n238409 );
not ( n239593 , n239114 );
or ( n239594 , n239592 , n239593 );
not ( n239595 , n237005 );
not ( n239596 , n219223 );
or ( n239597 , n239595 , n239596 );
not ( n239598 , n223156 );
not ( n239599 , n239598 );
nand ( n239600 , n219226 , n239599 );
nand ( n239601 , n239597 , n239600 );
nand ( n239602 , n239601 , n227294 );
nand ( n239603 , n239594 , n239602 );
not ( n239604 , n218232 );
not ( n239605 , n218205 );
not ( n239606 , n238728 );
or ( n239607 , n239605 , n239606 );
not ( n239608 , n227477 );
nand ( n239609 , n239608 , n234949 );
nand ( n239610 , n239607 , n239609 );
not ( n239611 , n239610 );
or ( n239612 , n239604 , n239611 );
nand ( n239613 , n239106 , n219461 );
nand ( n239614 , n239612 , n239613 );
xor ( n239615 , n239603 , n239614 );
not ( n239616 , n221933 );
not ( n239617 , n238835 );
and ( n239618 , n239617 , n226484 );
not ( n239619 , n239617 );
buf ( n239620 , n221938 );
and ( n239621 , n239619 , n239620 );
or ( n239622 , n239618 , n239621 );
not ( n239623 , n239622 );
or ( n239624 , n239616 , n239623 );
nand ( n239625 , n239208 , n219332 );
nand ( n239626 , n239624 , n239625 );
xor ( n239627 , n239615 , n239626 );
xor ( n239628 , n239591 , n239627 );
xor ( n239629 , n239628 , n239371 );
xor ( n239630 , n239591 , n239627 );
and ( n239631 , n239630 , n239371 );
and ( n239632 , n239591 , n239627 );
or ( n239633 , n239631 , n239632 );
not ( n239634 , n227260 );
not ( n239635 , n239241 );
or ( n239636 , n239634 , n239635 );
not ( n239637 , n226655 );
not ( n239638 , n39364 );
or ( n239639 , n239637 , n239638 );
nand ( n239640 , n237229 , n233053 );
nand ( n239641 , n239639 , n239640 );
nand ( n239642 , n239641 , n223949 );
nand ( n239643 , n239636 , n239642 );
not ( n239644 , n219501 );
not ( n239645 , n39089 );
not ( n239646 , n237203 );
and ( n239647 , n239645 , n239646 );
and ( n239648 , n238857 , n227599 );
nor ( n239649 , n239647 , n239648 );
not ( n239650 , n239649 );
not ( n239651 , n239650 );
or ( n239652 , n239644 , n239651 );
nand ( n239653 , n239250 , n225478 );
nand ( n239654 , n239652 , n239653 );
xor ( n239655 , n239643 , n239654 );
not ( n239656 , n234006 );
not ( n239657 , n239218 );
or ( n239658 , n239656 , n239657 );
not ( n239659 , n229261 );
not ( n239660 , n235516 );
or ( n239661 , n239659 , n239660 );
nand ( n239662 , n39747 , n234000 );
nand ( n239663 , n239661 , n239662 );
nand ( n239664 , n239663 , n229964 );
nand ( n239665 , n239658 , n239664 );
xor ( n239666 , n239655 , n239665 );
xor ( n239667 , n239666 , n239055 );
xor ( n239668 , n239428 , n239400 );
xor ( n239669 , n239668 , n239355 );
xor ( n239670 , n239667 , n239669 );
xor ( n239671 , n239666 , n239055 );
and ( n239672 , n239671 , n239669 );
and ( n239673 , n239666 , n239055 );
or ( n239674 , n239672 , n239673 );
xor ( n239675 , n239124 , n239061 );
xor ( n239676 , n239675 , n239434 );
xor ( n239677 , n239124 , n239061 );
and ( n239678 , n239677 , n239434 );
and ( n239679 , n239124 , n239061 );
or ( n239680 , n239678 , n239679 );
xor ( n239681 , n239260 , n239574 );
xor ( n239682 , n239681 , n239477 );
xor ( n239683 , n239260 , n239574 );
and ( n239684 , n239683 , n239477 );
and ( n239685 , n239260 , n239574 );
or ( n239686 , n239684 , n239685 );
xor ( n239687 , n239200 , n239629 );
xor ( n239688 , n239687 , n239291 );
xor ( n239689 , n239200 , n239629 );
and ( n239690 , n239689 , n239291 );
and ( n239691 , n239200 , n239629 );
or ( n239692 , n239690 , n239691 );
xor ( n239693 , n239670 , n239297 );
xor ( n239694 , n239693 , n239676 );
xor ( n239695 , n239670 , n239297 );
and ( n239696 , n239695 , n239676 );
and ( n239697 , n239670 , n239297 );
or ( n239698 , n239696 , n239697 );
xor ( n239699 , n239303 , n239682 );
xor ( n239700 , n239699 , n239309 );
xor ( n239701 , n239303 , n239682 );
and ( n239702 , n239701 , n239309 );
and ( n239703 , n239303 , n239682 );
or ( n239704 , n239702 , n239703 );
xor ( n239705 , n239494 , n239505 );
and ( n239706 , n239705 , n239519 );
and ( n239707 , n239494 , n239505 );
or ( n239708 , n239706 , n239707 );
xor ( n239709 , n239688 , n239315 );
xor ( n239710 , n239709 , n239694 );
xor ( n239711 , n239688 , n239315 );
and ( n239712 , n239711 , n239694 );
and ( n239713 , n239688 , n239315 );
or ( n239714 , n239712 , n239713 );
xor ( n239715 , n239700 , n239325 );
xor ( n239716 , n239715 , n239710 );
xor ( n239717 , n239700 , n239325 );
and ( n239718 , n239717 , n239710 );
and ( n239719 , n239700 , n239325 );
or ( n239720 , n239718 , n239719 );
xor ( n239721 , n239331 , n239716 );
xor ( n239722 , n239721 , n239337 );
xor ( n239723 , n239331 , n239716 );
and ( n239724 , n239723 , n239337 );
and ( n239725 , n239331 , n239716 );
or ( n239726 , n239724 , n239725 );
xor ( n239727 , n239532 , n239542 );
and ( n239728 , n239727 , n239554 );
and ( n239729 , n239532 , n239542 );
or ( n239730 , n239728 , n239729 );
xor ( n239731 , n239451 , n239462 );
and ( n239732 , n239731 , n239475 );
and ( n239733 , n239451 , n239462 );
or ( n239734 , n239732 , n239733 );
xor ( n239735 , n239603 , n239614 );
and ( n239736 , n239735 , n239626 );
and ( n239737 , n239603 , n239614 );
or ( n239738 , n239736 , n239737 );
xor ( n239739 , n239643 , n239654 );
and ( n239740 , n239739 , n239665 );
and ( n239741 , n239643 , n239654 );
or ( n239742 , n239740 , n239741 );
xor ( n239743 , n239559 , n239571 );
and ( n239744 , n239743 , n239013 );
and ( n239745 , n239559 , n239571 );
or ( n239746 , n239744 , n239745 );
xor ( n239747 , n239049 , n239589 );
and ( n239748 , n239747 , n239319 );
and ( n239749 , n239049 , n239589 );
or ( n239750 , n239748 , n239749 );
xor ( n239751 , n239428 , n239400 );
and ( n239752 , n239751 , n239355 );
and ( n239753 , n239428 , n239400 );
or ( n239754 , n239752 , n239753 );
or ( n239755 , n216204 , n219314 );
nand ( n239756 , n239755 , n219687 );
not ( n239757 , n239423 );
not ( n239758 , n232956 );
or ( n239759 , n239757 , n239758 );
not ( n239760 , n232493 );
not ( n239761 , n41165 );
or ( n239762 , n239760 , n239761 );
not ( n239763 , n219389 );
nand ( n239764 , n239763 , n229806 );
nand ( n239765 , n239762 , n239764 );
nand ( n239766 , n238776 , n239765 );
nand ( n239767 , n239759 , n239766 );
xor ( n239768 , n239756 , n239767 );
not ( n239769 , n237797 );
not ( n239770 , n239448 );
or ( n239771 , n239769 , n239770 );
and ( n239772 , n239001 , n234293 );
not ( n239773 , n239001 );
not ( n239774 , n238230 );
and ( n239775 , n239773 , n239774 );
nor ( n239776 , n239772 , n239775 );
or ( n239777 , n234896 , n239776 );
nand ( n239778 , n239771 , n239777 );
xor ( n239779 , n239768 , n239778 );
xor ( n239780 , n239756 , n239767 );
and ( n239781 , n239780 , n239778 );
and ( n239782 , n239756 , n239767 );
or ( n239783 , n239781 , n239782 );
not ( n239784 , n237810 );
not ( n239785 , n239379 );
or ( n239786 , n239784 , n239785 );
not ( n239787 , n233450 );
and ( n239788 , n239787 , n41250 );
and ( n239789 , n233450 , n217697 );
nor ( n239790 , n239788 , n239789 );
or ( n239791 , n228273 , n239790 );
nand ( n239792 , n239786 , n239791 );
not ( n239793 , n239388 );
not ( n239794 , n237038 );
not ( n239795 , n239794 );
or ( n239796 , n239793 , n239795 );
not ( n239797 , n234751 );
not ( n239798 , n228847 );
or ( n239799 , n239797 , n239798 );
nand ( n239800 , n228726 , n216500 );
nand ( n239801 , n239799 , n239800 );
nand ( n239802 , n228868 , n239801 );
nand ( n239803 , n239796 , n239802 );
xor ( n239804 , n239792 , n239803 );
buf ( n239805 , n231474 );
or ( n239806 , n239805 , n239397 );
not ( n239807 , n215616 );
not ( n239808 , n237014 );
or ( n239809 , n239807 , n239808 );
nand ( n239810 , n231480 , n236580 );
nand ( n239811 , n239809 , n239810 );
not ( n239812 , n239811 );
or ( n239813 , n231476 , n239812 );
nand ( n239814 , n239806 , n239813 );
xor ( n239815 , n239804 , n239814 );
xor ( n239816 , n239792 , n239803 );
and ( n239817 , n239816 , n239814 );
and ( n239818 , n239792 , n239803 );
or ( n239819 , n239817 , n239818 );
xor ( n239820 , n239708 , n239730 );
xor ( n239821 , n239820 , n239734 );
xor ( n239822 , n239708 , n239730 );
and ( n239823 , n239822 , n239734 );
and ( n239824 , n239708 , n239730 );
or ( n239825 , n239823 , n239824 );
xor ( n239826 , n239742 , n239746 );
xor ( n239827 , n239826 , n239750 );
xor ( n239828 , n239742 , n239746 );
and ( n239829 , n239828 , n239750 );
and ( n239830 , n239742 , n239746 );
or ( n239831 , n239829 , n239830 );
not ( n239832 , n220164 );
not ( n239833 , n239540 );
or ( n239834 , n239832 , n239833 );
not ( n239835 , n236768 );
not ( n239836 , n227004 );
or ( n239837 , n239835 , n239836 );
nand ( n239838 , n238362 , n222414 );
nand ( n239839 , n239837 , n239838 );
nand ( n239840 , n239839 , n219779 );
nand ( n239841 , n239834 , n239840 );
not ( n239842 , n221674 );
and ( n239843 , n220906 , n221712 );
not ( n239844 , n220906 );
and ( n239845 , n239844 , n236719 );
or ( n239846 , n239843 , n239845 );
not ( n239847 , n239846 );
or ( n239848 , n239842 , n239847 );
nand ( n239849 , n239550 , n235913 );
nand ( n239850 , n239848 , n239849 );
xor ( n239851 , n239841 , n239850 );
not ( n239852 , n221637 );
not ( n239853 , n222035 );
not ( n239854 , n226911 );
not ( n239855 , n239854 );
or ( n239856 , n239853 , n239855 );
nand ( n239857 , n40259 , n221612 );
nand ( n239858 , n239856 , n239857 );
not ( n239859 , n239858 );
or ( n239860 , n239852 , n239859 );
not ( n239861 , n222471 );
nand ( n239862 , n239861 , n239460 );
nand ( n239863 , n239860 , n239862 );
xor ( n239864 , n239851 , n239863 );
or ( n239865 , n239472 , n235644 );
not ( n239866 , n222430 );
not ( n239867 , n226921 );
or ( n239868 , n239866 , n239867 );
nand ( n239869 , n239080 , n238719 );
nand ( n239870 , n239868 , n239869 );
not ( n239871 , n239870 );
not ( n239872 , n237493 );
or ( n239873 , n239871 , n239872 );
nand ( n239874 , n239865 , n239873 );
xor ( n239875 , n239450 , n239874 );
not ( n239876 , n227294 );
not ( n239877 , n238681 );
not ( n239878 , n234108 );
or ( n239879 , n239877 , n239878 );
nand ( n239880 , n40625 , n238404 );
nand ( n239881 , n239879 , n239880 );
not ( n239882 , n239881 );
or ( n239883 , n239876 , n239882 );
nand ( n239884 , n239601 , n238409 );
nand ( n239885 , n239883 , n239884 );
xor ( n239886 , n239875 , n239885 );
xor ( n239887 , n239864 , n239886 );
not ( n239888 , n223665 );
not ( n239889 , n239517 );
or ( n239890 , n239888 , n239889 );
not ( n239891 , n221241 );
not ( n239892 , n226961 );
or ( n239893 , n239891 , n239892 );
nand ( n239894 , n39997 , n238363 );
nand ( n239895 , n239893 , n239894 );
nand ( n239896 , n239895 , n218843 );
nand ( n239897 , n239890 , n239896 );
not ( n239898 , n239495 );
not ( n239899 , n238672 );
not ( n239900 , n239899 );
not ( n239901 , n218912 );
or ( n239902 , n239900 , n239901 );
buf ( n239903 , n237129 );
nand ( n239904 , n236752 , n239903 );
nand ( n239905 , n239902 , n239904 );
not ( n239906 , n239905 );
or ( n239907 , n239898 , n239906 );
nand ( n239908 , n239501 , n224087 );
nand ( n239909 , n239907 , n239908 );
xor ( n239910 , n239897 , n239909 );
not ( n239911 , n220507 );
not ( n239912 , n239529 );
or ( n239913 , n239911 , n239912 );
and ( n239914 , n219797 , n237600 );
not ( n239915 , n219797 );
not ( n239916 , n40547 );
not ( n239917 , n239916 );
and ( n239918 , n239915 , n239917 );
or ( n239919 , n239914 , n239918 );
not ( n239920 , n239919 );
nand ( n239921 , n239920 , n239530 );
nand ( n239922 , n239913 , n239921 );
xor ( n239923 , n239910 , n239922 );
xor ( n239924 , n239887 , n239923 );
xor ( n239925 , n239864 , n239886 );
and ( n239926 , n239925 , n239923 );
and ( n239927 , n239864 , n239886 );
or ( n239928 , n239926 , n239927 );
or ( n239929 , n239649 , n225477 );
and ( n239930 , n233544 , n235962 );
not ( n239931 , n233544 );
not ( n239932 , n229704 );
and ( n239933 , n239931 , n239932 );
nor ( n239934 , n239930 , n239933 );
or ( n239935 , n239934 , n227121 );
nand ( n239936 , n239929 , n239935 );
not ( n239937 , n239663 );
not ( n239938 , n234006 );
or ( n239939 , n239937 , n239938 );
not ( n239940 , n229261 );
not ( n239941 , n226709 );
or ( n239942 , n239940 , n239941 );
nand ( n239943 , n235977 , n229262 );
nand ( n239944 , n239942 , n239943 );
not ( n239945 , n239944 );
not ( n239946 , n229964 );
or ( n239947 , n239945 , n239946 );
nand ( n239948 , n239939 , n239947 );
xor ( n239949 , n239936 , n239948 );
not ( n239950 , n239567 );
or ( n239951 , n239950 , n226942 );
buf ( n239952 , n209709 );
and ( n239953 , n227912 , n239952 );
not ( n239954 , n227912 );
and ( n239955 , n239954 , n235691 );
nor ( n239956 , n239953 , n239955 );
or ( n239957 , n239956 , n226940 );
nand ( n239958 , n239951 , n239957 );
xor ( n239959 , n239949 , n239958 );
xor ( n239960 , n239738 , n239959 );
xor ( n239961 , n239404 , n239432 );
not ( n239962 , n239587 );
or ( n239963 , n239962 , n227130 );
not ( n239964 , n233856 );
not ( n239965 , n231501 );
and ( n239966 , n239964 , n239965 );
and ( n239967 , n39714 , n234015 );
nor ( n239968 , n239966 , n239967 );
or ( n239969 , n239968 , n227138 );
nand ( n239970 , n239963 , n239969 );
xor ( n239971 , n239961 , n239970 );
xor ( n239972 , n239960 , n239971 );
xor ( n239973 , n239738 , n239959 );
and ( n239974 , n239973 , n239971 );
and ( n239975 , n239738 , n239959 );
or ( n239976 , n239974 , n239975 );
not ( n239977 , n219461 );
not ( n239978 , n239610 );
or ( n239979 , n239977 , n239978 );
not ( n239980 , n218775 );
not ( n239981 , n226724 );
or ( n239982 , n239980 , n239981 );
nand ( n239983 , n238323 , n234949 );
nand ( n239984 , n239982 , n239983 );
nand ( n239985 , n239984 , n218232 );
nand ( n239986 , n239979 , n239985 );
not ( n239987 , n219332 );
not ( n239988 , n239622 );
or ( n239989 , n239987 , n239988 );
not ( n239990 , n226484 );
not ( n239991 , n239186 );
or ( n239992 , n239990 , n239991 );
nand ( n239993 , n239185 , n221938 );
nand ( n239994 , n239992 , n239993 );
nand ( n239995 , n239994 , n221933 );
nand ( n239996 , n239989 , n239995 );
xor ( n239997 , n239986 , n239996 );
not ( n239998 , n223949 );
not ( n239999 , n226655 );
not ( n240000 , n238486 );
or ( n240001 , n239999 , n240000 );
nand ( n240002 , n236840 , n227927 );
nand ( n240003 , n240001 , n240002 );
not ( n240004 , n240003 );
or ( n240005 , n239998 , n240004 );
nand ( n240006 , n239641 , n227260 );
nand ( n240007 , n240005 , n240006 );
xor ( n240008 , n239997 , n240007 );
xor ( n240009 , n240008 , n239754 );
xor ( n240010 , n239815 , n239779 );
not ( n240011 , n239412 );
or ( n240012 , n230721 , n240011 );
xor ( n240013 , n225769 , n233885 );
not ( n240014 , n232402 );
or ( n240015 , n240013 , n240014 );
nand ( n240016 , n240012 , n240015 );
not ( n240017 , n231754 );
nor ( n240018 , n240017 , n226698 );
xor ( n240019 , n240016 , n240018 );
not ( n240020 , n236958 );
not ( n240021 , n240020 );
not ( n240022 , n219599 );
not ( n240023 , n237918 );
and ( n240024 , n240022 , n240023 );
and ( n240025 , n219599 , n237918 );
nor ( n240026 , n240024 , n240025 );
not ( n240027 , n240026 );
not ( n240028 , n240027 );
or ( n240029 , n240021 , n240028 );
nand ( n240030 , n239488 , n239492 );
nand ( n240031 , n240029 , n240030 );
xor ( n240032 , n240019 , n240031 );
xor ( n240033 , n240010 , n240032 );
xor ( n240034 , n240009 , n240033 );
xor ( n240035 , n240008 , n239754 );
and ( n240036 , n240035 , n240033 );
and ( n240037 , n240008 , n239754 );
or ( n240038 , n240036 , n240037 );
xor ( n240039 , n239438 , n239821 );
xor ( n240040 , n240039 , n239481 );
xor ( n240041 , n239438 , n239821 );
and ( n240042 , n240041 , n239481 );
and ( n240043 , n239438 , n239821 );
or ( n240044 , n240042 , n240043 );
xor ( n240045 , n239827 , n239924 );
xor ( n240046 , n240045 , n239633 );
xor ( n240047 , n239827 , n239924 );
and ( n240048 , n240047 , n239633 );
and ( n240049 , n239827 , n239924 );
or ( n240050 , n240048 , n240049 );
xor ( n240051 , n239578 , n239674 );
xor ( n240052 , n240051 , n239972 );
xor ( n240053 , n239578 , n239674 );
and ( n240054 , n240053 , n239972 );
and ( n240055 , n239578 , n239674 );
or ( n240056 , n240054 , n240055 );
xor ( n240057 , n239680 , n240034 );
xor ( n240058 , n240057 , n240040 );
xor ( n240059 , n239680 , n240034 );
and ( n240060 , n240059 , n240040 );
and ( n240061 , n239680 , n240034 );
or ( n240062 , n240060 , n240061 );
xor ( n240063 , n239686 , n240046 );
xor ( n240064 , n240063 , n240052 );
xor ( n240065 , n239686 , n240046 );
and ( n240066 , n240065 , n240052 );
and ( n240067 , n239686 , n240046 );
or ( n240068 , n240066 , n240067 );
xor ( n240069 , n240016 , n240018 );
and ( n240070 , n240069 , n240031 );
and ( n240071 , n240016 , n240018 );
or ( n240072 , n240070 , n240071 );
xor ( n240073 , n239692 , n239698 );
xor ( n240074 , n240073 , n240058 );
xor ( n240075 , n239692 , n239698 );
and ( n240076 , n240075 , n240058 );
and ( n240077 , n239692 , n239698 );
or ( n240078 , n240076 , n240077 );
xor ( n240079 , n240064 , n239704 );
xor ( n240080 , n240079 , n239714 );
xor ( n240081 , n240064 , n239704 );
and ( n240082 , n240081 , n239714 );
and ( n240083 , n240064 , n239704 );
or ( n240084 , n240082 , n240083 );
xor ( n240085 , n240074 , n240080 );
xor ( n240086 , n240085 , n239720 );
xor ( n240087 , n240074 , n240080 );
and ( n240088 , n240087 , n239720 );
and ( n240089 , n240074 , n240080 );
or ( n240090 , n240088 , n240089 );
xor ( n240091 , n239897 , n239909 );
and ( n240092 , n240091 , n239922 );
and ( n240093 , n239897 , n239909 );
or ( n240094 , n240092 , n240093 );
xor ( n240095 , n239841 , n239850 );
and ( n240096 , n240095 , n239863 );
and ( n240097 , n239841 , n239850 );
or ( n240098 , n240096 , n240097 );
xor ( n240099 , n239450 , n239874 );
and ( n240100 , n240099 , n239885 );
and ( n240101 , n239450 , n239874 );
or ( n240102 , n240100 , n240101 );
xor ( n240103 , n239986 , n239996 );
and ( n240104 , n240103 , n240007 );
and ( n240105 , n239986 , n239996 );
or ( n240106 , n240104 , n240105 );
xor ( n240107 , n239936 , n239948 );
and ( n240108 , n240107 , n239958 );
and ( n240109 , n239936 , n239948 );
or ( n240110 , n240108 , n240109 );
xor ( n240111 , n239404 , n239432 );
and ( n240112 , n240111 , n239970 );
and ( n240113 , n239404 , n239432 );
or ( n240114 , n240112 , n240113 );
xor ( n240115 , n239815 , n239779 );
and ( n240116 , n240115 , n240032 );
and ( n240117 , n239815 , n239779 );
or ( n240118 , n240116 , n240117 );
not ( n240119 , n239801 );
not ( n240120 , n237038 );
not ( n240121 , n240120 );
or ( n240122 , n240119 , n240121 );
not ( n240123 , n228850 );
not ( n240124 , n216307 );
or ( n240125 , n240123 , n240124 );
not ( n240126 , n233925 );
nand ( n240127 , n240126 , n41319 );
nand ( n240128 , n240125 , n240127 );
nand ( n240129 , n228868 , n240128 );
nand ( n240130 , n240122 , n240129 );
not ( n240131 , n239811 );
not ( n240132 , n234371 );
or ( n240133 , n240131 , n240132 );
not ( n240134 , n215796 );
not ( n240135 , n237014 );
or ( n240136 , n240134 , n240135 );
nand ( n240137 , n237017 , n216261 );
nand ( n240138 , n240136 , n240137 );
nand ( n240139 , n234378 , n240138 );
nand ( n240140 , n240133 , n240139 );
xor ( n240141 , n240130 , n240140 );
or ( n240142 , n239269 , n240013 );
not ( n240143 , n231754 );
not ( n240144 , n234256 );
and ( n240145 , n240143 , n240144 );
and ( n240146 , n231232 , n234256 );
nor ( n240147 , n240145 , n240146 );
not ( n240148 , n238274 );
or ( n240149 , n240147 , n240148 );
nand ( n240150 , n240142 , n240149 );
xor ( n240151 , n240141 , n240150 );
xor ( n240152 , n240130 , n240140 );
and ( n240153 , n240152 , n240150 );
and ( n240154 , n240130 , n240140 );
or ( n240155 , n240153 , n240154 );
buf ( n240156 , n232784 );
and ( n240157 , n240156 , n209437 );
not ( n240158 , n227852 );
not ( n240159 , n222984 );
not ( n240160 , n239774 );
or ( n240161 , n240159 , n240160 );
or ( n240162 , n229823 , n217330 );
nand ( n240163 , n240161 , n240162 );
not ( n240164 , n240163 );
or ( n240165 , n240158 , n240164 );
not ( n240166 , n239776 );
nand ( n240167 , n240166 , n237797 );
nand ( n240168 , n240165 , n240167 );
xor ( n240169 , n240157 , n240168 );
not ( n240170 , n238776 );
not ( n240171 , n232493 );
not ( n240172 , n238671 );
or ( n240173 , n240171 , n240172 );
or ( n240174 , n238671 , n232497 );
nand ( n240175 , n240173 , n240174 );
not ( n240176 , n240175 );
or ( n240177 , n240170 , n240176 );
nand ( n240178 , n232956 , n239765 );
nand ( n240179 , n240177 , n240178 );
xor ( n240180 , n240169 , n240179 );
xor ( n240181 , n240157 , n240168 );
and ( n240182 , n240181 , n240179 );
and ( n240183 , n240157 , n240168 );
or ( n240184 , n240182 , n240183 );
xor ( n240185 , n240102 , n240110 );
xor ( n240186 , n240185 , n240114 );
xor ( n240187 , n240102 , n240110 );
and ( n240188 , n240187 , n240114 );
and ( n240189 , n240102 , n240110 );
or ( n240190 , n240188 , n240189 );
not ( n240191 , n235913 );
not ( n240192 , n239846 );
or ( n240193 , n240191 , n240192 );
not ( n240194 , n220906 );
not ( n240195 , n236301 );
or ( n240196 , n240194 , n240195 );
nand ( n240197 , n236304 , n239548 );
nand ( n240198 , n240196 , n240197 );
nand ( n240199 , n240198 , n220930 );
nand ( n240200 , n240193 , n240199 );
not ( n240201 , n239790 );
not ( n240202 , n240201 );
not ( n240203 , n237810 );
or ( n240204 , n240202 , n240203 );
not ( n240205 , n233450 );
not ( n240206 , n40888 );
and ( n240207 , n240205 , n240206 );
and ( n240208 , n233450 , n40888 );
nor ( n240209 , n240207 , n240208 );
not ( n240210 , n240209 );
nand ( n240211 , n240210 , n238240 );
nand ( n240212 , n240204 , n240211 );
not ( n240213 , n240212 );
xor ( n240214 , n240200 , n240213 );
not ( n240215 , n239452 );
not ( n240216 , n239858 );
or ( n240217 , n240215 , n240216 );
not ( n240218 , n40397 );
not ( n240219 , n221612 );
or ( n240220 , n240218 , n240219 );
nand ( n240221 , n222121 , n222035 );
nand ( n240222 , n240220 , n240221 );
nand ( n240223 , n240222 , n221637 );
nand ( n240224 , n240217 , n240223 );
xor ( n240225 , n240214 , n240224 );
not ( n240226 , n237503 );
not ( n240227 , n239870 );
or ( n240228 , n240226 , n240227 );
buf ( n240229 , n222892 );
not ( n240230 , n240229 );
not ( n240231 , n220599 );
or ( n240232 , n240230 , n240231 );
not ( n240233 , n222892 );
nand ( n240234 , n240233 , n221956 );
nand ( n240235 , n240232 , n240234 );
nand ( n240236 , n240235 , n237493 );
nand ( n240237 , n240228 , n240236 );
not ( n240238 , n235172 );
not ( n240239 , n239881 );
or ( n240240 , n240238 , n240239 );
not ( n240241 , n239598 );
not ( n240242 , n40660 );
or ( n240243 , n240241 , n240242 );
nand ( n240244 , n235359 , n223156 );
nand ( n240245 , n240243 , n240244 );
nand ( n240246 , n240245 , n227294 );
nand ( n240247 , n240240 , n240246 );
xor ( n240248 , n240237 , n240247 );
not ( n240249 , n224087 );
not ( n240250 , n239905 );
or ( n240251 , n240249 , n240250 );
not ( n240252 , n237130 );
not ( n240253 , n40561 );
or ( n240254 , n240252 , n240253 );
not ( n240255 , n40560 );
nand ( n240256 , n240255 , n224095 );
nand ( n240257 , n240254 , n240256 );
nand ( n240258 , n240257 , n239495 );
nand ( n240259 , n240251 , n240258 );
xor ( n240260 , n240248 , n240259 );
xor ( n240261 , n240225 , n240260 );
not ( n240262 , n234878 );
not ( n240263 , n237948 );
or ( n240264 , n240262 , n240263 );
not ( n240265 , n40766 );
nand ( n240266 , n240265 , n235200 );
nand ( n240267 , n240264 , n240266 );
not ( n240268 , n240267 );
not ( n240269 , n237914 );
or ( n240270 , n240268 , n240269 );
buf ( n240271 , n227792 );
not ( n240272 , n240271 );
or ( n240273 , n240026 , n240272 );
nand ( n240274 , n240270 , n240273 );
or ( n240275 , n239919 , n219434 );
not ( n240276 , n223765 );
not ( n240277 , n219797 );
and ( n240278 , n240276 , n240277 );
not ( n240279 , n234503 );
and ( n240280 , n240279 , n219423 );
nor ( n240281 , n240278 , n240280 );
or ( n240282 , n240281 , n229612 );
nand ( n240283 , n240275 , n240282 );
xor ( n240284 , n240274 , n240283 );
not ( n240285 , n239839 );
or ( n240286 , n240285 , n237895 );
not ( n240287 , n236768 );
not ( n240288 , n222940 );
or ( n240289 , n240287 , n240288 );
not ( n240290 , n220151 );
nand ( n240291 , n240290 , n239527 );
nand ( n240292 , n240289 , n240291 );
not ( n240293 , n240292 );
or ( n240294 , n240293 , n224171 );
nand ( n240295 , n240286 , n240294 );
xor ( n240296 , n240284 , n240295 );
xor ( n240297 , n240261 , n240296 );
xor ( n240298 , n240225 , n240260 );
and ( n240299 , n240298 , n240296 );
and ( n240300 , n240225 , n240260 );
or ( n240301 , n240299 , n240300 );
not ( n240302 , n227260 );
not ( n240303 , n240003 );
or ( n240304 , n240302 , n240303 );
not ( n240305 , n226655 );
not ( n240306 , n237271 );
or ( n240307 , n240305 , n240306 );
not ( n240308 , n239562 );
nand ( n240309 , n240308 , n233053 );
nand ( n240310 , n240307 , n240309 );
nand ( n240311 , n240310 , n223949 );
nand ( n240312 , n240304 , n240311 );
xor ( n240313 , n239783 , n240312 );
xor ( n240314 , n240313 , n239819 );
xor ( n240315 , n240106 , n240314 );
not ( n240316 , n229964 );
not ( n240317 , n229261 );
not ( n240318 , n236382 );
or ( n240319 , n240317 , n240318 );
nand ( n240320 , n238857 , n234000 );
nand ( n240321 , n240319 , n240320 );
not ( n240322 , n240321 );
or ( n240323 , n240316 , n240322 );
nand ( n240324 , n239944 , n234006 );
nand ( n240325 , n240323 , n240324 );
not ( n240326 , n219332 );
not ( n240327 , n239994 );
or ( n240328 , n240326 , n240327 );
nand ( n240329 , n221933 , n226484 );
nand ( n240330 , n240328 , n240329 );
xor ( n240331 , n240325 , n240330 );
or ( n240332 , n239968 , n227130 );
and ( n240333 , n231501 , n235516 );
not ( n240334 , n231501 );
and ( n240335 , n240334 , n39747 );
or ( n240336 , n240333 , n240335 );
or ( n240337 , n240336 , n227138 );
nand ( n240338 , n240332 , n240337 );
xor ( n240339 , n240331 , n240338 );
xor ( n240340 , n240315 , n240339 );
xor ( n240341 , n240106 , n240314 );
and ( n240342 , n240341 , n240339 );
and ( n240343 , n240106 , n240314 );
or ( n240344 , n240342 , n240343 );
not ( n240345 , n218843 );
not ( n240346 , n221241 );
not ( n240347 , n227477 );
or ( n240348 , n240346 , n240347 );
nand ( n240349 , n39880 , n238363 );
nand ( n240350 , n240348 , n240349 );
not ( n240351 , n240350 );
or ( n240352 , n240345 , n240351 );
nand ( n240353 , n239895 , n239508 );
nand ( n240354 , n240352 , n240353 );
not ( n240355 , n226287 );
and ( n240356 , n229887 , n234579 );
not ( n240357 , n229887 );
not ( n240358 , n233611 );
and ( n240359 , n240357 , n240358 );
or ( n240360 , n240356 , n240359 );
not ( n240361 , n240360 );
not ( n240362 , n240361 );
or ( n240363 , n240355 , n240362 );
not ( n240364 , n239956 );
nand ( n240365 , n240364 , n226943 );
nand ( n240366 , n240363 , n240365 );
xor ( n240367 , n240354 , n240366 );
not ( n240368 , n229395 );
not ( n240369 , n239934 );
not ( n240370 , n240369 );
or ( n240371 , n240368 , n240370 );
buf ( n240372 , n230270 );
and ( n240373 , n237203 , n240372 );
not ( n240374 , n237203 );
not ( n240375 , n240372 );
and ( n240376 , n240374 , n240375 );
or ( n240377 , n240373 , n240376 );
not ( n240378 , n240377 );
nand ( n240379 , n240378 , n219501 );
nand ( n240380 , n240371 , n240379 );
xor ( n240381 , n240367 , n240380 );
xor ( n240382 , n240381 , n240118 );
xor ( n240383 , n240382 , n239825 );
xor ( n240384 , n240381 , n240118 );
and ( n240385 , n240384 , n239825 );
and ( n240386 , n240381 , n240118 );
or ( n240387 , n240385 , n240386 );
not ( n240388 , n219461 );
not ( n240389 , n239984 );
or ( n240390 , n240388 , n240389 );
not ( n240391 , n224497 );
not ( n240392 , n234350 );
or ( n240393 , n240391 , n240392 );
nand ( n240394 , n238819 , n238352 );
nand ( n240395 , n240393 , n240394 );
nand ( n240396 , n240395 , n218232 );
nand ( n240397 , n240390 , n240396 );
xor ( n240398 , n240397 , n240180 );
xor ( n240399 , n240398 , n240151 );
xor ( n240400 , n240399 , n239831 );
xor ( n240401 , n240400 , n239928 );
xor ( n240402 , n240399 , n239831 );
and ( n240403 , n240402 , n239928 );
and ( n240404 , n240399 , n239831 );
or ( n240405 , n240403 , n240404 );
xor ( n240406 , n240072 , n240094 );
xor ( n240407 , n240406 , n240098 );
xor ( n240408 , n240407 , n240297 );
xor ( n240409 , n240408 , n240186 );
xor ( n240410 , n240407 , n240297 );
and ( n240411 , n240410 , n240186 );
and ( n240412 , n240407 , n240297 );
or ( n240413 , n240411 , n240412 );
xor ( n240414 , n239976 , n240038 );
xor ( n240415 , n240414 , n240340 );
xor ( n240416 , n239976 , n240038 );
and ( n240417 , n240416 , n240340 );
and ( n240418 , n239976 , n240038 );
or ( n240419 , n240417 , n240418 );
xor ( n240420 , n240044 , n240383 );
xor ( n240421 , n240420 , n240401 );
xor ( n240422 , n240044 , n240383 );
and ( n240423 , n240422 , n240401 );
and ( n240424 , n240044 , n240383 );
or ( n240425 , n240423 , n240424 );
xor ( n240426 , n240050 , n240056 );
xor ( n240427 , n240426 , n240409 );
xor ( n240428 , n240050 , n240056 );
and ( n240429 , n240428 , n240409 );
and ( n240430 , n240050 , n240056 );
or ( n240431 , n240429 , n240430 );
xor ( n240432 , n240415 , n240421 );
xor ( n240433 , n240432 , n240062 );
xor ( n240434 , n240415 , n240421 );
and ( n240435 , n240434 , n240062 );
and ( n240436 , n240415 , n240421 );
or ( n240437 , n240435 , n240436 );
xor ( n240438 , n240274 , n240283 );
and ( n240439 , n240438 , n240295 );
and ( n240440 , n240274 , n240283 );
or ( n240441 , n240439 , n240440 );
xor ( n240442 , n240427 , n240068 );
xor ( n240443 , n240442 , n240078 );
xor ( n240444 , n240427 , n240068 );
and ( n240445 , n240444 , n240078 );
and ( n240446 , n240427 , n240068 );
or ( n240447 , n240445 , n240446 );
xor ( n240448 , n240433 , n240443 );
xor ( n240449 , n240448 , n240084 );
xor ( n240450 , n240433 , n240443 );
and ( n240451 , n240450 , n240084 );
and ( n240452 , n240433 , n240443 );
or ( n240453 , n240451 , n240452 );
xor ( n240454 , n240200 , n240213 );
and ( n240455 , n240454 , n240224 );
and ( n240456 , n240200 , n240213 );
or ( n240457 , n240455 , n240456 );
xor ( n240458 , n240237 , n240247 );
and ( n240459 , n240458 , n240259 );
and ( n240460 , n240237 , n240247 );
or ( n240461 , n240459 , n240460 );
xor ( n240462 , n240354 , n240366 );
and ( n240463 , n240462 , n240380 );
and ( n240464 , n240354 , n240366 );
or ( n240465 , n240463 , n240464 );
xor ( n240466 , n240325 , n240330 );
and ( n240467 , n240466 , n240338 );
and ( n240468 , n240325 , n240330 );
or ( n240469 , n240467 , n240468 );
xor ( n240470 , n239783 , n240312 );
and ( n240471 , n240470 , n239819 );
and ( n240472 , n239783 , n240312 );
or ( n240473 , n240471 , n240472 );
xor ( n240474 , n240397 , n240180 );
and ( n240475 , n240474 , n240151 );
and ( n240476 , n240397 , n240180 );
or ( n240477 , n240475 , n240476 );
xor ( n240478 , n240072 , n240094 );
and ( n240479 , n240478 , n240098 );
and ( n240480 , n240072 , n240094 );
or ( n240481 , n240479 , n240480 );
not ( n240482 , n221932 );
not ( n240483 , n234045 );
or ( n240484 , n240482 , n240483 );
nand ( n240485 , n240484 , n226484 );
not ( n240486 , n240163 );
not ( n240487 , n238225 );
or ( n240488 , n240486 , n240487 );
not ( n240489 , n226650 );
not ( n240490 , n238199 );
or ( n240491 , n240489 , n240490 );
not ( n240492 , n219389 );
nand ( n240493 , n240492 , n229823 );
nand ( n240494 , n240491 , n240493 );
nand ( n240495 , n226885 , n240494 );
nand ( n240496 , n240488 , n240495 );
xor ( n240497 , n240485 , n240496 );
or ( n240498 , n228270 , n240209 );
not ( n240499 , n238240 );
not ( n240500 , n237816 );
and ( n240501 , n239001 , n240500 );
not ( n240502 , n239001 );
and ( n240503 , n240502 , n237816 );
nor ( n240504 , n240501 , n240503 );
or ( n240505 , n240499 , n240504 );
nand ( n240506 , n240498 , n240505 );
xor ( n240507 , n240497 , n240506 );
xor ( n240508 , n240485 , n240496 );
and ( n240509 , n240508 , n240506 );
and ( n240510 , n240485 , n240496 );
or ( n240511 , n240509 , n240510 );
not ( n240512 , n240128 );
not ( n240513 , n228860 );
or ( n240514 , n240512 , n240513 );
not ( n240515 , n221016 );
not ( n240516 , n228727 );
or ( n240517 , n240515 , n240516 );
nand ( n240518 , n228726 , n220106 );
nand ( n240519 , n240517 , n240518 );
nand ( n240520 , n228868 , n240519 );
nand ( n240521 , n240514 , n240520 );
not ( n240522 , n240138 );
not ( n240523 , n234371 );
or ( n240524 , n240522 , n240523 );
not ( n240525 , n234751 );
not ( n240526 , n231477 );
or ( n240527 , n240525 , n240526 );
nand ( n240528 , n229761 , n215989 );
nand ( n240529 , n240527 , n240528 );
nand ( n240530 , n234378 , n240529 );
nand ( n240531 , n240524 , n240530 );
xor ( n240532 , n240521 , n240531 );
or ( n240533 , n239269 , n240147 );
not ( n240534 , n229629 );
not ( n240535 , n230725 );
or ( n240536 , n240534 , n240535 );
nand ( n240537 , n235279 , n211422 );
nand ( n240538 , n240536 , n240537 );
not ( n240539 , n240538 );
or ( n240540 , n238275 , n240539 );
nand ( n240541 , n240533 , n240540 );
xor ( n240542 , n240532 , n240541 );
xor ( n240543 , n240521 , n240531 );
and ( n240544 , n240543 , n240541 );
and ( n240545 , n240521 , n240531 );
or ( n240546 , n240544 , n240545 );
xor ( n240547 , n240461 , n240469 );
xor ( n240548 , n240547 , n240473 );
xor ( n240549 , n240461 , n240469 );
and ( n240550 , n240549 , n240473 );
and ( n240551 , n240461 , n240469 );
or ( n240552 , n240550 , n240551 );
not ( n240553 , n227294 );
not ( n240554 , n239598 );
not ( n240555 , n221725 );
or ( n240556 , n240554 , n240555 );
nand ( n240557 , n226922 , n223156 );
nand ( n240558 , n240556 , n240557 );
not ( n240559 , n240558 );
or ( n240560 , n240553 , n240559 );
nand ( n240561 , n240245 , n238409 );
nand ( n240562 , n240560 , n240561 );
not ( n240563 , n224087 );
not ( n240564 , n240257 );
or ( n240565 , n240563 , n240564 );
not ( n240566 , n40625 );
not ( n240567 , n224095 );
or ( n240568 , n240566 , n240567 );
nand ( n240569 , n221040 , n224096 );
nand ( n240570 , n240568 , n240569 );
nand ( n240571 , n240570 , n227782 );
nand ( n240572 , n240565 , n240571 );
xor ( n240573 , n240562 , n240572 );
not ( n240574 , n223665 );
not ( n240575 , n240350 );
or ( n240576 , n240574 , n240575 );
not ( n240577 , n221241 );
not ( n240578 , n235820 );
not ( n240579 , n240578 );
or ( n240580 , n240577 , n240579 );
not ( n240581 , n235817 );
nand ( n240582 , n240581 , n238363 );
nand ( n240583 , n240580 , n240582 );
nand ( n240584 , n240583 , n218843 );
nand ( n240585 , n240576 , n240584 );
xor ( n240586 , n240573 , n240585 );
not ( n240587 , n221637 );
not ( n240588 , n238705 );
buf ( n240589 , n40181 );
not ( n240590 , n240589 );
or ( n240591 , n240588 , n240590 );
not ( n240592 , n237937 );
nand ( n240593 , n240592 , n238377 );
nand ( n240594 , n240591 , n240593 );
not ( n240595 , n240594 );
or ( n240596 , n240587 , n240595 );
nand ( n240597 , n240222 , n221626 );
nand ( n240598 , n240596 , n240597 );
not ( n240599 , n237493 );
not ( n240600 , n222430 );
not ( n240601 , n238383 );
not ( n240602 , n240601 );
or ( n240603 , n240600 , n240602 );
nand ( n240604 , n40259 , n238719 );
nand ( n240605 , n240603 , n240604 );
not ( n240606 , n240605 );
or ( n240607 , n240599 , n240606 );
nand ( n240608 , n222454 , n240235 );
nand ( n240609 , n240607 , n240608 );
xor ( n240610 , n240598 , n240609 );
xor ( n240611 , n240610 , n240212 );
xor ( n240612 , n240586 , n240611 );
not ( n240613 , n237914 );
not ( n240614 , n234273 );
not ( n240615 , n218911 );
or ( n240616 , n240614 , n240615 );
buf ( n240617 , n234273 );
or ( n240618 , n240617 , n219533 );
nand ( n240619 , n240616 , n240618 );
not ( n240620 , n240619 );
or ( n240621 , n240613 , n240620 );
nand ( n240622 , n240267 , n239492 );
nand ( n240623 , n240621 , n240622 );
not ( n240624 , n220881 );
not ( n240625 , n220151 );
not ( n240626 , n237600 );
or ( n240627 , n240625 , n240626 );
nand ( n240628 , n235031 , n222414 );
nand ( n240629 , n240627 , n240628 );
not ( n240630 , n240629 );
or ( n240631 , n240624 , n240630 );
nand ( n240632 , n240292 , n220492 );
nand ( n240633 , n240631 , n240632 );
xor ( n240634 , n240623 , n240633 );
not ( n240635 , n220930 );
not ( n240636 , n220906 );
not ( n240637 , n238362 );
not ( n240638 , n240637 );
or ( n240639 , n240636 , n240638 );
nand ( n240640 , n40415 , n239066 );
nand ( n240641 , n240639 , n240640 );
not ( n240642 , n240641 );
or ( n240643 , n240635 , n240642 );
nand ( n240644 , n240198 , n235913 );
nand ( n240645 , n240643 , n240644 );
xor ( n240646 , n240634 , n240645 );
xor ( n240647 , n240612 , n240646 );
xor ( n240648 , n240586 , n240611 );
and ( n240649 , n240648 , n240646 );
and ( n240650 , n240586 , n240611 );
or ( n240651 , n240649 , n240650 );
and ( n240652 , n240156 , n225768 );
and ( n240653 , n218884 , n229806 );
not ( n240654 , n218884 );
and ( n240655 , n240654 , n229807 );
or ( n240656 , n240653 , n240655 );
not ( n240657 , n240656 );
or ( n240658 , n240657 , n238777 );
not ( n240659 , n238999 );
nand ( n240660 , n240659 , n240175 );
nand ( n240661 , n240658 , n240660 );
xor ( n240662 , n240652 , n240661 );
not ( n240663 , n239530 );
not ( n240664 , n219424 );
not ( n240665 , n39996 );
or ( n240666 , n240664 , n240665 );
buf ( n240667 , n225111 );
nand ( n240668 , n240667 , n219440 );
nand ( n240669 , n240666 , n240668 );
not ( n240670 , n240669 );
or ( n240671 , n240663 , n240670 );
or ( n240672 , n240281 , n219791 );
nand ( n240673 , n240671 , n240672 );
xor ( n240674 , n240662 , n240673 );
xor ( n240675 , n240674 , n240465 );
or ( n240676 , n240360 , n226942 );
not ( n240677 , n234094 );
not ( n240678 , n240677 );
not ( n240679 , n220038 );
and ( n240680 , n240678 , n240679 );
not ( n240681 , n238472 );
not ( n240682 , n240681 );
and ( n240683 , n240682 , n220038 );
nor ( n240684 , n240680 , n240683 );
or ( n240685 , n240684 , n226940 );
nand ( n240686 , n240676 , n240685 );
not ( n240687 , n229395 );
or ( n240688 , n240377 , n240687 );
xor ( n240689 , n227599 , n236840 );
or ( n240690 , n240689 , n227121 );
nand ( n240691 , n240688 , n240690 );
xor ( n240692 , n240686 , n240691 );
not ( n240693 , n240321 );
or ( n240694 , n240693 , n239938 );
not ( n240695 , n229261 );
not ( n240696 , n229704 );
or ( n240697 , n240695 , n240696 );
nand ( n240698 , n234792 , n234000 );
nand ( n240699 , n240697 , n240698 );
not ( n240700 , n240699 );
or ( n240701 , n240700 , n239946 );
nand ( n240702 , n240694 , n240701 );
xor ( n240703 , n240692 , n240702 );
xor ( n240704 , n240675 , n240703 );
xor ( n240705 , n240674 , n240465 );
and ( n240706 , n240705 , n240703 );
and ( n240707 , n240674 , n240465 );
or ( n240708 , n240706 , n240707 );
or ( n240709 , n240336 , n227130 );
not ( n240710 , n39607 );
and ( n240711 , n234015 , n240710 );
not ( n240712 , n234015 );
and ( n240713 , n240712 , n235977 );
or ( n240714 , n240711 , n240713 );
or ( n240715 , n240714 , n227138 );
nand ( n240716 , n240709 , n240715 );
xor ( n240717 , n240716 , n240155 );
not ( n240718 , n240310 );
not ( n240719 , n227260 );
or ( n240720 , n240718 , n240719 );
and ( n240721 , n233053 , n235691 );
not ( n240722 , n233053 );
and ( n240723 , n240722 , n209709 );
nor ( n240724 , n240721 , n240723 );
or ( n240725 , n240724 , n236271 );
nand ( n240726 , n240720 , n240725 );
xor ( n240727 , n240717 , n240726 );
xor ( n240728 , n240477 , n240727 );
xor ( n240729 , n240728 , n240481 );
xor ( n240730 , n240477 , n240727 );
and ( n240731 , n240730 , n240481 );
and ( n240732 , n240477 , n240727 );
or ( n240733 , n240731 , n240732 );
not ( n240734 , n219461 );
not ( n240735 , n240395 );
or ( n240736 , n240734 , n240735 );
not ( n240737 , n218775 );
not ( n240738 , n233856 );
not ( n240739 , n240738 );
or ( n240740 , n240737 , n240739 );
nand ( n240741 , n233856 , n238352 );
nand ( n240742 , n240740 , n240741 );
nand ( n240743 , n240742 , n218232 );
nand ( n240744 , n240736 , n240743 );
xor ( n240745 , n240744 , n240542 );
xor ( n240746 , n240745 , n240507 );
xor ( n240747 , n240746 , n240190 );
xor ( n240748 , n240747 , n240301 );
xor ( n240749 , n240746 , n240190 );
and ( n240750 , n240749 , n240301 );
and ( n240751 , n240746 , n240190 );
or ( n240752 , n240750 , n240751 );
xor ( n240753 , n240184 , n240441 );
xor ( n240754 , n240753 , n240457 );
xor ( n240755 , n240754 , n240344 );
xor ( n240756 , n240755 , n240704 );
xor ( n240757 , n240754 , n240344 );
and ( n240758 , n240757 , n240704 );
and ( n240759 , n240754 , n240344 );
or ( n240760 , n240758 , n240759 );
xor ( n240761 , n240647 , n240548 );
xor ( n240762 , n240761 , n240387 );
xor ( n240763 , n240647 , n240548 );
and ( n240764 , n240763 , n240387 );
and ( n240765 , n240647 , n240548 );
or ( n240766 , n240764 , n240765 );
xor ( n240767 , n240729 , n240405 );
xor ( n240768 , n240767 , n240413 );
xor ( n240769 , n240729 , n240405 );
and ( n240770 , n240769 , n240413 );
and ( n240771 , n240729 , n240405 );
or ( n240772 , n240770 , n240771 );
xor ( n240773 , n240748 , n240419 );
xor ( n240774 , n240773 , n240762 );
xor ( n240775 , n240748 , n240419 );
and ( n240776 , n240775 , n240762 );
and ( n240777 , n240748 , n240419 );
or ( n240778 , n240776 , n240777 );
xor ( n240779 , n240756 , n240768 );
xor ( n240780 , n240779 , n240425 );
xor ( n240781 , n240756 , n240768 );
and ( n240782 , n240781 , n240425 );
and ( n240783 , n240756 , n240768 );
or ( n240784 , n240782 , n240783 );
xor ( n240785 , n240652 , n240661 );
and ( n240786 , n240785 , n240673 );
and ( n240787 , n240652 , n240661 );
or ( n240788 , n240786 , n240787 );
xor ( n240789 , n240431 , n240774 );
xor ( n240790 , n240789 , n240437 );
xor ( n240791 , n240431 , n240774 );
and ( n240792 , n240791 , n240437 );
and ( n240793 , n240431 , n240774 );
or ( n240794 , n240792 , n240793 );
xor ( n240795 , n240780 , n240790 );
xor ( n240796 , n240795 , n240447 );
xor ( n240797 , n240780 , n240790 );
and ( n240798 , n240797 , n240447 );
and ( n240799 , n240780 , n240790 );
or ( n240800 , n240798 , n240799 );
xor ( n240801 , n240623 , n240633 );
and ( n240802 , n240801 , n240645 );
and ( n240803 , n240623 , n240633 );
or ( n240804 , n240802 , n240803 );
xor ( n240805 , n240598 , n240609 );
and ( n240806 , n240805 , n240212 );
and ( n240807 , n240598 , n240609 );
or ( n240808 , n240806 , n240807 );
xor ( n240809 , n240562 , n240572 );
and ( n240810 , n240809 , n240585 );
and ( n240811 , n240562 , n240572 );
or ( n240812 , n240810 , n240811 );
xor ( n240813 , n240686 , n240691 );
and ( n240814 , n240813 , n240702 );
and ( n240815 , n240686 , n240691 );
or ( n240816 , n240814 , n240815 );
xor ( n240817 , n240716 , n240155 );
and ( n240818 , n240817 , n240726 );
and ( n240819 , n240716 , n240155 );
or ( n240820 , n240818 , n240819 );
xor ( n240821 , n240744 , n240542 );
and ( n240822 , n240821 , n240507 );
and ( n240823 , n240744 , n240542 );
or ( n240824 , n240822 , n240823 );
xor ( n240825 , n240184 , n240441 );
and ( n240826 , n240825 , n240457 );
and ( n240827 , n240184 , n240441 );
or ( n240828 , n240826 , n240827 );
not ( n240829 , n240519 );
not ( n240830 , n228858 );
or ( n240831 , n240829 , n240830 );
not ( n240832 , n217318 );
not ( n240833 , n229249 );
or ( n240834 , n240832 , n240833 );
nand ( n240835 , n231943 , n217314 );
nand ( n240836 , n240834 , n240835 );
nand ( n240837 , n240836 , n229738 );
nand ( n240838 , n240831 , n240837 );
not ( n240839 , n240538 );
not ( n240840 , n230720 );
or ( n240841 , n240839 , n240840 );
not ( n240842 , n215796 );
not ( n240843 , n230725 );
or ( n240844 , n240842 , n240843 );
nand ( n240845 , n230991 , n216261 );
nand ( n240846 , n240844 , n240845 );
nand ( n240847 , n230708 , n240846 );
nand ( n240848 , n240841 , n240847 );
xor ( n240849 , n240838 , n240848 );
not ( n240850 , n240529 );
not ( n240851 , n229773 );
or ( n240852 , n240850 , n240851 );
not ( n240853 , n231476 );
not ( n240854 , n219902 );
not ( n240855 , n233399 );
or ( n240856 , n240854 , n240855 );
not ( n240857 , n231997 );
nand ( n240858 , n240857 , n208597 );
nand ( n240859 , n240856 , n240858 );
nand ( n240860 , n240853 , n240859 );
nand ( n240861 , n240852 , n240860 );
xor ( n240862 , n240849 , n240861 );
xor ( n240863 , n240838 , n240848 );
and ( n240864 , n240863 , n240861 );
and ( n240865 , n240838 , n240848 );
or ( n240866 , n240864 , n240865 );
and ( n240867 , n240156 , n226225 );
not ( n240868 , n226885 );
not ( n240869 , n239774 );
not ( n240870 , n217964 );
or ( n240871 , n240869 , n240870 );
nand ( n240872 , n208002 , n226650 );
nand ( n240873 , n240871 , n240872 );
not ( n240874 , n240873 );
or ( n240875 , n240868 , n240874 );
not ( n240876 , n234894 );
nand ( n240877 , n240876 , n240494 );
nand ( n240878 , n240875 , n240877 );
xor ( n240879 , n240867 , n240878 );
not ( n240880 , n238776 );
not ( n240881 , n229806 );
not ( n240882 , n40766 );
or ( n240883 , n240881 , n240882 );
nand ( n240884 , n221342 , n233962 );
nand ( n240885 , n240883 , n240884 );
not ( n240886 , n240885 );
or ( n240887 , n240880 , n240886 );
nand ( n240888 , n240656 , n239416 );
nand ( n240889 , n240887 , n240888 );
xor ( n240890 , n240879 , n240889 );
xor ( n240891 , n240867 , n240878 );
and ( n240892 , n240891 , n240889 );
and ( n240893 , n240867 , n240878 );
or ( n240894 , n240892 , n240893 );
not ( n240895 , n224087 );
not ( n240896 , n240570 );
or ( n240897 , n240895 , n240896 );
not ( n240898 , n237130 );
not ( n240899 , n40660 );
or ( n240900 , n240898 , n240899 );
nand ( n240901 , n207936 , n234764 );
nand ( n240902 , n240900 , n240901 );
nand ( n240903 , n240902 , n227782 );
nand ( n240904 , n240897 , n240903 );
not ( n240905 , n240619 );
not ( n240906 , n239492 );
or ( n240907 , n240905 , n240906 );
not ( n240908 , n233952 );
not ( n240909 , n219880 );
or ( n240910 , n240908 , n240909 );
nand ( n240911 , n219226 , n234273 );
nand ( n240912 , n240910 , n240911 );
nand ( n240913 , n240912 , n240020 );
nand ( n240914 , n240907 , n240913 );
xor ( n240915 , n240904 , n240914 );
not ( n240916 , n219076 );
not ( n240917 , n219797 );
not ( n240918 , n240917 );
not ( n240919 , n230280 );
or ( n240920 , n240918 , n240919 );
nand ( n240921 , n233525 , n219440 );
nand ( n240922 , n240920 , n240921 );
not ( n240923 , n240922 );
or ( n240924 , n240916 , n240923 );
nand ( n240925 , n240669 , n219792 );
nand ( n240926 , n240924 , n240925 );
xor ( n240927 , n240915 , n240926 );
not ( n240928 , n220164 );
not ( n240929 , n240629 );
or ( n240930 , n240928 , n240929 );
not ( n240931 , n221593 );
not ( n240932 , n230490 );
or ( n240933 , n240931 , n240932 );
nand ( n240934 , n234506 , n222414 );
nand ( n240935 , n240933 , n240934 );
nand ( n240936 , n240935 , n220881 );
nand ( n240937 , n240930 , n240936 );
not ( n240938 , n220930 );
not ( n240939 , n222399 );
not ( n240940 , n237971 );
or ( n240941 , n240939 , n240940 );
nand ( n240942 , n236290 , n236754 );
nand ( n240943 , n240941 , n240942 );
not ( n240944 , n240943 );
or ( n240945 , n240938 , n240944 );
nand ( n240946 , n240641 , n235913 );
nand ( n240947 , n240945 , n240946 );
xor ( n240948 , n240937 , n240947 );
not ( n240949 , n221626 );
not ( n240950 , n240594 );
or ( n240951 , n240949 , n240950 );
not ( n240952 , n238705 );
not ( n240953 , n224700 );
or ( n240954 , n240952 , n240953 );
nand ( n240955 , n236300 , n222586 );
nand ( n240956 , n240954 , n240955 );
nand ( n240957 , n240956 , n221637 );
nand ( n240958 , n240951 , n240957 );
xor ( n240959 , n240948 , n240958 );
xor ( n240960 , n240927 , n240959 );
xor ( n240961 , n240960 , n240820 );
xor ( n240962 , n240927 , n240959 );
and ( n240963 , n240962 , n240820 );
and ( n240964 , n240927 , n240959 );
or ( n240965 , n240963 , n240964 );
xor ( n240966 , n240812 , n240816 );
or ( n240967 , n240689 , n240687 );
not ( n240968 , n233544 );
not ( n240969 , n233362 );
or ( n240970 , n240968 , n240969 );
nand ( n240971 , n233363 , n227599 );
nand ( n240972 , n240970 , n240971 );
not ( n240973 , n240972 );
or ( n240974 , n240973 , n227121 );
nand ( n240975 , n240967 , n240974 );
xor ( n240976 , n240546 , n240975 );
not ( n240977 , n239508 );
not ( n240978 , n240583 );
or ( n240979 , n240977 , n240978 );
not ( n240980 , n221241 );
not ( n240981 , n234350 );
or ( n240982 , n240980 , n240981 );
nand ( n240983 , n238819 , n238755 );
nand ( n240984 , n240982 , n240983 );
nand ( n240985 , n240984 , n218843 );
nand ( n240986 , n240979 , n240985 );
xor ( n240987 , n240976 , n240986 );
xor ( n240988 , n240966 , n240987 );
xor ( n240989 , n240812 , n240816 );
and ( n240990 , n240989 , n240987 );
and ( n240991 , n240812 , n240816 );
or ( n240992 , n240990 , n240991 );
or ( n240993 , n240724 , n240719 );
not ( n240994 , n240358 );
not ( n240995 , n233053 );
and ( n240996 , n240994 , n240995 );
and ( n240997 , n240358 , n233053 );
nor ( n240998 , n240996 , n240997 );
or ( n240999 , n236271 , n240998 );
nand ( n241000 , n240993 , n240999 );
not ( n241001 , n229964 );
not ( n241002 , n229261 );
not ( n241003 , n230269 );
or ( n241004 , n241002 , n241003 );
nand ( n241005 , n39365 , n229262 );
nand ( n241006 , n241004 , n241005 );
not ( n241007 , n241006 );
or ( n241008 , n241001 , n241007 );
nand ( n241009 , n240699 , n234006 );
nand ( n241010 , n241008 , n241009 );
xor ( n241011 , n241000 , n241010 );
or ( n241012 , n240714 , n227130 );
not ( n241013 , n231500 );
not ( n241014 , n236382 );
or ( n241015 , n241013 , n241014 );
nand ( n241016 , n39089 , n234015 );
nand ( n241017 , n241015 , n241016 );
not ( n241018 , n241017 );
or ( n241019 , n241018 , n227138 );
nand ( n241020 , n241012 , n241019 );
xor ( n241021 , n241011 , n241020 );
xor ( n241022 , n241021 , n240824 );
not ( n241023 , n226287 );
not ( n241024 , n226292 );
or ( n241025 , n241023 , n241024 );
or ( n241026 , n240684 , n216730 );
nand ( n241027 , n241025 , n241026 );
not ( n241028 , n219461 );
not ( n241029 , n240742 );
or ( n241030 , n241028 , n241029 );
not ( n241031 , n218205 );
not ( n241032 , n230241 );
or ( n241033 , n241031 , n241032 );
nand ( n241034 , n238877 , n218226 );
nand ( n241035 , n241033 , n241034 );
nand ( n241036 , n241035 , n218232 );
nand ( n241037 , n241030 , n241036 );
xor ( n241038 , n241027 , n241037 );
xor ( n241039 , n241038 , n240511 );
xor ( n241040 , n241022 , n241039 );
xor ( n241041 , n241021 , n240824 );
and ( n241042 , n241041 , n241039 );
and ( n241043 , n241021 , n240824 );
or ( n241044 , n241042 , n241043 );
xor ( n241045 , n240804 , n240808 );
not ( n241046 , n240504 );
not ( n241047 , n241046 );
not ( n241048 , n237810 );
or ( n241049 , n241047 , n241048 );
not ( n241050 , n219201 );
not ( n241051 , n233451 );
or ( n241052 , n241050 , n241051 );
nand ( n241053 , n236188 , n231240 );
nand ( n241054 , n241052 , n241053 );
nand ( n241055 , n238240 , n241054 );
nand ( n241056 , n241049 , n241055 );
not ( n241057 , n241056 );
not ( n241058 , n222454 );
not ( n241059 , n240605 );
or ( n241060 , n241058 , n241059 );
not ( n241061 , n222892 );
not ( n241062 , n230511 );
or ( n241063 , n241061 , n241062 );
nand ( n241064 , n226505 , n222458 );
nand ( n241065 , n241063 , n241064 );
nand ( n241066 , n241065 , n237493 );
nand ( n241067 , n241060 , n241066 );
xor ( n241068 , n241057 , n241067 );
not ( n241069 , n238409 );
not ( n241070 , n240558 );
or ( n241071 , n241069 , n241070 );
not ( n241072 , n223156 );
not ( n241073 , n40410 );
or ( n241074 , n241072 , n241073 );
not ( n241075 , n239458 );
nand ( n241076 , n241075 , n239598 );
nand ( n241077 , n241074 , n241076 );
nand ( n241078 , n241077 , n222768 );
nand ( n241079 , n241071 , n241078 );
xor ( n241080 , n241068 , n241079 );
xor ( n241081 , n241045 , n241080 );
xor ( n241082 , n240828 , n241081 );
xor ( n241083 , n241082 , n240651 );
xor ( n241084 , n240828 , n241081 );
and ( n241085 , n241084 , n240651 );
and ( n241086 , n240828 , n241081 );
or ( n241087 , n241085 , n241086 );
xor ( n241088 , n240862 , n240890 );
xor ( n241089 , n241088 , n240788 );
xor ( n241090 , n240552 , n241089 );
xor ( n241091 , n241090 , n240708 );
xor ( n241092 , n240552 , n241089 );
and ( n241093 , n241092 , n240708 );
and ( n241094 , n240552 , n241089 );
or ( n241095 , n241093 , n241094 );
xor ( n241096 , n240988 , n240961 );
xor ( n241097 , n241096 , n241040 );
xor ( n241098 , n240988 , n240961 );
and ( n241099 , n241098 , n241040 );
and ( n241100 , n240988 , n240961 );
or ( n241101 , n241099 , n241100 );
xor ( n241102 , n240733 , n240752 );
xor ( n241103 , n241102 , n241091 );
xor ( n241104 , n240733 , n240752 );
and ( n241105 , n241104 , n241091 );
and ( n241106 , n240733 , n240752 );
or ( n241107 , n241105 , n241106 );
xor ( n241108 , n240760 , n241083 );
xor ( n241109 , n241108 , n241097 );
xor ( n241110 , n240760 , n241083 );
and ( n241111 , n241110 , n241097 );
and ( n241112 , n240760 , n241083 );
or ( n241113 , n241111 , n241112 );
xor ( n241114 , n240766 , n240772 );
xor ( n241115 , n241114 , n241103 );
xor ( n241116 , n240766 , n240772 );
and ( n241117 , n241116 , n241103 );
and ( n241118 , n240766 , n240772 );
or ( n241119 , n241117 , n241118 );
xor ( n241120 , n241109 , n240778 );
xor ( n241121 , n241120 , n240784 );
xor ( n241122 , n241109 , n240778 );
and ( n241123 , n241122 , n240784 );
and ( n241124 , n241109 , n240778 );
or ( n241125 , n241123 , n241124 );
xor ( n241126 , n240937 , n240947 );
and ( n241127 , n241126 , n240958 );
and ( n241128 , n240937 , n240947 );
or ( n241129 , n241127 , n241128 );
xor ( n241130 , n241115 , n241121 );
xor ( n241131 , n241130 , n240794 );
xor ( n241132 , n241115 , n241121 );
and ( n241133 , n241132 , n240794 );
and ( n241134 , n241115 , n241121 );
or ( n241135 , n241133 , n241134 );
xor ( n241136 , n241057 , n241067 );
and ( n241137 , n241136 , n241079 );
and ( n241138 , n241057 , n241067 );
or ( n241139 , n241137 , n241138 );
xor ( n241140 , n240904 , n240914 );
and ( n241141 , n241140 , n240926 );
and ( n241142 , n240904 , n240914 );
or ( n241143 , n241141 , n241142 );
xor ( n241144 , n241000 , n241010 );
and ( n241145 , n241144 , n241020 );
and ( n241146 , n241000 , n241010 );
or ( n241147 , n241145 , n241146 );
xor ( n241148 , n241027 , n241037 );
and ( n241149 , n241148 , n240511 );
and ( n241150 , n241027 , n241037 );
or ( n241151 , n241149 , n241150 );
xor ( n241152 , n240546 , n240975 );
and ( n241153 , n241152 , n240986 );
and ( n241154 , n240546 , n240975 );
or ( n241155 , n241153 , n241154 );
xor ( n241156 , n240862 , n240890 );
and ( n241157 , n241156 , n240788 );
and ( n241158 , n240862 , n240890 );
or ( n241159 , n241157 , n241158 );
xor ( n241160 , n240804 , n240808 );
and ( n241161 , n241160 , n241080 );
and ( n241162 , n240804 , n240808 );
or ( n241163 , n241161 , n241162 );
not ( n241164 , n220032 );
not ( n241165 , n216730 );
or ( n241166 , n241164 , n241165 );
nand ( n241167 , n241166 , n226292 );
not ( n241168 , n241054 );
not ( n241169 , n232440 );
or ( n241170 , n241168 , n241169 );
not ( n241171 , n233450 );
not ( n241172 , n219386 );
or ( n241173 , n241171 , n241172 );
nand ( n241174 , n234394 , n41165 );
nand ( n241175 , n241173 , n241174 );
nand ( n241176 , n227737 , n241175 );
nand ( n241177 , n241170 , n241176 );
xor ( n241178 , n241167 , n241177 );
not ( n241179 , n240836 );
or ( n241180 , n237038 , n241179 );
and ( n241181 , n231762 , n228847 );
not ( n241182 , n231762 );
and ( n241183 , n241182 , n228850 );
nor ( n241184 , n241181 , n241183 );
or ( n241185 , n237041 , n241184 );
nand ( n241186 , n241180 , n241185 );
xor ( n241187 , n241178 , n241186 );
xor ( n241188 , n241167 , n241177 );
and ( n241189 , n241188 , n241186 );
and ( n241190 , n241167 , n241177 );
or ( n241191 , n241189 , n241190 );
not ( n241192 , n240859 );
not ( n241193 , n234371 );
or ( n241194 , n241192 , n241193 );
not ( n241195 , n229761 );
not ( n241196 , n217147 );
and ( n241197 , n241195 , n241196 );
and ( n241198 , n231480 , n216520 );
nor ( n241199 , n241197 , n241198 );
not ( n241200 , n241199 );
nand ( n241201 , n241200 , n234378 );
nand ( n241202 , n241194 , n241201 );
not ( n241203 , n240846 );
not ( n241204 , n233879 );
or ( n241205 , n241203 , n241204 );
not ( n241206 , n234751 );
not ( n241207 , n232404 );
or ( n241208 , n241206 , n241207 );
nand ( n241209 , n234382 , n216500 );
nand ( n241210 , n241208 , n241209 );
nand ( n241211 , n232402 , n241210 );
nand ( n241212 , n241205 , n241211 );
xor ( n241213 , n241202 , n241212 );
and ( n241214 , n240156 , n41565 );
xor ( n241215 , n241213 , n241214 );
xor ( n241216 , n241202 , n241212 );
and ( n241217 , n241216 , n241214 );
and ( n241218 , n241202 , n241212 );
or ( n241219 , n241217 , n241218 );
not ( n241220 , n221266 );
not ( n241221 , n240943 );
or ( n241222 , n241220 , n241221 );
not ( n241223 , n222399 );
not ( n241224 , n239916 );
or ( n241225 , n241223 , n241224 );
nand ( n241226 , n40547 , n222400 );
nand ( n241227 , n241225 , n241226 );
nand ( n241228 , n241227 , n221674 );
nand ( n241229 , n241222 , n241228 );
not ( n241230 , n221637 );
not ( n241231 , n237937 );
not ( n241232 , n227004 );
or ( n241233 , n241231 , n241232 );
nand ( n241234 , n239139 , n221632 );
nand ( n241235 , n241233 , n241234 );
not ( n241236 , n241235 );
or ( n241237 , n241230 , n241236 );
nand ( n241238 , n240956 , n221626 );
nand ( n241239 , n241237 , n241238 );
xor ( n241240 , n241229 , n241239 );
xor ( n241241 , n241240 , n241056 );
not ( n241242 , n226885 );
not ( n241243 , n239774 );
not ( n241244 , n218884 );
or ( n241245 , n241243 , n241244 );
nand ( n241246 , n40710 , n238230 );
nand ( n241247 , n241245 , n241246 );
not ( n241248 , n241247 );
or ( n241249 , n241242 , n241248 );
nand ( n241250 , n240873 , n237797 );
nand ( n241251 , n241249 , n241250 );
not ( n241252 , n220492 );
not ( n241253 , n240935 );
or ( n241254 , n241252 , n241253 );
not ( n241255 , n221593 );
not ( n241256 , n39996 );
or ( n241257 , n241255 , n241256 );
nand ( n241258 , n226964 , n221257 );
nand ( n241259 , n241257 , n241258 );
nand ( n241260 , n241259 , n220881 );
nand ( n241261 , n241254 , n241260 );
xor ( n241262 , n241251 , n241261 );
not ( n241263 , n238776 );
not ( n241264 , n229806 );
not ( n241265 , n218912 );
or ( n241266 , n241264 , n241265 );
nand ( n241267 , n218911 , n229807 );
nand ( n241268 , n241266 , n241267 );
not ( n241269 , n241268 );
or ( n241270 , n241263 , n241269 );
nand ( n241271 , n240885 , n239416 );
nand ( n241272 , n241270 , n241271 );
xor ( n241273 , n241262 , n241272 );
xor ( n241274 , n241241 , n241273 );
xor ( n241275 , n241274 , n241155 );
xor ( n241276 , n241241 , n241273 );
and ( n241277 , n241276 , n241155 );
and ( n241278 , n241241 , n241273 );
or ( n241279 , n241277 , n241278 );
xor ( n241280 , n241143 , n241147 );
xor ( n241281 , n241280 , n241151 );
xor ( n241282 , n241143 , n241147 );
and ( n241283 , n241282 , n241151 );
and ( n241284 , n241143 , n241147 );
or ( n241285 , n241283 , n241284 );
not ( n241286 , n237914 );
not ( n241287 , n240617 );
not ( n241288 , n241287 );
not ( n241289 , n234108 );
or ( n241290 , n241288 , n241289 );
nand ( n241291 , n40625 , n235200 );
nand ( n241292 , n241290 , n241291 );
not ( n241293 , n241292 );
or ( n241294 , n241286 , n241293 );
nand ( n241295 , n240912 , n227792 );
nand ( n241296 , n241294 , n241295 );
not ( n241297 , n220507 );
not ( n241298 , n240922 );
or ( n241299 , n241297 , n241298 );
not ( n241300 , n219800 );
not ( n241301 , n226724 );
or ( n241302 , n241300 , n241301 );
not ( n241303 , n39927 );
nand ( n241304 , n241303 , n219440 );
nand ( n241305 , n241302 , n241304 );
nand ( n241306 , n241305 , n239530 );
nand ( n241307 , n241299 , n241306 );
xor ( n241308 , n241296 , n241307 );
not ( n241309 , n223949 );
not ( n241310 , n226655 );
not ( n241311 , n238473 );
or ( n241312 , n241310 , n241311 );
nand ( n241313 , n209964 , n233053 );
nand ( n241314 , n241312 , n241313 );
not ( n241315 , n241314 );
or ( n241316 , n241309 , n241315 );
not ( n241317 , n240998 );
nand ( n241318 , n241317 , n227260 );
nand ( n241319 , n241316 , n241318 );
xor ( n241320 , n241308 , n241319 );
not ( n241321 , n228237 );
not ( n241322 , n233544 );
not ( n241323 , n209709 );
or ( n241324 , n241322 , n241323 );
nand ( n241325 , n232856 , n227599 );
nand ( n241326 , n241324 , n241325 );
not ( n241327 , n241326 );
or ( n241328 , n241321 , n241327 );
nand ( n241329 , n240972 , n225478 );
nand ( n241330 , n241328 , n241329 );
xor ( n241331 , n240866 , n241330 );
not ( n241332 , n218843 );
not ( n241333 , n221241 );
not ( n241334 , n225792 );
or ( n241335 , n241333 , n241334 );
nand ( n241336 , n227696 , n238755 );
nand ( n241337 , n241335 , n241336 );
not ( n241338 , n241337 );
or ( n241339 , n241332 , n241338 );
nand ( n241340 , n240984 , n223665 );
nand ( n241341 , n241339 , n241340 );
xor ( n241342 , n241331 , n241341 );
xor ( n241343 , n241320 , n241342 );
not ( n241344 , n229974 );
not ( n241345 , n241006 );
or ( n241346 , n241344 , n241345 );
not ( n241347 , n229261 );
not ( n241348 , n233810 );
or ( n241349 , n241347 , n241348 );
nand ( n241350 , n39286 , n229262 );
nand ( n241351 , n241349 , n241350 );
nand ( n241352 , n241351 , n229964 );
nand ( n241353 , n241346 , n241352 );
not ( n241354 , n231018 );
not ( n241355 , n241017 );
or ( n241356 , n241354 , n241355 );
not ( n241357 , n217616 );
not ( n241358 , n235962 );
or ( n241359 , n241357 , n241358 );
nand ( n241360 , n234792 , n234015 );
nand ( n241361 , n241359 , n241360 );
nand ( n241362 , n241361 , n220067 );
nand ( n241363 , n241356 , n241362 );
xor ( n241364 , n241353 , n241363 );
not ( n241365 , n219461 );
not ( n241366 , n241035 );
or ( n241367 , n241365 , n241366 );
not ( n241368 , n233083 );
not ( n241369 , n39608 );
not ( n241370 , n241369 );
or ( n241371 , n241368 , n241370 );
nand ( n241372 , n39608 , n238352 );
nand ( n241373 , n241371 , n241372 );
nand ( n241374 , n241373 , n218232 );
nand ( n241375 , n241367 , n241374 );
xor ( n241376 , n241364 , n241375 );
xor ( n241377 , n241343 , n241376 );
xor ( n241378 , n241320 , n241342 );
and ( n241379 , n241378 , n241376 );
and ( n241380 , n241320 , n241342 );
or ( n241381 , n241379 , n241380 );
xor ( n241382 , n241215 , n241187 );
xor ( n241383 , n241382 , n240894 );
xor ( n241384 , n241159 , n241383 );
xor ( n241385 , n241384 , n240965 );
xor ( n241386 , n241159 , n241383 );
and ( n241387 , n241386 , n240965 );
and ( n241388 , n241159 , n241383 );
or ( n241389 , n241387 , n241388 );
xor ( n241390 , n241129 , n241139 );
not ( n241391 , n237503 );
not ( n241392 , n241065 );
or ( n241393 , n241391 , n241392 );
and ( n241394 , n222434 , n40181 );
not ( n241395 , n222434 );
and ( n241396 , n241395 , n236719 );
or ( n241397 , n241394 , n241396 );
nand ( n241398 , n241397 , n237493 );
nand ( n241399 , n241393 , n241398 );
not ( n241400 , n227294 );
not ( n241401 , n239598 );
not ( n241402 , n222552 );
or ( n241403 , n241401 , n241402 );
not ( n241404 , n237005 );
nand ( n241405 , n220970 , n241404 );
nand ( n241406 , n241403 , n241405 );
not ( n241407 , n241406 );
or ( n241408 , n241400 , n241407 );
nand ( n241409 , n238409 , n241077 );
nand ( n241410 , n241408 , n241409 );
xor ( n241411 , n241399 , n241410 );
not ( n241412 , n239495 );
not ( n241413 , n224096 );
not ( n241414 , n221725 );
or ( n241415 , n241413 , n241414 );
nand ( n241416 , n226922 , n238672 );
nand ( n241417 , n241415 , n241416 );
not ( n241418 , n241417 );
or ( n241419 , n241412 , n241418 );
nand ( n241420 , n240902 , n224087 );
nand ( n241421 , n241419 , n241420 );
xor ( n241422 , n241411 , n241421 );
xor ( n241423 , n241390 , n241422 );
xor ( n241424 , n241163 , n241423 );
xor ( n241425 , n241424 , n241044 );
xor ( n241426 , n241163 , n241423 );
and ( n241427 , n241426 , n241044 );
and ( n241428 , n241163 , n241423 );
or ( n241429 , n241427 , n241428 );
xor ( n241430 , n241281 , n240992 );
xor ( n241431 , n241430 , n241275 );
xor ( n241432 , n241281 , n240992 );
and ( n241433 , n241432 , n241275 );
and ( n241434 , n241281 , n240992 );
or ( n241435 , n241433 , n241434 );
xor ( n241436 , n241377 , n241087 );
xor ( n241437 , n241436 , n241385 );
xor ( n241438 , n241377 , n241087 );
and ( n241439 , n241438 , n241385 );
and ( n241440 , n241377 , n241087 );
or ( n241441 , n241439 , n241440 );
xor ( n241442 , n241095 , n241425 );
xor ( n241443 , n241442 , n241101 );
xor ( n241444 , n241095 , n241425 );
and ( n241445 , n241444 , n241101 );
and ( n241446 , n241095 , n241425 );
or ( n241447 , n241445 , n241446 );
xor ( n241448 , n241431 , n241107 );
xor ( n241449 , n241448 , n241437 );
xor ( n241450 , n241431 , n241107 );
and ( n241451 , n241450 , n241437 );
and ( n241452 , n241431 , n241107 );
or ( n241453 , n241451 , n241452 );
xor ( n241454 , n241443 , n241113 );
xor ( n241455 , n241454 , n241119 );
xor ( n241456 , n241443 , n241113 );
and ( n241457 , n241456 , n241119 );
and ( n241458 , n241443 , n241113 );
or ( n241459 , n241457 , n241458 );
xor ( n241460 , n241251 , n241261 );
and ( n241461 , n241460 , n241272 );
and ( n241462 , n241251 , n241261 );
or ( n241463 , n241461 , n241462 );
xor ( n241464 , n241449 , n241455 );
xor ( n241465 , n241464 , n241125 );
xor ( n241466 , n241449 , n241455 );
and ( n241467 , n241466 , n241125 );
and ( n241468 , n241449 , n241455 );
or ( n241469 , n241467 , n241468 );
xor ( n241470 , n241229 , n241239 );
and ( n241471 , n241470 , n241056 );
and ( n241472 , n241229 , n241239 );
or ( n241473 , n241471 , n241472 );
xor ( n241474 , n241399 , n241410 );
and ( n241475 , n241474 , n241421 );
and ( n241476 , n241399 , n241410 );
or ( n241477 , n241475 , n241476 );
xor ( n241478 , n241296 , n241307 );
and ( n241479 , n241478 , n241319 );
and ( n241480 , n241296 , n241307 );
or ( n241481 , n241479 , n241480 );
xor ( n241482 , n241353 , n241363 );
and ( n241483 , n241482 , n241375 );
and ( n241484 , n241353 , n241363 );
or ( n241485 , n241483 , n241484 );
xor ( n241486 , n240866 , n241330 );
and ( n241487 , n241486 , n241341 );
and ( n241488 , n240866 , n241330 );
or ( n241489 , n241487 , n241488 );
xor ( n241490 , n241215 , n241187 );
and ( n241491 , n241490 , n240894 );
and ( n241492 , n241215 , n241187 );
or ( n241493 , n241491 , n241492 );
xor ( n241494 , n241129 , n241139 );
and ( n241495 , n241494 , n241422 );
and ( n241496 , n241129 , n241139 );
or ( n241497 , n241495 , n241496 );
or ( n241498 , n231994 , n241199 );
and ( n241499 , n229762 , n223549 );
and ( n241500 , n234865 , n230171 );
nor ( n241501 , n241499 , n241500 );
or ( n241502 , n241501 , n231476 );
nand ( n241503 , n241498 , n241502 );
and ( n241504 , n233465 , n233279 );
xor ( n241505 , n241503 , n241504 );
not ( n241506 , n241210 );
not ( n241507 , n233105 );
or ( n241508 , n241506 , n241507 );
and ( n241509 , n41321 , n231753 );
not ( n241510 , n41321 );
and ( n241511 , n241510 , n231232 );
or ( n241512 , n241509 , n241511 );
nand ( n241513 , n241512 , n232402 );
nand ( n241514 , n241508 , n241513 );
xor ( n241515 , n241505 , n241514 );
xor ( n241516 , n241503 , n241504 );
and ( n241517 , n241516 , n241514 );
and ( n241518 , n241503 , n241504 );
or ( n241519 , n241517 , n241518 );
not ( n241520 , n241175 );
not ( n241521 , n233446 );
or ( n241522 , n241520 , n241521 );
not ( n241523 , n237816 );
not ( n241524 , n217964 );
or ( n241525 , n241523 , n241524 );
nand ( n241526 , n238671 , n240500 );
nand ( n241527 , n241525 , n241526 );
nand ( n241528 , n241527 , n238240 );
nand ( n241529 , n241522 , n241528 );
not ( n241530 , n227852 );
and ( n241531 , n219239 , n226650 );
not ( n241532 , n219239 );
and ( n241533 , n241532 , n239774 );
or ( n241534 , n241531 , n241533 );
not ( n241535 , n241534 );
or ( n241536 , n241530 , n241535 );
nand ( n241537 , n241247 , n239441 );
nand ( n241538 , n241536 , n241537 );
xor ( n241539 , n241529 , n241538 );
not ( n241540 , n221674 );
not ( n241541 , n220906 );
not ( n241542 , n230490 );
or ( n241543 , n241541 , n241542 );
nand ( n241544 , n223765 , n239066 );
nand ( n241545 , n241543 , n241544 );
not ( n241546 , n241545 );
or ( n241547 , n241540 , n241546 );
nand ( n241548 , n241227 , n235913 );
nand ( n241549 , n241547 , n241548 );
xor ( n241550 , n241539 , n241549 );
xor ( n241551 , n241529 , n241538 );
and ( n241552 , n241551 , n241549 );
and ( n241553 , n241529 , n241538 );
or ( n241554 , n241552 , n241553 );
xor ( n241555 , n241485 , n241481 );
not ( n241556 , n221626 );
not ( n241557 , n241235 );
or ( n241558 , n241556 , n241557 );
not ( n241559 , n222035 );
not ( n241560 , n237971 );
or ( n241561 , n241559 , n241560 );
nand ( n241562 , n236290 , n221612 );
nand ( n241563 , n241561 , n241562 );
nand ( n241564 , n241563 , n221637 );
nand ( n241565 , n241558 , n241564 );
not ( n241566 , n222454 );
not ( n241567 , n241397 );
or ( n241568 , n241566 , n241567 );
not ( n241569 , n222892 );
not ( n241570 , n235383 );
or ( n241571 , n241569 , n241570 );
nand ( n241572 , n222952 , n222429 );
nand ( n241573 , n241571 , n241572 );
nand ( n241574 , n241573 , n237493 );
nand ( n241575 , n241568 , n241574 );
xor ( n241576 , n241565 , n241575 );
not ( n241577 , n241184 );
not ( n241578 , n241577 );
not ( n241579 , n231421 );
or ( n241580 , n241578 , n241579 );
not ( n241581 , n217331 );
not ( n241582 , n228847 );
or ( n241583 , n241581 , n241582 );
not ( n241584 , n219201 );
nand ( n241585 , n241584 , n228850 );
nand ( n241586 , n241583 , n241585 );
nand ( n241587 , n228868 , n241586 );
nand ( n241588 , n241580 , n241587 );
not ( n241589 , n241588 );
xor ( n241590 , n241576 , n241589 );
xor ( n241591 , n241555 , n241590 );
xor ( n241592 , n241485 , n241481 );
and ( n241593 , n241592 , n241590 );
and ( n241594 , n241485 , n241481 );
or ( n241595 , n241593 , n241594 );
not ( n241596 , n239416 );
not ( n241597 , n241268 );
or ( n241598 , n241596 , n241597 );
not ( n241599 , n233962 );
not ( n241600 , n241599 );
not ( n241601 , n40560 );
or ( n241602 , n241600 , n241601 );
nand ( n241603 , n240255 , n233962 );
nand ( n241604 , n241602 , n241603 );
nand ( n241605 , n241604 , n238776 );
nand ( n241606 , n241598 , n241605 );
not ( n241607 , n219779 );
not ( n241608 , n221593 );
not ( n241609 , n39879 );
or ( n241610 , n241608 , n241609 );
nand ( n241611 , n235455 , n220147 );
nand ( n241612 , n241610 , n241611 );
not ( n241613 , n241612 );
or ( n241614 , n241607 , n241613 );
nand ( n241615 , n241259 , n220164 );
nand ( n241616 , n241614 , n241615 );
xor ( n241617 , n241606 , n241616 );
not ( n241618 , n229395 );
not ( n241619 , n241326 );
or ( n241620 , n241618 , n241619 );
not ( n241621 , n227599 );
not ( n241622 , n238835 );
or ( n241623 , n241621 , n241622 );
nand ( n241624 , n233611 , n229387 );
nand ( n241625 , n241623 , n241624 );
nand ( n241626 , n241625 , n219501 );
nand ( n241627 , n241620 , n241626 );
xor ( n241628 , n241617 , n241627 );
not ( n241629 , n229964 );
not ( n241630 , n229261 );
not ( n241631 , n233362 );
or ( n241632 , n241630 , n241631 );
nand ( n241633 , n229217 , n229262 );
nand ( n241634 , n241632 , n241633 );
not ( n241635 , n241634 );
or ( n241636 , n241629 , n241635 );
nand ( n241637 , n241351 , n219368 );
nand ( n241638 , n241636 , n241637 );
not ( n241639 , n239530 );
not ( n241640 , n219424 );
not ( n241641 , n234350 );
or ( n241642 , n241640 , n241641 );
nand ( n241643 , n227223 , n219440 );
nand ( n241644 , n241642 , n241643 );
not ( n241645 , n241644 );
or ( n241646 , n241639 , n241645 );
nand ( n241647 , n220507 , n241305 );
nand ( n241648 , n241646 , n241647 );
xor ( n241649 , n241638 , n241648 );
xor ( n241650 , n241649 , n241515 );
xor ( n241651 , n241628 , n241650 );
not ( n241652 , n220059 );
not ( n241653 , n241361 );
or ( n241654 , n241652 , n241653 );
not ( n241655 , n217616 );
not ( n241656 , n39366 );
or ( n241657 , n241655 , n241656 );
nand ( n241658 , n230273 , n234015 );
nand ( n241659 , n241657 , n241658 );
nand ( n241660 , n241659 , n220067 );
nand ( n241661 , n241654 , n241660 );
not ( n241662 , n218232 );
not ( n241663 , n218775 );
not ( n241664 , n236382 );
or ( n241665 , n241663 , n241664 );
nand ( n241666 , n39089 , n238352 );
nand ( n241667 , n241665 , n241666 );
not ( n241668 , n241667 );
or ( n241669 , n241662 , n241668 );
nand ( n241670 , n241373 , n219461 );
nand ( n241671 , n241669 , n241670 );
xor ( n241672 , n241661 , n241671 );
not ( n241673 , n227260 );
not ( n241674 , n241314 );
or ( n241675 , n241673 , n241674 );
nand ( n241676 , n223949 , n226655 );
nand ( n241677 , n241675 , n241676 );
xor ( n241678 , n241672 , n241677 );
xor ( n241679 , n241651 , n241678 );
xor ( n241680 , n241628 , n241650 );
and ( n241681 , n241680 , n241678 );
and ( n241682 , n241628 , n241650 );
or ( n241683 , n241681 , n241682 );
not ( n241684 , n239508 );
not ( n241685 , n241337 );
or ( n241686 , n241684 , n241685 );
not ( n241687 , n221241 );
not ( n241688 , n235516 );
or ( n241689 , n241687 , n241688 );
nand ( n241690 , n39747 , n238363 );
nand ( n241691 , n241689 , n241690 );
nand ( n241692 , n241691 , n218843 );
nand ( n241693 , n241686 , n241692 );
xor ( n241694 , n241191 , n241693 );
xor ( n241695 , n241694 , n241219 );
xor ( n241696 , n241695 , n241493 );
xor ( n241697 , n241696 , n241497 );
xor ( n241698 , n241695 , n241493 );
and ( n241699 , n241698 , n241497 );
and ( n241700 , n241695 , n241493 );
or ( n241701 , n241699 , n241700 );
xor ( n241702 , n241285 , n241279 );
xor ( n241703 , n241463 , n241473 );
xor ( n241704 , n241703 , n241477 );
xor ( n241705 , n241702 , n241704 );
xor ( n241706 , n241285 , n241279 );
and ( n241707 , n241706 , n241704 );
and ( n241708 , n241285 , n241279 );
or ( n241709 , n241707 , n241708 );
xor ( n241710 , n241381 , n241591 );
not ( n241711 , n227294 );
not ( n241712 , n236547 );
not ( n241713 , n241712 );
not ( n241714 , n222121 );
or ( n241715 , n241713 , n241714 );
nand ( n241716 , n226505 , n241404 );
nand ( n241717 , n241715 , n241716 );
not ( n241718 , n241717 );
or ( n241719 , n241711 , n241718 );
nand ( n241720 , n241406 , n235172 );
nand ( n241721 , n241719 , n241720 );
not ( n241722 , n224087 );
not ( n241723 , n241417 );
or ( n241724 , n241722 , n241723 );
not ( n241725 , n224096 );
not ( n241726 , n223786 );
or ( n241727 , n241725 , n241726 );
nand ( n241728 , n221956 , n238672 );
nand ( n241729 , n241727 , n241728 );
nand ( n241730 , n241729 , n227782 );
nand ( n241731 , n241724 , n241730 );
xor ( n241732 , n241721 , n241731 );
not ( n241733 , n240271 );
not ( n241734 , n241292 );
or ( n241735 , n241733 , n241734 );
not ( n241736 , n241287 );
not ( n241737 , n219742 );
or ( n241738 , n241736 , n241737 );
nand ( n241739 , n235359 , n235200 );
nand ( n241740 , n241738 , n241739 );
nand ( n241741 , n241740 , n240020 );
nand ( n241742 , n241735 , n241741 );
xor ( n241743 , n241732 , n241742 );
xor ( n241744 , n241489 , n241743 );
xor ( n241745 , n241744 , n241550 );
xor ( n241746 , n241710 , n241745 );
xor ( n241747 , n241381 , n241591 );
and ( n241748 , n241747 , n241745 );
and ( n241749 , n241381 , n241591 );
or ( n241750 , n241748 , n241749 );
xor ( n241751 , n241679 , n241389 );
xor ( n241752 , n241751 , n241697 );
xor ( n241753 , n241679 , n241389 );
and ( n241754 , n241753 , n241697 );
and ( n241755 , n241679 , n241389 );
or ( n241756 , n241754 , n241755 );
xor ( n241757 , n241705 , n241435 );
xor ( n241758 , n241757 , n241429 );
xor ( n241759 , n241705 , n241435 );
and ( n241760 , n241759 , n241429 );
and ( n241761 , n241705 , n241435 );
or ( n241762 , n241760 , n241761 );
xor ( n241763 , n241746 , n241441 );
xor ( n241764 , n241763 , n241752 );
xor ( n241765 , n241746 , n241441 );
and ( n241766 , n241765 , n241752 );
and ( n241767 , n241746 , n241441 );
or ( n241768 , n241766 , n241767 );
xor ( n241769 , n241758 , n241447 );
xor ( n241770 , n241769 , n241453 );
xor ( n241771 , n241758 , n241447 );
and ( n241772 , n241771 , n241453 );
and ( n241773 , n241758 , n241447 );
or ( n241774 , n241772 , n241773 );
xor ( n241775 , n241764 , n241770 );
xor ( n241776 , n241775 , n241459 );
xor ( n241777 , n241764 , n241770 );
and ( n241778 , n241777 , n241459 );
and ( n241779 , n241764 , n241770 );
or ( n241780 , n241778 , n241779 );
xor ( n241781 , n241565 , n241575 );
and ( n241782 , n241781 , n241589 );
and ( n241783 , n241565 , n241575 );
or ( n241784 , n241782 , n241783 );
xor ( n241785 , n241721 , n241731 );
and ( n241786 , n241785 , n241742 );
and ( n241787 , n241721 , n241731 );
or ( n241788 , n241786 , n241787 );
xor ( n241789 , n241606 , n241616 );
and ( n241790 , n241789 , n241627 );
and ( n241791 , n241606 , n241616 );
or ( n241792 , n241790 , n241791 );
xor ( n241793 , n241661 , n241671 );
and ( n241794 , n241793 , n241677 );
and ( n241795 , n241661 , n241671 );
or ( n241796 , n241794 , n241795 );
xor ( n241797 , n241191 , n241693 );
and ( n241798 , n241797 , n241219 );
and ( n241799 , n241191 , n241693 );
or ( n241800 , n241798 , n241799 );
xor ( n241801 , n241638 , n241648 );
and ( n241802 , n241801 , n241515 );
and ( n241803 , n241638 , n241648 );
or ( n241804 , n241802 , n241803 );
xor ( n241805 , n241463 , n241473 );
and ( n241806 , n241805 , n241477 );
and ( n241807 , n241463 , n241473 );
or ( n241808 , n241806 , n241807 );
xor ( n241809 , n241489 , n241743 );
and ( n241810 , n241809 , n241550 );
and ( n241811 , n241489 , n241743 );
or ( n241812 , n241810 , n241811 );
not ( n241813 , n236271 );
not ( n241814 , n240719 );
or ( n241815 , n241813 , n241814 );
nand ( n241816 , n241815 , n226655 );
not ( n241817 , n241586 );
not ( n241818 , n240120 );
or ( n241819 , n241817 , n241818 );
not ( n241820 , n238617 );
not ( n241821 , n41165 );
or ( n241822 , n241820 , n241821 );
not ( n241823 , n238199 );
nand ( n241824 , n241823 , n238619 );
nand ( n241825 , n241822 , n241824 );
nand ( n241826 , n228868 , n241825 );
nand ( n241827 , n241819 , n241826 );
xor ( n241828 , n241816 , n241827 );
or ( n241829 , n231474 , n241501 );
and ( n241830 , n237014 , n239001 );
and ( n241831 , n231480 , n231761 );
nor ( n241832 , n241830 , n241831 );
or ( n241833 , n231476 , n241832 );
nand ( n241834 , n241829 , n241833 );
xor ( n241835 , n241828 , n241834 );
xor ( n241836 , n241816 , n241827 );
and ( n241837 , n241836 , n241834 );
and ( n241838 , n241816 , n241827 );
or ( n241839 , n241837 , n241838 );
not ( n241840 , n241512 );
not ( n241841 , n233105 );
or ( n241842 , n241840 , n241841 );
and ( n241843 , n238218 , n231753 );
not ( n241844 , n238218 );
and ( n241845 , n241844 , n233885 );
or ( n241846 , n241843 , n241845 );
nand ( n241847 , n238274 , n241846 );
nand ( n241848 , n241842 , n241847 );
and ( n241849 , n239281 , n234751 );
xor ( n241850 , n241848 , n241849 );
not ( n241851 , n238240 );
not ( n241852 , n237816 );
not ( n241853 , n218884 );
or ( n241854 , n241852 , n241853 );
nand ( n241855 , n235908 , n234394 );
nand ( n241856 , n241854 , n241855 );
not ( n241857 , n241856 );
or ( n241858 , n241851 , n241857 );
nand ( n241859 , n237810 , n241527 );
nand ( n241860 , n241858 , n241859 );
xor ( n241861 , n241850 , n241860 );
xor ( n241862 , n241848 , n241849 );
and ( n241863 , n241862 , n241860 );
and ( n241864 , n241848 , n241849 );
or ( n241865 , n241863 , n241864 );
not ( n241866 , n227782 );
not ( n241867 , n239899 );
not ( n241868 , n40258 );
or ( n241869 , n241867 , n241868 );
nand ( n241870 , n221743 , n224095 );
nand ( n241871 , n241869 , n241870 );
not ( n241872 , n241871 );
or ( n241873 , n241866 , n241872 );
nand ( n241874 , n224087 , n241729 );
nand ( n241875 , n241873 , n241874 );
not ( n241876 , n237914 );
not ( n241877 , n230966 );
not ( n241878 , n241287 );
or ( n241879 , n241877 , n241878 );
nand ( n241880 , n239080 , n235200 );
nand ( n241881 , n241879 , n241880 );
not ( n241882 , n241881 );
or ( n241883 , n241876 , n241882 );
nand ( n241884 , n241740 , n239492 );
nand ( n241885 , n241883 , n241884 );
xor ( n241886 , n241875 , n241885 );
not ( n241887 , n228775 );
not ( n241888 , n229806 );
not ( n241889 , n234108 );
or ( n241890 , n241888 , n241889 );
not ( n241891 , n234108 );
nand ( n241892 , n232493 , n241891 );
nand ( n241893 , n241890 , n241892 );
not ( n241894 , n241893 );
or ( n241895 , n241887 , n241894 );
nand ( n241896 , n241604 , n232956 );
nand ( n241897 , n241895 , n241896 );
xor ( n241898 , n241886 , n241897 );
not ( n241899 , n235913 );
not ( n241900 , n241545 );
or ( n241901 , n241899 , n241900 );
not ( n241902 , n220906 );
not ( n241903 , n235921 );
or ( n241904 , n241902 , n241903 );
nand ( n241905 , n39997 , n238301 );
nand ( n241906 , n241904 , n241905 );
nand ( n241907 , n241906 , n220930 );
nand ( n241908 , n241901 , n241907 );
not ( n241909 , n227852 );
not ( n241910 , n226651 );
not ( n241911 , n237588 );
or ( n241912 , n241910 , n241911 );
nand ( n241913 , n236752 , n226650 );
nand ( n241914 , n241912 , n241913 );
not ( n241915 , n241914 );
or ( n241916 , n241909 , n241915 );
nand ( n241917 , n241534 , n237797 );
nand ( n241918 , n241916 , n241917 );
xor ( n241919 , n241908 , n241918 );
not ( n241920 , n221637 );
not ( n241921 , n222035 );
not ( n241922 , n237600 );
or ( n241923 , n241921 , n241922 );
nand ( n241924 , n239917 , n221778 );
nand ( n241925 , n241923 , n241924 );
not ( n241926 , n241925 );
or ( n241927 , n241920 , n241926 );
nand ( n241928 , n241563 , n221626 );
nand ( n241929 , n241927 , n241928 );
xor ( n241930 , n241919 , n241929 );
xor ( n241931 , n241898 , n241930 );
xor ( n241932 , n241931 , n241800 );
xor ( n241933 , n241898 , n241930 );
and ( n241934 , n241933 , n241800 );
and ( n241935 , n241898 , n241930 );
or ( n241936 , n241934 , n241935 );
not ( n241937 , n220881 );
not ( n241938 , n220151 );
not ( n241939 , n226724 );
or ( n241940 , n241938 , n241939 );
nand ( n241941 , n233018 , n220147 );
nand ( n241942 , n241940 , n241941 );
not ( n241943 , n241942 );
or ( n241944 , n241937 , n241943 );
nand ( n241945 , n241612 , n220492 );
nand ( n241946 , n241944 , n241945 );
not ( n241947 , n228237 );
not ( n241948 , n229387 );
not ( n241949 , n209964 );
not ( n241950 , n241949 );
or ( n241951 , n241948 , n241950 );
nand ( n241952 , n239185 , n227599 );
nand ( n241953 , n241951 , n241952 );
not ( n241954 , n241953 );
or ( n241955 , n241947 , n241954 );
nand ( n241956 , n241625 , n225478 );
nand ( n241957 , n241955 , n241956 );
xor ( n241958 , n241946 , n241957 );
not ( n241959 , n220067 );
not ( n241960 , n217616 );
not ( n241961 , n238486 );
or ( n241962 , n241960 , n241961 );
nand ( n241963 , n236840 , n231501 );
nand ( n241964 , n241962 , n241963 );
not ( n241965 , n241964 );
or ( n241966 , n241959 , n241965 );
nand ( n241967 , n241659 , n231018 );
nand ( n241968 , n241966 , n241967 );
xor ( n241969 , n241958 , n241968 );
xor ( n241970 , n241796 , n241969 );
not ( n241971 , n229964 );
not ( n241972 , n229261 );
not ( n241973 , n238449 );
or ( n241974 , n241972 , n241973 );
nand ( n241975 , n209710 , n234000 );
nand ( n241976 , n241974 , n241975 );
not ( n241977 , n241976 );
or ( n241978 , n241971 , n241977 );
nand ( n241979 , n241634 , n234006 );
nand ( n241980 , n241978 , n241979 );
not ( n241981 , n239530 );
not ( n241982 , n219800 );
not ( n241983 , n233856 );
not ( n241984 , n241983 );
or ( n241985 , n241982 , n241984 );
nand ( n241986 , n225795 , n219440 );
nand ( n241987 , n241985 , n241986 );
not ( n241988 , n241987 );
or ( n241989 , n241981 , n241988 );
nand ( n241990 , n241644 , n220507 );
nand ( n241991 , n241989 , n241990 );
xor ( n241992 , n241980 , n241991 );
xor ( n241993 , n241992 , n241835 );
xor ( n241994 , n241970 , n241993 );
xor ( n241995 , n241796 , n241969 );
and ( n241996 , n241995 , n241993 );
and ( n241997 , n241796 , n241969 );
or ( n241998 , n241996 , n241997 );
not ( n241999 , n219461 );
not ( n242000 , n241667 );
or ( n242001 , n241999 , n242000 );
not ( n242002 , n224497 );
not ( n242003 , n229704 );
or ( n242004 , n242002 , n242003 );
nand ( n242005 , n234792 , n218256 );
nand ( n242006 , n242004 , n242005 );
nand ( n242007 , n242006 , n218232 );
nand ( n242008 , n242001 , n242007 );
xor ( n242009 , n242008 , n241519 );
not ( n242010 , n218843 );
not ( n242011 , n221241 );
not ( n242012 , n232842 );
or ( n242013 , n242011 , n242012 );
nand ( n242014 , n39608 , n238363 );
nand ( n242015 , n242013 , n242014 );
not ( n242016 , n242015 );
or ( n242017 , n242010 , n242016 );
nand ( n242018 , n241691 , n239508 );
nand ( n242019 , n242017 , n242018 );
xor ( n242020 , n242009 , n242019 );
xor ( n242021 , n242020 , n241804 );
xor ( n242022 , n242021 , n241808 );
xor ( n242023 , n242020 , n241804 );
and ( n242024 , n242023 , n241808 );
and ( n242025 , n242020 , n241804 );
or ( n242026 , n242024 , n242025 );
xor ( n242027 , n241812 , n241595 );
xor ( n242028 , n241861 , n241554 );
xor ( n242029 , n242028 , n241784 );
xor ( n242030 , n242027 , n242029 );
xor ( n242031 , n241812 , n241595 );
and ( n242032 , n242031 , n242029 );
and ( n242033 , n241812 , n241595 );
or ( n242034 , n242032 , n242033 );
xor ( n242035 , n241683 , n241932 );
xor ( n242036 , n241788 , n241792 );
not ( n242037 , n237493 );
not ( n242038 , n222434 );
not ( n242039 , n227004 );
or ( n242040 , n242038 , n242039 );
nand ( n242041 , n238362 , n238719 );
nand ( n242042 , n242040 , n242041 );
not ( n242043 , n242042 );
or ( n242044 , n242037 , n242043 );
nand ( n242045 , n241573 , n237503 );
nand ( n242046 , n242044 , n242045 );
xor ( n242047 , n242046 , n241588 );
not ( n242048 , n227294 );
not ( n242049 , n239598 );
not ( n242050 , n221712 );
or ( n242051 , n242049 , n242050 );
not ( n242052 , n237005 );
nand ( n242053 , n242052 , n40182 );
nand ( n242054 , n242051 , n242053 );
not ( n242055 , n242054 );
or ( n242056 , n242048 , n242055 );
nand ( n242057 , n241717 , n235172 );
nand ( n242058 , n242056 , n242057 );
xor ( n242059 , n242047 , n242058 );
xor ( n242060 , n242036 , n242059 );
xor ( n242061 , n242035 , n242060 );
xor ( n242062 , n241683 , n241932 );
and ( n242063 , n242062 , n242060 );
and ( n242064 , n241683 , n241932 );
or ( n242065 , n242063 , n242064 );
xor ( n242066 , n242022 , n241994 );
xor ( n242067 , n242066 , n241709 );
xor ( n242068 , n242022 , n241994 );
and ( n242069 , n242068 , n241709 );
and ( n242070 , n242022 , n241994 );
or ( n242071 , n242069 , n242070 );
xor ( n242072 , n241701 , n242030 );
xor ( n242073 , n242072 , n241750 );
xor ( n242074 , n241701 , n242030 );
and ( n242075 , n242074 , n241750 );
and ( n242076 , n241701 , n242030 );
or ( n242077 , n242075 , n242076 );
xor ( n242078 , n242061 , n241756 );
xor ( n242079 , n242078 , n242067 );
xor ( n242080 , n242061 , n241756 );
and ( n242081 , n242080 , n242067 );
and ( n242082 , n242061 , n241756 );
or ( n242083 , n242081 , n242082 );
xor ( n242084 , n241762 , n242073 );
xor ( n242085 , n242084 , n242079 );
xor ( n242086 , n241762 , n242073 );
and ( n242087 , n242086 , n242079 );
and ( n242088 , n241762 , n242073 );
or ( n242089 , n242087 , n242088 );
xor ( n242090 , n241768 , n242085 );
xor ( n242091 , n242090 , n241774 );
xor ( n242092 , n241768 , n242085 );
and ( n242093 , n242092 , n241774 );
and ( n242094 , n241768 , n242085 );
or ( n242095 , n242093 , n242094 );
xor ( n242096 , n241908 , n241918 );
and ( n242097 , n242096 , n241929 );
and ( n242098 , n241908 , n241918 );
or ( n242099 , n242097 , n242098 );
xor ( n242100 , n242046 , n241588 );
and ( n242101 , n242100 , n242058 );
and ( n242102 , n242046 , n241588 );
or ( n242103 , n242101 , n242102 );
xor ( n242104 , n241875 , n241885 );
and ( n242105 , n242104 , n241897 );
and ( n242106 , n241875 , n241885 );
or ( n242107 , n242105 , n242106 );
xor ( n242108 , n241946 , n241957 );
and ( n242109 , n242108 , n241968 );
and ( n242110 , n241946 , n241957 );
or ( n242111 , n242109 , n242110 );
xor ( n242112 , n242008 , n241519 );
and ( n242113 , n242112 , n242019 );
and ( n242114 , n242008 , n241519 );
or ( n242115 , n242113 , n242114 );
xor ( n242116 , n241980 , n241991 );
and ( n242117 , n242116 , n241835 );
and ( n242118 , n241980 , n241991 );
or ( n242119 , n242117 , n242118 );
xor ( n242120 , n241861 , n241554 );
and ( n242121 , n242120 , n241784 );
and ( n242122 , n241861 , n241554 );
or ( n242123 , n242121 , n242122 );
xor ( n242124 , n241788 , n241792 );
and ( n242125 , n242124 , n242059 );
and ( n242126 , n241788 , n241792 );
or ( n242127 , n242125 , n242126 );
not ( n242128 , n241846 );
not ( n242129 , n233105 );
or ( n242130 , n242128 , n242129 );
xor ( n242131 , n216859 , n234382 );
nand ( n242132 , n238274 , n242131 );
nand ( n242133 , n242130 , n242132 );
and ( n242134 , n231754 , n41321 );
xor ( n242135 , n242133 , n242134 );
not ( n242136 , n228868 );
and ( n242137 , n238671 , n238617 );
not ( n242138 , n238671 );
and ( n242139 , n242138 , n238619 );
or ( n242140 , n242137 , n242139 );
not ( n242141 , n242140 );
or ( n242142 , n242136 , n242141 );
nand ( n242143 , n239794 , n241825 );
nand ( n242144 , n242142 , n242143 );
xor ( n242145 , n242135 , n242144 );
xor ( n242146 , n242133 , n242134 );
and ( n242147 , n242146 , n242144 );
and ( n242148 , n242133 , n242134 );
or ( n242149 , n242147 , n242148 );
not ( n242150 , n238240 );
not ( n242151 , n236188 );
not ( n242152 , n219235 );
or ( n242153 , n242151 , n242152 );
nand ( n242154 , n220568 , n239787 );
nand ( n242155 , n242153 , n242154 );
not ( n242156 , n242155 );
or ( n242157 , n242150 , n242156 );
not ( n242158 , n228270 );
nand ( n242159 , n242158 , n241856 );
nand ( n242160 , n242157 , n242159 );
not ( n242161 , n221626 );
not ( n242162 , n241925 );
or ( n242163 , n242161 , n242162 );
not ( n242164 , n237937 );
not ( n242165 , n230490 );
or ( n242166 , n242164 , n242165 );
nand ( n242167 , n240279 , n221778 );
nand ( n242168 , n242166 , n242167 );
nand ( n242169 , n242168 , n221637 );
nand ( n242170 , n242163 , n242169 );
xor ( n242171 , n242160 , n242170 );
not ( n242172 , n222454 );
not ( n242173 , n242042 );
or ( n242174 , n242172 , n242173 );
not ( n242175 , n240229 );
not ( n242176 , n223717 );
or ( n242177 , n242175 , n242176 );
nand ( n242178 , n239527 , n238719 );
nand ( n242179 , n242177 , n242178 );
nand ( n242180 , n242179 , n237493 );
nand ( n242181 , n242174 , n242180 );
xor ( n242182 , n242171 , n242181 );
xor ( n242183 , n242160 , n242170 );
and ( n242184 , n242183 , n242181 );
and ( n242185 , n242160 , n242170 );
or ( n242186 , n242184 , n242185 );
not ( n242187 , n219076 );
not ( n242188 , n240917 );
not ( n242189 , n230241 );
or ( n242190 , n242188 , n242189 );
nand ( n242191 , n238877 , n219797 );
nand ( n242192 , n242190 , n242191 );
not ( n242193 , n242192 );
or ( n242194 , n242187 , n242193 );
nand ( n242195 , n241987 , n220507 );
nand ( n242196 , n242194 , n242195 );
not ( n242197 , n220067 );
not ( n242198 , n231500 );
not ( n242199 , n237271 );
or ( n242200 , n242198 , n242199 );
nand ( n242201 , n240308 , n231501 );
nand ( n242202 , n242200 , n242201 );
not ( n242203 , n242202 );
or ( n242204 , n242197 , n242203 );
nand ( n242205 , n241964 , n231018 );
nand ( n242206 , n242204 , n242205 );
xor ( n242207 , n242196 , n242206 );
not ( n242208 , n219779 );
not ( n242209 , n236768 );
not ( n242210 , n227223 );
not ( n242211 , n242210 );
or ( n242212 , n242209 , n242211 );
nand ( n242213 , n238819 , n222414 );
nand ( n242214 , n242212 , n242213 );
not ( n242215 , n242214 );
or ( n242216 , n242208 , n242215 );
nand ( n242217 , n241942 , n220164 );
nand ( n242218 , n242216 , n242217 );
xor ( n242219 , n242207 , n242218 );
xor ( n242220 , n242115 , n242219 );
xor ( n242221 , n242220 , n242119 );
xor ( n242222 , n242115 , n242219 );
and ( n242223 , n242222 , n242119 );
and ( n242224 , n242115 , n242219 );
or ( n242225 , n242223 , n242224 );
not ( n242226 , n218843 );
not ( n242227 , n221241 );
not ( n242228 , n227201 );
or ( n242229 , n242227 , n242228 );
nand ( n242230 , n39089 , n238363 );
nand ( n242231 , n242229 , n242230 );
not ( n242232 , n242231 );
or ( n242233 , n242226 , n242232 );
nand ( n242234 , n223665 , n242015 );
nand ( n242235 , n242233 , n242234 );
not ( n242236 , n229395 );
not ( n242237 , n241953 );
or ( n242238 , n242236 , n242237 );
nand ( n242239 , n219501 , n229387 );
nand ( n242240 , n242238 , n242239 );
xor ( n242241 , n242235 , n242240 );
xor ( n242242 , n242241 , n241839 );
not ( n242243 , n221674 );
not ( n242244 , n220906 );
not ( n242245 , n238728 );
or ( n242246 , n242244 , n242245 );
not ( n242247 , n235452 );
nand ( n242248 , n242247 , n239066 );
nand ( n242249 , n242246 , n242248 );
not ( n242250 , n242249 );
or ( n242251 , n242243 , n242250 );
nand ( n242252 , n241906 , n235913 );
nand ( n242253 , n242251 , n242252 );
not ( n242254 , n229964 );
not ( n242255 , n229261 );
not ( n242256 , n239617 );
or ( n242257 , n242255 , n242256 );
nand ( n242258 , n233614 , n234000 );
nand ( n242259 , n242257 , n242258 );
not ( n242260 , n242259 );
or ( n242261 , n242254 , n242260 );
nand ( n242262 , n241976 , n234006 );
nand ( n242263 , n242261 , n242262 );
xor ( n242264 , n242253 , n242263 );
not ( n242265 , n218232 );
not ( n242266 , n233083 );
not ( n242267 , n39366 );
or ( n242268 , n242266 , n242267 );
nand ( n242269 , n39365 , n238352 );
nand ( n242270 , n242268 , n242269 );
not ( n242271 , n242270 );
or ( n242272 , n242265 , n242271 );
nand ( n242273 , n242006 , n219461 );
nand ( n242274 , n242272 , n242273 );
xor ( n242275 , n242264 , n242274 );
xor ( n242276 , n242242 , n242275 );
xor ( n242277 , n242276 , n242123 );
xor ( n242278 , n242242 , n242275 );
and ( n242279 , n242278 , n242123 );
and ( n242280 , n242242 , n242275 );
or ( n242281 , n242279 , n242280 );
xor ( n242282 , n242103 , n242107 );
not ( n242283 , n242054 );
not ( n242284 , n238409 );
or ( n242285 , n242283 , n242284 );
not ( n242286 , n239598 );
not ( n242287 , n224700 );
or ( n242288 , n242286 , n242287 );
nand ( n242289 , n236300 , n241404 );
nand ( n242290 , n242288 , n242289 );
nand ( n242291 , n242290 , n227294 );
nand ( n242292 , n242285 , n242291 );
not ( n242293 , n231474 );
not ( n242294 , n241832 );
and ( n242295 , n242293 , n242294 );
and ( n242296 , n231480 , n238640 );
not ( n242297 , n231480 );
and ( n242298 , n242297 , n219201 );
or ( n242299 , n242296 , n242298 );
not ( n242300 , n242299 );
nor ( n242301 , n242300 , n237013 );
nor ( n242302 , n242295 , n242301 );
xor ( n242303 , n242292 , n242302 );
not ( n242304 , n224087 );
not ( n242305 , n241871 );
or ( n242306 , n242304 , n242305 );
not ( n242307 , n237130 );
not ( n242308 , n238786 );
or ( n242309 , n242307 , n242308 );
nand ( n242310 , n230514 , n224095 );
nand ( n242311 , n242309 , n242310 );
nand ( n242312 , n242311 , n227782 );
nand ( n242313 , n242306 , n242312 );
xor ( n242314 , n242303 , n242313 );
xor ( n242315 , n242282 , n242314 );
xor ( n242316 , n242315 , n241936 );
xor ( n242317 , n242316 , n242127 );
xor ( n242318 , n242315 , n241936 );
and ( n242319 , n242318 , n242127 );
and ( n242320 , n242315 , n241936 );
or ( n242321 , n242319 , n242320 );
xor ( n242322 , n242145 , n241865 );
xor ( n242323 , n242322 , n242099 );
xor ( n242324 , n242323 , n241998 );
not ( n242325 , n240271 );
not ( n242326 , n241881 );
or ( n242327 , n242325 , n242326 );
not ( n242328 , n234878 );
not ( n242329 , n220599 );
or ( n242330 , n242328 , n242329 );
nand ( n242331 , n221956 , n240617 );
nand ( n242332 , n242330 , n242331 );
nand ( n242333 , n242332 , n237914 );
nand ( n242334 , n242327 , n242333 );
buf ( n242335 , n232956 );
not ( n242336 , n242335 );
not ( n242337 , n241893 );
or ( n242338 , n242336 , n242337 );
not ( n242339 , n232494 );
not ( n242340 , n40660 );
or ( n242341 , n242339 , n242340 );
nand ( n242342 , n239470 , n232493 );
nand ( n242343 , n242341 , n242342 );
nand ( n242344 , n242343 , n238776 );
nand ( n242345 , n242338 , n242344 );
xor ( n242346 , n242334 , n242345 );
not ( n242347 , n237797 );
not ( n242348 , n241914 );
or ( n242349 , n242347 , n242348 );
and ( n242350 , n239774 , n219223 );
not ( n242351 , n239774 );
and ( n242352 , n242351 , n219226 );
or ( n242353 , n242350 , n242352 );
nand ( n242354 , n242353 , n227852 );
nand ( n242355 , n242349 , n242354 );
xor ( n242356 , n242346 , n242355 );
xor ( n242357 , n242356 , n242182 );
xor ( n242358 , n242357 , n242111 );
xor ( n242359 , n242324 , n242358 );
xor ( n242360 , n242323 , n241998 );
and ( n242361 , n242360 , n242358 );
and ( n242362 , n242323 , n241998 );
or ( n242363 , n242361 , n242362 );
xor ( n242364 , n242277 , n242221 );
xor ( n242365 , n242364 , n242026 );
xor ( n242366 , n242277 , n242221 );
and ( n242367 , n242366 , n242026 );
and ( n242368 , n242277 , n242221 );
or ( n242369 , n242367 , n242368 );
xor ( n242370 , n242034 , n242065 );
xor ( n242371 , n242370 , n242317 );
xor ( n242372 , n242034 , n242065 );
and ( n242373 , n242372 , n242317 );
and ( n242374 , n242034 , n242065 );
or ( n242375 , n242373 , n242374 );
xor ( n242376 , n242359 , n242071 );
xor ( n242377 , n242376 , n242365 );
xor ( n242378 , n242359 , n242071 );
and ( n242379 , n242378 , n242365 );
and ( n242380 , n242359 , n242071 );
or ( n242381 , n242379 , n242380 );
xor ( n242382 , n242077 , n242371 );
xor ( n242383 , n242382 , n242083 );
xor ( n242384 , n242077 , n242371 );
and ( n242385 , n242384 , n242083 );
and ( n242386 , n242077 , n242371 );
or ( n242387 , n242385 , n242386 );
xor ( n242388 , n242377 , n242383 );
xor ( n242389 , n242388 , n242089 );
xor ( n242390 , n242377 , n242383 );
and ( n242391 , n242390 , n242089 );
and ( n242392 , n242377 , n242383 );
or ( n242393 , n242391 , n242392 );
xor ( n242394 , n242292 , n242302 );
and ( n242395 , n242394 , n242313 );
and ( n242396 , n242292 , n242302 );
or ( n242397 , n242395 , n242396 );
xor ( n242398 , n242334 , n242345 );
and ( n242399 , n242398 , n242355 );
and ( n242400 , n242334 , n242345 );
or ( n242401 , n242399 , n242400 );
xor ( n242402 , n242253 , n242263 );
and ( n242403 , n242402 , n242274 );
and ( n242404 , n242253 , n242263 );
or ( n242405 , n242403 , n242404 );
xor ( n242406 , n242235 , n242240 );
and ( n242407 , n242406 , n241839 );
and ( n242408 , n242235 , n242240 );
or ( n242409 , n242407 , n242408 );
xor ( n242410 , n242196 , n242206 );
and ( n242411 , n242410 , n242218 );
and ( n242412 , n242196 , n242206 );
or ( n242413 , n242411 , n242412 );
xor ( n242414 , n242145 , n241865 );
and ( n242415 , n242414 , n242099 );
and ( n242416 , n242145 , n241865 );
or ( n242417 , n242415 , n242416 );
xor ( n242418 , n242103 , n242107 );
and ( n242419 , n242418 , n242314 );
and ( n242420 , n242103 , n242107 );
or ( n242421 , n242419 , n242420 );
xor ( n242422 , n242356 , n242182 );
and ( n242423 , n242422 , n242111 );
and ( n242424 , n242356 , n242182 );
or ( n242425 , n242423 , n242424 );
not ( n242426 , n227121 );
not ( n242427 , n225477 );
or ( n242428 , n242426 , n242427 );
nand ( n242429 , n242428 , n229387 );
not ( n242430 , n242299 );
not ( n242431 , n234371 );
or ( n242432 , n242430 , n242431 );
not ( n242433 , n237014 );
not ( n242434 , n238199 );
or ( n242435 , n242433 , n242434 );
not ( n242436 , n219389 );
nand ( n242437 , n242436 , n231480 );
nand ( n242438 , n242435 , n242437 );
nand ( n242439 , n234378 , n242438 );
nand ( n242440 , n242432 , n242439 );
xor ( n242441 , n242429 , n242440 );
not ( n242442 , n242131 );
or ( n242443 , n239269 , n242442 );
and ( n242444 , n231753 , n239001 );
and ( n242445 , n239281 , n231761 );
nor ( n242446 , n242444 , n242445 );
or ( n242447 , n242446 , n238275 );
nand ( n242448 , n242443 , n242447 );
xor ( n242449 , n242441 , n242448 );
xor ( n242450 , n242429 , n242440 );
and ( n242451 , n242450 , n242448 );
and ( n242452 , n242429 , n242440 );
or ( n242453 , n242451 , n242452 );
and ( n242454 , n239281 , n41250 );
not ( n242455 , n228868 );
not ( n242456 , n238619 );
not ( n242457 , n237496 );
or ( n242458 , n242456 , n242457 );
nand ( n242459 , n235908 , n236643 );
nand ( n242460 , n242458 , n242459 );
not ( n242461 , n242460 );
or ( n242462 , n242455 , n242461 );
not ( n242463 , n237038 );
nand ( n242464 , n242463 , n242140 );
nand ( n242465 , n242462 , n242464 );
xor ( n242466 , n242454 , n242465 );
not ( n242467 , n221626 );
not ( n242468 , n242168 );
or ( n242469 , n242467 , n242468 );
not ( n242470 , n238705 );
buf ( n242471 , n235012 );
not ( n242472 , n242471 );
not ( n242473 , n242472 );
or ( n242474 , n242470 , n242473 );
nand ( n242475 , n229928 , n221778 );
nand ( n242476 , n242474 , n242475 );
nand ( n242477 , n242476 , n221637 );
nand ( n242478 , n242469 , n242477 );
xor ( n242479 , n242466 , n242478 );
xor ( n242480 , n242454 , n242465 );
and ( n242481 , n242480 , n242478 );
and ( n242482 , n242454 , n242465 );
or ( n242483 , n242481 , n242482 );
xor ( n242484 , n242405 , n242413 );
not ( n242485 , n228775 );
and ( n242486 , n233962 , n239077 );
not ( n242487 , n233962 );
and ( n242488 , n242487 , n226922 );
nor ( n242489 , n242486 , n242488 );
not ( n242490 , n242489 );
or ( n242491 , n242485 , n242490 );
nand ( n242492 , n242343 , n242335 );
nand ( n242493 , n242491 , n242492 );
not ( n242494 , n242353 );
not ( n242495 , n237797 );
or ( n242496 , n242494 , n242495 );
not ( n242497 , n239774 );
not ( n242498 , n234108 );
or ( n242499 , n242497 , n242498 );
nand ( n242500 , n241891 , n234293 );
nand ( n242501 , n242499 , n242500 );
nand ( n242502 , n242501 , n227852 );
nand ( n242503 , n242496 , n242502 );
xor ( n242504 , n242493 , n242503 );
not ( n242505 , n235913 );
not ( n242506 , n242249 );
or ( n242507 , n242505 , n242506 );
not ( n242508 , n222399 );
not ( n242509 , n39927 );
or ( n242510 , n242508 , n242509 );
nand ( n242511 , n239173 , n239548 );
nand ( n242512 , n242510 , n242511 );
nand ( n242513 , n242512 , n220930 );
nand ( n242514 , n242507 , n242513 );
xor ( n242515 , n242504 , n242514 );
xor ( n242516 , n242484 , n242515 );
xor ( n242517 , n242405 , n242413 );
and ( n242518 , n242517 , n242515 );
and ( n242519 , n242405 , n242413 );
or ( n242520 , n242518 , n242519 );
not ( n242521 , n219076 );
not ( n242522 , n240917 );
not ( n242523 , n240710 );
or ( n242524 , n242522 , n242523 );
nand ( n242525 , n235977 , n219797 );
nand ( n242526 , n242524 , n242525 );
not ( n242527 , n242526 );
or ( n242528 , n242521 , n242527 );
nand ( n242529 , n242192 , n220507 );
nand ( n242530 , n242528 , n242529 );
not ( n242531 , n231018 );
not ( n242532 , n242202 );
or ( n242533 , n242531 , n242532 );
not ( n242534 , n217616 );
not ( n242535 , n209709 );
or ( n242536 , n242534 , n242535 );
nand ( n242537 , n235691 , n234015 );
nand ( n242538 , n242536 , n242537 );
nand ( n242539 , n242538 , n220067 );
nand ( n242540 , n242533 , n242539 );
xor ( n242541 , n242530 , n242540 );
not ( n242542 , n220881 );
not ( n242543 , n236768 );
not ( n242544 , n240738 );
or ( n242545 , n242543 , n242544 );
nand ( n242546 , n227696 , n222414 );
nand ( n242547 , n242545 , n242546 );
not ( n242548 , n242547 );
or ( n242549 , n242542 , n242548 );
nand ( n242550 , n242214 , n220164 );
nand ( n242551 , n242549 , n242550 );
xor ( n242552 , n242541 , n242551 );
not ( n242553 , n229964 );
not ( n242554 , n229261 );
not ( n242555 , n241949 );
or ( n242556 , n242554 , n242555 );
nand ( n242557 , n239185 , n234000 );
nand ( n242558 , n242556 , n242557 );
not ( n242559 , n242558 );
or ( n242560 , n242553 , n242559 );
nand ( n242561 , n242259 , n234006 );
nand ( n242562 , n242560 , n242561 );
not ( n242563 , n219461 );
not ( n242564 , n242270 );
or ( n242565 , n242563 , n242564 );
not ( n242566 , n233083 );
not ( n242567 , n39287 );
or ( n242568 , n242566 , n242567 );
nand ( n242569 , n236840 , n238352 );
nand ( n242570 , n242568 , n242569 );
nand ( n242571 , n242570 , n218232 );
nand ( n242572 , n242565 , n242571 );
xor ( n242573 , n242562 , n242572 );
not ( n242574 , n239508 );
not ( n242575 , n242231 );
or ( n242576 , n242574 , n242575 );
not ( n242577 , n221241 );
not ( n242578 , n229704 );
or ( n242579 , n242577 , n242578 );
nand ( n242580 , n38532 , n238363 );
nand ( n242581 , n242579 , n242580 );
nand ( n242582 , n242581 , n218843 );
nand ( n242583 , n242576 , n242582 );
xor ( n242584 , n242573 , n242583 );
xor ( n242585 , n242552 , n242584 );
xor ( n242586 , n242585 , n242417 );
xor ( n242587 , n242552 , n242584 );
and ( n242588 , n242587 , n242417 );
and ( n242589 , n242552 , n242584 );
or ( n242590 , n242588 , n242589 );
xor ( n242591 , n242449 , n242149 );
xor ( n242592 , n242591 , n242186 );
xor ( n242593 , n242592 , n242425 );
xor ( n242594 , n242397 , n242401 );
not ( n242595 , n238240 );
not ( n242596 , n239787 );
not ( n242597 , n242596 );
not ( n242598 , n237588 );
or ( n242599 , n242597 , n242598 );
nand ( n242600 , n236752 , n239787 );
nand ( n242601 , n242599 , n242600 );
not ( n242602 , n242601 );
or ( n242603 , n242595 , n242602 );
nand ( n242604 , n242155 , n233446 );
nand ( n242605 , n242603 , n242604 );
not ( n242606 , n237493 );
not ( n242607 , n222430 );
not ( n242608 , n237600 );
or ( n242609 , n242607 , n242608 );
nand ( n242610 , n239917 , n238719 );
nand ( n242611 , n242609 , n242610 );
not ( n242612 , n242611 );
or ( n242613 , n242606 , n242612 );
nand ( n242614 , n242179 , n222454 );
nand ( n242615 , n242613 , n242614 );
xor ( n242616 , n242605 , n242615 );
not ( n242617 , n242302 );
xor ( n242618 , n242616 , n242617 );
xor ( n242619 , n242594 , n242618 );
xor ( n242620 , n242593 , n242619 );
xor ( n242621 , n242592 , n242425 );
and ( n242622 , n242621 , n242619 );
and ( n242623 , n242592 , n242425 );
or ( n242624 , n242622 , n242623 );
xor ( n242625 , n242421 , n242225 );
xor ( n242626 , n242625 , n242516 );
xor ( n242627 , n242421 , n242225 );
and ( n242628 , n242627 , n242516 );
and ( n242629 , n242421 , n242225 );
or ( n242630 , n242628 , n242629 );
not ( n242631 , n227294 );
not ( n242632 , n241712 );
not ( n242633 , n240637 );
or ( n242634 , n242632 , n242633 );
nand ( n242635 , n40415 , n239599 );
nand ( n242636 , n242634 , n242635 );
not ( n242637 , n242636 );
or ( n242638 , n242631 , n242637 );
nand ( n242639 , n242290 , n235172 );
nand ( n242640 , n242638 , n242639 );
not ( n242641 , n227782 );
not ( n242642 , n237130 );
not ( n242643 , n221712 );
or ( n242644 , n242642 , n242643 );
nand ( n242645 , n236719 , n237129 );
nand ( n242646 , n242644 , n242645 );
not ( n242647 , n242646 );
or ( n242648 , n242641 , n242647 );
nand ( n242649 , n242311 , n224087 );
nand ( n242650 , n242648 , n242649 );
xor ( n242651 , n242640 , n242650 );
not ( n242652 , n240020 );
not ( n242653 , n234273 );
not ( n242654 , n242653 );
not ( n242655 , n220971 );
or ( n242656 , n242654 , n242655 );
nand ( n242657 , n226911 , n240617 );
nand ( n242658 , n242656 , n242657 );
not ( n242659 , n242658 );
or ( n242660 , n242652 , n242659 );
nand ( n242661 , n240271 , n242332 );
nand ( n242662 , n242660 , n242661 );
xor ( n242663 , n242651 , n242662 );
xor ( n242664 , n242663 , n242479 );
xor ( n242665 , n242664 , n242409 );
xor ( n242666 , n242665 , n242586 );
xor ( n242667 , n242666 , n242281 );
xor ( n242668 , n242665 , n242586 );
and ( n242669 , n242668 , n242281 );
and ( n242670 , n242665 , n242586 );
or ( n242671 , n242669 , n242670 );
xor ( n242672 , n242321 , n242620 );
xor ( n242673 , n242672 , n242363 );
xor ( n242674 , n242321 , n242620 );
and ( n242675 , n242674 , n242363 );
and ( n242676 , n242321 , n242620 );
or ( n242677 , n242675 , n242676 );
xor ( n242678 , n242626 , n242369 );
xor ( n242679 , n242678 , n242667 );
xor ( n242680 , n242626 , n242369 );
and ( n242681 , n242680 , n242667 );
and ( n242682 , n242626 , n242369 );
or ( n242683 , n242681 , n242682 );
xor ( n242684 , n242375 , n242673 );
xor ( n242685 , n242684 , n242381 );
xor ( n242686 , n242375 , n242673 );
and ( n242687 , n242686 , n242381 );
and ( n242688 , n242375 , n242673 );
or ( n242689 , n242687 , n242688 );
xor ( n242690 , n242679 , n242685 );
xor ( n242691 , n242690 , n242387 );
xor ( n242692 , n242679 , n242685 );
and ( n242693 , n242692 , n242387 );
and ( n242694 , n242679 , n242685 );
or ( n242695 , n242693 , n242694 );
xor ( n242696 , n242605 , n242615 );
and ( n242697 , n242696 , n242617 );
and ( n242698 , n242605 , n242615 );
or ( n242699 , n242697 , n242698 );
xor ( n242700 , n242640 , n242650 );
and ( n242701 , n242700 , n242662 );
and ( n242702 , n242640 , n242650 );
or ( n242703 , n242701 , n242702 );
xor ( n242704 , n242493 , n242503 );
and ( n242705 , n242704 , n242514 );
and ( n242706 , n242493 , n242503 );
or ( n242707 , n242705 , n242706 );
xor ( n242708 , n242562 , n242572 );
and ( n242709 , n242708 , n242583 );
and ( n242710 , n242562 , n242572 );
or ( n242711 , n242709 , n242710 );
xor ( n242712 , n242530 , n242540 );
and ( n242713 , n242712 , n242551 );
and ( n242714 , n242530 , n242540 );
or ( n242715 , n242713 , n242714 );
xor ( n242716 , n242449 , n242149 );
and ( n242717 , n242716 , n242186 );
and ( n242718 , n242449 , n242149 );
or ( n242719 , n242717 , n242718 );
xor ( n242720 , n242397 , n242401 );
and ( n242721 , n242720 , n242618 );
and ( n242722 , n242397 , n242401 );
or ( n242723 , n242721 , n242722 );
xor ( n242724 , n242663 , n242479 );
and ( n242725 , n242724 , n242409 );
and ( n242726 , n242663 , n242479 );
or ( n242727 , n242725 , n242726 );
and ( n242728 , n216859 , n234382 );
not ( n242729 , n242438 );
not ( n242730 , n234371 );
or ( n242731 , n242729 , n242730 );
not ( n242732 , n239393 );
not ( n242733 , n217964 );
or ( n242734 , n242732 , n242733 );
nand ( n242735 , n238671 , n237014 );
nand ( n242736 , n242734 , n242735 );
buf ( n242737 , n234378 );
nand ( n242738 , n242736 , n242737 );
nand ( n242739 , n242731 , n242738 );
xor ( n242740 , n242728 , n242739 );
not ( n242741 , n230721 );
not ( n242742 , n242446 );
and ( n242743 , n242741 , n242742 );
not ( n242744 , n238641 );
not ( n242745 , n231753 );
or ( n242746 , n242744 , n242745 );
nand ( n242747 , n234382 , n41070 );
nand ( n242748 , n242746 , n242747 );
not ( n242749 , n242748 );
nor ( n242750 , n242749 , n238275 );
nor ( n242751 , n242743 , n242750 );
xor ( n242752 , n242740 , n242751 );
xor ( n242753 , n242728 , n242739 );
and ( n242754 , n242753 , n242751 );
and ( n242755 , n242728 , n242739 );
or ( n242756 , n242754 , n242755 );
not ( n242757 , n228868 );
not ( n242758 , n228850 );
not ( n242759 , n219235 );
or ( n242760 , n242758 , n242759 );
nand ( n242761 , n220568 , n236643 );
nand ( n242762 , n242760 , n242761 );
not ( n242763 , n242762 );
or ( n242764 , n242757 , n242763 );
nand ( n242765 , n242460 , n240120 );
nand ( n242766 , n242764 , n242765 );
not ( n242767 , n237503 );
not ( n242768 , n242611 );
or ( n242769 , n242767 , n242768 );
not ( n242770 , n222430 );
not ( n242771 , n230490 );
or ( n242772 , n242770 , n242771 );
nand ( n242773 , n237963 , n238719 );
nand ( n242774 , n242772 , n242773 );
nand ( n242775 , n242774 , n237493 );
nand ( n242776 , n242769 , n242775 );
xor ( n242777 , n242766 , n242776 );
not ( n242778 , n235172 );
not ( n242779 , n242636 );
or ( n242780 , n242778 , n242779 );
not ( n242781 , n241712 );
not ( n242782 , n237971 );
or ( n242783 , n242781 , n242782 );
nand ( n242784 , n239527 , n223156 );
nand ( n242785 , n242783 , n242784 );
nand ( n242786 , n242785 , n227294 );
nand ( n242787 , n242780 , n242786 );
xor ( n242788 , n242777 , n242787 );
xor ( n242789 , n242766 , n242776 );
and ( n242790 , n242789 , n242787 );
and ( n242791 , n242766 , n242776 );
or ( n242792 , n242790 , n242791 );
not ( n242793 , n234006 );
not ( n242794 , n242558 );
or ( n242795 , n242793 , n242794 );
nand ( n242796 , n229964 , n229261 );
nand ( n242797 , n242795 , n242796 );
xor ( n242798 , n242453 , n242797 );
not ( n242799 , n219779 );
and ( n242800 , n220151 , n238877 );
not ( n242801 , n220151 );
and ( n242802 , n242801 , n235516 );
nor ( n242803 , n242800 , n242802 );
not ( n242804 , n242803 );
or ( n242805 , n242799 , n242804 );
nand ( n242806 , n242547 , n220164 );
nand ( n242807 , n242805 , n242806 );
xor ( n242808 , n242798 , n242807 );
not ( n242809 , n231018 );
not ( n242810 , n242538 );
or ( n242811 , n242809 , n242810 );
not ( n242812 , n217616 );
not ( n242813 , n234579 );
or ( n242814 , n242812 , n242813 );
nand ( n242815 , n240358 , n231501 );
nand ( n242816 , n242814 , n242815 );
nand ( n242817 , n242816 , n220067 );
nand ( n242818 , n242811 , n242817 );
not ( n242819 , n239508 );
not ( n242820 , n242581 );
or ( n242821 , n242819 , n242820 );
not ( n242822 , n221241 );
not ( n242823 , n228165 );
or ( n242824 , n242822 , n242823 );
nand ( n242825 , n237229 , n238363 );
nand ( n242826 , n242824 , n242825 );
nand ( n242827 , n242826 , n218843 );
nand ( n242828 , n242821 , n242827 );
xor ( n242829 , n242818 , n242828 );
not ( n242830 , n239530 );
not ( n242831 , n240917 );
not ( n242832 , n227201 );
or ( n242833 , n242831 , n242832 );
nand ( n242834 , n39089 , n219420 );
nand ( n242835 , n242833 , n242834 );
not ( n242836 , n242835 );
or ( n242837 , n242830 , n242836 );
nand ( n242838 , n242526 , n220507 );
nand ( n242839 , n242837 , n242838 );
xor ( n242840 , n242829 , n242839 );
xor ( n242841 , n242808 , n242840 );
not ( n242842 , n219461 );
not ( n242843 , n242570 );
or ( n242844 , n242842 , n242843 );
not ( n242845 , n224497 );
not ( n242846 , n239562 );
or ( n242847 , n242845 , n242846 );
nand ( n242848 , n238887 , n238352 );
nand ( n242849 , n242847 , n242848 );
nand ( n242850 , n242849 , n218232 );
nand ( n242851 , n242844 , n242850 );
not ( n242852 , n235913 );
not ( n242853 , n242512 );
or ( n242854 , n242852 , n242853 );
not ( n242855 , n222399 );
not ( n242856 , n234347 );
or ( n242857 , n242855 , n242856 );
not ( n242858 , n234350 );
nand ( n242859 , n242858 , n239548 );
nand ( n242860 , n242857 , n242859 );
nand ( n242861 , n242860 , n221674 );
nand ( n242862 , n242854 , n242861 );
xor ( n242863 , n242851 , n242862 );
xor ( n242864 , n242863 , n242752 );
xor ( n242865 , n242841 , n242864 );
xor ( n242866 , n242808 , n242840 );
and ( n242867 , n242866 , n242864 );
and ( n242868 , n242808 , n242840 );
or ( n242869 , n242867 , n242868 );
xor ( n242870 , n242719 , n242520 );
xor ( n242871 , n242483 , n242699 );
xor ( n242872 , n242871 , n242703 );
xor ( n242873 , n242870 , n242872 );
xor ( n242874 , n242719 , n242520 );
and ( n242875 , n242874 , n242872 );
and ( n242876 , n242719 , n242520 );
or ( n242877 , n242875 , n242876 );
xor ( n242878 , n242727 , n242723 );
xor ( n242879 , n242707 , n242711 );
not ( n242880 , n239441 );
not ( n242881 , n242501 );
or ( n242882 , n242880 , n242881 );
not ( n242883 , n239774 );
not ( n242884 , n219742 );
or ( n242885 , n242883 , n242884 );
nand ( n242886 , n239470 , n234293 );
nand ( n242887 , n242885 , n242886 );
buf ( n242888 , n227852 );
nand ( n242889 , n242887 , n242888 );
nand ( n242890 , n242882 , n242889 );
not ( n242891 , n237810 );
not ( n242892 , n242601 );
or ( n242893 , n242891 , n242892 );
not ( n242894 , n237816 );
not ( n242895 , n227448 );
or ( n242896 , n242894 , n242895 );
nand ( n242897 , n240255 , n234394 );
nand ( n242898 , n242896 , n242897 );
nand ( n242899 , n242898 , n238240 );
nand ( n242900 , n242893 , n242899 );
xor ( n242901 , n242890 , n242900 );
not ( n242902 , n221637 );
not ( n242903 , n237937 );
not ( n242904 , n233525 );
not ( n242905 , n242904 );
or ( n242906 , n242903 , n242905 );
nand ( n242907 , n233525 , n221778 );
nand ( n242908 , n242906 , n242907 );
not ( n242909 , n242908 );
or ( n242910 , n242902 , n242909 );
nand ( n242911 , n242476 , n239452 );
nand ( n242912 , n242910 , n242911 );
xor ( n242913 , n242901 , n242912 );
xor ( n242914 , n242879 , n242913 );
xor ( n242915 , n242878 , n242914 );
xor ( n242916 , n242727 , n242723 );
and ( n242917 , n242916 , n242914 );
and ( n242918 , n242727 , n242723 );
or ( n242919 , n242917 , n242918 );
not ( n242920 , n224087 );
not ( n242921 , n242646 );
or ( n242922 , n242920 , n242921 );
not ( n242923 , n239899 );
not ( n242924 , n224700 );
or ( n242925 , n242923 , n242924 );
nand ( n242926 , n236304 , n238672 );
nand ( n242927 , n242925 , n242926 );
nand ( n242928 , n242927 , n239495 );
nand ( n242929 , n242922 , n242928 );
not ( n242930 , n239492 );
not ( n242931 , n242658 );
or ( n242932 , n242930 , n242931 );
not ( n242933 , n241287 );
not ( n242934 , n233546 );
or ( n242935 , n242933 , n242934 );
nand ( n242936 , n40397 , n234273 );
nand ( n242937 , n242935 , n242936 );
nand ( n242938 , n242937 , n240020 );
nand ( n242939 , n242932 , n242938 );
xor ( n242940 , n242929 , n242939 );
not ( n242941 , n242335 );
not ( n242942 , n242489 );
or ( n242943 , n242941 , n242942 );
not ( n242944 , n225952 );
not ( n242945 , n221330 );
or ( n242946 , n242944 , n242945 );
nand ( n242947 , n221956 , n233962 );
nand ( n242948 , n242946 , n242947 );
nand ( n242949 , n242948 , n228775 );
nand ( n242950 , n242943 , n242949 );
xor ( n242951 , n242940 , n242950 );
xor ( n242952 , n242788 , n242951 );
xor ( n242953 , n242952 , n242715 );
xor ( n242954 , n242953 , n242590 );
xor ( n242955 , n242954 , n242865 );
xor ( n242956 , n242953 , n242590 );
and ( n242957 , n242956 , n242865 );
and ( n242958 , n242953 , n242590 );
or ( n242959 , n242957 , n242958 );
xor ( n242960 , n242624 , n242873 );
xor ( n242961 , n242960 , n242630 );
xor ( n242962 , n242624 , n242873 );
and ( n242963 , n242962 , n242630 );
and ( n242964 , n242624 , n242873 );
or ( n242965 , n242963 , n242964 );
xor ( n242966 , n242915 , n242671 );
xor ( n242967 , n242966 , n242955 );
xor ( n242968 , n242915 , n242671 );
and ( n242969 , n242968 , n242955 );
and ( n242970 , n242915 , n242671 );
or ( n242971 , n242969 , n242970 );
xor ( n242972 , n242677 , n242961 );
xor ( n242973 , n242972 , n242683 );
xor ( n242974 , n242677 , n242961 );
and ( n242975 , n242974 , n242683 );
and ( n242976 , n242677 , n242961 );
or ( n242977 , n242975 , n242976 );
xor ( n242978 , n242967 , n242973 );
xor ( n242979 , n242978 , n242689 );
xor ( n242980 , n242967 , n242973 );
and ( n242981 , n242980 , n242689 );
and ( n242982 , n242967 , n242973 );
or ( n242983 , n242981 , n242982 );
xor ( n242984 , n242929 , n242939 );
and ( n242985 , n242984 , n242950 );
and ( n242986 , n242929 , n242939 );
or ( n242987 , n242985 , n242986 );
xor ( n242988 , n242890 , n242900 );
and ( n242989 , n242988 , n242912 );
and ( n242990 , n242890 , n242900 );
or ( n242991 , n242989 , n242990 );
xor ( n242992 , n242818 , n242828 );
and ( n242993 , n242992 , n242839 );
and ( n242994 , n242818 , n242828 );
or ( n242995 , n242993 , n242994 );
xor ( n242996 , n242453 , n242797 );
and ( n242997 , n242996 , n242807 );
and ( n242998 , n242453 , n242797 );
or ( n242999 , n242997 , n242998 );
xor ( n243000 , n242851 , n242862 );
and ( n243001 , n243000 , n242752 );
and ( n243002 , n242851 , n242862 );
or ( n243003 , n243001 , n243002 );
xor ( n243004 , n242483 , n242699 );
and ( n243005 , n243004 , n242703 );
and ( n243006 , n242483 , n242699 );
or ( n243007 , n243005 , n243006 );
xor ( n243008 , n242788 , n242951 );
and ( n243009 , n243008 , n242715 );
and ( n243010 , n242788 , n242951 );
or ( n243011 , n243009 , n243010 );
xor ( n243012 , n242707 , n242711 );
and ( n243013 , n243012 , n242913 );
and ( n243014 , n242707 , n242711 );
or ( n243015 , n243013 , n243014 );
not ( n243016 , n239946 );
not ( n243017 , n229973 );
or ( n243018 , n243016 , n243017 );
nand ( n243019 , n243018 , n229261 );
not ( n243020 , n242748 );
not ( n243021 , n232399 );
or ( n243022 , n243020 , n243021 );
xor ( n243023 , n238199 , n233885 );
nand ( n243024 , n238274 , n243023 );
nand ( n243025 , n243022 , n243024 );
xor ( n243026 , n243019 , n243025 );
and ( n243027 , n234382 , n239001 );
xor ( n243028 , n243026 , n243027 );
xor ( n243029 , n243019 , n243025 );
and ( n243030 , n243029 , n243027 );
and ( n243031 , n243019 , n243025 );
or ( n243032 , n243030 , n243031 );
not ( n243033 , n242737 );
not ( n243034 , n231480 );
not ( n243035 , n219596 );
or ( n243036 , n243034 , n243035 );
nand ( n243037 , n238403 , n233399 );
nand ( n243038 , n243036 , n243037 );
not ( n243039 , n243038 );
or ( n243040 , n243033 , n243039 );
nand ( n243041 , n234371 , n242736 );
nand ( n243042 , n243040 , n243041 );
not ( n243043 , n222454 );
not ( n243044 , n242774 );
or ( n243045 , n243043 , n243044 );
not ( n243046 , n222430 );
not ( n243047 , n226961 );
or ( n243048 , n243046 , n243047 );
nand ( n243049 , n242471 , n238719 );
nand ( n243050 , n243048 , n243049 );
nand ( n243051 , n243050 , n237493 );
nand ( n243052 , n243045 , n243051 );
xor ( n243053 , n243042 , n243052 );
not ( n243054 , n228868 );
not ( n243055 , n228850 );
not ( n243056 , n218912 );
or ( n243057 , n243055 , n243056 );
not ( n243058 , n228850 );
nand ( n243059 , n236752 , n243058 );
nand ( n243060 , n243057 , n243059 );
not ( n243061 , n243060 );
or ( n243062 , n243054 , n243061 );
not ( n243063 , n237038 );
nand ( n243064 , n242762 , n243063 );
nand ( n243065 , n243062 , n243064 );
xor ( n243066 , n243053 , n243065 );
xor ( n243067 , n243042 , n243052 );
and ( n243068 , n243067 , n243065 );
and ( n243069 , n243042 , n243052 );
or ( n243070 , n243068 , n243069 );
not ( n243071 , n218232 );
and ( n243072 , n218205 , n235691 );
not ( n243073 , n218205 );
and ( n243074 , n243073 , n209709 );
nor ( n243075 , n243072 , n243074 );
not ( n243076 , n243075 );
or ( n243077 , n243071 , n243076 );
nand ( n243078 , n242849 , n219461 );
nand ( n243079 , n243077 , n243078 );
not ( n243080 , n220930 );
not ( n243081 , n222399 );
not ( n243082 , n239214 );
or ( n243083 , n243081 , n243082 );
nand ( n243084 , n239548 , n39714 );
nand ( n243085 , n243083 , n243084 );
not ( n243086 , n243085 );
or ( n243087 , n243080 , n243086 );
nand ( n243088 , n242860 , n235913 );
nand ( n243089 , n243087 , n243088 );
xor ( n243090 , n243079 , n243089 );
xor ( n243091 , n243090 , n243028 );
not ( n243092 , n218843 );
not ( n243093 , n221241 );
not ( n243094 , n238486 );
or ( n243095 , n243093 , n243094 );
nand ( n243096 , n236840 , n238363 );
nand ( n243097 , n243095 , n243096 );
not ( n243098 , n243097 );
or ( n243099 , n243092 , n243098 );
nand ( n243100 , n242826 , n223665 );
nand ( n243101 , n243099 , n243100 );
not ( n243102 , n220507 );
not ( n243103 , n242835 );
or ( n243104 , n243102 , n243103 );
not ( n243105 , n240917 );
not ( n243106 , n235962 );
or ( n243107 , n243105 , n243106 );
nand ( n243108 , n38532 , n219797 );
nand ( n243109 , n243107 , n243108 );
nand ( n243110 , n243109 , n239530 );
nand ( n243111 , n243104 , n243110 );
xor ( n243112 , n243101 , n243111 );
not ( n243113 , n220164 );
not ( n243114 , n242803 );
or ( n243115 , n243113 , n243114 );
not ( n243116 , n236768 );
not ( n243117 , n232842 );
or ( n243118 , n243116 , n243117 );
nand ( n243119 , n39608 , n221257 );
nand ( n243120 , n243118 , n243119 );
nand ( n243121 , n243120 , n220881 );
nand ( n243122 , n243115 , n243121 );
xor ( n243123 , n243112 , n243122 );
xor ( n243124 , n243091 , n243123 );
not ( n243125 , n233446 );
not ( n243126 , n242898 );
or ( n243127 , n243125 , n243126 );
not ( n243128 , n236188 );
not ( n243129 , n219518 );
or ( n243130 , n243128 , n243129 );
nand ( n243131 , n40625 , n234394 );
nand ( n243132 , n243130 , n243131 );
nand ( n243133 , n243132 , n238240 );
nand ( n243134 , n243127 , n243133 );
not ( n243135 , n221626 );
not ( n243136 , n242908 );
or ( n243137 , n243135 , n243136 );
not ( n243138 , n237937 );
not ( n243139 , n226724 );
or ( n243140 , n243138 , n243139 );
nand ( n243141 , n238323 , n221778 );
nand ( n243142 , n243140 , n243141 );
nand ( n243143 , n243142 , n221637 );
nand ( n243144 , n243137 , n243143 );
xor ( n243145 , n243134 , n243144 );
not ( n243146 , n220067 );
and ( n243147 , n231501 , n240681 );
not ( n243148 , n231501 );
and ( n243149 , n243148 , n238472 );
nor ( n243150 , n243147 , n243149 );
not ( n243151 , n243150 );
or ( n243152 , n243146 , n243151 );
nand ( n243153 , n242816 , n231018 );
nand ( n243154 , n243152 , n243153 );
xor ( n243155 , n243145 , n243154 );
xor ( n243156 , n243124 , n243155 );
xor ( n243157 , n243091 , n243123 );
and ( n243158 , n243157 , n243155 );
and ( n243159 , n243091 , n243123 );
or ( n243160 , n243158 , n243159 );
xor ( n243161 , n243007 , n243003 );
xor ( n243162 , n243161 , n243015 );
xor ( n243163 , n243007 , n243003 );
and ( n243164 , n243163 , n243015 );
and ( n243165 , n243007 , n243003 );
or ( n243166 , n243164 , n243165 );
xor ( n243167 , n242756 , n242792 );
xor ( n243168 , n243167 , n242987 );
xor ( n243169 , n243011 , n243168 );
not ( n243170 , n227294 );
not ( n243171 , n238681 );
not ( n243172 , n239916 );
or ( n243173 , n243171 , n243172 );
nand ( n243174 , n236547 , n40547 );
nand ( n243175 , n243173 , n243174 );
not ( n243176 , n243175 );
or ( n243177 , n243170 , n243176 );
nand ( n243178 , n242785 , n238409 );
nand ( n243179 , n243177 , n243178 );
not ( n243180 , n242751 );
xor ( n243181 , n243179 , n243180 );
not ( n243182 , n239495 );
not ( n243183 , n224096 );
not ( n243184 , n227004 );
or ( n243185 , n243183 , n243184 );
nand ( n243186 , n40415 , n224095 );
nand ( n243187 , n243185 , n243186 );
not ( n243188 , n243187 );
or ( n243189 , n243182 , n243188 );
nand ( n243190 , n242927 , n224087 );
nand ( n243191 , n243189 , n243190 );
xor ( n243192 , n243181 , n243191 );
xor ( n243193 , n243066 , n243192 );
xor ( n243194 , n243193 , n242991 );
xor ( n243195 , n243169 , n243194 );
xor ( n243196 , n243011 , n243168 );
and ( n243197 , n243196 , n243194 );
and ( n243198 , n243011 , n243168 );
or ( n243199 , n243197 , n243198 );
xor ( n243200 , n242995 , n242999 );
not ( n243201 , n240020 );
not ( n243202 , n241287 );
not ( n243203 , n221712 );
or ( n243204 , n243202 , n243203 );
nand ( n243205 , n40182 , n234273 );
nand ( n243206 , n243204 , n243205 );
not ( n243207 , n243206 );
or ( n243208 , n243201 , n243207 );
nand ( n243209 , n242937 , n239492 );
nand ( n243210 , n243208 , n243209 );
not ( n243211 , n228775 );
not ( n243212 , n225952 );
not ( n243213 , n40258 );
or ( n243214 , n243212 , n243213 );
nand ( n243215 , n220970 , n233962 );
nand ( n243216 , n243214 , n243215 );
not ( n243217 , n243216 );
or ( n243218 , n243211 , n243217 );
nand ( n243219 , n242335 , n242948 );
nand ( n243220 , n243218 , n243219 );
xor ( n243221 , n243210 , n243220 );
not ( n243222 , n227852 );
not ( n243223 , n226651 );
not ( n243224 , n221725 );
or ( n243225 , n243223 , n243224 );
nand ( n243226 , n234014 , n234293 );
nand ( n243227 , n243225 , n243226 );
not ( n243228 , n243227 );
or ( n243229 , n243222 , n243228 );
nand ( n243230 , n242887 , n237797 );
nand ( n243231 , n243229 , n243230 );
xor ( n243232 , n243221 , n243231 );
xor ( n243233 , n243200 , n243232 );
xor ( n243234 , n243233 , n243156 );
xor ( n243235 , n243234 , n242869 );
xor ( n243236 , n243233 , n243156 );
and ( n243237 , n243236 , n242869 );
and ( n243238 , n243233 , n243156 );
or ( n243239 , n243237 , n243238 );
xor ( n243240 , n242877 , n243162 );
xor ( n243241 , n243240 , n242919 );
xor ( n243242 , n242877 , n243162 );
and ( n243243 , n243242 , n242919 );
and ( n243244 , n242877 , n243162 );
or ( n243245 , n243243 , n243244 );
xor ( n243246 , n243195 , n242959 );
xor ( n243247 , n243246 , n243235 );
xor ( n243248 , n243195 , n242959 );
and ( n243249 , n243248 , n243235 );
and ( n243250 , n243195 , n242959 );
or ( n243251 , n243249 , n243250 );
xor ( n243252 , n243241 , n242965 );
xor ( n243253 , n243252 , n242971 );
xor ( n243254 , n243241 , n242965 );
and ( n243255 , n243254 , n242971 );
and ( n243256 , n243241 , n242965 );
or ( n243257 , n243255 , n243256 );
xor ( n243258 , n243247 , n243253 );
xor ( n243259 , n243258 , n242977 );
xor ( n243260 , n243247 , n243253 );
and ( n243261 , n243260 , n242977 );
and ( n243262 , n243247 , n243253 );
or ( n243263 , n243261 , n243262 );
xor ( n243264 , n243179 , n243180 );
and ( n243265 , n243264 , n243191 );
and ( n243266 , n243179 , n243180 );
or ( n243267 , n243265 , n243266 );
xor ( n243268 , n243210 , n243220 );
and ( n243269 , n243268 , n243231 );
and ( n243270 , n243210 , n243220 );
or ( n243271 , n243269 , n243270 );
xor ( n243272 , n243134 , n243144 );
and ( n243273 , n243272 , n243154 );
and ( n243274 , n243134 , n243144 );
or ( n243275 , n243273 , n243274 );
xor ( n243276 , n243101 , n243111 );
and ( n243277 , n243276 , n243122 );
and ( n243278 , n243101 , n243111 );
or ( n243279 , n243277 , n243278 );
xor ( n243280 , n243079 , n243089 );
and ( n243281 , n243280 , n243028 );
and ( n243282 , n243079 , n243089 );
or ( n243283 , n243281 , n243282 );
xor ( n243284 , n242756 , n242792 );
and ( n243285 , n243284 , n242987 );
and ( n243286 , n242756 , n242792 );
or ( n243287 , n243285 , n243286 );
xor ( n243288 , n243066 , n243192 );
and ( n243289 , n243288 , n242991 );
and ( n243290 , n243066 , n243192 );
or ( n243291 , n243289 , n243290 );
xor ( n243292 , n242995 , n242999 );
and ( n243293 , n243292 , n243232 );
and ( n243294 , n242995 , n242999 );
or ( n243295 , n243293 , n243294 );
not ( n243296 , n238274 );
not ( n243297 , n234382 );
not ( n243298 , n243297 );
not ( n243299 , n40724 );
or ( n243300 , n243298 , n243299 );
not ( n243301 , n238671 );
nand ( n243302 , n243301 , n239281 );
nand ( n243303 , n243300 , n243302 );
not ( n243304 , n243303 );
or ( n243305 , n243296 , n243304 );
nand ( n243306 , n233105 , n243023 );
nand ( n243307 , n243305 , n243306 );
not ( n243308 , n234371 );
not ( n243309 , n243038 );
or ( n243310 , n243308 , n243309 );
not ( n243311 , n231480 );
not ( n243312 , n237948 );
or ( n243313 , n243311 , n243312 );
not ( n243314 , n231480 );
nand ( n243315 , n220568 , n243314 );
nand ( n243316 , n243313 , n243315 );
nand ( n243317 , n243316 , n242737 );
nand ( n243318 , n243310 , n243317 );
xor ( n243319 , n243307 , n243318 );
not ( n243320 , n238409 );
not ( n243321 , n243175 );
or ( n243322 , n243320 , n243321 );
not ( n243323 , n223182 );
not ( n243324 , n230490 );
or ( n243325 , n243323 , n243324 );
not ( n243326 , n238681 );
nand ( n243327 , n237963 , n243326 );
nand ( n243328 , n243325 , n243327 );
nand ( n243329 , n243328 , n227294 );
nand ( n243330 , n243322 , n243329 );
xor ( n243331 , n243319 , n243330 );
xor ( n243332 , n243307 , n243318 );
and ( n243333 , n243332 , n243330 );
and ( n243334 , n243307 , n243318 );
or ( n243335 , n243333 , n243334 );
not ( n243336 , n224087 );
not ( n243337 , n243187 );
or ( n243338 , n243336 , n243337 );
not ( n243339 , n224096 );
not ( n243340 , n237971 );
or ( n243341 , n243339 , n243340 );
nand ( n243342 , n239527 , n237129 );
nand ( n243343 , n243341 , n243342 );
nand ( n243344 , n243343 , n227782 );
nand ( n243345 , n243338 , n243344 );
nand ( n243346 , n240156 , n41071 );
xor ( n243347 , n243345 , n243346 );
not ( n243348 , n240020 );
and ( n243349 , n241287 , n222101 );
not ( n243350 , n241287 );
and ( n243351 , n243350 , n224700 );
nor ( n243352 , n243349 , n243351 );
not ( n243353 , n243352 );
or ( n243354 , n243348 , n243353 );
nand ( n243355 , n243206 , n240271 );
nand ( n243356 , n243354 , n243355 );
xor ( n243357 , n243347 , n243356 );
xor ( n243358 , n243345 , n243346 );
and ( n243359 , n243358 , n243356 );
and ( n243360 , n243345 , n243346 );
or ( n243361 , n243359 , n243360 );
not ( n243362 , n220507 );
not ( n243363 , n243109 );
or ( n243364 , n243362 , n243363 );
not ( n243365 , n219424 );
not ( n243366 , n39366 );
or ( n243367 , n243365 , n243366 );
not ( n243368 , n240917 );
nand ( n243369 , n243368 , n237229 );
nand ( n243370 , n243367 , n243369 );
nand ( n243371 , n243370 , n219076 );
nand ( n243372 , n243364 , n243371 );
not ( n243373 , n220164 );
not ( n243374 , n243120 );
or ( n243375 , n243373 , n243374 );
not ( n243376 , n220151 );
not ( n243377 , n227201 );
or ( n243378 , n243376 , n243377 );
nand ( n243379 , n39089 , n221257 );
nand ( n243380 , n243378 , n243379 );
nand ( n243381 , n243380 , n220881 );
nand ( n243382 , n243375 , n243381 );
xor ( n243383 , n243372 , n243382 );
xor ( n243384 , n243383 , n243032 );
xor ( n243385 , n243384 , n243287 );
not ( n243386 , n239452 );
not ( n243387 , n243142 );
or ( n243388 , n243386 , n243387 );
not ( n243389 , n238705 );
not ( n243390 , n234350 );
or ( n243391 , n243389 , n243390 );
not ( n243392 , n242210 );
nand ( n243393 , n243392 , n221778 );
nand ( n243394 , n243391 , n243393 );
nand ( n243395 , n243394 , n221637 );
nand ( n243396 , n243388 , n243395 );
xor ( n243397 , n243396 , n243070 );
xor ( n243398 , n243397 , n243267 );
xor ( n243399 , n243385 , n243398 );
xor ( n243400 , n243384 , n243287 );
and ( n243401 , n243400 , n243398 );
and ( n243402 , n243384 , n243287 );
or ( n243403 , n243401 , n243402 );
xor ( n243404 , n243295 , n243291 );
xor ( n243405 , n243404 , n243160 );
xor ( n243406 , n243295 , n243291 );
and ( n243407 , n243406 , n243160 );
and ( n243408 , n243295 , n243291 );
or ( n243409 , n243407 , n243408 );
xor ( n243410 , n243271 , n243331 );
xor ( n243411 , n243410 , n243357 );
xor ( n243412 , n243275 , n243279 );
not ( n243413 , n228775 );
not ( n243414 , n225952 );
not ( n243415 , n238786 );
or ( n243416 , n243414 , n243415 );
nand ( n243417 , n226505 , n232493 );
nand ( n243418 , n243416 , n243417 );
not ( n243419 , n243418 );
or ( n243420 , n243413 , n243419 );
nand ( n243421 , n243216 , n242335 );
nand ( n243422 , n243420 , n243421 );
not ( n243423 , n237797 );
not ( n243424 , n243227 );
or ( n243425 , n243423 , n243424 );
and ( n243426 , n220599 , n226651 );
not ( n243427 , n220599 );
and ( n243428 , n243427 , n226650 );
or ( n243429 , n243426 , n243428 );
nand ( n243430 , n243429 , n242888 );
nand ( n243431 , n243425 , n243430 );
xor ( n243432 , n243422 , n243431 );
not ( n243433 , n238240 );
not ( n243434 , n237816 );
not ( n243435 , n219742 );
or ( n243436 , n243434 , n243435 );
nand ( n243437 , n239470 , n227596 );
nand ( n243438 , n243436 , n243437 );
not ( n243439 , n243438 );
or ( n243440 , n243433 , n243439 );
nand ( n243441 , n243132 , n237810 );
nand ( n243442 , n243440 , n243441 );
xor ( n243443 , n243432 , n243442 );
xor ( n243444 , n243412 , n243443 );
xor ( n243445 , n243411 , n243444 );
not ( n243446 , n220059 );
not ( n243447 , n243150 );
or ( n243448 , n243446 , n243447 );
nand ( n243449 , n220067 , n231500 );
nand ( n243450 , n243448 , n243449 );
not ( n243451 , n235913 );
not ( n243452 , n243085 );
or ( n243453 , n243451 , n243452 );
not ( n243454 , n222399 );
not ( n243455 , n234324 );
or ( n243456 , n243454 , n243455 );
not ( n243457 , n220906 );
not ( n243458 , n234324 );
nand ( n243459 , n243457 , n243458 );
nand ( n243460 , n243456 , n243459 );
nand ( n243461 , n243460 , n221674 );
nand ( n243462 , n243453 , n243461 );
xor ( n243463 , n243450 , n243462 );
not ( n243464 , n223665 );
not ( n243465 , n243097 );
or ( n243466 , n243464 , n243465 );
not ( n243467 , n221241 );
not ( n243468 , n237271 );
or ( n243469 , n243467 , n243468 );
nand ( n243470 , n237272 , n238363 );
nand ( n243471 , n243469 , n243470 );
nand ( n243472 , n243471 , n218843 );
nand ( n243473 , n243466 , n243472 );
xor ( n243474 , n243463 , n243473 );
xor ( n243475 , n243474 , n243283 );
not ( n243476 , n243063 );
not ( n243477 , n243060 );
or ( n243478 , n243476 , n243477 );
not ( n243479 , n228850 );
not ( n243480 , n219880 );
or ( n243481 , n243479 , n243480 );
nand ( n243482 , n219226 , n238617 );
nand ( n243483 , n243481 , n243482 );
nand ( n243484 , n243483 , n228868 );
nand ( n243485 , n243478 , n243484 );
not ( n243486 , n237493 );
and ( n243487 , n222430 , n235452 );
not ( n243488 , n222430 );
and ( n243489 , n243488 , n39880 );
or ( n243490 , n243487 , n243489 );
not ( n243491 , n243490 );
or ( n243492 , n243486 , n243491 );
nand ( n243493 , n243050 , n222454 );
nand ( n243494 , n243492 , n243493 );
xor ( n243495 , n243485 , n243494 );
not ( n243496 , n219461 );
not ( n243497 , n243075 );
or ( n243498 , n243496 , n243497 );
not ( n243499 , n224497 );
not ( n243500 , n239617 );
or ( n243501 , n243499 , n243500 );
nand ( n243502 , n238835 , n218256 );
nand ( n243503 , n243501 , n243502 );
nand ( n243504 , n243503 , n218232 );
nand ( n243505 , n243498 , n243504 );
xor ( n243506 , n243495 , n243505 );
xor ( n243507 , n243475 , n243506 );
xor ( n243508 , n243445 , n243507 );
xor ( n243509 , n243411 , n243444 );
and ( n243510 , n243509 , n243507 );
and ( n243511 , n243411 , n243444 );
or ( n243512 , n243510 , n243511 );
xor ( n243513 , n243399 , n243166 );
xor ( n243514 , n243513 , n243199 );
xor ( n243515 , n243399 , n243166 );
and ( n243516 , n243515 , n243199 );
and ( n243517 , n243399 , n243166 );
or ( n243518 , n243516 , n243517 );
xor ( n243519 , n243405 , n243239 );
xor ( n243520 , n243519 , n243508 );
xor ( n243521 , n243405 , n243239 );
and ( n243522 , n243521 , n243508 );
and ( n243523 , n243405 , n243239 );
or ( n243524 , n243522 , n243523 );
xor ( n243525 , n243514 , n243245 );
xor ( n243526 , n243525 , n243251 );
xor ( n243527 , n243514 , n243245 );
and ( n243528 , n243527 , n243251 );
and ( n243529 , n243514 , n243245 );
or ( n243530 , n243528 , n243529 );
xor ( n243531 , n243520 , n243526 );
xor ( n243532 , n243531 , n243257 );
xor ( n243533 , n243520 , n243526 );
and ( n243534 , n243533 , n243257 );
and ( n243535 , n243520 , n243526 );
or ( n243536 , n243534 , n243535 );
xor ( n243537 , n243422 , n243431 );
and ( n243538 , n243537 , n243442 );
and ( n243539 , n243422 , n243431 );
or ( n243540 , n243538 , n243539 );
xor ( n243541 , n243485 , n243494 );
and ( n243542 , n243541 , n243505 );
and ( n243543 , n243485 , n243494 );
or ( n243544 , n243542 , n243543 );
xor ( n243545 , n243372 , n243382 );
and ( n243546 , n243545 , n243032 );
and ( n243547 , n243372 , n243382 );
or ( n243548 , n243546 , n243547 );
xor ( n243549 , n243450 , n243462 );
and ( n243550 , n243549 , n243473 );
and ( n243551 , n243450 , n243462 );
or ( n243552 , n243550 , n243551 );
xor ( n243553 , n243396 , n243070 );
and ( n243554 , n243553 , n243267 );
and ( n243555 , n243396 , n243070 );
or ( n243556 , n243554 , n243555 );
xor ( n243557 , n243271 , n243331 );
and ( n243558 , n243557 , n243357 );
and ( n243559 , n243271 , n243331 );
or ( n243560 , n243558 , n243559 );
xor ( n243561 , n243275 , n243279 );
and ( n243562 , n243561 , n243443 );
and ( n243563 , n243275 , n243279 );
or ( n243564 , n243562 , n243563 );
xor ( n243565 , n243474 , n243283 );
and ( n243566 , n243565 , n243506 );
and ( n243567 , n243474 , n243283 );
or ( n243568 , n243566 , n243567 );
not ( n243569 , n227138 );
not ( n243570 , n227130 );
or ( n243571 , n243569 , n243570 );
nand ( n243572 , n243571 , n217616 );
and ( n243573 , n238199 , n233885 );
xor ( n243574 , n243572 , n243573 );
not ( n243575 , n238409 );
not ( n243576 , n243328 );
or ( n243577 , n243575 , n243576 );
not ( n243578 , n223182 );
not ( n243579 , n242472 );
or ( n243580 , n243578 , n243579 );
nand ( n243581 , n229928 , n238404 );
nand ( n243582 , n243580 , n243581 );
nand ( n243583 , n243582 , n227294 );
nand ( n243584 , n243577 , n243583 );
xor ( n243585 , n243574 , n243584 );
xor ( n243586 , n243572 , n243573 );
and ( n243587 , n243586 , n243584 );
and ( n243588 , n243572 , n243573 );
or ( n243589 , n243587 , n243588 );
not ( n243590 , n238274 );
not ( n243591 , n239281 );
not ( n243592 , n219596 );
or ( n243593 , n243591 , n243592 );
nand ( n243594 , n238403 , n231753 );
nand ( n243595 , n243593 , n243594 );
not ( n243596 , n243595 );
or ( n243597 , n243590 , n243596 );
nand ( n243598 , n243303 , n233105 );
nand ( n243599 , n243597 , n243598 );
not ( n243600 , n234378 );
not ( n243601 , n239393 );
not ( n243602 , n218912 );
or ( n243603 , n243601 , n243602 );
nand ( n243604 , n218911 , n243314 );
nand ( n243605 , n243603 , n243604 );
not ( n243606 , n243605 );
or ( n243607 , n243600 , n243606 );
nand ( n243608 , n243316 , n234371 );
nand ( n243609 , n243607 , n243608 );
xor ( n243610 , n243599 , n243609 );
not ( n243611 , n243346 );
xor ( n243612 , n243610 , n243611 );
xor ( n243613 , n243599 , n243609 );
and ( n243614 , n243613 , n243611 );
and ( n243615 , n243599 , n243609 );
or ( n243616 , n243614 , n243615 );
not ( n243617 , n237493 );
not ( n243618 , n222430 );
not ( n243619 , n233018 );
not ( n243620 , n243619 );
or ( n243621 , n243618 , n243620 );
nand ( n243622 , n238323 , n238719 );
nand ( n243623 , n243621 , n243622 );
not ( n243624 , n243623 );
or ( n243625 , n243617 , n243624 );
nand ( n243626 , n243490 , n222454 );
nand ( n243627 , n243625 , n243626 );
not ( n243628 , n219461 );
not ( n243629 , n243503 );
or ( n243630 , n243628 , n243629 );
not ( n243631 , n224497 );
not ( n243632 , n239186 );
or ( n243633 , n243631 , n243632 );
nand ( n243634 , n239185 , n234949 );
nand ( n243635 , n243633 , n243634 );
nand ( n243636 , n243635 , n218232 );
nand ( n243637 , n243630 , n243636 );
xor ( n243638 , n243627 , n243637 );
not ( n243639 , n239530 );
not ( n243640 , n219424 );
not ( n243641 , n238486 );
or ( n243642 , n243640 , n243641 );
nand ( n243643 , n39288 , n219423 );
nand ( n243644 , n243642 , n243643 );
not ( n243645 , n243644 );
or ( n243646 , n243639 , n243645 );
nand ( n243647 , n220507 , n243370 );
nand ( n243648 , n243646 , n243647 );
xor ( n243649 , n243638 , n243648 );
xor ( n243650 , n243649 , n243556 );
xor ( n243651 , n243650 , n243564 );
xor ( n243652 , n243649 , n243556 );
and ( n243653 , n243652 , n243564 );
and ( n243654 , n243649 , n243556 );
or ( n243655 , n243653 , n243654 );
xor ( n243656 , n243361 , n243540 );
xor ( n243657 , n243656 , n243612 );
xor ( n243658 , n243560 , n243657 );
not ( n243659 , n221637 );
and ( n243660 , n237937 , n39714 );
not ( n243661 , n237937 );
and ( n243662 , n243661 , n240738 );
nor ( n243663 , n243660 , n243662 );
not ( n243664 , n243663 );
or ( n243665 , n243659 , n243664 );
nand ( n243666 , n243394 , n239452 );
nand ( n243667 , n243665 , n243666 );
xor ( n243668 , n243667 , n243585 );
xor ( n243669 , n243668 , n243335 );
xor ( n243670 , n243658 , n243669 );
xor ( n243671 , n243560 , n243657 );
and ( n243672 , n243671 , n243669 );
and ( n243673 , n243560 , n243657 );
or ( n243674 , n243672 , n243673 );
not ( n243675 , n242888 );
not ( n243676 , n234295 );
not ( n243677 , n240601 );
or ( n243678 , n243676 , n243677 );
nand ( n243679 , n40259 , n226650 );
nand ( n243680 , n243678 , n243679 );
not ( n243681 , n243680 );
or ( n243682 , n243675 , n243681 );
nand ( n243683 , n237797 , n243429 );
nand ( n243684 , n243682 , n243683 );
not ( n243685 , n238240 );
not ( n243686 , n236188 );
not ( n243687 , n239077 );
or ( n243688 , n243686 , n243687 );
nand ( n243689 , n239080 , n227596 );
nand ( n243690 , n243688 , n243689 );
not ( n243691 , n243690 );
or ( n243692 , n243685 , n243691 );
nand ( n243693 , n243438 , n237810 );
nand ( n243694 , n243692 , n243693 );
xor ( n243695 , n243684 , n243694 );
not ( n243696 , n239794 );
not ( n243697 , n243483 );
or ( n243698 , n243696 , n243697 );
not ( n243699 , n228850 );
not ( n243700 , n234108 );
or ( n243701 , n243699 , n243700 );
nand ( n243702 , n40625 , n238617 );
nand ( n243703 , n243701 , n243702 );
nand ( n243704 , n243703 , n228868 );
nand ( n243705 , n243698 , n243704 );
xor ( n243706 , n243695 , n243705 );
not ( n243707 , n239495 );
not ( n243708 , n239899 );
not ( n243709 , n237600 );
or ( n243710 , n243708 , n243709 );
nand ( n243711 , n239917 , n239903 );
nand ( n243712 , n243710 , n243711 );
not ( n243713 , n243712 );
or ( n243714 , n243707 , n243713 );
nand ( n243715 , n243343 , n224087 );
nand ( n243716 , n243714 , n243715 );
not ( n243717 , n239492 );
not ( n243718 , n243352 );
or ( n243719 , n243717 , n243718 );
not ( n243720 , n234878 );
not ( n243721 , n240637 );
or ( n243722 , n243720 , n243721 );
nand ( n243723 , n238362 , n240617 );
nand ( n243724 , n243722 , n243723 );
nand ( n243725 , n243724 , n240020 );
nand ( n243726 , n243719 , n243725 );
xor ( n243727 , n243716 , n243726 );
not ( n243728 , n242335 );
not ( n243729 , n243418 );
or ( n243730 , n243728 , n243729 );
not ( n243731 , n232494 );
not ( n243732 , n229936 );
or ( n243733 , n243731 , n243732 );
buf ( n243734 , n236719 );
nand ( n243735 , n243734 , n229807 );
nand ( n243736 , n243733 , n243735 );
nand ( n243737 , n243736 , n238776 );
nand ( n243738 , n243730 , n243737 );
xor ( n243739 , n243727 , n243738 );
xor ( n243740 , n243706 , n243739 );
not ( n243741 , n220164 );
not ( n243742 , n243380 );
or ( n243743 , n243741 , n243742 );
not ( n243744 , n220151 );
not ( n243745 , n235962 );
or ( n243746 , n243744 , n243745 );
nand ( n243747 , n38532 , n221257 );
nand ( n243748 , n243746 , n243747 );
nand ( n243749 , n243748 , n219779 );
nand ( n243750 , n243743 , n243749 );
not ( n243751 , n220930 );
and ( n243752 , n222399 , n39608 );
not ( n243753 , n222399 );
not ( n243754 , n39608 );
and ( n243755 , n243753 , n243754 );
nor ( n243756 , n243752 , n243755 );
not ( n243757 , n243756 );
or ( n243758 , n243751 , n243757 );
nand ( n243759 , n243460 , n235913 );
nand ( n243760 , n243758 , n243759 );
xor ( n243761 , n243750 , n243760 );
not ( n243762 , n218843 );
not ( n243763 , n221241 );
buf ( n243764 , n235691 );
not ( n243765 , n243764 );
not ( n243766 , n243765 );
or ( n243767 , n243763 , n243766 );
nand ( n243768 , n243764 , n238363 );
nand ( n243769 , n243767 , n243768 );
not ( n243770 , n243769 );
or ( n243771 , n243762 , n243770 );
nand ( n243772 , n243471 , n239508 );
nand ( n243773 , n243771 , n243772 );
xor ( n243774 , n243761 , n243773 );
xor ( n243775 , n243740 , n243774 );
xor ( n243776 , n243568 , n243775 );
xor ( n243777 , n243544 , n243548 );
xor ( n243778 , n243777 , n243552 );
xor ( n243779 , n243776 , n243778 );
xor ( n243780 , n243568 , n243775 );
and ( n243781 , n243780 , n243778 );
and ( n243782 , n243568 , n243775 );
or ( n243783 , n243781 , n243782 );
xor ( n243784 , n243403 , n243651 );
xor ( n243785 , n243784 , n243670 );
xor ( n243786 , n243403 , n243651 );
and ( n243787 , n243786 , n243670 );
and ( n243788 , n243403 , n243651 );
or ( n243789 , n243787 , n243788 );
xor ( n243790 , n243409 , n243512 );
xor ( n243791 , n243790 , n243779 );
xor ( n243792 , n243409 , n243512 );
and ( n243793 , n243792 , n243779 );
and ( n243794 , n243409 , n243512 );
or ( n243795 , n243793 , n243794 );
xor ( n243796 , n243785 , n243518 );
xor ( n243797 , n243796 , n243524 );
xor ( n243798 , n243785 , n243518 );
and ( n243799 , n243798 , n243524 );
and ( n243800 , n243785 , n243518 );
or ( n243801 , n243799 , n243800 );
xor ( n243802 , n243791 , n243797 );
xor ( n243803 , n243802 , n243530 );
xor ( n243804 , n243791 , n243797 );
and ( n243805 , n243804 , n243530 );
and ( n243806 , n243791 , n243797 );
or ( n243807 , n243805 , n243806 );
xor ( n243808 , n243716 , n243726 );
and ( n243809 , n243808 , n243738 );
and ( n243810 , n243716 , n243726 );
or ( n243811 , n243809 , n243810 );
xor ( n243812 , n243684 , n243694 );
and ( n243813 , n243812 , n243705 );
and ( n243814 , n243684 , n243694 );
or ( n243815 , n243813 , n243814 );
xor ( n243816 , n243627 , n243637 );
and ( n243817 , n243816 , n243648 );
and ( n243818 , n243627 , n243637 );
or ( n243819 , n243817 , n243818 );
xor ( n243820 , n243750 , n243760 );
and ( n243821 , n243820 , n243773 );
and ( n243822 , n243750 , n243760 );
or ( n243823 , n243821 , n243822 );
xor ( n243824 , n243667 , n243585 );
and ( n243825 , n243824 , n243335 );
and ( n243826 , n243667 , n243585 );
or ( n243827 , n243825 , n243826 );
xor ( n243828 , n243361 , n243540 );
and ( n243829 , n243828 , n243612 );
and ( n243830 , n243361 , n243540 );
or ( n243831 , n243829 , n243830 );
xor ( n243832 , n243544 , n243548 );
and ( n243833 , n243832 , n243552 );
and ( n243834 , n243544 , n243548 );
or ( n243835 , n243833 , n243834 );
xor ( n243836 , n243706 , n243739 );
and ( n243837 , n243836 , n243774 );
and ( n243838 , n243706 , n243739 );
or ( n243839 , n243837 , n243838 );
not ( n243840 , n224087 );
not ( n243841 , n243712 );
or ( n243842 , n243840 , n243841 );
not ( n243843 , n224096 );
not ( n243844 , n230490 );
or ( n243845 , n243843 , n243844 );
nand ( n243846 , n239515 , n224095 );
nand ( n243847 , n243845 , n243846 );
nand ( n243848 , n243847 , n239495 );
nand ( n243849 , n243842 , n243848 );
not ( n243850 , n238274 );
xor ( n243851 , n233891 , n208046 );
not ( n243852 , n243851 );
or ( n243853 , n243850 , n243852 );
nand ( n243854 , n243595 , n233105 );
nand ( n243855 , n243853 , n243854 );
xor ( n243856 , n243849 , n243855 );
not ( n243857 , n239492 );
not ( n243858 , n243724 );
or ( n243859 , n243857 , n243858 );
not ( n243860 , n242653 );
not ( n243861 , n222940 );
or ( n243862 , n243860 , n243861 );
nand ( n243863 , n236290 , n240617 );
nand ( n243864 , n243862 , n243863 );
nand ( n243865 , n243864 , n240020 );
nand ( n243866 , n243859 , n243865 );
xor ( n243867 , n243856 , n243866 );
xor ( n243868 , n243849 , n243855 );
and ( n243869 , n243868 , n243866 );
and ( n243870 , n243849 , n243855 );
or ( n243871 , n243869 , n243870 );
not ( n243872 , n242335 );
not ( n243873 , n243736 );
or ( n243874 , n243872 , n243873 );
not ( n243875 , n232494 );
not ( n243876 , n235383 );
or ( n243877 , n243875 , n243876 );
nand ( n243878 , n236304 , n232497 );
nand ( n243879 , n243877 , n243878 );
nand ( n243880 , n243879 , n238776 );
nand ( n243881 , n243874 , n243880 );
not ( n243882 , n242888 );
not ( n243883 , n226651 );
not ( n243884 , n222121 );
or ( n243885 , n243883 , n243884 );
nand ( n243886 , n40397 , n238230 );
nand ( n243887 , n243885 , n243886 );
not ( n243888 , n243887 );
or ( n243889 , n243882 , n243888 );
nand ( n243890 , n243680 , n237797 );
nand ( n243891 , n243889 , n243890 );
xor ( n243892 , n243881 , n243891 );
not ( n243893 , n237810 );
not ( n243894 , n243690 );
or ( n243895 , n243893 , n243894 );
not ( n243896 , n233450 );
not ( n243897 , n220599 );
or ( n243898 , n243896 , n243897 );
nand ( n243899 , n221956 , n234394 );
nand ( n243900 , n243898 , n243899 );
nand ( n243901 , n243900 , n238240 );
nand ( n243902 , n243895 , n243901 );
xor ( n243903 , n243892 , n243902 );
xor ( n243904 , n243881 , n243891 );
and ( n243905 , n243904 , n243902 );
and ( n243906 , n243881 , n243891 );
or ( n243907 , n243905 , n243906 );
xor ( n243908 , n243616 , n243811 );
xor ( n243909 , n243908 , n243815 );
xor ( n243910 , n243831 , n243909 );
xor ( n243911 , n243910 , n243835 );
xor ( n243912 , n243831 , n243909 );
and ( n243913 , n243912 , n243835 );
and ( n243914 , n243831 , n243909 );
or ( n243915 , n243913 , n243914 );
not ( n243916 , n228868 );
not ( n243917 , n228850 );
not ( n243918 , n219742 );
or ( n243919 , n243917 , n243918 );
nand ( n243920 , n239470 , n228847 );
nand ( n243921 , n243919 , n243920 );
not ( n243922 , n243921 );
or ( n243923 , n243916 , n243922 );
nand ( n243924 , n243703 , n243063 );
nand ( n243925 , n243923 , n243924 );
not ( n243926 , n239393 );
not ( n243927 , n227448 );
or ( n243928 , n243926 , n243927 );
not ( n243929 , n40561 );
nand ( n243930 , n243929 , n243314 );
nand ( n243931 , n243928 , n243930 );
nand ( n243932 , n243931 , n242737 );
nand ( n243933 , n234371 , n243605 );
nand ( n243934 , n243932 , n243933 );
xor ( n243935 , n243925 , n243934 );
nand ( n243936 , n40724 , n239281 );
xor ( n243937 , n243935 , n243936 );
xor ( n243938 , n243937 , n243903 );
not ( n243939 , n235913 );
not ( n243940 , n243756 );
or ( n243941 , n243939 , n243940 );
not ( n243942 , n222399 );
not ( n243943 , n236382 );
or ( n243944 , n243942 , n243943 );
nand ( n243945 , n238857 , n239548 );
nand ( n243946 , n243944 , n243945 );
nand ( n243947 , n243946 , n220930 );
nand ( n243948 , n243941 , n243947 );
not ( n243949 , n219461 );
not ( n243950 , n243635 );
or ( n243951 , n243949 , n243950 );
nand ( n243952 , n218232 , n224497 );
nand ( n243953 , n243951 , n243952 );
xor ( n243954 , n243948 , n243953 );
not ( n243955 , n221626 );
not ( n243956 , n243663 );
or ( n243957 , n243955 , n243956 );
not ( n243958 , n237937 );
not ( n243959 , n234324 );
or ( n243960 , n243958 , n243959 );
nand ( n243961 , n243458 , n221612 );
nand ( n243962 , n243960 , n243961 );
nand ( n243963 , n243962 , n221637 );
nand ( n243964 , n243957 , n243963 );
xor ( n243965 , n243954 , n243964 );
xor ( n243966 , n243938 , n243965 );
xor ( n243967 , n243966 , n243839 );
xor ( n243968 , n243867 , n243819 );
xor ( n243969 , n243968 , n243823 );
xor ( n243970 , n243967 , n243969 );
xor ( n243971 , n243966 , n243839 );
and ( n243972 , n243971 , n243969 );
and ( n243973 , n243966 , n243839 );
or ( n243974 , n243972 , n243973 );
xor ( n243975 , n243674 , n243655 );
not ( n243976 , n227294 );
not ( n243977 , n238681 );
not ( n243978 , n238728 );
or ( n243979 , n243977 , n243978 );
nand ( n243980 , n39880 , n243326 );
nand ( n243981 , n243979 , n243980 );
not ( n243982 , n243981 );
or ( n243983 , n243976 , n243982 );
nand ( n243984 , n243582 , n238409 );
nand ( n243985 , n243983 , n243984 );
not ( n243986 , n239508 );
not ( n243987 , n243769 );
or ( n243988 , n243986 , n243987 );
not ( n243989 , n221241 );
not ( n243990 , n239617 );
or ( n243991 , n243989 , n243990 );
nand ( n243992 , n209866 , n238363 );
nand ( n243993 , n243991 , n243992 );
nand ( n243994 , n243993 , n218843 );
nand ( n243995 , n243988 , n243994 );
xor ( n243996 , n243985 , n243995 );
not ( n243997 , n219779 );
not ( n243998 , n236768 );
not ( n243999 , n228165 );
or ( n244000 , n243998 , n243999 );
nand ( n244001 , n39365 , n222414 );
nand ( n244002 , n244000 , n244001 );
not ( n244003 , n244002 );
or ( n244004 , n243997 , n244003 );
nand ( n244005 , n243748 , n220164 );
nand ( n244006 , n244004 , n244005 );
xor ( n244007 , n243996 , n244006 );
not ( n244008 , n220507 );
not ( n244009 , n243644 );
or ( n244010 , n244008 , n244009 );
not ( n244011 , n240917 );
not ( n244012 , n237271 );
or ( n244013 , n244011 , n244012 );
nand ( n244014 , n240308 , n219420 );
nand ( n244015 , n244013 , n244014 );
nand ( n244016 , n244015 , n239530 );
nand ( n244017 , n244010 , n244016 );
not ( n244018 , n237503 );
not ( n244019 , n243623 );
or ( n244020 , n244018 , n244019 );
not ( n244021 , n222430 );
not ( n244022 , n242210 );
or ( n244023 , n244021 , n244022 );
not ( n244024 , n240229 );
nand ( n244025 , n242858 , n244024 );
nand ( n244026 , n244023 , n244025 );
nand ( n244027 , n244026 , n237493 );
nand ( n244028 , n244020 , n244027 );
xor ( n244029 , n244017 , n244028 );
xor ( n244030 , n244029 , n243589 );
xor ( n244031 , n244007 , n244030 );
xor ( n244032 , n244031 , n243827 );
xor ( n244033 , n243975 , n244032 );
xor ( n244034 , n243674 , n243655 );
and ( n244035 , n244034 , n244032 );
and ( n244036 , n243674 , n243655 );
or ( n244037 , n244035 , n244036 );
xor ( n244038 , n243911 , n243783 );
xor ( n244039 , n244038 , n243970 );
xor ( n244040 , n243911 , n243783 );
and ( n244041 , n244040 , n243970 );
and ( n244042 , n243911 , n243783 );
or ( n244043 , n244041 , n244042 );
xor ( n244044 , n244033 , n243789 );
xor ( n244045 , n244044 , n244039 );
xor ( n244046 , n244033 , n243789 );
and ( n244047 , n244046 , n244039 );
and ( n244048 , n244033 , n243789 );
or ( n244049 , n244047 , n244048 );
xor ( n244050 , n243795 , n244045 );
xor ( n244051 , n244050 , n243801 );
xor ( n244052 , n243795 , n244045 );
and ( n244053 , n244052 , n243801 );
and ( n244054 , n243795 , n244045 );
or ( n244055 , n244053 , n244054 );
xor ( n244056 , n243925 , n243934 );
and ( n244057 , n244056 , n243936 );
and ( n244058 , n243925 , n243934 );
or ( n244059 , n244057 , n244058 );
xor ( n244060 , n243985 , n243995 );
and ( n244061 , n244060 , n244006 );
and ( n244062 , n243985 , n243995 );
or ( n244063 , n244061 , n244062 );
xor ( n244064 , n243948 , n243953 );
and ( n244065 , n244064 , n243964 );
and ( n244066 , n243948 , n243953 );
or ( n244067 , n244065 , n244066 );
xor ( n244068 , n244017 , n244028 );
and ( n244069 , n244068 , n243589 );
and ( n244070 , n244017 , n244028 );
or ( n244071 , n244069 , n244070 );
xor ( n244072 , n243616 , n243811 );
and ( n244073 , n244072 , n243815 );
and ( n244074 , n243616 , n243811 );
or ( n244075 , n244073 , n244074 );
xor ( n244076 , n243867 , n243819 );
and ( n244077 , n244076 , n243823 );
and ( n244078 , n243867 , n243819 );
or ( n244079 , n244077 , n244078 );
xor ( n244080 , n243937 , n243903 );
and ( n244081 , n244080 , n243965 );
and ( n244082 , n243937 , n243903 );
or ( n244083 , n244081 , n244082 );
xor ( n244084 , n244007 , n244030 );
and ( n244085 , n244084 , n243827 );
and ( n244086 , n244007 , n244030 );
or ( n244087 , n244085 , n244086 );
not ( n244088 , n218232 );
not ( n244089 , n244088 );
not ( n244090 , n222002 );
or ( n244091 , n244089 , n244090 );
nand ( n244092 , n244091 , n224497 );
not ( n244093 , n224087 );
not ( n244094 , n243847 );
or ( n244095 , n244093 , n244094 );
not ( n244096 , n239903 );
not ( n244097 , n244096 );
not ( n244098 , n226961 );
or ( n244099 , n244097 , n244098 );
nand ( n244100 , n242471 , n239903 );
nand ( n244101 , n244099 , n244100 );
nand ( n244102 , n244101 , n227782 );
nand ( n244103 , n244095 , n244102 );
xor ( n244104 , n244092 , n244103 );
not ( n244105 , n238274 );
xor ( n244106 , n233465 , n236752 );
not ( n244107 , n244106 );
or ( n244108 , n244105 , n244107 );
nand ( n244109 , n243851 , n239270 );
nand ( n244110 , n244108 , n244109 );
xor ( n244111 , n244104 , n244110 );
xor ( n244112 , n244092 , n244103 );
and ( n244113 , n244112 , n244110 );
and ( n244114 , n244092 , n244103 );
or ( n244115 , n244113 , n244114 );
and ( n244116 , n238403 , n233891 );
not ( n244117 , n240020 );
not ( n244118 , n234878 );
not ( n244119 , n237600 );
or ( n244120 , n244118 , n244119 );
not ( n244121 , n234878 );
nand ( n244122 , n235031 , n244121 );
nand ( n244123 , n244120 , n244122 );
not ( n244124 , n244123 );
or ( n244125 , n244117 , n244124 );
nand ( n244126 , n243864 , n239492 );
nand ( n244127 , n244125 , n244126 );
xor ( n244128 , n244116 , n244127 );
not ( n244129 , n238776 );
not ( n244130 , n232494 );
not ( n244131 , n40415 );
not ( n244132 , n244131 );
or ( n244133 , n244130 , n244132 );
nand ( n244134 , n238362 , n229807 );
nand ( n244135 , n244133 , n244134 );
not ( n244136 , n244135 );
or ( n244137 , n244129 , n244136 );
not ( n244138 , n238999 );
nand ( n244139 , n243879 , n244138 );
nand ( n244140 , n244137 , n244139 );
xor ( n244141 , n244128 , n244140 );
xor ( n244142 , n244116 , n244127 );
and ( n244143 , n244142 , n244140 );
and ( n244144 , n244116 , n244127 );
or ( n244145 , n244143 , n244144 );
xor ( n244146 , n244071 , n244079 );
xor ( n244147 , n243871 , n243907 );
xor ( n244148 , n244147 , n244111 );
xor ( n244149 , n244146 , n244148 );
xor ( n244150 , n244071 , n244079 );
and ( n244151 , n244150 , n244148 );
and ( n244152 , n244071 , n244079 );
or ( n244153 , n244151 , n244152 );
not ( n244154 , n227852 );
and ( n244155 , n234293 , n221712 );
not ( n244156 , n234293 );
and ( n244157 , n244156 , n236719 );
nor ( n244158 , n244155 , n244157 );
not ( n244159 , n244158 );
or ( n244160 , n244154 , n244159 );
nand ( n244161 , n243887 , n239441 );
nand ( n244162 , n244160 , n244161 );
not ( n244163 , n238240 );
not ( n244164 , n236188 );
not ( n244165 , n220971 );
or ( n244166 , n244164 , n244165 );
nand ( n244167 , n40259 , n234394 );
nand ( n244168 , n244166 , n244167 );
not ( n244169 , n244168 );
or ( n244170 , n244163 , n244169 );
nand ( n244171 , n233446 , n243900 );
nand ( n244172 , n244170 , n244171 );
xor ( n244173 , n244162 , n244172 );
not ( n244174 , n228868 );
not ( n244175 , n238619 );
not ( n244176 , n221725 );
or ( n244177 , n244175 , n244176 );
nand ( n244178 , n234014 , n243058 );
nand ( n244179 , n244177 , n244178 );
not ( n244180 , n244179 );
or ( n244181 , n244174 , n244180 );
nand ( n244182 , n243921 , n243063 );
nand ( n244183 , n244181 , n244182 );
xor ( n244184 , n244173 , n244183 );
xor ( n244185 , n244184 , n244141 );
not ( n244186 , n243962 );
not ( n244187 , n221626 );
or ( n244188 , n244186 , n244187 );
and ( n244189 , n221778 , n235977 );
not ( n244190 , n221778 );
and ( n244191 , n244190 , n241369 );
or ( n244192 , n244189 , n244191 );
nand ( n244193 , n244192 , n221637 );
nand ( n244194 , n244188 , n244193 );
not ( n244195 , n220507 );
not ( n244196 , n244015 );
or ( n244197 , n244195 , n244196 );
and ( n244198 , n240917 , n243764 );
not ( n244199 , n240917 );
and ( n244200 , n244199 , n209709 );
nor ( n244201 , n244198 , n244200 );
nand ( n244202 , n244201 , n239530 );
nand ( n244203 , n244197 , n244202 );
xor ( n244204 , n244194 , n244203 );
not ( n244205 , n237503 );
not ( n244206 , n244026 );
or ( n244207 , n244205 , n244206 );
not ( n244208 , n240229 );
not ( n244209 , n241983 );
or ( n244210 , n244208 , n244209 );
nand ( n244211 , n225795 , n238719 );
nand ( n244212 , n244210 , n244211 );
nand ( n244213 , n244212 , n237493 );
nand ( n244214 , n244207 , n244213 );
xor ( n244215 , n244204 , n244214 );
xor ( n244216 , n244185 , n244215 );
xor ( n244217 , n244083 , n244216 );
xor ( n244218 , n244059 , n244063 );
xor ( n244219 , n244218 , n244067 );
xor ( n244220 , n244217 , n244219 );
xor ( n244221 , n244083 , n244216 );
and ( n244222 , n244221 , n244219 );
and ( n244223 , n244083 , n244216 );
or ( n244224 , n244222 , n244223 );
not ( n244225 , n242737 );
not ( n244226 , n239393 );
not ( n244227 , n234108 );
or ( n244228 , n244226 , n244227 );
nand ( n244229 , n40625 , n243314 );
nand ( n244230 , n244228 , n244229 );
not ( n244231 , n244230 );
or ( n244232 , n244225 , n244231 );
nand ( n244233 , n243931 , n234371 );
nand ( n244234 , n244232 , n244233 );
not ( n244235 , n238409 );
not ( n244236 , n243981 );
or ( n244237 , n244235 , n244236 );
nand ( n244238 , n239173 , n243326 );
not ( n244239 , n244238 );
not ( n244240 , n240581 );
nand ( n244241 , n244240 , n223182 );
not ( n244242 , n244241 );
or ( n244243 , n244239 , n244242 );
nand ( n244244 , n244243 , n227294 );
nand ( n244245 , n244237 , n244244 );
xor ( n244246 , n244234 , n244245 );
not ( n244247 , n239508 );
not ( n244248 , n243993 );
or ( n244249 , n244247 , n244248 );
and ( n244250 , n238363 , n239185 );
not ( n244251 , n238363 );
and ( n244252 , n244251 , n239186 );
nor ( n244253 , n244250 , n244252 );
not ( n244254 , n244253 );
nand ( n244255 , n244254 , n218843 );
nand ( n244256 , n244249 , n244255 );
xor ( n244257 , n244246 , n244256 );
not ( n244258 , n220164 );
not ( n244259 , n244002 );
or ( n244260 , n244258 , n244259 );
not ( n244261 , n236768 );
not ( n244262 , n238486 );
or ( n244263 , n244261 , n244262 );
nand ( n244264 , n236840 , n222414 );
nand ( n244265 , n244263 , n244264 );
nand ( n244266 , n244265 , n220881 );
nand ( n244267 , n244260 , n244266 );
not ( n244268 , n243936 );
xor ( n244269 , n244267 , n244268 );
not ( n244270 , n221674 );
not ( n244271 , n220906 );
not ( n244272 , n229704 );
or ( n244273 , n244271 , n244272 );
nand ( n244274 , n38532 , n239548 );
nand ( n244275 , n244273 , n244274 );
not ( n244276 , n244275 );
or ( n244277 , n244270 , n244276 );
nand ( n244278 , n243946 , n235913 );
nand ( n244279 , n244277 , n244278 );
xor ( n244280 , n244269 , n244279 );
xor ( n244281 , n244257 , n244280 );
xor ( n244282 , n244281 , n244075 );
xor ( n244283 , n244282 , n244087 );
xor ( n244284 , n244283 , n243915 );
xor ( n244285 , n244282 , n244087 );
and ( n244286 , n244285 , n243915 );
and ( n244287 , n244282 , n244087 );
or ( n244288 , n244286 , n244287 );
xor ( n244289 , n244149 , n243974 );
xor ( n244290 , n244289 , n244220 );
xor ( n244291 , n244149 , n243974 );
and ( n244292 , n244291 , n244220 );
and ( n244293 , n244149 , n243974 );
or ( n244294 , n244292 , n244293 );
xor ( n244295 , n244037 , n244284 );
xor ( n244296 , n244295 , n244290 );
xor ( n244297 , n244037 , n244284 );
and ( n244298 , n244297 , n244290 );
and ( n244299 , n244037 , n244284 );
or ( n244300 , n244298 , n244299 );
xor ( n244301 , n244043 , n244296 );
xor ( n244302 , n244301 , n244049 );
xor ( n244303 , n244043 , n244296 );
and ( n244304 , n244303 , n244049 );
and ( n244305 , n244043 , n244296 );
or ( n244306 , n244304 , n244305 );
xor ( n244307 , n244162 , n244172 );
and ( n244308 , n244307 , n244183 );
and ( n244309 , n244162 , n244172 );
or ( n244310 , n244308 , n244309 );
xor ( n244311 , n244234 , n244245 );
and ( n244312 , n244311 , n244256 );
and ( n244313 , n244234 , n244245 );
or ( n244314 , n244312 , n244313 );
xor ( n244315 , n244267 , n244268 );
and ( n244316 , n244315 , n244279 );
and ( n244317 , n244267 , n244268 );
or ( n244318 , n244316 , n244317 );
xor ( n244319 , n244194 , n244203 );
and ( n244320 , n244319 , n244214 );
and ( n244321 , n244194 , n244203 );
or ( n244322 , n244320 , n244321 );
xor ( n244323 , n243871 , n243907 );
and ( n244324 , n244323 , n244111 );
and ( n244325 , n243871 , n243907 );
or ( n244326 , n244324 , n244325 );
xor ( n244327 , n244059 , n244063 );
and ( n244328 , n244327 , n244067 );
and ( n244329 , n244059 , n244063 );
or ( n244330 , n244328 , n244329 );
xor ( n244331 , n244184 , n244141 );
and ( n244332 , n244331 , n244215 );
and ( n244333 , n244184 , n244141 );
or ( n244334 , n244332 , n244333 );
xor ( n244335 , n244257 , n244280 );
and ( n244336 , n244335 , n244075 );
and ( n244337 , n244257 , n244280 );
or ( n244338 , n244336 , n244337 );
not ( n244339 , n244138 );
not ( n244340 , n244135 );
or ( n244341 , n244339 , n244340 );
not ( n244342 , n229806 );
not ( n244343 , n238752 );
or ( n244344 , n244342 , n244343 );
nand ( n244345 , n239527 , n233962 );
nand ( n244346 , n244344 , n244345 );
nand ( n244347 , n244346 , n238776 );
nand ( n244348 , n244341 , n244347 );
and ( n244349 , n233891 , n208046 );
xor ( n244350 , n244348 , n244349 );
not ( n244351 , n237797 );
not ( n244352 , n244158 );
or ( n244353 , n244351 , n244352 );
not ( n244354 , n239774 );
not ( n244355 , n236301 );
or ( n244356 , n244354 , n244355 );
nand ( n244357 , n236304 , n234293 );
nand ( n244358 , n244356 , n244357 );
nand ( n244359 , n244358 , n242888 );
nand ( n244360 , n244353 , n244359 );
xor ( n244361 , n244350 , n244360 );
xor ( n244362 , n244348 , n244349 );
and ( n244363 , n244362 , n244360 );
and ( n244364 , n244348 , n244349 );
or ( n244365 , n244363 , n244364 );
not ( n244366 , n233446 );
not ( n244367 , n244168 );
or ( n244368 , n244366 , n244367 );
not ( n244369 , n236188 );
not ( n244370 , n226504 );
or ( n244371 , n244369 , n244370 );
nand ( n244372 , n230514 , n239787 );
nand ( n244373 , n244371 , n244372 );
nand ( n244374 , n238240 , n244373 );
nand ( n244375 , n244368 , n244374 );
not ( n244376 , n239794 );
not ( n244377 , n244179 );
or ( n244378 , n244376 , n244377 );
not ( n244379 , n228850 );
not ( n244380 , n223786 );
or ( n244381 , n244379 , n244380 );
nand ( n244382 , n221956 , n243058 );
nand ( n244383 , n244381 , n244382 );
nand ( n244384 , n228868 , n244383 );
nand ( n244385 , n244378 , n244384 );
xor ( n244386 , n244375 , n244385 );
buf ( n244387 , n234371 );
not ( n244388 , n244387 );
not ( n244389 , n244230 );
or ( n244390 , n244388 , n244389 );
not ( n244391 , n231480 );
not ( n244392 , n219742 );
or ( n244393 , n244391 , n244392 );
nand ( n244394 , n239470 , n233399 );
nand ( n244395 , n244393 , n244394 );
nand ( n244396 , n244395 , n234378 );
nand ( n244397 , n244390 , n244396 );
xor ( n244398 , n244386 , n244397 );
xor ( n244399 , n244375 , n244385 );
and ( n244400 , n244399 , n244397 );
and ( n244401 , n244375 , n244385 );
or ( n244402 , n244400 , n244401 );
xor ( n244403 , n244310 , n244314 );
xor ( n244404 , n244403 , n244318 );
xor ( n244405 , n244322 , n244398 );
xor ( n244406 , n244405 , n244361 );
xor ( n244407 , n244404 , n244406 );
xor ( n244408 , n244407 , n244334 );
xor ( n244409 , n244404 , n244406 );
and ( n244410 , n244409 , n244334 );
and ( n244411 , n244404 , n244406 );
or ( n244412 , n244410 , n244411 );
not ( n244413 , n222454 );
not ( n244414 , n244212 );
or ( n244415 , n244413 , n244414 );
not ( n244416 , n222430 );
not ( n244417 , n234324 );
or ( n244418 , n244416 , n244417 );
nand ( n244419 , n238877 , n238719 );
nand ( n244420 , n244418 , n244419 );
nand ( n244421 , n244420 , n237493 );
nand ( n244422 , n244415 , n244421 );
not ( n244423 , n220164 );
not ( n244424 , n244265 );
or ( n244425 , n244423 , n244424 );
not ( n244426 , n236768 );
not ( n244427 , n237271 );
or ( n244428 , n244426 , n244427 );
nand ( n244429 , n237272 , n222414 );
nand ( n244430 , n244428 , n244429 );
nand ( n244431 , n219779 , n244430 );
nand ( n244432 , n244425 , n244431 );
xor ( n244433 , n244422 , n244432 );
not ( n244434 , n238409 );
nand ( n244435 , n244238 , n244241 );
not ( n244436 , n244435 );
or ( n244437 , n244434 , n244436 );
not ( n244438 , n237005 );
not ( n244439 , n227224 );
or ( n244440 , n244438 , n244439 );
nand ( n244441 , n227223 , n243326 );
nand ( n244442 , n244440 , n244441 );
nand ( n244443 , n244442 , n222768 );
nand ( n244444 , n244437 , n244443 );
xor ( n244445 , n244433 , n244444 );
not ( n244446 , n239270 );
not ( n244447 , n244106 );
or ( n244448 , n244446 , n244447 );
xor ( n244449 , n240156 , n40562 );
nand ( n244450 , n238274 , n244449 );
nand ( n244451 , n244448 , n244450 );
not ( n244452 , n239495 );
not ( n244453 , n239899 );
not ( n244454 , n238728 );
or ( n244455 , n244453 , n244454 );
nand ( n244456 , n239608 , n239903 );
nand ( n244457 , n244455 , n244456 );
not ( n244458 , n244457 );
or ( n244459 , n244452 , n244458 );
nand ( n244460 , n244101 , n224087 );
nand ( n244461 , n244459 , n244460 );
xor ( n244462 , n244451 , n244461 );
not ( n244463 , n220507 );
not ( n244464 , n244201 );
or ( n244465 , n244463 , n244464 );
not ( n244466 , n236241 );
not ( n244467 , n234579 );
or ( n244468 , n244466 , n244467 );
nand ( n244469 , n209865 , n219420 );
nand ( n244470 , n244468 , n244469 );
nand ( n244471 , n244470 , n239530 );
nand ( n244472 , n244465 , n244471 );
xor ( n244473 , n244462 , n244472 );
xor ( n244474 , n244445 , n244473 );
not ( n244475 , n235913 );
not ( n244476 , n244275 );
or ( n244477 , n244475 , n244476 );
not ( n244478 , n222399 );
not ( n244479 , n39366 );
or ( n244480 , n244478 , n244479 );
not ( n244481 , n39364 );
nand ( n244482 , n244481 , n239548 );
nand ( n244483 , n244480 , n244482 );
nand ( n244484 , n244483 , n220930 );
nand ( n244485 , n244477 , n244484 );
not ( n244486 , n221637 );
not ( n244487 , n221608 );
not ( n244488 , n236382 );
or ( n244489 , n244487 , n244488 );
nand ( n244490 , n39089 , n221612 );
nand ( n244491 , n244489 , n244490 );
not ( n244492 , n244491 );
or ( n244493 , n244486 , n244492 );
nand ( n244494 , n244192 , n221626 );
nand ( n244495 , n244493 , n244494 );
xor ( n244496 , n244485 , n244495 );
or ( n244497 , n244253 , n239507 );
or ( n244498 , n221237 , n238363 );
nand ( n244499 , n244497 , n244498 );
xor ( n244500 , n244496 , n244499 );
xor ( n244501 , n244474 , n244500 );
xor ( n244502 , n244338 , n244501 );
xor ( n244503 , n244502 , n244153 );
xor ( n244504 , n244338 , n244501 );
and ( n244505 , n244504 , n244153 );
and ( n244506 , n244338 , n244501 );
or ( n244507 , n244505 , n244506 );
not ( n244508 , n239492 );
not ( n244509 , n244123 );
or ( n244510 , n244508 , n244509 );
not ( n244511 , n241287 );
not ( n244512 , n234503 );
or ( n244513 , n244511 , n244512 );
nand ( n244514 , n234506 , n234273 );
nand ( n244515 , n244513 , n244514 );
nand ( n244516 , n244515 , n240020 );
nand ( n244517 , n244510 , n244516 );
not ( n244518 , n244517 );
xor ( n244519 , n244518 , n244115 );
xor ( n244520 , n244519 , n244145 );
xor ( n244521 , n244330 , n244520 );
xor ( n244522 , n244521 , n244326 );
xor ( n244523 , n244224 , n244522 );
xor ( n244524 , n244523 , n244408 );
xor ( n244525 , n244224 , n244522 );
and ( n244526 , n244525 , n244408 );
and ( n244527 , n244224 , n244522 );
or ( n244528 , n244526 , n244527 );
xor ( n244529 , n244503 , n244288 );
xor ( n244530 , n244529 , n244294 );
xor ( n244531 , n244503 , n244288 );
and ( n244532 , n244531 , n244294 );
and ( n244533 , n244503 , n244288 );
or ( n244534 , n244532 , n244533 );
xor ( n244535 , n244524 , n244530 );
xor ( n244536 , n244535 , n244300 );
xor ( n244537 , n244524 , n244530 );
and ( n244538 , n244537 , n244300 );
and ( n244539 , n244524 , n244530 );
or ( n244540 , n244538 , n244539 );
xor ( n244541 , n244451 , n244461 );
and ( n244542 , n244541 , n244472 );
and ( n244543 , n244451 , n244461 );
or ( n244544 , n244542 , n244543 );
xor ( n244545 , n244485 , n244495 );
and ( n244546 , n244545 , n244499 );
and ( n244547 , n244485 , n244495 );
or ( n244548 , n244546 , n244547 );
xor ( n244549 , n244422 , n244432 );
and ( n244550 , n244549 , n244444 );
and ( n244551 , n244422 , n244432 );
or ( n244552 , n244550 , n244551 );
xor ( n244553 , n244518 , n244115 );
and ( n244554 , n244553 , n244145 );
and ( n244555 , n244518 , n244115 );
or ( n244556 , n244554 , n244555 );
xor ( n244557 , n244310 , n244314 );
and ( n244558 , n244557 , n244318 );
and ( n244559 , n244310 , n244314 );
or ( n244560 , n244558 , n244559 );
xor ( n244561 , n244322 , n244398 );
and ( n244562 , n244561 , n244361 );
and ( n244563 , n244322 , n244398 );
or ( n244564 , n244562 , n244563 );
xor ( n244565 , n244445 , n244473 );
and ( n244566 , n244565 , n244500 );
and ( n244567 , n244445 , n244473 );
or ( n244568 , n244566 , n244567 );
xor ( n244569 , n244330 , n244520 );
and ( n244570 , n244569 , n244326 );
and ( n244571 , n244330 , n244520 );
or ( n244572 , n244570 , n244571 );
not ( n244573 , n221237 );
not ( n244574 , n232421 );
or ( n244575 , n244573 , n244574 );
nand ( n244576 , n244575 , n221241 );
not ( n244577 , n240271 );
not ( n244578 , n244515 );
or ( n244579 , n244577 , n244578 );
not ( n244580 , n242653 );
not ( n244581 , n226961 );
or ( n244582 , n244580 , n244581 );
nand ( n244583 , n226964 , n244121 );
nand ( n244584 , n244582 , n244583 );
nand ( n244585 , n244584 , n240020 );
nand ( n244586 , n244579 , n244585 );
xor ( n244587 , n244576 , n244586 );
and ( n244588 , n233465 , n236752 );
xor ( n244589 , n244587 , n244588 );
xor ( n244590 , n244576 , n244586 );
and ( n244591 , n244590 , n244588 );
and ( n244592 , n244576 , n244586 );
or ( n244593 , n244591 , n244592 );
not ( n244594 , n228775 );
not ( n244595 , n225952 );
not ( n244596 , n237600 );
or ( n244597 , n244595 , n244596 );
nand ( n244598 , n40547 , n233962 );
nand ( n244599 , n244597 , n244598 );
not ( n244600 , n244599 );
or ( n244601 , n244594 , n244600 );
nand ( n244602 , n244346 , n244138 );
nand ( n244603 , n244601 , n244602 );
not ( n244604 , n242888 );
not ( n244605 , n239774 );
not ( n244606 , n244131 );
or ( n244607 , n244605 , n244606 );
nand ( n244608 , n239139 , n234293 );
nand ( n244609 , n244607 , n244608 );
not ( n244610 , n244609 );
or ( n244611 , n244604 , n244610 );
nand ( n244612 , n244358 , n237797 );
nand ( n244613 , n244611 , n244612 );
xor ( n244614 , n244603 , n244613 );
not ( n244615 , n238240 );
not ( n244616 , n236188 );
not ( n244617 , n221712 );
or ( n244618 , n244616 , n244617 );
nand ( n244619 , n238377 , n239787 );
nand ( n244620 , n244618 , n244619 );
not ( n244621 , n244620 );
or ( n244622 , n244615 , n244621 );
nand ( n244623 , n244373 , n237810 );
nand ( n244624 , n244622 , n244623 );
xor ( n244625 , n244614 , n244624 );
xor ( n244626 , n244603 , n244613 );
and ( n244627 , n244626 , n244624 );
and ( n244628 , n244603 , n244613 );
or ( n244629 , n244627 , n244628 );
xor ( n244630 , n244560 , n244568 );
xor ( n244631 , n244402 , n244589 );
xor ( n244632 , n244631 , n244544 );
xor ( n244633 , n244630 , n244632 );
xor ( n244634 , n244560 , n244568 );
and ( n244635 , n244634 , n244632 );
and ( n244636 , n244560 , n244568 );
or ( n244637 , n244635 , n244636 );
xor ( n244638 , n244548 , n244552 );
not ( n244639 , n228868 );
not ( n244640 , n228850 );
not ( n244641 , n239854 );
or ( n244642 , n244640 , n244641 );
not ( n244643 , n238619 );
nand ( n244644 , n40259 , n244643 );
nand ( n244645 , n244642 , n244644 );
not ( n244646 , n244645 );
or ( n244647 , n244639 , n244646 );
nand ( n244648 , n240120 , n244383 );
nand ( n244649 , n244647 , n244648 );
not ( n244650 , n234378 );
not ( n244651 , n239393 );
not ( n244652 , n239077 );
or ( n244653 , n244651 , n244652 );
not ( n244654 , n239393 );
nand ( n244655 , n239080 , n244654 );
nand ( n244656 , n244653 , n244655 );
not ( n244657 , n244656 );
or ( n244658 , n244650 , n244657 );
nand ( n244659 , n244395 , n234371 );
nand ( n244660 , n244658 , n244659 );
xor ( n244661 , n244649 , n244660 );
not ( n244662 , n239270 );
not ( n244663 , n244449 );
or ( n244664 , n244662 , n244663 );
xor ( n244665 , n233465 , n241891 );
nand ( n244666 , n244665 , n238274 );
nand ( n244667 , n244664 , n244666 );
xor ( n244668 , n244661 , n244667 );
xor ( n244669 , n244638 , n244668 );
not ( n244670 , n244491 );
not ( n244671 , n221626 );
or ( n244672 , n244670 , n244671 );
not ( n244673 , n221608 );
not ( n244674 , n235962 );
or ( n244675 , n244673 , n244674 );
nand ( n244676 , n38532 , n221612 );
nand ( n244677 , n244675 , n244676 );
nand ( n244678 , n244677 , n221637 );
nand ( n244679 , n244672 , n244678 );
not ( n244680 , n237493 );
and ( n244681 , n238719 , n243754 );
not ( n244682 , n238719 );
and ( n244683 , n244682 , n39608 );
nor ( n244684 , n244681 , n244683 );
not ( n244685 , n244684 );
or ( n244686 , n244680 , n244685 );
nand ( n244687 , n244420 , n237503 );
nand ( n244688 , n244686 , n244687 );
xor ( n244689 , n244679 , n244688 );
not ( n244690 , n220164 );
not ( n244691 , n244430 );
or ( n244692 , n244690 , n244691 );
not ( n244693 , n221593 );
not ( n244694 , n209709 );
or ( n244695 , n244693 , n244694 );
nand ( n244696 , n209710 , n222414 );
nand ( n244697 , n244695 , n244696 );
nand ( n244698 , n244697 , n219779 );
nand ( n244699 , n244692 , n244698 );
xor ( n244700 , n244689 , n244699 );
xor ( n244701 , n244625 , n244700 );
not ( n244702 , n219076 );
not ( n244703 , n236241 );
not ( n244704 , n234094 );
or ( n244705 , n244703 , n244704 );
nand ( n244706 , n209964 , n219420 );
nand ( n244707 , n244705 , n244706 );
not ( n244708 , n244707 );
or ( n244709 , n244702 , n244708 );
nand ( n244710 , n244470 , n220507 );
nand ( n244711 , n244709 , n244710 );
not ( n244712 , n224087 );
not ( n244713 , n244457 );
or ( n244714 , n244712 , n244713 );
and ( n244715 , n233018 , n239903 );
not ( n244716 , n233018 );
and ( n244717 , n244716 , n224096 );
or ( n244718 , n244715 , n244717 );
nand ( n244719 , n244718 , n227782 );
nand ( n244720 , n244714 , n244719 );
xor ( n244721 , n244711 , n244720 );
not ( n244722 , n220930 );
and ( n244723 , n236840 , n239066 );
not ( n244724 , n236840 );
and ( n244725 , n244724 , n220906 );
or ( n244726 , n244723 , n244725 );
not ( n244727 , n244726 );
or ( n244728 , n244722 , n244727 );
nand ( n244729 , n244483 , n235913 );
nand ( n244730 , n244728 , n244729 );
xor ( n244731 , n244721 , n244730 );
xor ( n244732 , n244701 , n244731 );
xor ( n244733 , n244669 , n244732 );
not ( n244734 , n222768 );
not ( n244735 , n238681 );
not ( n244736 , n210823 );
or ( n244737 , n244735 , n244736 );
nand ( n244738 , n227696 , n236547 );
nand ( n244739 , n244737 , n244738 );
not ( n244740 , n244739 );
or ( n244741 , n244734 , n244740 );
nand ( n244742 , n244442 , n238409 );
nand ( n244743 , n244741 , n244742 );
xor ( n244744 , n244743 , n244517 );
xor ( n244745 , n244744 , n244365 );
xor ( n244746 , n244745 , n244556 );
xor ( n244747 , n244746 , n244564 );
xor ( n244748 , n244733 , n244747 );
xor ( n244749 , n244669 , n244732 );
and ( n244750 , n244749 , n244747 );
and ( n244751 , n244669 , n244732 );
or ( n244752 , n244750 , n244751 );
xor ( n244753 , n244572 , n244412 );
xor ( n244754 , n244753 , n244633 );
xor ( n244755 , n244572 , n244412 );
and ( n244756 , n244755 , n244633 );
and ( n244757 , n244572 , n244412 );
or ( n244758 , n244756 , n244757 );
xor ( n244759 , n244748 , n244507 );
xor ( n244760 , n244759 , n244528 );
xor ( n244761 , n244748 , n244507 );
and ( n244762 , n244761 , n244528 );
and ( n244763 , n244748 , n244507 );
or ( n244764 , n244762 , n244763 );
xor ( n244765 , n244754 , n244760 );
xor ( n244766 , n244765 , n244534 );
xor ( n244767 , n244754 , n244760 );
and ( n244768 , n244767 , n244534 );
and ( n244769 , n244754 , n244760 );
or ( n244770 , n244768 , n244769 );
xor ( n244771 , n244649 , n244660 );
and ( n244772 , n244771 , n244667 );
and ( n244773 , n244649 , n244660 );
or ( n244774 , n244772 , n244773 );
xor ( n244775 , n244711 , n244720 );
and ( n244776 , n244775 , n244730 );
and ( n244777 , n244711 , n244720 );
or ( n244778 , n244776 , n244777 );
xor ( n244779 , n244679 , n244688 );
and ( n244780 , n244779 , n244699 );
and ( n244781 , n244679 , n244688 );
or ( n244782 , n244780 , n244781 );
xor ( n244783 , n244743 , n244517 );
and ( n244784 , n244783 , n244365 );
and ( n244785 , n244743 , n244517 );
or ( n244786 , n244784 , n244785 );
xor ( n244787 , n244402 , n244589 );
and ( n244788 , n244787 , n244544 );
and ( n244789 , n244402 , n244589 );
or ( n244790 , n244788 , n244789 );
xor ( n244791 , n244548 , n244552 );
and ( n244792 , n244791 , n244668 );
and ( n244793 , n244548 , n244552 );
or ( n244794 , n244792 , n244793 );
xor ( n244795 , n244625 , n244700 );
and ( n244796 , n244795 , n244731 );
and ( n244797 , n244625 , n244700 );
or ( n244798 , n244796 , n244797 );
xor ( n244799 , n244745 , n244556 );
and ( n244800 , n244799 , n244564 );
and ( n244801 , n244745 , n244556 );
or ( n244802 , n244800 , n244801 );
not ( n244803 , n237797 );
not ( n244804 , n244609 );
or ( n244805 , n244803 , n244804 );
not ( n244806 , n226651 );
not ( n244807 , n238752 );
or ( n244808 , n244806 , n244807 );
nand ( n244809 , n239527 , n226650 );
nand ( n244810 , n244808 , n244809 );
nand ( n244811 , n244810 , n227852 );
nand ( n244812 , n244805 , n244811 );
not ( n244813 , n237810 );
not ( n244814 , n244620 );
or ( n244815 , n244813 , n244814 );
not ( n244816 , n236188 );
not ( n244817 , n236301 );
or ( n244818 , n244816 , n244817 );
nand ( n244819 , n236304 , n239787 );
nand ( n244820 , n244818 , n244819 );
nand ( n244821 , n244820 , n238240 );
nand ( n244822 , n244815 , n244821 );
xor ( n244823 , n244812 , n244822 );
not ( n244824 , n239794 );
not ( n244825 , n244645 );
or ( n244826 , n244824 , n244825 );
not ( n244827 , n238617 );
not ( n244828 , n244827 );
not ( n244829 , n233546 );
or ( n244830 , n244828 , n244829 );
nand ( n244831 , n238789 , n244643 );
nand ( n244832 , n244830 , n244831 );
nand ( n244833 , n244832 , n228868 );
nand ( n244834 , n244826 , n244833 );
xor ( n244835 , n244823 , n244834 );
xor ( n244836 , n244812 , n244822 );
and ( n244837 , n244836 , n244834 );
and ( n244838 , n244812 , n244822 );
or ( n244839 , n244837 , n244838 );
not ( n244840 , n244387 );
not ( n244841 , n244656 );
or ( n244842 , n244840 , n244841 );
and ( n244843 , n239458 , n243314 );
not ( n244844 , n239458 );
and ( n244845 , n244844 , n231480 );
or ( n244846 , n244843 , n244845 );
nand ( n244847 , n244846 , n234378 );
nand ( n244848 , n244842 , n244847 );
not ( n244849 , n238274 );
xor ( n244850 , n233465 , n239470 );
not ( n244851 , n244850 );
or ( n244852 , n244849 , n244851 );
nand ( n244853 , n244665 , n239270 );
nand ( n244854 , n244852 , n244853 );
xor ( n244855 , n244848 , n244854 );
and ( n244856 , n240156 , n40562 );
xor ( n244857 , n244855 , n244856 );
xor ( n244858 , n244848 , n244854 );
and ( n244859 , n244858 , n244856 );
and ( n244860 , n244848 , n244854 );
or ( n244861 , n244859 , n244860 );
not ( n244862 , n235913 );
not ( n244863 , n244726 );
or ( n244864 , n244862 , n244863 );
not ( n244865 , n220906 );
not ( n244866 , n237271 );
or ( n244867 , n244865 , n244866 );
nand ( n244868 , n237272 , n239066 );
nand ( n244869 , n244867 , n244868 );
nand ( n244870 , n244869 , n221674 );
nand ( n244871 , n244864 , n244870 );
not ( n244872 , n239495 );
not ( n244873 , n244096 );
not ( n244874 , n234350 );
or ( n244875 , n244873 , n244874 );
nand ( n244876 , n227223 , n239903 );
nand ( n244877 , n244875 , n244876 );
not ( n244878 , n244877 );
or ( n244879 , n244872 , n244878 );
nand ( n244880 , n244718 , n224087 );
nand ( n244881 , n244879 , n244880 );
xor ( n244882 , n244871 , n244881 );
and ( n244883 , n244599 , n242335 );
not ( n244884 , n241599 );
not ( n244885 , n237963 );
not ( n244886 , n244885 );
or ( n244887 , n244884 , n244886 );
nand ( n244888 , n237963 , n232497 );
nand ( n244889 , n244887 , n244888 );
and ( n244890 , n244889 , n228775 );
nor ( n244891 , n244883 , n244890 );
xor ( n244892 , n244882 , n244891 );
xor ( n244893 , n244835 , n244892 );
not ( n244894 , n237503 );
not ( n244895 , n244684 );
or ( n244896 , n244894 , n244895 );
not ( n244897 , n222430 );
not ( n244898 , n236382 );
or ( n244899 , n244897 , n244898 );
nand ( n244900 , n39089 , n238719 );
nand ( n244901 , n244899 , n244900 );
nand ( n244902 , n244901 , n237493 );
nand ( n244903 , n244896 , n244902 );
not ( n244904 , n220507 );
not ( n244905 , n244707 );
or ( n244906 , n244904 , n244905 );
not ( n244907 , n219423 );
nand ( n244908 , n244907 , n239530 );
nand ( n244909 , n244906 , n244908 );
xor ( n244910 , n244903 , n244909 );
not ( n244911 , n238409 );
not ( n244912 , n244739 );
or ( n244913 , n244911 , n244912 );
not ( n244914 , n241712 );
not ( n244915 , n230241 );
or ( n244916 , n244914 , n244915 );
nand ( n244917 , n39747 , n243326 );
nand ( n244918 , n244916 , n244917 );
nand ( n244919 , n244918 , n222768 );
nand ( n244920 , n244913 , n244919 );
xor ( n244921 , n244910 , n244920 );
xor ( n244922 , n244893 , n244921 );
xor ( n244923 , n244798 , n244922 );
xor ( n244924 , n244923 , n244802 );
xor ( n244925 , n244798 , n244922 );
and ( n244926 , n244925 , n244802 );
and ( n244927 , n244798 , n244922 );
or ( n244928 , n244926 , n244927 );
not ( n244929 , n219779 );
not ( n244930 , n221593 );
not ( n244931 , n234579 );
or ( n244932 , n244930 , n244931 );
nand ( n244933 , n240358 , n222414 );
nand ( n244934 , n244932 , n244933 );
not ( n244935 , n244934 );
or ( n244936 , n244929 , n244935 );
nand ( n244937 , n244697 , n220164 );
nand ( n244938 , n244936 , n244937 );
not ( n244939 , n240020 );
and ( n244940 , n240617 , n235452 );
not ( n244941 , n240617 );
and ( n244942 , n244941 , n233525 );
nor ( n244943 , n244940 , n244942 );
not ( n244944 , n244943 );
or ( n244945 , n244939 , n244944 );
nand ( n244946 , n244584 , n240271 );
nand ( n244947 , n244945 , n244946 );
xor ( n244948 , n244938 , n244947 );
not ( n244949 , n239452 );
not ( n244950 , n244677 );
or ( n244951 , n244949 , n244950 );
not ( n244952 , n237937 );
not ( n244953 , n240372 );
or ( n244954 , n244952 , n244953 );
or ( n244955 , n240372 , n237937 );
nand ( n244956 , n244954 , n244955 );
nand ( n244957 , n244956 , n221637 );
nand ( n244958 , n244951 , n244957 );
xor ( n244959 , n244948 , n244958 );
xor ( n244960 , n244959 , n244786 );
xor ( n244961 , n244960 , n244794 );
xor ( n244962 , n244961 , n244637 );
xor ( n244963 , n244593 , n244629 );
xor ( n244964 , n244963 , n244774 );
xor ( n244965 , n244964 , n244790 );
xor ( n244966 , n244778 , n244782 );
xor ( n244967 , n244966 , n244857 );
xor ( n244968 , n244965 , n244967 );
xor ( n244969 , n244962 , n244968 );
xor ( n244970 , n244961 , n244637 );
and ( n244971 , n244970 , n244968 );
and ( n244972 , n244961 , n244637 );
or ( n244973 , n244971 , n244972 );
xor ( n244974 , n244752 , n244924 );
xor ( n244975 , n244974 , n244969 );
xor ( n244976 , n244752 , n244924 );
and ( n244977 , n244976 , n244969 );
and ( n244978 , n244752 , n244924 );
or ( n244979 , n244977 , n244978 );
xor ( n244980 , n244758 , n244975 );
xor ( n244981 , n244980 , n244764 );
xor ( n244982 , n244758 , n244975 );
and ( n244983 , n244982 , n244764 );
and ( n244984 , n244758 , n244975 );
or ( n244985 , n244983 , n244984 );
xor ( n244986 , n244938 , n244947 );
and ( n244987 , n244986 , n244958 );
and ( n244988 , n244938 , n244947 );
or ( n244989 , n244987 , n244988 );
xor ( n244990 , n244903 , n244909 );
and ( n244991 , n244990 , n244920 );
and ( n244992 , n244903 , n244909 );
or ( n244993 , n244991 , n244992 );
xor ( n244994 , n244871 , n244881 );
and ( n244995 , n244994 , n244891 );
and ( n244996 , n244871 , n244881 );
or ( n244997 , n244995 , n244996 );
xor ( n244998 , n244593 , n244629 );
and ( n244999 , n244998 , n244774 );
and ( n245000 , n244593 , n244629 );
or ( n245001 , n244999 , n245000 );
xor ( n245002 , n244778 , n244782 );
and ( n245003 , n245002 , n244857 );
and ( n245004 , n244778 , n244782 );
or ( n245005 , n245003 , n245004 );
xor ( n245006 , n244835 , n244892 );
and ( n245007 , n245006 , n244921 );
and ( n245008 , n244835 , n244892 );
or ( n245009 , n245007 , n245008 );
xor ( n245010 , n244959 , n244786 );
and ( n245011 , n245010 , n244794 );
and ( n245012 , n244959 , n244786 );
or ( n245013 , n245011 , n245012 );
xor ( n245014 , n244964 , n244790 );
and ( n245015 , n245014 , n244967 );
and ( n245016 , n244964 , n244790 );
or ( n245017 , n245015 , n245016 );
not ( n245018 , n229612 );
not ( n245019 , n219791 );
or ( n245020 , n245018 , n245019 );
nand ( n245021 , n245020 , n219800 );
not ( n245022 , n242335 );
not ( n245023 , n244889 );
or ( n245024 , n245022 , n245023 );
not ( n245025 , n241599 );
not ( n245026 , n242472 );
or ( n245027 , n245025 , n245026 );
nand ( n245028 , n242471 , n232497 );
nand ( n245029 , n245027 , n245028 );
nand ( n245030 , n245029 , n238776 );
nand ( n245031 , n245024 , n245030 );
xor ( n245032 , n245021 , n245031 );
not ( n245033 , n242888 );
not ( n245034 , n234295 );
not ( n245035 , n237600 );
or ( n245036 , n245034 , n245035 );
nand ( n245037 , n40547 , n226650 );
nand ( n245038 , n245036 , n245037 );
not ( n245039 , n245038 );
or ( n245040 , n245033 , n245039 );
nand ( n245041 , n244810 , n237797 );
nand ( n245042 , n245040 , n245041 );
xor ( n245043 , n245032 , n245042 );
xor ( n245044 , n245021 , n245031 );
and ( n245045 , n245044 , n245042 );
and ( n245046 , n245021 , n245031 );
or ( n245047 , n245045 , n245046 );
not ( n245048 , n237810 );
not ( n245049 , n244820 );
or ( n245050 , n245048 , n245049 );
not ( n245051 , n236188 );
not ( n245052 , n240637 );
or ( n245053 , n245051 , n245052 );
nand ( n245054 , n40415 , n239787 );
nand ( n245055 , n245053 , n245054 );
nand ( n245056 , n245055 , n238240 );
nand ( n245057 , n245050 , n245056 );
not ( n245058 , n228868 );
and ( n245059 , n244643 , n221712 );
not ( n245060 , n244643 );
and ( n245061 , n245060 , n40182 );
nor ( n245062 , n245059 , n245061 );
not ( n245063 , n245062 );
or ( n245064 , n245058 , n245063 );
nand ( n245065 , n244832 , n243063 );
nand ( n245066 , n245064 , n245065 );
xor ( n245067 , n245057 , n245066 );
not ( n245068 , n242737 );
not ( n245069 , n239393 );
not ( n245070 , n40258 );
or ( n245071 , n245069 , n245070 );
nand ( n245072 , n40259 , n244654 );
nand ( n245073 , n245071 , n245072 );
not ( n245074 , n245073 );
or ( n245075 , n245068 , n245074 );
nand ( n245076 , n244387 , n244846 );
nand ( n245077 , n245075 , n245076 );
xor ( n245078 , n245067 , n245077 );
xor ( n245079 , n245057 , n245066 );
and ( n245080 , n245079 , n245077 );
and ( n245081 , n245057 , n245066 );
or ( n245082 , n245080 , n245081 );
not ( n245083 , n238274 );
not ( n245084 , n221725 );
xor ( n245085 , n240156 , n245084 );
not ( n245086 , n245085 );
or ( n245087 , n245083 , n245086 );
nand ( n245088 , n244850 , n239270 );
nand ( n245089 , n245087 , n245088 );
and ( n245090 , n233465 , n241891 );
xor ( n245091 , n245089 , n245090 );
not ( n245092 , n219779 );
buf ( n245093 , n237643 );
and ( n245094 , n221593 , n245093 );
not ( n245095 , n221593 );
and ( n245096 , n245095 , n239186 );
nor ( n245097 , n245094 , n245096 );
not ( n245098 , n245097 );
or ( n245099 , n245092 , n245098 );
nand ( n245100 , n244934 , n220164 );
nand ( n245101 , n245099 , n245100 );
xor ( n245102 , n245091 , n245101 );
xor ( n245103 , n244989 , n245102 );
xor ( n245104 , n245103 , n244993 );
xor ( n245105 , n245043 , n245078 );
not ( n245106 , n227294 );
and ( n245107 , n243326 , n243754 );
not ( n245108 , n243326 );
and ( n245109 , n245108 , n235977 );
nor ( n245110 , n245107 , n245109 );
not ( n245111 , n245110 );
or ( n245112 , n245106 , n245111 );
nand ( n245113 , n244918 , n238409 );
nand ( n245114 , n245112 , n245113 );
not ( n245115 , n220930 );
not ( n245116 , n222399 );
not ( n245117 , n239952 );
or ( n245118 , n245116 , n245117 );
nand ( n245119 , n243764 , n239548 );
nand ( n245120 , n245118 , n245119 );
not ( n245121 , n245120 );
or ( n245122 , n245115 , n245121 );
nand ( n245123 , n244869 , n235913 );
nand ( n245124 , n245122 , n245123 );
xor ( n245125 , n245114 , n245124 );
not ( n245126 , n239495 );
not ( n245127 , n244096 );
not ( n245128 , n240738 );
or ( n245129 , n245127 , n245128 );
nand ( n245130 , n227696 , n239903 );
nand ( n245131 , n245129 , n245130 );
not ( n245132 , n245131 );
or ( n245133 , n245126 , n245132 );
nand ( n245134 , n244877 , n224087 );
nand ( n245135 , n245133 , n245134 );
xor ( n245136 , n245125 , n245135 );
xor ( n245137 , n245105 , n245136 );
xor ( n245138 , n245104 , n245137 );
not ( n245139 , n226724 );
nand ( n245140 , n245139 , n242653 );
not ( n245141 , n245140 );
not ( n245142 , n242653 );
not ( n245143 , n240581 );
and ( n245144 , n245142 , n245143 );
nor ( n245145 , n245144 , n236958 );
not ( n245146 , n245145 );
or ( n245147 , n245141 , n245146 );
nand ( n245148 , n244943 , n239492 );
nand ( n245149 , n245147 , n245148 );
not ( n245150 , n244956 );
not ( n245151 , n221626 );
or ( n245152 , n245150 , n245151 );
not ( n245153 , n237937 );
not ( n245154 , n238486 );
or ( n245155 , n245153 , n245154 );
nand ( n245156 , n236840 , n221612 );
nand ( n245157 , n245155 , n245156 );
nand ( n245158 , n245157 , n221637 );
nand ( n245159 , n245152 , n245158 );
xor ( n245160 , n245149 , n245159 );
not ( n245161 , n237493 );
not ( n245162 , n222430 );
not ( n245163 , n235962 );
or ( n245164 , n245162 , n245163 );
nand ( n245165 , n38532 , n244024 );
nand ( n245166 , n245164 , n245165 );
not ( n245167 , n245166 );
or ( n245168 , n245161 , n245167 );
nand ( n245169 , n244901 , n222454 );
nand ( n245170 , n245168 , n245169 );
xor ( n245171 , n245160 , n245170 );
xor ( n245172 , n245171 , n244997 );
xor ( n245173 , n245172 , n245001 );
xor ( n245174 , n245138 , n245173 );
xor ( n245175 , n245104 , n245137 );
and ( n245176 , n245175 , n245173 );
and ( n245177 , n245104 , n245137 );
or ( n245178 , n245176 , n245177 );
xor ( n245179 , n245013 , n245017 );
not ( n245180 , n244891 );
xor ( n245181 , n245180 , n244839 );
xor ( n245182 , n245181 , n244861 );
xor ( n245183 , n245005 , n245182 );
xor ( n245184 , n245183 , n245009 );
xor ( n245185 , n245179 , n245184 );
xor ( n245186 , n245013 , n245017 );
and ( n245187 , n245186 , n245184 );
and ( n245188 , n245013 , n245017 );
or ( n245189 , n245187 , n245188 );
xor ( n245190 , n245174 , n244928 );
xor ( n245191 , n245190 , n244973 );
xor ( n245192 , n245174 , n244928 );
and ( n245193 , n245192 , n244973 );
and ( n245194 , n245174 , n244928 );
or ( n245195 , n245193 , n245194 );
xor ( n245196 , n245185 , n245191 );
xor ( n245197 , n245196 , n244979 );
xor ( n245198 , n245185 , n245191 );
and ( n245199 , n245198 , n244979 );
and ( n245200 , n245185 , n245191 );
or ( n245201 , n245199 , n245200 );
xor ( n245202 , n245089 , n245090 );
and ( n245203 , n245202 , n245101 );
and ( n245204 , n245089 , n245090 );
or ( n245205 , n245203 , n245204 );
xor ( n245206 , n245149 , n245159 );
and ( n245207 , n245206 , n245170 );
and ( n245208 , n245149 , n245159 );
or ( n245209 , n245207 , n245208 );
xor ( n245210 , n245114 , n245124 );
and ( n245211 , n245210 , n245135 );
and ( n245212 , n245114 , n245124 );
or ( n245213 , n245211 , n245212 );
xor ( n245214 , n245180 , n244839 );
and ( n245215 , n245214 , n244861 );
and ( n245216 , n245180 , n244839 );
or ( n245217 , n245215 , n245216 );
xor ( n245218 , n244989 , n245102 );
and ( n245219 , n245218 , n244993 );
and ( n245220 , n244989 , n245102 );
or ( n245221 , n245219 , n245220 );
xor ( n245222 , n245043 , n245078 );
and ( n245223 , n245222 , n245136 );
and ( n245224 , n245043 , n245078 );
or ( n245225 , n245223 , n245224 );
xor ( n245226 , n245171 , n244997 );
and ( n245227 , n245226 , n245001 );
and ( n245228 , n245171 , n244997 );
or ( n245229 , n245227 , n245228 );
xor ( n245230 , n245005 , n245182 );
and ( n245231 , n245230 , n245009 );
and ( n245232 , n245005 , n245182 );
or ( n245233 , n245231 , n245232 );
not ( n245234 , n239794 );
not ( n245235 , n245062 );
or ( n245236 , n245234 , n245235 );
not ( n245237 , n244827 );
not ( n245238 , n224700 );
or ( n245239 , n245237 , n245238 );
not ( n245240 , n236301 );
nand ( n245241 , n245240 , n238617 );
nand ( n245242 , n245239 , n245241 );
nand ( n245243 , n245242 , n228868 );
nand ( n245244 , n245236 , n245243 );
not ( n245245 , n237797 );
not ( n245246 , n245038 );
or ( n245247 , n245245 , n245246 );
not ( n245248 , n239774 );
not ( n245249 , n244885 );
or ( n245250 , n245248 , n245249 );
nand ( n245251 , n237963 , n238230 );
nand ( n245252 , n245250 , n245251 );
nand ( n245253 , n245252 , n242888 );
nand ( n245254 , n245247 , n245253 );
xor ( n245255 , n245244 , n245254 );
not ( n245256 , n239270 );
not ( n245257 , n245085 );
or ( n245258 , n245256 , n245257 );
xor ( n245259 , n239458 , n239281 );
nand ( n245260 , n245259 , n238274 );
nand ( n245261 , n245258 , n245260 );
xor ( n245262 , n245255 , n245261 );
xor ( n245263 , n245244 , n245254 );
and ( n245264 , n245263 , n245261 );
and ( n245265 , n245244 , n245254 );
or ( n245266 , n245264 , n245265 );
not ( n245267 , n244387 );
not ( n245268 , n245073 );
or ( n245269 , n245267 , n245268 );
not ( n245270 , n239393 );
not ( n245271 , n230511 );
or ( n245272 , n245270 , n245271 );
buf ( n245273 , n226505 );
nand ( n245274 , n245273 , n244654 );
nand ( n245275 , n245272 , n245274 );
nand ( n245276 , n245275 , n242737 );
nand ( n245277 , n245269 , n245276 );
and ( n245278 , n233465 , n239470 );
xor ( n245279 , n245277 , n245278 );
not ( n245280 , n221674 );
not ( n245281 , n222399 );
not ( n245282 , n209866 );
not ( n245283 , n245282 );
or ( n245284 , n245281 , n245283 );
nand ( n245285 , n209866 , n239548 );
nand ( n245286 , n245284 , n245285 );
not ( n245287 , n245286 );
or ( n245288 , n245280 , n245287 );
nand ( n245289 , n245120 , n235913 );
nand ( n245290 , n245288 , n245289 );
xor ( n245291 , n245279 , n245290 );
xor ( n245292 , n245277 , n245278 );
and ( n245293 , n245292 , n245290 );
and ( n245294 , n245277 , n245278 );
or ( n245295 , n245293 , n245294 );
not ( n245296 , n220164 );
not ( n245297 , n245097 );
or ( n245298 , n245296 , n245297 );
nand ( n245299 , n220881 , n236768 );
nand ( n245300 , n245298 , n245299 );
not ( n245301 , n224087 );
not ( n245302 , n245131 );
or ( n245303 , n245301 , n245302 );
not ( n245304 , n239899 );
not ( n245305 , n235516 );
or ( n245306 , n245304 , n245305 );
nand ( n245307 , n39747 , n238672 );
nand ( n245308 , n245306 , n245307 );
nand ( n245309 , n245308 , n239495 );
nand ( n245310 , n245303 , n245309 );
xor ( n245311 , n245300 , n245310 );
not ( n245312 , n221637 );
not ( n245313 , n237937 );
not ( n245314 , n237271 );
or ( n245315 , n245313 , n245314 );
nand ( n245316 , n237272 , n221778 );
nand ( n245317 , n245315 , n245316 );
not ( n245318 , n245317 );
or ( n245319 , n245312 , n245318 );
nand ( n245320 , n245157 , n239452 );
nand ( n245321 , n245319 , n245320 );
xor ( n245322 , n245311 , n245321 );
not ( n245323 , n238776 );
not ( n245324 , n232494 );
not ( n245325 , n242904 );
or ( n245326 , n245324 , n245325 );
nand ( n245327 , n39880 , n232493 );
nand ( n245328 , n245326 , n245327 );
not ( n245329 , n245328 );
or ( n245330 , n245323 , n245329 );
nand ( n245331 , n245029 , n242335 );
nand ( n245332 , n245330 , n245331 );
not ( n245333 , n222454 );
not ( n245334 , n245166 );
or ( n245335 , n245333 , n245334 );
not ( n245336 , n240229 );
not ( n245337 , n240372 );
or ( n245338 , n245336 , n245337 );
nand ( n245339 , n240375 , n244024 );
nand ( n245340 , n245338 , n245339 );
nand ( n245341 , n245340 , n237493 );
nand ( n245342 , n245335 , n245341 );
xor ( n245343 , n245332 , n245342 );
not ( n245344 , n245110 );
not ( n245345 , n238409 );
or ( n245346 , n245344 , n245345 );
not ( n245347 , n241712 );
not ( n245348 , n227201 );
or ( n245349 , n245347 , n245348 );
nand ( n245350 , n238857 , n236547 );
nand ( n245351 , n245349 , n245350 );
nand ( n245352 , n245351 , n227294 );
nand ( n245353 , n245346 , n245352 );
xor ( n245354 , n245343 , n245353 );
xor ( n245355 , n245322 , n245354 );
and ( n245356 , n242653 , n239173 );
not ( n245357 , n242653 );
and ( n245358 , n245357 , n244240 );
nor ( n245359 , n245356 , n245358 );
nand ( n245360 , n245359 , n239492 );
and ( n245361 , n234878 , n242210 );
not ( n245362 , n234878 );
and ( n245363 , n245362 , n242858 );
or ( n245364 , n245361 , n245363 );
nand ( n245365 , n245364 , n240020 );
nand ( n245366 , n245360 , n245365 );
not ( n245367 , n237810 );
not ( n245368 , n245055 );
or ( n245369 , n245367 , n245368 );
not ( n245370 , n242596 );
not ( n245371 , n238752 );
or ( n245372 , n245370 , n245371 );
nand ( n245373 , n239527 , n240500 );
nand ( n245374 , n245372 , n245373 );
nand ( n245375 , n245374 , n238240 );
nand ( n245376 , n245369 , n245375 );
not ( n245377 , n245376 );
xor ( n245378 , n245366 , n245377 );
xor ( n245379 , n245378 , n245047 );
xor ( n245380 , n245355 , n245379 );
xor ( n245381 , n245380 , n245233 );
xor ( n245382 , n245217 , n245221 );
xor ( n245383 , n245082 , n245209 );
xor ( n245384 , n245383 , n245205 );
xor ( n245385 , n245382 , n245384 );
xor ( n245386 , n245381 , n245385 );
xor ( n245387 , n245380 , n245233 );
and ( n245388 , n245387 , n245385 );
and ( n245389 , n245380 , n245233 );
or ( n245390 , n245388 , n245389 );
xor ( n245391 , n245213 , n245291 );
xor ( n245392 , n245391 , n245262 );
xor ( n245393 , n245392 , n245225 );
xor ( n245394 , n245393 , n245229 );
xor ( n245395 , n245178 , n245394 );
xor ( n245396 , n245395 , n245189 );
xor ( n245397 , n245178 , n245394 );
and ( n245398 , n245397 , n245189 );
and ( n245399 , n245178 , n245394 );
or ( n245400 , n245398 , n245399 );
xor ( n245401 , n245386 , n245396 );
xor ( n245402 , n245401 , n245195 );
xor ( n245403 , n245386 , n245396 );
and ( n245404 , n245403 , n245195 );
and ( n245405 , n245386 , n245396 );
or ( n245406 , n245404 , n245405 );
xor ( n245407 , n245332 , n245342 );
and ( n245408 , n245407 , n245353 );
and ( n245409 , n245332 , n245342 );
or ( n245410 , n245408 , n245409 );
xor ( n245411 , n245300 , n245310 );
and ( n245412 , n245411 , n245321 );
and ( n245413 , n245300 , n245310 );
or ( n245414 , n245412 , n245413 );
xor ( n245415 , n245366 , n245377 );
and ( n245416 , n245415 , n245047 );
and ( n245417 , n245366 , n245377 );
or ( n245418 , n245416 , n245417 );
xor ( n245419 , n245082 , n245209 );
and ( n245420 , n245419 , n245205 );
and ( n245421 , n245082 , n245209 );
or ( n245422 , n245420 , n245421 );
xor ( n245423 , n245213 , n245291 );
and ( n245424 , n245423 , n245262 );
and ( n245425 , n245213 , n245291 );
or ( n245426 , n245424 , n245425 );
xor ( n245427 , n245322 , n245354 );
and ( n245428 , n245427 , n245379 );
and ( n245429 , n245322 , n245354 );
or ( n245430 , n245428 , n245429 );
xor ( n245431 , n245217 , n245221 );
and ( n245432 , n245431 , n245384 );
and ( n245433 , n245217 , n245221 );
or ( n245434 , n245432 , n245433 );
xor ( n245435 , n245392 , n245225 );
and ( n245436 , n245435 , n245229 );
and ( n245437 , n245392 , n245225 );
or ( n245438 , n245436 , n245437 );
not ( n245439 , n224171 );
not ( n245440 , n237895 );
or ( n245441 , n245439 , n245440 );
nand ( n245442 , n245441 , n236768 );
not ( n245443 , n239441 );
not ( n245444 , n245252 );
or ( n245445 , n245443 , n245444 );
not ( n245446 , n226651 );
not ( n245447 , n242472 );
or ( n245448 , n245446 , n245447 );
nand ( n245449 , n242471 , n238230 );
nand ( n245450 , n245448 , n245449 );
nand ( n245451 , n245450 , n242888 );
nand ( n245452 , n245445 , n245451 );
xor ( n245453 , n245442 , n245452 );
not ( n245454 , n238240 );
not ( n245455 , n242596 );
not ( n245456 , n237600 );
or ( n245457 , n245455 , n245456 );
not ( n245458 , n237816 );
nand ( n245459 , n235031 , n245458 );
nand ( n245460 , n245457 , n245459 );
not ( n245461 , n245460 );
or ( n245462 , n245454 , n245461 );
nand ( n245463 , n245374 , n237810 );
nand ( n245464 , n245462 , n245463 );
xor ( n245465 , n245453 , n245464 );
xor ( n245466 , n245442 , n245452 );
and ( n245467 , n245466 , n245464 );
and ( n245468 , n245442 , n245452 );
or ( n245469 , n245467 , n245468 );
not ( n245470 , n243063 );
not ( n245471 , n245242 );
or ( n245472 , n245470 , n245471 );
not ( n245473 , n238619 );
not ( n245474 , n244131 );
or ( n245475 , n245473 , n245474 );
nand ( n245476 , n40415 , n231940 );
nand ( n245477 , n245475 , n245476 );
nand ( n245478 , n245477 , n228868 );
nand ( n245479 , n245472 , n245478 );
not ( n245480 , n244387 );
not ( n245481 , n245275 );
or ( n245482 , n245480 , n245481 );
not ( n245483 , n231480 );
not ( n245484 , n240589 );
or ( n245485 , n245483 , n245484 );
nand ( n245486 , n236719 , n243314 );
nand ( n245487 , n245485 , n245486 );
nand ( n245488 , n245487 , n242737 );
nand ( n245489 , n245482 , n245488 );
xor ( n245490 , n245479 , n245489 );
not ( n245491 , n238274 );
xor ( n245492 , n234382 , n40259 );
not ( n245493 , n245492 );
or ( n245494 , n245491 , n245493 );
nand ( n245495 , n239270 , n245259 );
nand ( n245496 , n245494 , n245495 );
xor ( n245497 , n245490 , n245496 );
xor ( n245498 , n245479 , n245489 );
and ( n245499 , n245498 , n245496 );
and ( n245500 , n245479 , n245489 );
or ( n245501 , n245499 , n245500 );
not ( n245502 , n221637 );
not ( n245503 , n237937 );
not ( n245504 , n238449 );
or ( n245505 , n245503 , n245504 );
nand ( n245506 , n209710 , n221778 );
nand ( n245507 , n245505 , n245506 );
not ( n245508 , n245507 );
or ( n245509 , n245502 , n245508 );
nand ( n245510 , n245317 , n239452 );
nand ( n245511 , n245509 , n245510 );
not ( n245512 , n240020 );
not ( n245513 , n234878 );
not ( n245514 , n210823 );
or ( n245515 , n245513 , n245514 );
nand ( n245516 , n227696 , n244121 );
nand ( n245517 , n245515 , n245516 );
not ( n245518 , n245517 );
or ( n245519 , n245512 , n245518 );
nand ( n245520 , n245364 , n240271 );
nand ( n245521 , n245519 , n245520 );
xor ( n245522 , n245511 , n245521 );
xor ( n245523 , n245522 , n245376 );
and ( n245524 , n240156 , n245084 );
not ( n245525 , n221674 );
not ( n245526 , n222399 );
not ( n245527 , n209965 );
or ( n245528 , n245526 , n245527 );
not ( n245529 , n209965 );
nand ( n245530 , n245529 , n239548 );
nand ( n245531 , n245528 , n245530 );
not ( n245532 , n245531 );
or ( n245533 , n245525 , n245532 );
nand ( n245534 , n245286 , n235913 );
nand ( n245535 , n245533 , n245534 );
xor ( n245536 , n245524 , n245535 );
not ( n245537 , n244138 );
not ( n245538 , n245328 );
or ( n245539 , n245537 , n245538 );
not ( n245540 , n232494 );
not ( n245541 , n39928 );
or ( n245542 , n245540 , n245541 );
nand ( n245543 , n39929 , n232493 );
nand ( n245544 , n245542 , n245543 );
nand ( n245545 , n245544 , n238776 );
nand ( n245546 , n245539 , n245545 );
xor ( n245547 , n245536 , n245546 );
xor ( n245548 , n245523 , n245547 );
not ( n245549 , n237493 );
not ( n245550 , n240229 );
not ( n245551 , n238486 );
or ( n245552 , n245550 , n245551 );
nand ( n245553 , n39288 , n244024 );
nand ( n245554 , n245552 , n245553 );
not ( n245555 , n245554 );
or ( n245556 , n245549 , n245555 );
nand ( n245557 , n245340 , n237503 );
nand ( n245558 , n245556 , n245557 );
not ( n245559 , n227294 );
not ( n245560 , n235962 );
not ( n245561 , n238681 );
or ( n245562 , n245560 , n245561 );
nand ( n245563 , n38532 , n236547 );
nand ( n245564 , n245562 , n245563 );
not ( n245565 , n245564 );
or ( n245566 , n245559 , n245565 );
nand ( n245567 , n245351 , n238409 );
nand ( n245568 , n245566 , n245567 );
xor ( n245569 , n245558 , n245568 );
not ( n245570 , n239495 );
not ( n245571 , n244096 );
not ( n245572 , n243754 );
or ( n245573 , n245571 , n245572 );
nand ( n245574 , n39608 , n238672 );
nand ( n245575 , n245573 , n245574 );
not ( n245576 , n245575 );
or ( n245577 , n245570 , n245576 );
nand ( n245578 , n245308 , n224087 );
nand ( n245579 , n245577 , n245578 );
xor ( n245580 , n245569 , n245579 );
xor ( n245581 , n245548 , n245580 );
xor ( n245582 , n245581 , n245434 );
xor ( n245583 , n245418 , n245426 );
xor ( n245584 , n245583 , n245422 );
xor ( n245585 , n245582 , n245584 );
xor ( n245586 , n245581 , n245434 );
and ( n245587 , n245586 , n245584 );
and ( n245588 , n245581 , n245434 );
or ( n245589 , n245587 , n245588 );
xor ( n245590 , n245266 , n245410 );
xor ( n245591 , n245590 , n245295 );
xor ( n245592 , n245497 , n245414 );
xor ( n245593 , n245592 , n245465 );
xor ( n245594 , n245591 , n245593 );
xor ( n245595 , n245594 , n245430 );
xor ( n245596 , n245595 , n245438 );
xor ( n245597 , n245596 , n245390 );
xor ( n245598 , n245595 , n245438 );
and ( n245599 , n245598 , n245390 );
and ( n245600 , n245595 , n245438 );
or ( n245601 , n245599 , n245600 );
xor ( n245602 , n245585 , n245597 );
xor ( n245603 , n245602 , n245400 );
xor ( n245604 , n245585 , n245597 );
and ( n245605 , n245604 , n245400 );
and ( n245606 , n245585 , n245597 );
or ( n245607 , n245605 , n245606 );
xor ( n245608 , n245524 , n245535 );
and ( n245609 , n245608 , n245546 );
and ( n245610 , n245524 , n245535 );
or ( n245611 , n245609 , n245610 );
xor ( n245612 , n245558 , n245568 );
and ( n245613 , n245612 , n245579 );
and ( n245614 , n245558 , n245568 );
or ( n245615 , n245613 , n245614 );
xor ( n245616 , n245511 , n245521 );
and ( n245617 , n245616 , n245376 );
and ( n245618 , n245511 , n245521 );
or ( n245619 , n245617 , n245618 );
xor ( n245620 , n245266 , n245410 );
and ( n245621 , n245620 , n245295 );
and ( n245622 , n245266 , n245410 );
or ( n245623 , n245621 , n245622 );
xor ( n245624 , n245497 , n245414 );
and ( n245625 , n245624 , n245465 );
and ( n245626 , n245497 , n245414 );
or ( n245627 , n245625 , n245626 );
xor ( n245628 , n245523 , n245547 );
and ( n245629 , n245628 , n245580 );
and ( n245630 , n245523 , n245547 );
or ( n245631 , n245629 , n245630 );
xor ( n245632 , n245418 , n245426 );
and ( n245633 , n245632 , n245422 );
and ( n245634 , n245418 , n245426 );
or ( n245635 , n245633 , n245634 );
xor ( n245636 , n245591 , n245593 );
and ( n245637 , n245636 , n245430 );
and ( n245638 , n245591 , n245593 );
or ( n245639 , n245637 , n245638 );
not ( n245640 , n244387 );
not ( n245641 , n245487 );
or ( n245642 , n245640 , n245641 );
not ( n245643 , n243314 );
not ( n245644 , n222101 );
or ( n245645 , n245643 , n245644 );
nand ( n245646 , n231480 , n235383 );
nand ( n245647 , n245645 , n245646 );
nand ( n245648 , n245647 , n234378 );
nand ( n245649 , n245642 , n245648 );
not ( n245650 , n237810 );
not ( n245651 , n245460 );
or ( n245652 , n245650 , n245651 );
not ( n245653 , n242596 );
not ( n245654 , n244885 );
or ( n245655 , n245653 , n245654 );
nand ( n245656 , n237963 , n240500 );
nand ( n245657 , n245655 , n245656 );
nand ( n245658 , n245657 , n238240 );
nand ( n245659 , n245652 , n245658 );
xor ( n245660 , n245649 , n245659 );
and ( n245661 , n239458 , n239281 );
xor ( n245662 , n245660 , n245661 );
xor ( n245663 , n245649 , n245659 );
and ( n245664 , n245663 , n245661 );
and ( n245665 , n245649 , n245659 );
or ( n245666 , n245664 , n245665 );
not ( n245667 , n239270 );
not ( n245668 , n245492 );
or ( n245669 , n245667 , n245668 );
xor ( n245670 , n236615 , n226505 );
nand ( n245671 , n245670 , n238274 );
nand ( n245672 , n245669 , n245671 );
not ( n245673 , n221637 );
and ( n245674 , n222035 , n209865 );
not ( n245675 , n222035 );
and ( n245676 , n245675 , n239617 );
nor ( n245677 , n245674 , n245676 );
not ( n245678 , n245677 );
or ( n245679 , n245673 , n245678 );
nand ( n245680 , n245507 , n239452 );
nand ( n245681 , n245679 , n245680 );
xor ( n245682 , n245672 , n245681 );
not ( n245683 , n242888 );
not ( n245684 , n226651 );
not ( n245685 , n242904 );
or ( n245686 , n245684 , n245685 );
nand ( n245687 , n39880 , n238230 );
nand ( n245688 , n245686 , n245687 );
not ( n245689 , n245688 );
or ( n245690 , n245683 , n245689 );
nand ( n245691 , n245450 , n239441 );
nand ( n245692 , n245690 , n245691 );
xor ( n245693 , n245682 , n245692 );
xor ( n245694 , n245672 , n245681 );
and ( n245695 , n245694 , n245692 );
and ( n245696 , n245672 , n245681 );
or ( n245697 , n245695 , n245696 );
xor ( n245698 , n245623 , n245631 );
xor ( n245699 , n245611 , n245662 );
xor ( n245700 , n245699 , n245615 );
xor ( n245701 , n245698 , n245700 );
xor ( n245702 , n245639 , n245701 );
not ( n245703 , n240271 );
not ( n245704 , n245517 );
or ( n245705 , n245703 , n245704 );
not ( n245706 , n234878 );
not ( n245707 , n39748 );
or ( n245708 , n245706 , n245707 );
nand ( n245709 , n238877 , n244121 );
nand ( n245710 , n245708 , n245709 );
nand ( n245711 , n245710 , n240020 );
nand ( n245712 , n245705 , n245711 );
not ( n245713 , n222454 );
not ( n245714 , n245554 );
or ( n245715 , n245713 , n245714 );
not ( n245716 , n240229 );
not ( n245717 , n237271 );
or ( n245718 , n245716 , n245717 );
nand ( n245719 , n237272 , n244024 );
nand ( n245720 , n245718 , n245719 );
nand ( n245721 , n245720 , n237493 );
nand ( n245722 , n245715 , n245721 );
xor ( n245723 , n245712 , n245722 );
not ( n245724 , n244138 );
not ( n245725 , n245544 );
or ( n245726 , n245724 , n245725 );
not ( n245727 , n232494 );
not ( n245728 , n242210 );
or ( n245729 , n245727 , n245728 );
nand ( n245730 , n242858 , n232493 );
nand ( n245731 , n245729 , n245730 );
nand ( n245732 , n245731 , n238776 );
nand ( n245733 , n245726 , n245732 );
xor ( n245734 , n245723 , n245733 );
xor ( n245735 , n245734 , n245693 );
not ( n245736 , n223182 );
not ( n245737 , n240372 );
or ( n245738 , n245736 , n245737 );
nand ( n245739 , n240375 , n243326 );
nand ( n245740 , n245738 , n245739 );
not ( n245741 , n245740 );
not ( n245742 , n227294 );
or ( n245743 , n245741 , n245742 );
nand ( n245744 , n245564 , n238409 );
nand ( n245745 , n245743 , n245744 );
not ( n245746 , n224087 );
not ( n245747 , n245575 );
or ( n245748 , n245746 , n245747 );
not ( n245749 , n239899 );
not ( n245750 , n227201 );
or ( n245751 , n245749 , n245750 );
nand ( n245752 , n238857 , n238672 );
nand ( n245753 , n245751 , n245752 );
nand ( n245754 , n245753 , n239495 );
nand ( n245755 , n245748 , n245754 );
xor ( n245756 , n245745 , n245755 );
not ( n245757 , n221674 );
not ( n245758 , n222399 );
or ( n245759 , n245757 , n245758 );
not ( n245760 , n245531 );
not ( n245761 , n235913 );
or ( n245762 , n245760 , n245761 );
nand ( n245763 , n245759 , n245762 );
xor ( n245764 , n245756 , n245763 );
xor ( n245765 , n245735 , n245764 );
xor ( n245766 , n245765 , n245635 );
not ( n245767 , n228868 );
xnor ( n245768 , n238619 , n238752 );
not ( n245769 , n245768 );
or ( n245770 , n245767 , n245769 );
nand ( n245771 , n245477 , n239794 );
nand ( n245772 , n245770 , n245771 );
not ( n245773 , n245772 );
xor ( n245774 , n245773 , n245501 );
xor ( n245775 , n245774 , n245469 );
xor ( n245776 , n245619 , n245775 );
xor ( n245777 , n245776 , n245627 );
xor ( n245778 , n245766 , n245777 );
xor ( n245779 , n245702 , n245778 );
xor ( n245780 , n245639 , n245701 );
and ( n245781 , n245780 , n245778 );
and ( n245782 , n245639 , n245701 );
or ( n245783 , n245781 , n245782 );
xor ( n245784 , n245589 , n245779 );
xor ( n245785 , n245784 , n245601 );
xor ( n245786 , n245589 , n245779 );
and ( n245787 , n245786 , n245601 );
and ( n245788 , n245589 , n245779 );
or ( n245789 , n245787 , n245788 );
xor ( n245790 , n245745 , n245755 );
and ( n245791 , n245790 , n245763 );
and ( n245792 , n245745 , n245755 );
or ( n245793 , n245791 , n245792 );
xor ( n245794 , n245712 , n245722 );
and ( n245795 , n245794 , n245733 );
and ( n245796 , n245712 , n245722 );
or ( n245797 , n245795 , n245796 );
xor ( n245798 , n245773 , n245501 );
and ( n245799 , n245798 , n245469 );
and ( n245800 , n245773 , n245501 );
or ( n245801 , n245799 , n245800 );
xor ( n245802 , n245611 , n245662 );
and ( n245803 , n245802 , n245615 );
and ( n245804 , n245611 , n245662 );
or ( n245805 , n245803 , n245804 );
xor ( n245806 , n245734 , n245693 );
and ( n245807 , n245806 , n245764 );
and ( n245808 , n245734 , n245693 );
or ( n245809 , n245807 , n245808 );
xor ( n245810 , n245619 , n245775 );
and ( n245811 , n245810 , n245627 );
and ( n245812 , n245619 , n245775 );
or ( n245813 , n245811 , n245812 );
xor ( n245814 , n245623 , n245631 );
and ( n245815 , n245814 , n245700 );
and ( n245816 , n245623 , n245631 );
or ( n245817 , n245815 , n245816 );
xor ( n245818 , n245765 , n245635 );
and ( n245819 , n245818 , n245777 );
and ( n245820 , n245765 , n245635 );
or ( n245821 , n245819 , n245820 );
not ( n245822 , n220930 );
not ( n245823 , n245822 );
not ( n245824 , n245761 );
or ( n245825 , n245823 , n245824 );
nand ( n245826 , n245825 , n222399 );
not ( n245827 , n237810 );
not ( n245828 , n245657 );
or ( n245829 , n245827 , n245828 );
and ( n245830 , n237816 , n226961 );
not ( n245831 , n237816 );
and ( n245832 , n245831 , n242471 );
or ( n245833 , n245830 , n245832 );
nand ( n245834 , n245833 , n238240 );
nand ( n245835 , n245829 , n245834 );
xor ( n245836 , n245826 , n245835 );
not ( n245837 , n228868 );
not ( n245838 , n228850 );
not ( n245839 , n237600 );
or ( n245840 , n245838 , n245839 );
not ( n245841 , n238619 );
nand ( n245842 , n245841 , n235031 );
nand ( n245843 , n245840 , n245842 );
not ( n245844 , n245843 );
or ( n245845 , n245837 , n245844 );
nand ( n245846 , n245768 , n243063 );
nand ( n245847 , n245845 , n245846 );
xor ( n245848 , n245836 , n245847 );
xor ( n245849 , n245826 , n245835 );
and ( n245850 , n245849 , n245847 );
and ( n245851 , n245826 , n245835 );
or ( n245852 , n245850 , n245851 );
not ( n245853 , n242737 );
not ( n245854 , n239393 );
not ( n245855 , n244131 );
or ( n245856 , n245854 , n245855 );
nand ( n245857 , n239139 , n244654 );
nand ( n245858 , n245856 , n245857 );
not ( n245859 , n245858 );
or ( n245860 , n245853 , n245859 );
nand ( n245861 , n245647 , n244387 );
nand ( n245862 , n245860 , n245861 );
not ( n245863 , n239270 );
not ( n245864 , n245670 );
or ( n245865 , n245863 , n245864 );
xor ( n245866 , n233465 , n236719 );
nand ( n245867 , n245866 , n238274 );
nand ( n245868 , n245865 , n245867 );
xor ( n245869 , n245862 , n245868 );
and ( n245870 , n234382 , n40259 );
xor ( n245871 , n245869 , n245870 );
xor ( n245872 , n245862 , n245868 );
and ( n245873 , n245872 , n245870 );
and ( n245874 , n245862 , n245868 );
or ( n245875 , n245873 , n245874 );
xor ( n245876 , n245805 , n245809 );
xor ( n245877 , n245871 , n245848 );
not ( n245878 , n221626 );
not ( n245879 , n245677 );
or ( n245880 , n245878 , n245879 );
and ( n245881 , n221612 , n239186 );
not ( n245882 , n221612 );
and ( n245883 , n245882 , n245093 );
nor ( n245884 , n245881 , n245883 );
nand ( n245885 , n245884 , n221637 );
nand ( n245886 , n245880 , n245885 );
not ( n245887 , n239441 );
not ( n245888 , n245688 );
or ( n245889 , n245887 , n245888 );
and ( n245890 , n226723 , n226650 );
not ( n245891 , n226723 );
and ( n245892 , n245891 , n226651 );
or ( n245893 , n245890 , n245892 );
nand ( n245894 , n245893 , n242888 );
nand ( n245895 , n245889 , n245894 );
xor ( n245896 , n245886 , n245895 );
not ( n245897 , n227294 );
not ( n245898 , n223182 );
not ( n245899 , n238486 );
or ( n245900 , n245898 , n245899 );
nand ( n245901 , n236840 , n243326 );
nand ( n245902 , n245900 , n245901 );
not ( n245903 , n245902 );
or ( n245904 , n245897 , n245903 );
nand ( n245905 , n245740 , n238409 );
nand ( n245906 , n245904 , n245905 );
xor ( n245907 , n245896 , n245906 );
xor ( n245908 , n245877 , n245907 );
xor ( n245909 , n245876 , n245908 );
xor ( n245910 , n245817 , n245909 );
xor ( n245911 , n245697 , n245793 );
xor ( n245912 , n245911 , n245797 );
xor ( n245913 , n245912 , n245813 );
not ( n245914 , n239495 );
not ( n245915 , n239899 );
not ( n245916 , n235962 );
or ( n245917 , n245915 , n245916 );
nand ( n245918 , n239932 , n239903 );
nand ( n245919 , n245917 , n245918 );
not ( n245920 , n245919 );
or ( n245921 , n245914 , n245920 );
nand ( n245922 , n245753 , n224087 );
nand ( n245923 , n245921 , n245922 );
not ( n245924 , n240020 );
and ( n245925 , n244121 , n240710 );
not ( n245926 , n244121 );
and ( n245927 , n245926 , n235977 );
nor ( n245928 , n245925 , n245927 );
not ( n245929 , n245928 );
or ( n245930 , n245924 , n245929 );
nand ( n245931 , n245710 , n240271 );
nand ( n245932 , n245930 , n245931 );
xor ( n245933 , n245923 , n245932 );
not ( n245934 , n237503 );
not ( n245935 , n245720 );
or ( n245936 , n245934 , n245935 );
not ( n245937 , n222430 );
not ( n245938 , n243765 );
or ( n245939 , n245937 , n245938 );
nand ( n245940 , n243764 , n238719 );
nand ( n245941 , n245939 , n245940 );
nand ( n245942 , n245941 , n237493 );
nand ( n245943 , n245936 , n245942 );
xor ( n245944 , n245933 , n245943 );
not ( n245945 , n238776 );
and ( n245946 , n241599 , n227696 );
not ( n245947 , n241599 );
and ( n245948 , n245947 , n239214 );
nor ( n245949 , n245946 , n245948 );
not ( n245950 , n245949 );
or ( n245951 , n245945 , n245950 );
nand ( n245952 , n245731 , n244138 );
nand ( n245953 , n245951 , n245952 );
xor ( n245954 , n245953 , n245772 );
xor ( n245955 , n245954 , n245666 );
xor ( n245956 , n245944 , n245955 );
xor ( n245957 , n245956 , n245801 );
xor ( n245958 , n245913 , n245957 );
xor ( n245959 , n245910 , n245958 );
xor ( n245960 , n245817 , n245909 );
and ( n245961 , n245960 , n245958 );
and ( n245962 , n245817 , n245909 );
or ( n245963 , n245961 , n245962 );
xor ( n245964 , n245821 , n245959 );
xor ( n245965 , n245964 , n245783 );
xor ( n245966 , n245821 , n245959 );
and ( n245967 , n245966 , n245783 );
and ( n245968 , n245821 , n245959 );
or ( n245969 , n245967 , n245968 );
xor ( n245970 , n245886 , n245895 );
and ( n245971 , n245970 , n245906 );
and ( n245972 , n245886 , n245895 );
or ( n245973 , n245971 , n245972 );
xor ( n245974 , n245923 , n245932 );
and ( n245975 , n245974 , n245943 );
and ( n245976 , n245923 , n245932 );
or ( n245977 , n245975 , n245976 );
xor ( n245978 , n245953 , n245772 );
and ( n245979 , n245978 , n245666 );
and ( n245980 , n245953 , n245772 );
or ( n245981 , n245979 , n245980 );
xor ( n245982 , n245697 , n245793 );
and ( n245983 , n245982 , n245797 );
and ( n245984 , n245697 , n245793 );
or ( n245985 , n245983 , n245984 );
xor ( n245986 , n245871 , n245848 );
and ( n245987 , n245986 , n245907 );
and ( n245988 , n245871 , n245848 );
or ( n245989 , n245987 , n245988 );
xor ( n245990 , n245944 , n245955 );
and ( n245991 , n245990 , n245801 );
and ( n245992 , n245944 , n245955 );
or ( n245993 , n245991 , n245992 );
xor ( n245994 , n245805 , n245809 );
and ( n245995 , n245994 , n245908 );
and ( n245996 , n245805 , n245809 );
or ( n245997 , n245995 , n245996 );
xor ( n245998 , n245912 , n245813 );
and ( n245999 , n245998 , n245957 );
and ( n246000 , n245912 , n245813 );
or ( n246001 , n245999 , n246000 );
not ( n246002 , n239270 );
not ( n246003 , n245866 );
or ( n246004 , n246002 , n246003 );
xor ( n246005 , n233465 , n236300 );
nand ( n246006 , n246005 , n238274 );
nand ( n246007 , n246004 , n246006 );
not ( n246008 , n239794 );
not ( n246009 , n245843 );
or ( n246010 , n246008 , n246009 );
not ( n246011 , n238619 );
not ( n246012 , n230490 );
or ( n246013 , n246011 , n246012 );
nand ( n246014 , n237963 , n243058 );
nand ( n246015 , n246013 , n246014 );
nand ( n246016 , n246015 , n228868 );
nand ( n246017 , n246010 , n246016 );
xor ( n246018 , n246007 , n246017 );
and ( n246019 , n236615 , n226505 );
xor ( n246020 , n246018 , n246019 );
xor ( n246021 , n246007 , n246017 );
and ( n246022 , n246021 , n246019 );
and ( n246023 , n246007 , n246017 );
or ( n246024 , n246022 , n246023 );
not ( n246025 , n222454 );
not ( n246026 , n245941 );
or ( n246027 , n246025 , n246026 );
not ( n246028 , n222430 );
not ( n246029 , n239617 );
or ( n246030 , n246028 , n246029 );
nand ( n246031 , n209866 , n238719 );
nand ( n246032 , n246030 , n246031 );
nand ( n246033 , n246032 , n237493 );
nand ( n246034 , n246027 , n246033 );
not ( n246035 , n238240 );
not ( n246036 , n242596 );
not ( n246037 , n242904 );
or ( n246038 , n246036 , n246037 );
nand ( n246039 , n39880 , n239787 );
nand ( n246040 , n246038 , n246039 );
not ( n246041 , n246040 );
or ( n246042 , n246035 , n246041 );
nand ( n246043 , n245833 , n237810 );
nand ( n246044 , n246042 , n246043 );
xor ( n246045 , n246034 , n246044 );
not ( n246046 , n224087 );
not ( n246047 , n245919 );
or ( n246048 , n246046 , n246047 );
not ( n246049 , n244096 );
not ( n246050 , n240372 );
or ( n246051 , n246049 , n246050 );
nand ( n246052 , n240375 , n239903 );
nand ( n246053 , n246051 , n246052 );
nand ( n246054 , n246053 , n239495 );
nand ( n246055 , n246048 , n246054 );
xor ( n246056 , n246045 , n246055 );
xor ( n246057 , n246034 , n246044 );
and ( n246058 , n246057 , n246055 );
and ( n246059 , n246034 , n246044 );
or ( n246060 , n246058 , n246059 );
xor ( n246061 , n245852 , n245875 );
xor ( n246062 , n246061 , n246020 );
xor ( n246063 , n245985 , n246062 );
xor ( n246064 , n246063 , n245989 );
xor ( n246065 , n246064 , n245997 );
xor ( n246066 , n245973 , n245977 );
not ( n246067 , n240271 );
not ( n246068 , n245928 );
or ( n246069 , n246067 , n246068 );
not ( n246070 , n242653 );
not ( n246071 , n236382 );
or ( n246072 , n246070 , n246071 );
nand ( n246073 , n39089 , n234273 );
nand ( n246074 , n246072 , n246073 );
nand ( n246075 , n246074 , n240020 );
nand ( n246076 , n246069 , n246075 );
not ( n246077 , n239452 );
not ( n246078 , n245884 );
or ( n246079 , n246077 , n246078 );
not ( n246080 , n221612 );
nand ( n246081 , n246080 , n221637 );
nand ( n246082 , n246079 , n246081 );
xor ( n246083 , n246076 , n246082 );
not ( n246084 , n244138 );
not ( n246085 , n245949 );
or ( n246086 , n246084 , n246085 );
not ( n246087 , n241599 );
not ( n246088 , n39748 );
or ( n246089 , n246087 , n246088 );
nand ( n246090 , n39747 , n233962 );
nand ( n246091 , n246089 , n246090 );
nand ( n246092 , n246091 , n238776 );
nand ( n246093 , n246086 , n246092 );
xor ( n246094 , n246083 , n246093 );
xor ( n246095 , n246066 , n246094 );
not ( n246096 , n238409 );
not ( n246097 , n245902 );
or ( n246098 , n246096 , n246097 );
not ( n246099 , n237005 );
not ( n246100 , n237271 );
or ( n246101 , n246099 , n246100 );
nand ( n246102 , n238887 , n243326 );
nand ( n246103 , n246101 , n246102 );
nand ( n246104 , n246103 , n227294 );
nand ( n246105 , n246098 , n246104 );
not ( n246106 , n239441 );
not ( n246107 , n245893 );
or ( n246108 , n246106 , n246107 );
not ( n246109 , n226651 );
not ( n246110 , n227224 );
or ( n246111 , n246109 , n246110 );
nand ( n246112 , n242858 , n234293 );
nand ( n246113 , n246111 , n246112 );
nand ( n246114 , n246113 , n242888 );
nand ( n246115 , n246108 , n246114 );
xor ( n246116 , n246105 , n246115 );
not ( n246117 , n244387 );
not ( n246118 , n245858 );
or ( n246119 , n246117 , n246118 );
not ( n246120 , n239393 );
not ( n246121 , n222940 );
or ( n246122 , n246120 , n246121 );
nand ( n246123 , n236290 , n243314 );
nand ( n246124 , n246122 , n246123 );
nand ( n246125 , n246124 , n234378 );
nand ( n246126 , n246119 , n246125 );
not ( n246127 , n246126 );
xor ( n246128 , n246116 , n246127 );
xor ( n246129 , n246056 , n246128 );
xor ( n246130 , n246129 , n245981 );
xor ( n246131 , n246095 , n246130 );
xor ( n246132 , n246131 , n245993 );
xor ( n246133 , n246065 , n246132 );
xor ( n246134 , n246001 , n246133 );
xor ( n246135 , n246134 , n245963 );
xor ( n246136 , n246001 , n246133 );
and ( n246137 , n246136 , n245963 );
and ( n246138 , n246001 , n246133 );
or ( n246139 , n246137 , n246138 );
xor ( n246140 , n246076 , n246082 );
and ( n246141 , n246140 , n246093 );
and ( n246142 , n246076 , n246082 );
or ( n246143 , n246141 , n246142 );
xor ( n246144 , n246105 , n246115 );
and ( n246145 , n246144 , n246127 );
and ( n246146 , n246105 , n246115 );
or ( n246147 , n246145 , n246146 );
xor ( n246148 , n245852 , n245875 );
and ( n246149 , n246148 , n246020 );
and ( n246150 , n245852 , n245875 );
or ( n246151 , n246149 , n246150 );
xor ( n246152 , n245973 , n245977 );
and ( n246153 , n246152 , n246094 );
and ( n246154 , n245973 , n245977 );
or ( n246155 , n246153 , n246154 );
xor ( n246156 , n246056 , n246128 );
and ( n246157 , n246156 , n245981 );
and ( n246158 , n246056 , n246128 );
or ( n246159 , n246157 , n246158 );
xor ( n246160 , n245985 , n246062 );
and ( n246161 , n246160 , n245989 );
and ( n246162 , n245985 , n246062 );
or ( n246163 , n246161 , n246162 );
xor ( n246164 , n246095 , n246130 );
and ( n246165 , n246164 , n245993 );
and ( n246166 , n246095 , n246130 );
or ( n246167 , n246165 , n246166 );
xor ( n246168 , n246064 , n245997 );
and ( n246169 , n246168 , n246132 );
and ( n246170 , n246064 , n245997 );
or ( n246171 , n246169 , n246170 );
not ( n246172 , n221636 );
not ( n246173 , n222471 );
or ( n246174 , n246172 , n246173 );
nand ( n246175 , n246174 , n238705 );
not ( n246176 , n239794 );
not ( n246177 , n246015 );
or ( n246178 , n246176 , n246177 );
not ( n246179 , n228850 );
not ( n246180 , n226961 );
or ( n246181 , n246179 , n246180 );
not ( n246182 , n238619 );
nand ( n246183 , n246182 , n242471 );
nand ( n246184 , n246181 , n246183 );
nand ( n246185 , n246184 , n228868 );
nand ( n246186 , n246178 , n246185 );
xor ( n246187 , n246175 , n246186 );
not ( n246188 , n242737 );
not ( n246189 , n239393 );
not ( n246190 , n237600 );
or ( n246191 , n246189 , n246190 );
nand ( n246192 , n235031 , n244654 );
nand ( n246193 , n246191 , n246192 );
not ( n246194 , n246193 );
or ( n246195 , n246188 , n246194 );
nand ( n246196 , n246124 , n244387 );
nand ( n246197 , n246195 , n246196 );
xor ( n246198 , n246187 , n246197 );
xor ( n246199 , n246175 , n246186 );
and ( n246200 , n246199 , n246197 );
and ( n246201 , n246175 , n246186 );
or ( n246202 , n246200 , n246201 );
not ( n246203 , n238274 );
xor ( n246204 , n234382 , n239139 );
not ( n246205 , n246204 );
or ( n246206 , n246203 , n246205 );
nand ( n246207 , n246005 , n233105 );
nand ( n246208 , n246206 , n246207 );
and ( n246209 , n233465 , n236719 );
xor ( n246210 , n246208 , n246209 );
not ( n246211 , n237493 );
not ( n246212 , n222430 );
not ( n246213 , n239186 );
or ( n246214 , n246212 , n246213 );
nand ( n246215 , n245093 , n238719 );
nand ( n246216 , n246214 , n246215 );
not ( n246217 , n246216 );
or ( n246218 , n246211 , n246217 );
nand ( n246219 , n246032 , n237503 );
nand ( n246220 , n246218 , n246219 );
xor ( n246221 , n246210 , n246220 );
xor ( n246222 , n246208 , n246209 );
and ( n246223 , n246222 , n246220 );
and ( n246224 , n246208 , n246209 );
or ( n246225 , n246223 , n246224 );
xor ( n246226 , n246221 , n246198 );
xor ( n246227 , n246226 , n246060 );
xor ( n246228 , n246227 , n246159 );
not ( n246229 , n222768 );
and ( n246230 , n238681 , n209710 );
not ( n246231 , n238681 );
and ( n246232 , n246231 , n238449 );
nor ( n246233 , n246230 , n246232 );
not ( n246234 , n246233 );
or ( n246235 , n246229 , n246234 );
nand ( n246236 , n246103 , n238409 );
nand ( n246237 , n246235 , n246236 );
not ( n246238 , n238776 );
and ( n246239 , n233962 , n243754 );
not ( n246240 , n233962 );
and ( n246241 , n246240 , n235977 );
nor ( n246242 , n246239 , n246241 );
not ( n246243 , n246242 );
or ( n246244 , n246238 , n246243 );
nand ( n246245 , n246091 , n242335 );
nand ( n246246 , n246244 , n246245 );
xor ( n246247 , n246237 , n246246 );
not ( n246248 , n242888 );
not ( n246249 , n239774 );
not ( n246250 , n210823 );
or ( n246251 , n246249 , n246250 );
nand ( n246252 , n227696 , n238230 );
nand ( n246253 , n246251 , n246252 );
not ( n246254 , n246253 );
or ( n246255 , n246248 , n246254 );
nand ( n246256 , n246113 , n239441 );
nand ( n246257 , n246255 , n246256 );
xor ( n246258 , n246247 , n246257 );
xor ( n246259 , n246147 , n246258 );
not ( n246260 , n237810 );
not ( n246261 , n246040 );
or ( n246262 , n246260 , n246261 );
and ( n246263 , n239787 , n226723 );
not ( n246264 , n239787 );
and ( n246265 , n246264 , n240578 );
or ( n246266 , n246263 , n246265 );
nand ( n246267 , n246266 , n238240 );
nand ( n246268 , n246262 , n246267 );
not ( n246269 , n224087 );
not ( n246270 , n246053 );
or ( n246271 , n246269 , n246270 );
not ( n246272 , n239899 );
not ( n246273 , n238486 );
or ( n246274 , n246272 , n246273 );
not ( n246275 , n244096 );
nand ( n246276 , n246275 , n39288 );
nand ( n246277 , n246274 , n246276 );
nand ( n246278 , n246277 , n239495 );
nand ( n246279 , n246271 , n246278 );
xor ( n246280 , n246268 , n246279 );
not ( n246281 , n240020 );
not ( n246282 , n234878 );
not ( n246283 , n229704 );
or ( n246284 , n246282 , n246283 );
nand ( n246285 , n239932 , n237918 );
nand ( n246286 , n246284 , n246285 );
not ( n246287 , n246286 );
or ( n246288 , n246281 , n246287 );
nand ( n246289 , n246074 , n239492 );
nand ( n246290 , n246288 , n246289 );
xor ( n246291 , n246280 , n246290 );
xor ( n246292 , n246259 , n246291 );
xor ( n246293 , n246228 , n246292 );
xor ( n246294 , n246126 , n246024 );
xor ( n246295 , n246294 , n246143 );
xor ( n246296 , n246295 , n246151 );
xor ( n246297 , n246296 , n246155 );
xor ( n246298 , n246297 , n246163 );
xor ( n246299 , n246298 , n246167 );
xor ( n246300 , n246293 , n246299 );
xor ( n246301 , n246300 , n246171 );
xor ( n246302 , n246293 , n246299 );
and ( n246303 , n246302 , n246171 );
and ( n246304 , n246293 , n246299 );
or ( n246305 , n246303 , n246304 );
xor ( n246306 , n246268 , n246279 );
and ( n246307 , n246306 , n246290 );
and ( n246308 , n246268 , n246279 );
or ( n246309 , n246307 , n246308 );
xor ( n246310 , n246237 , n246246 );
and ( n246311 , n246310 , n246257 );
and ( n246312 , n246237 , n246246 );
or ( n246313 , n246311 , n246312 );
xor ( n246314 , n246126 , n246024 );
and ( n246315 , n246314 , n246143 );
and ( n246316 , n246126 , n246024 );
or ( n246317 , n246315 , n246316 );
xor ( n246318 , n246221 , n246198 );
and ( n246319 , n246318 , n246060 );
and ( n246320 , n246221 , n246198 );
or ( n246321 , n246319 , n246320 );
xor ( n246322 , n246147 , n246258 );
and ( n246323 , n246322 , n246291 );
and ( n246324 , n246147 , n246258 );
or ( n246325 , n246323 , n246324 );
xor ( n246326 , n246295 , n246151 );
and ( n246327 , n246326 , n246155 );
and ( n246328 , n246295 , n246151 );
or ( n246329 , n246327 , n246328 );
xor ( n246330 , n246227 , n246159 );
and ( n246331 , n246330 , n246292 );
and ( n246332 , n246227 , n246159 );
or ( n246333 , n246331 , n246332 );
xor ( n246334 , n246297 , n246163 );
and ( n246335 , n246334 , n246167 );
and ( n246336 , n246297 , n246163 );
or ( n246337 , n246335 , n246336 );
and ( n246338 , n233465 , n236300 );
and ( n246339 , n230490 , n239393 );
not ( n246340 , n230490 );
and ( n246341 , n246340 , n244654 );
or ( n246342 , n246339 , n246341 );
not ( n246343 , n246342 );
not ( n246344 , n242737 );
or ( n246345 , n246343 , n246344 );
nand ( n246346 , n244387 , n246193 );
nand ( n246347 , n246345 , n246346 );
xor ( n246348 , n246338 , n246347 );
not ( n246349 , n238409 );
not ( n246350 , n246233 );
or ( n246351 , n246349 , n246350 );
not ( n246352 , n237005 );
not ( n246353 , n245282 );
or ( n246354 , n246352 , n246353 );
nand ( n246355 , n209866 , n236547 );
nand ( n246356 , n246354 , n246355 );
nand ( n246357 , n246356 , n227294 );
nand ( n246358 , n246351 , n246357 );
xor ( n246359 , n246348 , n246358 );
xor ( n246360 , n246338 , n246347 );
and ( n246361 , n246360 , n246358 );
and ( n246362 , n246338 , n246347 );
or ( n246363 , n246361 , n246362 );
not ( n246364 , n228868 );
not ( n246365 , n238619 );
not ( n246366 , n242904 );
or ( n246367 , n246365 , n246366 );
nand ( n246368 , n233525 , n244643 );
nand ( n246369 , n246367 , n246368 );
not ( n246370 , n246369 );
or ( n246371 , n246364 , n246370 );
nand ( n246372 , n246184 , n243063 );
nand ( n246373 , n246371 , n246372 );
not ( n246374 , n240020 );
and ( n246375 , n244121 , n39367 );
not ( n246376 , n244121 );
not ( n246377 , n39367 );
and ( n246378 , n246376 , n246377 );
nor ( n246379 , n246375 , n246378 );
not ( n246380 , n246379 );
or ( n246381 , n246374 , n246380 );
nand ( n246382 , n246286 , n239492 );
nand ( n246383 , n246381 , n246382 );
xor ( n246384 , n246373 , n246383 );
not ( n246385 , n244138 );
not ( n246386 , n246242 );
or ( n246387 , n246385 , n246386 );
not ( n246388 , n232494 );
not ( n246389 , n227201 );
or ( n246390 , n246388 , n246389 );
nand ( n246391 , n238857 , n232493 );
nand ( n246392 , n246390 , n246391 );
nand ( n246393 , n246392 , n238776 );
nand ( n246394 , n246387 , n246393 );
xor ( n246395 , n246384 , n246394 );
xor ( n246396 , n246373 , n246383 );
and ( n246397 , n246396 , n246394 );
and ( n246398 , n246373 , n246383 );
or ( n246399 , n246397 , n246398 );
not ( n246400 , n222454 );
not ( n246401 , n246216 );
or ( n246402 , n246400 , n246401 );
nand ( n246403 , n237493 , n240229 );
nand ( n246404 , n246402 , n246403 );
not ( n246405 , n224087 );
not ( n246406 , n246277 );
or ( n246407 , n246405 , n246406 );
not ( n246408 , n239899 );
not ( n246409 , n237271 );
or ( n246410 , n246408 , n246409 );
nand ( n246411 , n237272 , n238672 );
nand ( n246412 , n246410 , n246411 );
nand ( n246413 , n246412 , n239495 );
nand ( n246414 , n246407 , n246413 );
xor ( n246415 , n246404 , n246414 );
not ( n246416 , n242888 );
not ( n246417 , n238230 );
not ( n246418 , n246417 );
not ( n246419 , n226243 );
or ( n246420 , n246418 , n246419 );
nand ( n246421 , n39747 , n238230 );
nand ( n246422 , n246420 , n246421 );
not ( n246423 , n246422 );
or ( n246424 , n246416 , n246423 );
nand ( n246425 , n246253 , n239441 );
nand ( n246426 , n246424 , n246425 );
xor ( n246427 , n246415 , n246426 );
xor ( n246428 , n246404 , n246414 );
and ( n246429 , n246428 , n246426 );
and ( n246430 , n246404 , n246414 );
or ( n246431 , n246429 , n246430 );
not ( n246432 , n237810 );
not ( n246433 , n246266 );
or ( n246434 , n246432 , n246433 );
not ( n246435 , n237816 );
not ( n246436 , n234350 );
or ( n246437 , n246435 , n246436 );
nand ( n246438 , n243392 , n245458 );
nand ( n246439 , n246437 , n246438 );
nand ( n246440 , n246439 , n238240 );
nand ( n246441 , n246434 , n246440 );
not ( n246442 , n239270 );
not ( n246443 , n246204 );
or ( n246444 , n246442 , n246443 );
xor ( n246445 , n239281 , n239527 );
nand ( n246446 , n246445 , n238274 );
nand ( n246447 , n246444 , n246446 );
not ( n246448 , n246447 );
xor ( n246449 , n246441 , n246448 );
xor ( n246450 , n246449 , n246202 );
xor ( n246451 , n246441 , n246448 );
and ( n246452 , n246451 , n246202 );
and ( n246453 , n246441 , n246448 );
or ( n246454 , n246452 , n246453 );
xor ( n246455 , n246313 , n246359 );
xor ( n246456 , n246455 , n246309 );
xor ( n246457 , n246313 , n246359 );
and ( n246458 , n246457 , n246309 );
and ( n246459 , n246313 , n246359 );
or ( n246460 , n246458 , n246459 );
xor ( n246461 , n246225 , n246395 );
xor ( n246462 , n246461 , n246427 );
xor ( n246463 , n246225 , n246395 );
and ( n246464 , n246463 , n246427 );
and ( n246465 , n246225 , n246395 );
or ( n246466 , n246464 , n246465 );
xor ( n246467 , n246450 , n246317 );
xor ( n246468 , n246467 , n246321 );
xor ( n246469 , n246450 , n246317 );
and ( n246470 , n246469 , n246321 );
and ( n246471 , n246450 , n246317 );
or ( n246472 , n246470 , n246471 );
xor ( n246473 , n246325 , n246456 );
xor ( n246474 , n246473 , n246462 );
xor ( n246475 , n246325 , n246456 );
and ( n246476 , n246475 , n246462 );
and ( n246477 , n246325 , n246456 );
or ( n246478 , n246476 , n246477 );
xor ( n246479 , n246329 , n246468 );
xor ( n246480 , n246479 , n246333 );
xor ( n246481 , n246329 , n246468 );
and ( n246482 , n246481 , n246333 );
and ( n246483 , n246329 , n246468 );
or ( n246484 , n246482 , n246483 );
xor ( n246485 , n246474 , n246480 );
xor ( n246486 , n246485 , n246337 );
xor ( n246487 , n246474 , n246480 );
and ( n246488 , n246487 , n246337 );
and ( n246489 , n246474 , n246480 );
or ( n246490 , n246488 , n246489 );
not ( n246491 , n239872 );
not ( n246492 , n235644 );
or ( n246493 , n246491 , n246492 );
nand ( n246494 , n246493 , n240229 );
not ( n246495 , n244387 );
not ( n246496 , n246342 );
or ( n246497 , n246495 , n246496 );
not ( n246498 , n239393 );
not ( n246499 , n226961 );
or ( n246500 , n246498 , n246499 );
nand ( n246501 , n242471 , n244654 );
nand ( n246502 , n246500 , n246501 );
nand ( n246503 , n246502 , n242737 );
nand ( n246504 , n246497 , n246503 );
xor ( n246505 , n246494 , n246504 );
not ( n246506 , n238274 );
xor ( n246507 , n233465 , n235031 );
not ( n246508 , n246507 );
or ( n246509 , n246506 , n246508 );
nand ( n246510 , n246445 , n239270 );
nand ( n246511 , n246509 , n246510 );
xor ( n246512 , n246505 , n246511 );
xor ( n246513 , n246494 , n246504 );
and ( n246514 , n246513 , n246511 );
and ( n246515 , n246494 , n246504 );
or ( n246516 , n246514 , n246515 );
and ( n246517 , n234382 , n239139 );
not ( n246518 , n227294 );
not ( n246519 , n237005 );
not ( n246520 , n245529 );
not ( n246521 , n246520 );
or ( n246522 , n246519 , n246521 );
nand ( n246523 , n209966 , n241404 );
nand ( n246524 , n246522 , n246523 );
not ( n246525 , n246524 );
or ( n246526 , n246518 , n246525 );
nand ( n246527 , n246356 , n238409 );
nand ( n246528 , n246526 , n246527 );
xor ( n246529 , n246517 , n246528 );
not ( n246530 , n239794 );
not ( n246531 , n246369 );
or ( n246532 , n246530 , n246531 );
not ( n246533 , n238619 );
not ( n246534 , n39928 );
or ( n246535 , n246533 , n246534 );
nand ( n246536 , n39929 , n244643 );
nand ( n246537 , n246535 , n246536 );
nand ( n246538 , n246537 , n228868 );
nand ( n246539 , n246532 , n246538 );
xor ( n246540 , n246529 , n246539 );
xor ( n246541 , n246517 , n246528 );
and ( n246542 , n246541 , n246539 );
and ( n246543 , n246517 , n246528 );
or ( n246544 , n246542 , n246543 );
not ( n246545 , n240271 );
not ( n246546 , n246379 );
or ( n246547 , n246545 , n246546 );
not ( n246548 , n234878 );
not ( n246549 , n238486 );
or ( n246550 , n246548 , n246549 );
nand ( n246551 , n39288 , n244121 );
nand ( n246552 , n246550 , n246551 );
nand ( n246553 , n246552 , n240020 );
nand ( n246554 , n246547 , n246553 );
not ( n246555 , n238776 );
not ( n246556 , n239932 );
and ( n246557 , n232493 , n246556 );
not ( n246558 , n232493 );
and ( n246559 , n246558 , n239932 );
nor ( n246560 , n246557 , n246559 );
not ( n246561 , n246560 );
or ( n246562 , n246555 , n246561 );
nand ( n246563 , n246392 , n242335 );
nand ( n246564 , n246562 , n246563 );
xor ( n246565 , n246554 , n246564 );
not ( n246566 , n239495 );
not ( n246567 , n239899 );
not ( n246568 , n243765 );
or ( n246569 , n246567 , n246568 );
nand ( n246570 , n243764 , n238672 );
nand ( n246571 , n246569 , n246570 );
not ( n246572 , n246571 );
or ( n246573 , n246566 , n246572 );
nand ( n246574 , n246412 , n224087 );
nand ( n246575 , n246573 , n246574 );
xor ( n246576 , n246565 , n246575 );
xor ( n246577 , n246554 , n246564 );
and ( n246578 , n246577 , n246575 );
and ( n246579 , n246554 , n246564 );
or ( n246580 , n246578 , n246579 );
not ( n246581 , n242888 );
and ( n246582 , n238230 , n243754 );
not ( n246583 , n238230 );
and ( n246584 , n246583 , n39608 );
nor ( n246585 , n246582 , n246584 );
not ( n246586 , n246585 );
or ( n246587 , n246581 , n246586 );
nand ( n246588 , n246422 , n239441 );
nand ( n246589 , n246587 , n246588 );
buf ( n246590 , n238240 );
not ( n246591 , n246590 );
not ( n246592 , n237816 );
not ( n246593 , n210823 );
or ( n246594 , n246592 , n246593 );
nand ( n246595 , n239787 , n39714 );
nand ( n246596 , n246594 , n246595 );
not ( n246597 , n246596 );
or ( n246598 , n246591 , n246597 );
nand ( n246599 , n246439 , n237810 );
nand ( n246600 , n246598 , n246599 );
xor ( n246601 , n246589 , n246600 );
xor ( n246602 , n246601 , n246447 );
xor ( n246603 , n246589 , n246600 );
and ( n246604 , n246603 , n246447 );
and ( n246605 , n246589 , n246600 );
or ( n246606 , n246604 , n246605 );
xor ( n246607 , n246512 , n246431 );
xor ( n246608 , n246607 , n246363 );
xor ( n246609 , n246512 , n246431 );
and ( n246610 , n246609 , n246363 );
and ( n246611 , n246512 , n246431 );
or ( n246612 , n246610 , n246611 );
xor ( n246613 , n246399 , n246540 );
xor ( n246614 , n246613 , n246576 );
xor ( n246615 , n246399 , n246540 );
and ( n246616 , n246615 , n246576 );
and ( n246617 , n246399 , n246540 );
or ( n246618 , n246616 , n246617 );
xor ( n246619 , n246602 , n246454 );
xor ( n246620 , n246619 , n246460 );
xor ( n246621 , n246602 , n246454 );
and ( n246622 , n246621 , n246460 );
and ( n246623 , n246602 , n246454 );
or ( n246624 , n246622 , n246623 );
xor ( n246625 , n246466 , n246608 );
xor ( n246626 , n246625 , n246614 );
xor ( n246627 , n246466 , n246608 );
and ( n246628 , n246627 , n246614 );
and ( n246629 , n246466 , n246608 );
or ( n246630 , n246628 , n246629 );
xor ( n246631 , n246472 , n246620 );
xor ( n246632 , n246631 , n246478 );
xor ( n246633 , n246472 , n246620 );
and ( n246634 , n246633 , n246478 );
and ( n246635 , n246472 , n246620 );
or ( n246636 , n246634 , n246635 );
xor ( n246637 , n246626 , n246632 );
xor ( n246638 , n246637 , n246484 );
xor ( n246639 , n246626 , n246632 );
and ( n246640 , n246639 , n246484 );
and ( n246641 , n246626 , n246632 );
or ( n246642 , n246640 , n246641 );
and ( n246643 , n239281 , n239527 );
not ( n246644 , n224087 );
not ( n246645 , n246571 );
or ( n246646 , n246644 , n246645 );
not ( n246647 , n239899 );
not ( n246648 , n245282 );
or ( n246649 , n246647 , n246648 );
nand ( n246650 , n209866 , n238672 );
nand ( n246651 , n246649 , n246650 );
nand ( n246652 , n246651 , n239495 );
nand ( n246653 , n246646 , n246652 );
xor ( n246654 , n246643 , n246653 );
not ( n246655 , n242737 );
not ( n246656 , n239393 );
not ( n246657 , n39879 );
or ( n246658 , n246656 , n246657 );
nand ( n246659 , n39880 , n244654 );
nand ( n246660 , n246658 , n246659 );
not ( n246661 , n246660 );
or ( n246662 , n246655 , n246661 );
nand ( n246663 , n246502 , n244387 );
nand ( n246664 , n246662 , n246663 );
xor ( n246665 , n246654 , n246664 );
xor ( n246666 , n246643 , n246653 );
and ( n246667 , n246666 , n246664 );
and ( n246668 , n246643 , n246653 );
or ( n246669 , n246667 , n246668 );
not ( n246670 , n242335 );
not ( n246671 , n246560 );
or ( n246672 , n246670 , n246671 );
not ( n246673 , n232494 );
not ( n246674 , n39367 );
or ( n246675 , n246673 , n246674 );
nand ( n246676 , n246377 , n232493 );
nand ( n246677 , n246675 , n246676 );
nand ( n246678 , n246677 , n238776 );
nand ( n246679 , n246672 , n246678 );
not ( n246680 , n239441 );
not ( n246681 , n246585 );
or ( n246682 , n246680 , n246681 );
and ( n246683 , n227201 , n246417 );
not ( n246684 , n227201 );
and ( n246685 , n246684 , n238230 );
or ( n246686 , n246683 , n246685 );
nand ( n246687 , n246686 , n242888 );
nand ( n246688 , n246682 , n246687 );
xor ( n246689 , n246679 , n246688 );
not ( n246690 , n238409 );
not ( n246691 , n246524 );
or ( n246692 , n246690 , n246691 );
nand ( n246693 , n227294 , n237005 );
nand ( n246694 , n246692 , n246693 );
xor ( n246695 , n246689 , n246694 );
xor ( n246696 , n246679 , n246688 );
and ( n246697 , n246696 , n246694 );
and ( n246698 , n246679 , n246688 );
or ( n246699 , n246697 , n246698 );
not ( n246700 , n240271 );
not ( n246701 , n246552 );
or ( n246702 , n246700 , n246701 );
not ( n246703 , n234878 );
not ( n246704 , n237271 );
or ( n246705 , n246703 , n246704 );
nand ( n246706 , n237272 , n237918 );
nand ( n246707 , n246705 , n246706 );
nand ( n246708 , n246707 , n240020 );
nand ( n246709 , n246702 , n246708 );
not ( n246710 , n237810 );
not ( n246711 , n246596 );
or ( n246712 , n246710 , n246711 );
not ( n246713 , n242596 );
not ( n246714 , n39748 );
or ( n246715 , n246713 , n246714 );
not ( n246716 , n226243 );
nand ( n246717 , n246716 , n245458 );
nand ( n246718 , n246715 , n246717 );
nand ( n246719 , n246718 , n246590 );
nand ( n246720 , n246712 , n246719 );
xor ( n246721 , n246709 , n246720 );
not ( n246722 , n239794 );
not ( n246723 , n246537 );
or ( n246724 , n246722 , n246723 );
not ( n246725 , n238619 );
not ( n246726 , n242210 );
or ( n246727 , n246725 , n246726 );
nand ( n246728 , n243392 , n244643 );
nand ( n246729 , n246727 , n246728 );
nand ( n246730 , n246729 , n228868 );
nand ( n246731 , n246724 , n246730 );
xor ( n246732 , n246721 , n246731 );
xor ( n246733 , n246709 , n246720 );
and ( n246734 , n246733 , n246731 );
and ( n246735 , n246709 , n246720 );
or ( n246736 , n246734 , n246735 );
not ( n246737 , n239270 );
not ( n246738 , n246507 );
or ( n246739 , n246737 , n246738 );
and ( n246740 , n239281 , n244885 );
not ( n246741 , n239281 );
and ( n246742 , n246741 , n237963 );
or ( n246743 , n246740 , n246742 );
nand ( n246744 , n246743 , n238274 );
nand ( n246745 , n246739 , n246744 );
not ( n246746 , n246745 );
xor ( n246747 , n246746 , n246516 );
xor ( n246748 , n246747 , n246544 );
xor ( n246749 , n246746 , n246516 );
and ( n246750 , n246749 , n246544 );
and ( n246751 , n246746 , n246516 );
or ( n246752 , n246750 , n246751 );
xor ( n246753 , n246580 , n246665 );
xor ( n246754 , n246753 , n246695 );
xor ( n246755 , n246580 , n246665 );
and ( n246756 , n246755 , n246695 );
and ( n246757 , n246580 , n246665 );
or ( n246758 , n246756 , n246757 );
xor ( n246759 , n246732 , n246606 );
xor ( n246760 , n246759 , n246612 );
xor ( n246761 , n246732 , n246606 );
and ( n246762 , n246761 , n246612 );
and ( n246763 , n246732 , n246606 );
or ( n246764 , n246762 , n246763 );
xor ( n246765 , n246748 , n246618 );
xor ( n246766 , n246765 , n246754 );
xor ( n246767 , n246748 , n246618 );
and ( n246768 , n246767 , n246754 );
and ( n246769 , n246748 , n246618 );
or ( n246770 , n246768 , n246769 );
xor ( n246771 , n246760 , n246624 );
xor ( n246772 , n246771 , n246630 );
xor ( n246773 , n246760 , n246624 );
and ( n246774 , n246773 , n246630 );
and ( n246775 , n246760 , n246624 );
or ( n246776 , n246774 , n246775 );
xor ( n246777 , n246766 , n246772 );
xor ( n246778 , n246777 , n246636 );
xor ( n246779 , n246766 , n246772 );
and ( n246780 , n246779 , n246636 );
and ( n246781 , n246766 , n246772 );
or ( n246782 , n246780 , n246781 );
not ( n246783 , n225376 );
not ( n246784 , n236338 );
or ( n246785 , n246783 , n246784 );
nand ( n246786 , n246785 , n237005 );
not ( n246787 , n239270 );
not ( n246788 , n246743 );
or ( n246789 , n246787 , n246788 );
xor ( n246790 , n240156 , n229928 );
nand ( n246791 , n246790 , n238274 );
nand ( n246792 , n246789 , n246791 );
xor ( n246793 , n246786 , n246792 );
and ( n246794 , n233465 , n235031 );
xor ( n246795 , n246793 , n246794 );
xor ( n246796 , n246786 , n246792 );
and ( n246797 , n246796 , n246794 );
and ( n246798 , n246786 , n246792 );
or ( n246799 , n246797 , n246798 );
not ( n246800 , n239495 );
not ( n246801 , n239899 );
not ( n246802 , n246520 );
or ( n246803 , n246801 , n246802 );
buf ( n246804 , n245093 );
nand ( n246805 , n246804 , n238672 );
nand ( n246806 , n246803 , n246805 );
not ( n246807 , n246806 );
or ( n246808 , n246800 , n246807 );
nand ( n246809 , n246651 , n224087 );
nand ( n246810 , n246808 , n246809 );
not ( n246811 , n244387 );
not ( n246812 , n246660 );
or ( n246813 , n246811 , n246812 );
and ( n246814 , n239393 , n39928 );
not ( n246815 , n239393 );
and ( n246816 , n246815 , n39929 );
or ( n246817 , n246814 , n246816 );
nand ( n246818 , n246817 , n242737 );
nand ( n246819 , n246813 , n246818 );
xor ( n246820 , n246810 , n246819 );
not ( n246821 , n238776 );
not ( n246822 , n232494 );
not ( n246823 , n39287 );
or ( n246824 , n246822 , n246823 );
nand ( n246825 , n39288 , n232493 );
nand ( n246826 , n246824 , n246825 );
not ( n246827 , n246826 );
or ( n246828 , n246821 , n246827 );
nand ( n246829 , n246677 , n242335 );
nand ( n246830 , n246828 , n246829 );
xor ( n246831 , n246820 , n246830 );
xor ( n246832 , n246810 , n246819 );
and ( n246833 , n246832 , n246830 );
and ( n246834 , n246810 , n246819 );
or ( n246835 , n246833 , n246834 );
not ( n246836 , n242888 );
and ( n246837 , n238230 , n246556 );
not ( n246838 , n238230 );
and ( n246839 , n246838 , n239932 );
nor ( n246840 , n246837 , n246839 );
not ( n246841 , n246840 );
or ( n246842 , n246836 , n246841 );
nand ( n246843 , n246686 , n239441 );
nand ( n246844 , n246842 , n246843 );
not ( n246845 , n240020 );
and ( n246846 , n237918 , n243765 );
not ( n246847 , n237918 );
and ( n246848 , n246847 , n243764 );
nor ( n246849 , n246846 , n246848 );
not ( n246850 , n246849 );
or ( n246851 , n246845 , n246850 );
nand ( n246852 , n246707 , n240271 );
nand ( n246853 , n246851 , n246852 );
xor ( n246854 , n246844 , n246853 );
not ( n246855 , n246590 );
not ( n246856 , n237816 );
not ( n246857 , n39608 );
not ( n246858 , n246857 );
or ( n246859 , n246856 , n246858 );
nand ( n246860 , n39608 , n245458 );
nand ( n246861 , n246859 , n246860 );
not ( n246862 , n246861 );
or ( n246863 , n246855 , n246862 );
nand ( n246864 , n246718 , n237810 );
nand ( n246865 , n246863 , n246864 );
xor ( n246866 , n246854 , n246865 );
xor ( n246867 , n246844 , n246853 );
and ( n246868 , n246867 , n246865 );
and ( n246869 , n246844 , n246853 );
or ( n246870 , n246868 , n246869 );
not ( n246871 , n228868 );
and ( n246872 , n238619 , n39714 );
not ( n246873 , n238619 );
and ( n246874 , n246873 , n210823 );
nor ( n246875 , n246872 , n246874 );
not ( n246876 , n246875 );
or ( n246877 , n246871 , n246876 );
nand ( n246878 , n246729 , n239794 );
nand ( n246879 , n246877 , n246878 );
xor ( n246880 , n246879 , n246745 );
xor ( n246881 , n246880 , n246795 );
xor ( n246882 , n246879 , n246745 );
and ( n246883 , n246882 , n246795 );
and ( n246884 , n246879 , n246745 );
or ( n246885 , n246883 , n246884 );
xor ( n246886 , n246669 , n246699 );
xor ( n246887 , n246886 , n246736 );
xor ( n246888 , n246669 , n246699 );
and ( n246889 , n246888 , n246736 );
and ( n246890 , n246669 , n246699 );
or ( n246891 , n246889 , n246890 );
xor ( n246892 , n246866 , n246831 );
xor ( n246893 , n246892 , n246752 );
xor ( n246894 , n246866 , n246831 );
and ( n246895 , n246894 , n246752 );
and ( n246896 , n246866 , n246831 );
or ( n246897 , n246895 , n246896 );
xor ( n246898 , n246881 , n246887 );
xor ( n246899 , n246898 , n246758 );
xor ( n246900 , n246881 , n246887 );
and ( n246901 , n246900 , n246758 );
and ( n246902 , n246881 , n246887 );
or ( n246903 , n246901 , n246902 );
xor ( n246904 , n246893 , n246764 );
xor ( n246905 , n246904 , n246770 );
xor ( n246906 , n246893 , n246764 );
and ( n246907 , n246906 , n246770 );
and ( n246908 , n246893 , n246764 );
or ( n246909 , n246907 , n246908 );
xor ( n246910 , n246899 , n246905 );
xor ( n246911 , n246910 , n246776 );
xor ( n246912 , n246899 , n246905 );
and ( n246913 , n246912 , n246776 );
and ( n246914 , n246899 , n246905 );
or ( n246915 , n246913 , n246914 );
not ( n246916 , n240271 );
not ( n246917 , n246849 );
or ( n246918 , n246916 , n246917 );
not ( n246919 , n234878 );
not ( n246920 , n245282 );
or ( n246921 , n246919 , n246920 );
not ( n246922 , n245282 );
nand ( n246923 , n246922 , n237918 );
nand ( n246924 , n246921 , n246923 );
nand ( n246925 , n246924 , n240020 );
nand ( n246926 , n246918 , n246925 );
not ( n246927 , n238274 );
xor ( n246928 , n233891 , n39880 );
not ( n246929 , n246928 );
or ( n246930 , n246927 , n246929 );
nand ( n246931 , n246790 , n239270 );
nand ( n246932 , n246930 , n246931 );
xor ( n246933 , n246926 , n246932 );
not ( n246934 , n239441 );
not ( n246935 , n246840 );
or ( n246936 , n246934 , n246935 );
not ( n246937 , n246417 );
not ( n246938 , n39367 );
or ( n246939 , n246937 , n246938 );
nand ( n246940 , n246377 , n238230 );
nand ( n246941 , n246939 , n246940 );
nand ( n246942 , n246941 , n242888 );
nand ( n246943 , n246936 , n246942 );
xor ( n246944 , n246933 , n246943 );
xor ( n246945 , n246926 , n246932 );
and ( n246946 , n246945 , n246943 );
and ( n246947 , n246926 , n246932 );
or ( n246948 , n246946 , n246947 );
not ( n246949 , n224087 );
not ( n246950 , n246806 );
or ( n246951 , n246949 , n246950 );
nand ( n246952 , n239495 , n239899 );
nand ( n246953 , n246951 , n246952 );
not ( n246954 , n237810 );
not ( n246955 , n246861 );
or ( n246956 , n246954 , n246955 );
and ( n246957 , n242596 , n238857 );
not ( n246958 , n242596 );
and ( n246959 , n246958 , n227201 );
nor ( n246960 , n246957 , n246959 );
nand ( n246961 , n246960 , n246590 );
nand ( n246962 , n246956 , n246961 );
xor ( n246963 , n246953 , n246962 );
not ( n246964 , n242335 );
not ( n246965 , n246826 );
or ( n246966 , n246964 , n246965 );
not ( n246967 , n232494 );
not ( n246968 , n237271 );
or ( n246969 , n246967 , n246968 );
nand ( n246970 , n237272 , n232493 );
nand ( n246971 , n246969 , n246970 );
not ( n246972 , n246971 );
or ( n246973 , n246972 , n238777 );
nand ( n246974 , n246966 , n246973 );
xor ( n246975 , n246963 , n246974 );
xor ( n246976 , n246953 , n246962 );
and ( n246977 , n246976 , n246974 );
and ( n246978 , n246953 , n246962 );
or ( n246979 , n246977 , n246978 );
not ( n246980 , n239794 );
not ( n246981 , n246875 );
or ( n246982 , n246980 , n246981 );
not ( n246983 , n238619 );
not ( n246984 , n39748 );
or ( n246985 , n246983 , n246984 );
nand ( n246986 , n39749 , n244643 );
nand ( n246987 , n246985 , n246986 );
nand ( n246988 , n246987 , n228868 );
nand ( n246989 , n246982 , n246988 );
not ( n246990 , n244387 );
not ( n246991 , n246817 );
or ( n246992 , n246990 , n246991 );
and ( n246993 , n239393 , n243392 );
not ( n246994 , n239393 );
and ( n246995 , n246994 , n242210 );
nor ( n246996 , n246993 , n246995 );
nand ( n246997 , n246996 , n242737 );
nand ( n246998 , n246992 , n246997 );
xor ( n246999 , n246989 , n246998 );
nand ( n247000 , n237963 , n234382 );
xor ( n247001 , n246999 , n247000 );
xor ( n247002 , n246989 , n246998 );
and ( n247003 , n247002 , n247000 );
and ( n247004 , n246989 , n246998 );
or ( n247005 , n247003 , n247004 );
xor ( n247006 , n246799 , n246835 );
xor ( n247007 , n247006 , n246870 );
xor ( n247008 , n246799 , n246835 );
and ( n247009 , n247008 , n246870 );
and ( n247010 , n246799 , n246835 );
or ( n247011 , n247009 , n247010 );
xor ( n247012 , n246944 , n247001 );
xor ( n247013 , n247012 , n246975 );
xor ( n247014 , n246944 , n247001 );
and ( n247015 , n247014 , n246975 );
and ( n247016 , n246944 , n247001 );
or ( n247017 , n247015 , n247016 );
xor ( n247018 , n246891 , n246885 );
xor ( n247019 , n247018 , n247007 );
xor ( n247020 , n246891 , n246885 );
and ( n247021 , n247020 , n247007 );
and ( n247022 , n246891 , n246885 );
or ( n247023 , n247021 , n247022 );
xor ( n247024 , n247013 , n246897 );
xor ( n247025 , n247024 , n246903 );
xor ( n247026 , n247013 , n246897 );
and ( n247027 , n247026 , n246903 );
and ( n247028 , n247013 , n246897 );
or ( n247029 , n247027 , n247028 );
xor ( n247030 , n247019 , n247025 );
xor ( n247031 , n247030 , n246909 );
xor ( n247032 , n247019 , n247025 );
and ( n247033 , n247032 , n246909 );
and ( n247034 , n247019 , n247025 );
or ( n247035 , n247033 , n247034 );
or ( n247036 , n239495 , n224087 );
nand ( n247037 , n247036 , n239899 );
and ( n247038 , n240156 , n229928 );
xor ( n247039 , n247037 , n247038 );
not ( n247040 , n240020 );
not ( n247041 , n234878 );
not ( n247042 , n246520 );
or ( n247043 , n247041 , n247042 );
nand ( n247044 , n246804 , n237918 );
nand ( n247045 , n247043 , n247044 );
not ( n247046 , n247045 );
or ( n247047 , n247040 , n247046 );
nand ( n247048 , n246924 , n240271 );
nand ( n247049 , n247047 , n247048 );
xor ( n247050 , n247039 , n247049 );
xor ( n247051 , n247037 , n247038 );
and ( n247052 , n247051 , n247049 );
and ( n247053 , n247037 , n247038 );
or ( n247054 , n247052 , n247053 );
not ( n247055 , n239270 );
not ( n247056 , n246928 );
or ( n247057 , n247055 , n247056 );
xor ( n247058 , n233891 , n210919 );
nand ( n247059 , n247058 , n238274 );
nand ( n247060 , n247057 , n247059 );
not ( n247061 , n239441 );
not ( n247062 , n246941 );
or ( n247063 , n247061 , n247062 );
not ( n247064 , n246417 );
not ( n247065 , n39287 );
or ( n247066 , n247064 , n247065 );
nand ( n247067 , n238230 , n39288 );
nand ( n247068 , n247066 , n247067 );
nand ( n247069 , n247068 , n242888 );
nand ( n247070 , n247063 , n247069 );
xor ( n247071 , n247060 , n247070 );
not ( n247072 , n237810 );
not ( n247073 , n246960 );
or ( n247074 , n247072 , n247073 );
and ( n247075 , n239787 , n239932 );
not ( n247076 , n239787 );
and ( n247077 , n247076 , n246556 );
nor ( n247078 , n247075 , n247077 );
not ( n247079 , n246590 );
or ( n247080 , n247078 , n247079 );
nand ( n247081 , n247074 , n247080 );
xor ( n247082 , n247071 , n247081 );
xor ( n247083 , n247060 , n247070 );
and ( n247084 , n247083 , n247081 );
and ( n247085 , n247060 , n247070 );
or ( n247086 , n247084 , n247085 );
not ( n247087 , n238776 );
not ( n247088 , n232494 );
not ( n247089 , n243765 );
or ( n247090 , n247088 , n247089 );
nand ( n247091 , n243764 , n232493 );
nand ( n247092 , n247090 , n247091 );
not ( n247093 , n247092 );
or ( n247094 , n247087 , n247093 );
nand ( n247095 , n246971 , n242335 );
nand ( n247096 , n247094 , n247095 );
not ( n247097 , n239794 );
not ( n247098 , n246987 );
or ( n247099 , n247097 , n247098 );
not ( n247100 , n238619 );
not ( n247101 , n246857 );
or ( n247102 , n247100 , n247101 );
nand ( n247103 , n244643 , n39608 );
nand ( n247104 , n247102 , n247103 );
nand ( n247105 , n247104 , n228868 );
nand ( n247106 , n247099 , n247105 );
xor ( n247107 , n247096 , n247106 );
not ( n247108 , n244387 );
not ( n247109 , n246996 );
or ( n247110 , n247108 , n247109 );
and ( n247111 , n239393 , n210823 );
not ( n247112 , n239393 );
and ( n247113 , n247112 , n39714 );
nor ( n247114 , n247111 , n247113 );
not ( n247115 , n247114 );
nand ( n247116 , n247115 , n242737 );
nand ( n247117 , n247110 , n247116 );
xor ( n247118 , n247107 , n247117 );
xor ( n247119 , n247096 , n247106 );
and ( n247120 , n247119 , n247117 );
and ( n247121 , n247096 , n247106 );
or ( n247122 , n247120 , n247121 );
not ( n247123 , n247000 );
xor ( n247124 , n247123 , n247050 );
xor ( n247125 , n247124 , n246948 );
xor ( n247126 , n247123 , n247050 );
and ( n247127 , n247126 , n246948 );
and ( n247128 , n247123 , n247050 );
or ( n247129 , n247127 , n247128 );
xor ( n247130 , n246979 , n247118 );
xor ( n247131 , n247130 , n247005 );
xor ( n247132 , n246979 , n247118 );
and ( n247133 , n247132 , n247005 );
and ( n247134 , n246979 , n247118 );
or ( n247135 , n247133 , n247134 );
xor ( n247136 , n247082 , n247011 );
xor ( n247137 , n247136 , n247125 );
xor ( n247138 , n247082 , n247011 );
and ( n247139 , n247138 , n247125 );
and ( n247140 , n247082 , n247011 );
or ( n247141 , n247139 , n247140 );
xor ( n247142 , n247017 , n247131 );
xor ( n247143 , n247142 , n247137 );
xor ( n247144 , n247017 , n247131 );
and ( n247145 , n247144 , n247137 );
and ( n247146 , n247017 , n247131 );
or ( n247147 , n247145 , n247146 );
xor ( n247148 , n247023 , n247143 );
xor ( n247149 , n247148 , n247029 );
xor ( n247150 , n247023 , n247143 );
and ( n247151 , n247150 , n247029 );
and ( n247152 , n247023 , n247143 );
or ( n247153 , n247151 , n247152 );
not ( n247154 , n242335 );
not ( n247155 , n247092 );
or ( n247156 , n247154 , n247155 );
not ( n247157 , n232494 );
not ( n247158 , n245282 );
or ( n247159 , n247157 , n247158 );
nand ( n247160 , n246922 , n232493 );
nand ( n247161 , n247159 , n247160 );
nand ( n247162 , n247161 , n238776 );
nand ( n247163 , n247156 , n247162 );
and ( n247164 , n233891 , n39880 );
xor ( n247165 , n247163 , n247164 );
not ( n247166 , n246590 );
and ( n247167 , n242596 , n246377 );
not ( n247168 , n242596 );
and ( n247169 , n247168 , n39367 );
nor ( n247170 , n247167 , n247169 );
not ( n247171 , n247170 );
or ( n247172 , n247166 , n247171 );
not ( n247173 , n247078 );
nand ( n247174 , n247173 , n237810 );
nand ( n247175 , n247172 , n247174 );
xor ( n247176 , n247165 , n247175 );
xor ( n247177 , n247163 , n247164 );
and ( n247178 , n247177 , n247175 );
and ( n247179 , n247163 , n247164 );
or ( n247180 , n247178 , n247179 );
not ( n247181 , n239794 );
not ( n247182 , n247104 );
or ( n247183 , n247181 , n247182 );
not ( n247184 , n238619 );
not ( n247185 , n227201 );
or ( n247186 , n247184 , n247185 );
nand ( n247187 , n238857 , n244643 );
nand ( n247188 , n247186 , n247187 );
nand ( n247189 , n247188 , n228868 );
nand ( n247190 , n247183 , n247189 );
not ( n247191 , n239441 );
not ( n247192 , n247068 );
or ( n247193 , n247191 , n247192 );
not ( n247194 , n246417 );
not ( n247195 , n237271 );
or ( n247196 , n247194 , n247195 );
nand ( n247197 , n237272 , n238230 );
nand ( n247198 , n247196 , n247197 );
nand ( n247199 , n247198 , n242888 );
nand ( n247200 , n247193 , n247199 );
xor ( n247201 , n247190 , n247200 );
not ( n247202 , n242737 );
not ( n247203 , n239393 );
not ( n247204 , n39748 );
or ( n247205 , n247203 , n247204 );
nand ( n247206 , n39749 , n244654 );
nand ( n247207 , n247205 , n247206 );
not ( n247208 , n247207 );
or ( n247209 , n247202 , n247208 );
buf ( n247210 , n239805 );
or ( n247211 , n247114 , n247210 );
nand ( n247212 , n247209 , n247211 );
xor ( n247213 , n247201 , n247212 );
xor ( n247214 , n247190 , n247200 );
and ( n247215 , n247214 , n247212 );
and ( n247216 , n247190 , n247200 );
or ( n247217 , n247215 , n247216 );
not ( n247218 , n239270 );
not ( n247219 , n247058 );
or ( n247220 , n247218 , n247219 );
xor ( n247221 , n233891 , n243392 );
nand ( n247222 , n247221 , n238274 );
nand ( n247223 , n247220 , n247222 );
not ( n247224 , n236958 );
not ( n247225 , n237918 );
and ( n247226 , n247224 , n247225 );
and ( n247227 , n247045 , n240271 );
nor ( n247228 , n247226 , n247227 );
xor ( n247229 , n247223 , n247228 );
xor ( n247230 , n247229 , n247054 );
xor ( n247231 , n247223 , n247228 );
and ( n247232 , n247231 , n247054 );
and ( n247233 , n247223 , n247228 );
or ( n247234 , n247232 , n247233 );
xor ( n247235 , n247086 , n247122 );
xor ( n247236 , n247235 , n247213 );
xor ( n247237 , n247086 , n247122 );
and ( n247238 , n247237 , n247213 );
and ( n247239 , n247086 , n247122 );
or ( n247240 , n247238 , n247239 );
xor ( n247241 , n247176 , n247230 );
xor ( n247242 , n247241 , n247129 );
xor ( n247243 , n247176 , n247230 );
and ( n247244 , n247243 , n247129 );
and ( n247245 , n247176 , n247230 );
or ( n247246 , n247244 , n247245 );
xor ( n247247 , n247236 , n247135 );
xor ( n247248 , n247247 , n247242 );
xor ( n247249 , n247236 , n247135 );
and ( n247250 , n247249 , n247242 );
and ( n247251 , n247236 , n247135 );
or ( n247252 , n247250 , n247251 );
xor ( n247253 , n247141 , n247248 );
xor ( n247254 , n247253 , n247147 );
xor ( n247255 , n247141 , n247248 );
and ( n247256 , n247255 , n247147 );
and ( n247257 , n247141 , n247248 );
or ( n247258 , n247256 , n247257 );
not ( n247259 , n236958 );
not ( n247260 , n240272 );
or ( n247261 , n247259 , n247260 );
nand ( n247262 , n247261 , n234878 );
not ( n247263 , n238776 );
not ( n247264 , n246804 );
and ( n247265 , n232494 , n247264 );
not ( n247266 , n232494 );
and ( n247267 , n247266 , n209967 );
nor ( n247268 , n247265 , n247267 );
not ( n247269 , n247268 );
not ( n247270 , n247269 );
or ( n247271 , n247263 , n247270 );
nand ( n247272 , n247161 , n242335 );
nand ( n247273 , n247271 , n247272 );
xor ( n247274 , n247262 , n247273 );
not ( n247275 , n246590 );
not ( n247276 , n242596 );
not ( n247277 , n39287 );
or ( n247278 , n247276 , n247277 );
nand ( n247279 , n39288 , n239787 );
nand ( n247280 , n247278 , n247279 );
not ( n247281 , n247280 );
or ( n247282 , n247275 , n247281 );
nand ( n247283 , n247170 , n237810 );
nand ( n247284 , n247282 , n247283 );
xor ( n247285 , n247274 , n247284 );
xor ( n247286 , n247262 , n247273 );
and ( n247287 , n247286 , n247284 );
and ( n247288 , n247262 , n247273 );
or ( n247289 , n247287 , n247288 );
and ( n247290 , n233891 , n210919 );
not ( n247291 , n228868 );
and ( n247292 , n244643 , n246556 );
not ( n247293 , n244643 );
and ( n247294 , n247293 , n239932 );
nor ( n247295 , n247292 , n247294 );
not ( n247296 , n247295 );
or ( n247297 , n247291 , n247296 );
nand ( n247298 , n247188 , n239794 );
nand ( n247299 , n247297 , n247298 );
xor ( n247300 , n247290 , n247299 );
not ( n247301 , n242888 );
and ( n247302 , n246417 , n243764 );
not ( n247303 , n246417 );
and ( n247304 , n247303 , n243765 );
nor ( n247305 , n247302 , n247304 );
not ( n247306 , n247305 );
or ( n247307 , n247301 , n247306 );
not ( n247308 , n247198 );
not ( n247309 , n239441 );
or ( n247310 , n247308 , n247309 );
nand ( n247311 , n247307 , n247310 );
xor ( n247312 , n247300 , n247311 );
xor ( n247313 , n247290 , n247299 );
and ( n247314 , n247313 , n247311 );
and ( n247315 , n247290 , n247299 );
or ( n247316 , n247314 , n247315 );
not ( n247317 , n242737 );
buf ( n247318 , n239393 );
and ( n247319 , n247318 , n39608 );
not ( n247320 , n247318 );
and ( n247321 , n247320 , n246857 );
nor ( n247322 , n247319 , n247321 );
not ( n247323 , n247322 );
or ( n247324 , n247317 , n247323 );
nand ( n247325 , n247207 , n244387 );
nand ( n247326 , n247324 , n247325 );
not ( n247327 , n238274 );
xor ( n247328 , n233891 , n39714 );
not ( n247329 , n247328 );
or ( n247330 , n247327 , n247329 );
nand ( n247331 , n247221 , n239270 );
nand ( n247332 , n247330 , n247331 );
xor ( n247333 , n247326 , n247332 );
not ( n247334 , n247228 );
xor ( n247335 , n247333 , n247334 );
xor ( n247336 , n247326 , n247332 );
and ( n247337 , n247336 , n247334 );
and ( n247338 , n247326 , n247332 );
or ( n247339 , n247337 , n247338 );
xor ( n247340 , n247217 , n247180 );
xor ( n247341 , n247340 , n247285 );
xor ( n247342 , n247217 , n247180 );
and ( n247343 , n247342 , n247285 );
and ( n247344 , n247217 , n247180 );
or ( n247345 , n247343 , n247344 );
xor ( n247346 , n247312 , n247335 );
xor ( n247347 , n247346 , n247234 );
xor ( n247348 , n247312 , n247335 );
and ( n247349 , n247348 , n247234 );
and ( n247350 , n247312 , n247335 );
or ( n247351 , n247349 , n247350 );
xor ( n247352 , n247341 , n247240 );
xor ( n247353 , n247352 , n247246 );
xor ( n247354 , n247341 , n247240 );
and ( n247355 , n247354 , n247246 );
and ( n247356 , n247341 , n247240 );
or ( n247357 , n247355 , n247356 );
xor ( n247358 , n247347 , n247353 );
xor ( n247359 , n247358 , n247252 );
xor ( n247360 , n247347 , n247353 );
and ( n247361 , n247360 , n247252 );
and ( n247362 , n247347 , n247353 );
or ( n247363 , n247361 , n247362 );
not ( n247364 , n239441 );
not ( n247365 , n247305 );
or ( n247366 , n247364 , n247365 );
and ( n247367 , n238230 , n246922 );
not ( n247368 , n238230 );
and ( n247369 , n247368 , n245282 );
nor ( n247370 , n247367 , n247369 );
not ( n247371 , n247370 );
nand ( n247372 , n247371 , n242888 );
nand ( n247373 , n247366 , n247372 );
not ( n247374 , n228868 );
and ( n247375 , n238619 , n246377 );
not ( n247376 , n238619 );
and ( n247377 , n247376 , n39367 );
nor ( n247378 , n247375 , n247377 );
not ( n247379 , n247378 );
or ( n247380 , n247374 , n247379 );
nand ( n247381 , n247295 , n239794 );
nand ( n247382 , n247380 , n247381 );
xor ( n247383 , n247373 , n247382 );
not ( n247384 , n247322 );
or ( n247385 , n247384 , n247210 );
and ( n247386 , n244654 , n238857 );
not ( n247387 , n244654 );
and ( n247388 , n247387 , n227201 );
nor ( n247389 , n247386 , n247388 );
or ( n247390 , n247389 , n237013 );
nand ( n247391 , n247385 , n247390 );
xor ( n247392 , n247383 , n247391 );
xor ( n247393 , n247373 , n247382 );
and ( n247394 , n247393 , n247391 );
and ( n247395 , n247373 , n247382 );
or ( n247396 , n247394 , n247395 );
not ( n247397 , n237810 );
not ( n247398 , n247280 );
or ( n247399 , n247397 , n247398 );
not ( n247400 , n242596 );
not ( n247401 , n237271 );
or ( n247402 , n247400 , n247401 );
nand ( n247403 , n237272 , n245458 );
nand ( n247404 , n247402 , n247403 );
nand ( n247405 , n247404 , n246590 );
nand ( n247406 , n247399 , n247405 );
not ( n247407 , n239270 );
not ( n247408 , n247328 );
or ( n247409 , n247407 , n247408 );
xor ( n247410 , n234382 , n246716 );
nand ( n247411 , n247410 , n238274 );
nand ( n247412 , n247409 , n247411 );
xor ( n247413 , n247406 , n247412 );
and ( n247414 , n233891 , n243392 );
xor ( n247415 , n247413 , n247414 );
xor ( n247416 , n247406 , n247412 );
and ( n247417 , n247416 , n247414 );
and ( n247418 , n247406 , n247412 );
or ( n247419 , n247417 , n247418 );
not ( n247420 , n247268 );
not ( n247421 , n242335 );
not ( n247422 , n247421 );
and ( n247423 , n247420 , n247422 );
and ( n247424 , n238776 , n232494 );
nor ( n247425 , n247423 , n247424 );
xor ( n247426 , n247425 , n247289 );
xor ( n247427 , n247426 , n247316 );
xor ( n247428 , n247425 , n247289 );
and ( n247429 , n247428 , n247316 );
and ( n247430 , n247425 , n247289 );
or ( n247431 , n247429 , n247430 );
xor ( n247432 , n247415 , n247392 );
xor ( n247433 , n247432 , n247339 );
xor ( n247434 , n247415 , n247392 );
and ( n247435 , n247434 , n247339 );
and ( n247436 , n247415 , n247392 );
or ( n247437 , n247435 , n247436 );
xor ( n247438 , n247427 , n247345 );
xor ( n247439 , n247438 , n247433 );
xor ( n247440 , n247427 , n247345 );
and ( n247441 , n247440 , n247433 );
and ( n247442 , n247427 , n247345 );
or ( n247443 , n247441 , n247442 );
xor ( n247444 , n247351 , n247439 );
xor ( n247445 , n247444 , n247357 );
xor ( n247446 , n247351 , n247439 );
and ( n247447 , n247446 , n247357 );
and ( n247448 , n247351 , n247439 );
or ( n247449 , n247447 , n247448 );
or ( n247450 , n242335 , n238776 );
nand ( n247451 , n247450 , n232494 );
or ( n247452 , n247370 , n247309 );
and ( n247453 , n246417 , n247264 );
not ( n247454 , n246417 );
not ( n247455 , n247264 );
and ( n247456 , n247454 , n247455 );
nor ( n247457 , n247453 , n247456 );
not ( n247458 , n242888 );
or ( n247459 , n247457 , n247458 );
nand ( n247460 , n247452 , n247459 );
xor ( n247461 , n247451 , n247460 );
not ( n247462 , n239794 );
not ( n247463 , n247378 );
or ( n247464 , n247462 , n247463 );
and ( n247465 , n244643 , n39288 );
and ( n247466 , n39287 , n238619 );
nor ( n247467 , n247465 , n247466 );
or ( n247468 , n247467 , n237041 );
nand ( n247469 , n247464 , n247468 );
xor ( n247470 , n247461 , n247469 );
xor ( n247471 , n247451 , n247460 );
and ( n247472 , n247471 , n247469 );
and ( n247473 , n247451 , n247460 );
or ( n247474 , n247472 , n247473 );
not ( n247475 , n244387 );
not ( n247476 , n247389 );
not ( n247477 , n247476 );
or ( n247478 , n247475 , n247477 );
and ( n247479 , n239932 , n244654 );
and ( n247480 , n246556 , n247318 );
nor ( n247481 , n247479 , n247480 );
or ( n247482 , n247481 , n237013 );
nand ( n247483 , n247478 , n247482 );
not ( n247484 , n246590 );
and ( n247485 , n245458 , n243764 );
not ( n247486 , n245458 );
and ( n247487 , n247486 , n243765 );
nor ( n247488 , n247485 , n247487 );
not ( n247489 , n247488 );
not ( n247490 , n247489 );
or ( n247491 , n247484 , n247490 );
not ( n247492 , n247404 );
or ( n247493 , n247492 , n239784 );
nand ( n247494 , n247491 , n247493 );
xor ( n247495 , n247483 , n247494 );
not ( n247496 , n247410 );
not ( n247497 , n239270 );
or ( n247498 , n247496 , n247497 );
and ( n247499 , n39608 , n243297 );
and ( n247500 , n246857 , n234382 );
nor ( n247501 , n247499 , n247500 );
or ( n247502 , n247501 , n240148 );
nand ( n247503 , n247498 , n247502 );
xor ( n247504 , n247495 , n247503 );
xor ( n247505 , n247483 , n247494 );
and ( n247506 , n247505 , n247503 );
and ( n247507 , n247483 , n247494 );
or ( n247508 , n247506 , n247507 );
and ( n247509 , n233891 , n39714 );
not ( n247510 , n247425 );
xor ( n247511 , n247509 , n247510 );
xor ( n247512 , n247511 , n247396 );
xor ( n247513 , n247509 , n247510 );
and ( n247514 , n247513 , n247396 );
and ( n247515 , n247509 , n247510 );
or ( n247516 , n247514 , n247515 );
xor ( n247517 , n247419 , n247504 );
xor ( n247518 , n247517 , n247470 );
xor ( n247519 , n247419 , n247504 );
and ( n247520 , n247519 , n247470 );
and ( n247521 , n247419 , n247504 );
or ( n247522 , n247520 , n247521 );
xor ( n247523 , n247512 , n247431 );
xor ( n247524 , n247523 , n247437 );
xor ( n247525 , n247512 , n247431 );
and ( n247526 , n247525 , n247437 );
and ( n247527 , n247512 , n247431 );
or ( n247528 , n247526 , n247527 );
xor ( n247529 , n247518 , n247524 );
xor ( n247530 , n247529 , n247443 );
xor ( n247531 , n247518 , n247524 );
and ( n247532 , n247531 , n247443 );
and ( n247533 , n247518 , n247524 );
or ( n247534 , n247532 , n247533 );
or ( n247535 , n247481 , n247210 );
and ( n247536 , n246377 , n244654 );
not ( n247537 , n246377 );
and ( n247538 , n247537 , n239393 );
nor ( n247539 , n247536 , n247538 );
or ( n247540 , n247539 , n237013 );
nand ( n247541 , n247535 , n247540 );
or ( n247542 , n247501 , n247497 );
and ( n247543 , n234382 , n227201 );
not ( n247544 , n234382 );
and ( n247545 , n247544 , n238857 );
nor ( n247546 , n247543 , n247545 );
or ( n247547 , n247546 , n240148 );
nand ( n247548 , n247542 , n247547 );
xor ( n247549 , n247541 , n247548 );
or ( n247550 , n247457 , n247309 );
or ( n247551 , n247458 , n238230 );
nand ( n247552 , n247550 , n247551 );
xor ( n247553 , n247549 , n247552 );
xor ( n247554 , n247541 , n247548 );
and ( n247555 , n247554 , n247552 );
and ( n247556 , n247541 , n247548 );
or ( n247557 , n247555 , n247556 );
and ( n247558 , n234382 , n246716 );
not ( n247559 , n239794 );
or ( n247560 , n247467 , n247559 );
and ( n247561 , n237271 , n238619 );
not ( n247562 , n237271 );
and ( n247563 , n247562 , n244643 );
nor ( n247564 , n247561 , n247563 );
or ( n247565 , n247564 , n237041 );
nand ( n247566 , n247560 , n247565 );
xor ( n247567 , n247558 , n247566 );
or ( n247568 , n247488 , n239784 );
and ( n247569 , n209866 , n239787 );
and ( n247570 , n245282 , n242596 );
nor ( n247571 , n247569 , n247570 );
or ( n247572 , n247571 , n247079 );
nand ( n247573 , n247568 , n247572 );
not ( n247574 , n247573 );
xor ( n247575 , n247567 , n247574 );
xor ( n247576 , n247558 , n247566 );
and ( n247577 , n247576 , n247574 );
and ( n247578 , n247558 , n247566 );
or ( n247579 , n247577 , n247578 );
xor ( n247580 , n247508 , n247474 );
xor ( n247581 , n247580 , n247553 );
xor ( n247582 , n247508 , n247474 );
and ( n247583 , n247582 , n247553 );
and ( n247584 , n247508 , n247474 );
or ( n247585 , n247583 , n247584 );
xor ( n247586 , n247575 , n247516 );
xor ( n247587 , n247586 , n247522 );
xor ( n247588 , n247575 , n247516 );
and ( n247589 , n247588 , n247522 );
and ( n247590 , n247575 , n247516 );
or ( n247591 , n247589 , n247590 );
xor ( n247592 , n247581 , n247587 );
xor ( n247593 , n247592 , n247528 );
xor ( n247594 , n247581 , n247587 );
and ( n247595 , n247594 , n247528 );
and ( n247596 , n247581 , n247587 );
or ( n247597 , n247595 , n247596 );
or ( n247598 , n239441 , n242888 );
nand ( n247599 , n247598 , n246417 );
or ( n247600 , n247571 , n239784 );
and ( n247601 , n242596 , n209968 );
not ( n247602 , n242596 );
and ( n247603 , n247602 , n247455 );
nor ( n247604 , n247601 , n247603 );
or ( n247605 , n247604 , n247079 );
nand ( n247606 , n247600 , n247605 );
xor ( n247607 , n247599 , n247606 );
or ( n247608 , n247539 , n247210 );
and ( n247609 , n39288 , n244654 );
and ( n247610 , n39287 , n247318 );
nor ( n247611 , n247609 , n247610 );
or ( n247612 , n247611 , n237013 );
nand ( n247613 , n247608 , n247612 );
xor ( n247614 , n247607 , n247613 );
xor ( n247615 , n247599 , n247606 );
and ( n247616 , n247615 , n247613 );
and ( n247617 , n247599 , n247606 );
or ( n247618 , n247616 , n247617 );
and ( n247619 , n234382 , n246556 );
not ( n247620 , n234382 );
and ( n247621 , n247620 , n239932 );
nor ( n247622 , n247619 , n247621 );
not ( n247623 , n247622 );
not ( n247624 , n247623 );
not ( n247625 , n238274 );
or ( n247626 , n247624 , n247625 );
or ( n247627 , n247546 , n247497 );
nand ( n247628 , n247626 , n247627 );
or ( n247629 , n247564 , n247559 );
and ( n247630 , n243764 , n244643 );
and ( n247631 , n243765 , n238619 );
nor ( n247632 , n247630 , n247631 );
or ( n247633 , n247632 , n237041 );
nand ( n247634 , n247629 , n247633 );
xor ( n247635 , n247628 , n247634 );
nor ( n247636 , n243754 , n243297 );
xor ( n247637 , n247635 , n247636 );
xor ( n247638 , n247628 , n247634 );
and ( n247639 , n247638 , n247636 );
and ( n247640 , n247628 , n247634 );
or ( n247641 , n247639 , n247640 );
xor ( n247642 , n247573 , n247557 );
xor ( n247643 , n247642 , n247637 );
xor ( n247644 , n247573 , n247557 );
and ( n247645 , n247644 , n247637 );
and ( n247646 , n247573 , n247557 );
or ( n247647 , n247645 , n247646 );
xor ( n247648 , n247614 , n247579 );
xor ( n247649 , n247648 , n247643 );
xor ( n247650 , n247614 , n247579 );
and ( n247651 , n247650 , n247643 );
and ( n247652 , n247614 , n247579 );
or ( n247653 , n247651 , n247652 );
xor ( n247654 , n247585 , n247649 );
xor ( n247655 , n247654 , n247591 );
xor ( n247656 , n247585 , n247649 );
and ( n247657 , n247656 , n247591 );
and ( n247658 , n247585 , n247649 );
or ( n247659 , n247657 , n247658 );
or ( n247660 , n247622 , n239269 );
and ( n247661 , n39368 , n243297 );
and ( n247662 , n39367 , n234382 );
nor ( n247663 , n247661 , n247662 );
or ( n247664 , n247663 , n240148 );
nand ( n247665 , n247660 , n247664 );
not ( n247666 , n243297 );
and ( n247667 , n238857 , n247666 );
xor ( n247668 , n247665 , n247667 );
not ( n247669 , n242596 );
not ( n247670 , n246590 );
or ( n247671 , n247669 , n247670 );
or ( n247672 , n247604 , n239784 );
nand ( n247673 , n247671 , n247672 );
xor ( n247674 , n247668 , n247673 );
xor ( n247675 , n247665 , n247667 );
and ( n247676 , n247675 , n247673 );
and ( n247677 , n247665 , n247667 );
or ( n247678 , n247676 , n247677 );
or ( n247679 , n247611 , n247210 );
not ( n247680 , n237271 );
and ( n247681 , n247680 , n244654 );
and ( n247682 , n237271 , n247318 );
nor ( n247683 , n247681 , n247682 );
or ( n247684 , n247683 , n237013 );
nand ( n247685 , n247679 , n247684 );
or ( n247686 , n247632 , n247559 );
and ( n247687 , n238619 , n245282 );
not ( n247688 , n238619 );
and ( n247689 , n247688 , n246922 );
nor ( n247690 , n247687 , n247689 );
or ( n247691 , n247690 , n237041 );
nand ( n247692 , n247686 , n247691 );
not ( n247693 , n247692 );
xor ( n247694 , n247685 , n247693 );
xor ( n247695 , n247694 , n247641 );
xor ( n247696 , n247685 , n247693 );
and ( n247697 , n247696 , n247641 );
and ( n247698 , n247685 , n247693 );
or ( n247699 , n247697 , n247698 );
xor ( n247700 , n247618 , n247674 );
xor ( n247701 , n247700 , n247695 );
xor ( n247702 , n247618 , n247674 );
and ( n247703 , n247702 , n247695 );
and ( n247704 , n247618 , n247674 );
or ( n247705 , n247703 , n247704 );
xor ( n247706 , n247647 , n247701 );
xor ( n247707 , n247706 , n247653 );
xor ( n247708 , n247647 , n247701 );
and ( n247709 , n247708 , n247653 );
and ( n247710 , n247647 , n247701 );
or ( n247711 , n247709 , n247710 );
or ( n247712 , n237810 , n246590 );
nand ( n247713 , n247712 , n242596 );
not ( n247714 , n239794 );
not ( n247715 , n247690 );
not ( n247716 , n247715 );
or ( n247717 , n247714 , n247716 );
not ( n247718 , n209969 );
and ( n247719 , n247718 , n244643 );
and ( n247720 , n209969 , n238619 );
nor ( n247721 , n247719 , n247720 );
or ( n247722 , n247721 , n237041 );
nand ( n247723 , n247717 , n247722 );
xor ( n247724 , n247713 , n247723 );
or ( n247725 , n247663 , n239269 );
and ( n247726 , n39288 , n243297 );
and ( n247727 , n39287 , n234382 );
nor ( n247728 , n247726 , n247727 );
or ( n247729 , n247728 , n240148 );
nand ( n247730 , n247725 , n247729 );
xor ( n247731 , n247724 , n247730 );
xor ( n247732 , n247713 , n247723 );
and ( n247733 , n247732 , n247730 );
and ( n247734 , n247713 , n247723 );
or ( n247735 , n247733 , n247734 );
not ( n247736 , n239932 );
nor ( n247737 , n247736 , n243297 );
or ( n247738 , n247683 , n247210 );
and ( n247739 , n247318 , n243765 );
not ( n247740 , n247318 );
and ( n247741 , n247740 , n243764 );
nor ( n247742 , n247739 , n247741 );
or ( n247743 , n247742 , n237013 );
nand ( n247744 , n247738 , n247743 );
xor ( n247745 , n247737 , n247744 );
xor ( n247746 , n247745 , n247692 );
xor ( n247747 , n247737 , n247744 );
and ( n247748 , n247747 , n247692 );
and ( n247749 , n247737 , n247744 );
or ( n247750 , n247748 , n247749 );
xor ( n247751 , n247678 , n247731 );
xor ( n247752 , n247751 , n247746 );
xor ( n247753 , n247678 , n247731 );
and ( n247754 , n247753 , n247746 );
and ( n247755 , n247678 , n247731 );
or ( n247756 , n247754 , n247755 );
xor ( n247757 , n247699 , n247752 );
xor ( n247758 , n247757 , n247705 );
xor ( n247759 , n247699 , n247752 );
and ( n247760 , n247759 , n247705 );
and ( n247761 , n247699 , n247752 );
or ( n247762 , n247760 , n247761 );
nor ( n247763 , n39367 , n243297 );
or ( n247764 , n247742 , n247210 );
and ( n247765 , n209866 , n244654 );
and ( n247766 , n245282 , n247318 );
nor ( n247767 , n247765 , n247766 );
or ( n247768 , n247767 , n237013 );
nand ( n247769 , n247764 , n247768 );
xor ( n247770 , n247763 , n247769 );
or ( n247771 , n247728 , n247497 );
and ( n247772 , n247680 , n243297 );
and ( n247773 , n237271 , n247666 );
nor ( n247774 , n247772 , n247773 );
or ( n247775 , n247774 , n240148 );
nand ( n247776 , n247771 , n247775 );
xor ( n247777 , n247770 , n247776 );
xor ( n247778 , n247763 , n247769 );
and ( n247779 , n247778 , n247776 );
and ( n247780 , n247763 , n247769 );
or ( n247781 , n247779 , n247780 );
or ( n247782 , n247721 , n247559 );
or ( n247783 , n237041 , n244643 );
nand ( n247784 , n247782 , n247783 );
not ( n247785 , n247784 );
xor ( n247786 , n247785 , n247735 );
xor ( n247787 , n247786 , n247777 );
xor ( n247788 , n247785 , n247735 );
and ( n247789 , n247788 , n247777 );
and ( n247790 , n247785 , n247735 );
or ( n247791 , n247789 , n247790 );
xor ( n247792 , n247750 , n247787 );
xor ( n247793 , n247792 , n247756 );
xor ( n247794 , n247750 , n247787 );
and ( n247795 , n247794 , n247756 );
and ( n247796 , n247750 , n247787 );
or ( n247797 , n247795 , n247796 );
or ( n247798 , n239794 , n228868 );
nand ( n247799 , n247798 , n238619 );
not ( n247800 , n242737 );
or ( n247801 , n209970 , n239393 );
not ( n247802 , n209970 );
or ( n247803 , n247802 , n244654 );
nand ( n247804 , n247801 , n247803 );
not ( n247805 , n247804 );
or ( n247806 , n247800 , n247805 );
or ( n247807 , n247767 , n247210 );
nand ( n247808 , n247806 , n247807 );
xor ( n247809 , n247799 , n247808 );
nor ( n247810 , n39287 , n243297 );
xor ( n247811 , n247809 , n247810 );
xor ( n247812 , n247799 , n247808 );
and ( n247813 , n247812 , n247810 );
and ( n247814 , n247799 , n247808 );
or ( n247815 , n247813 , n247814 );
or ( n247816 , n247774 , n247497 );
and ( n247817 , n243764 , n243297 );
and ( n247818 , n243765 , n234382 );
nor ( n247819 , n247817 , n247818 );
or ( n247820 , n247819 , n240148 );
nand ( n247821 , n247816 , n247820 );
xor ( n247822 , n247821 , n247784 );
xor ( n247823 , n247822 , n247781 );
xor ( n247824 , n247821 , n247784 );
and ( n247825 , n247824 , n247781 );
and ( n247826 , n247821 , n247784 );
or ( n247827 , n247825 , n247826 );
xor ( n247828 , n247811 , n247823 );
xor ( n247829 , n247828 , n247791 );
xor ( n247830 , n247811 , n247823 );
and ( n247831 , n247830 , n247791 );
and ( n247832 , n247811 , n247823 );
or ( n247833 , n247831 , n247832 );
or ( n247834 , n247819 , n247497 );
and ( n247835 , n209867 , n243297 );
not ( n247836 , n209867 );
and ( n247837 , n247836 , n247666 );
nor ( n247838 , n247835 , n247837 );
or ( n247839 , n247838 , n240148 );
nand ( n247840 , n247834 , n247839 );
not ( n247841 , n247680 );
nor ( n247842 , n247841 , n243297 );
xor ( n247843 , n247840 , n247842 );
and ( n247844 , n247804 , n244387 );
and ( n247845 , n242737 , n239393 );
nor ( n247846 , n247844 , n247845 );
xor ( n247847 , n247843 , n247846 );
xor ( n247848 , n247840 , n247842 );
and ( n247849 , n247848 , n247846 );
and ( n247850 , n247840 , n247842 );
or ( n247851 , n247849 , n247850 );
xor ( n247852 , n247815 , n247847 );
xor ( n247853 , n247852 , n247827 );
xor ( n247854 , n247815 , n247847 );
and ( n247855 , n247854 , n247827 );
and ( n247856 , n247815 , n247847 );
or ( n247857 , n247855 , n247856 );
or ( n247858 , n244387 , n242737 );
nand ( n247859 , n247858 , n239393 );
or ( n247860 , n247838 , n247497 );
xnor ( n247861 , n209971 , n243297 );
or ( n247862 , n247861 , n240148 );
nand ( n247863 , n247860 , n247862 );
xor ( n247864 , n247859 , n247863 );
nor ( n247865 , n243765 , n243297 );
xor ( n247866 , n247864 , n247865 );
xor ( n247867 , n247859 , n247863 );
and ( n247868 , n247867 , n247865 );
and ( n247869 , n247859 , n247863 );
or ( n247870 , n247868 , n247869 );
not ( n247871 , n247846 );
xor ( n247872 , n247871 , n247866 );
xor ( n247873 , n247872 , n247851 );
xor ( n247874 , n247871 , n247866 );
and ( n247875 , n247874 , n247851 );
and ( n247876 , n247871 , n247866 );
or ( n247877 , n247875 , n247876 );
or ( n247878 , n247861 , n247497 );
nand ( n247879 , n238274 , n247666 );
nand ( n247880 , n247878 , n247879 );
nand ( n247881 , n209867 , n247666 );
xor ( n247882 , n247880 , n247881 );
xor ( n247883 , n247882 , n247870 );
xor ( n247884 , n247880 , n247881 );
and ( n247885 , n247884 , n247870 );
and ( n247886 , n247880 , n247881 );
or ( n247887 , n247885 , n247886 );
or ( n247888 , n247762 , n247793 );
not ( n247889 , n247888 );
nor ( n247890 , n245197 , n244985 );
nor ( n247891 , n245402 , n245201 );
nor ( n247892 , n247890 , n247891 );
not ( n247893 , n245603 );
not ( n247894 , n245406 );
nand ( n247895 , n247893 , n247894 );
buf ( n247896 , n247895 );
or ( n247897 , n245607 , n245785 );
and ( n247898 , n247892 , n247896 , n247897 );
not ( n247899 , n247898 );
nor ( n247900 , n245969 , n246135 );
not ( n247901 , n247900 );
or ( n247902 , n246139 , n246301 );
nand ( n247903 , n247901 , n247902 );
nor ( n247904 , n245789 , n245965 );
nor ( n247905 , n247903 , n247904 );
buf ( n247906 , n247905 );
nor ( n247907 , n246486 , n246305 );
nor ( n247908 , n246490 , n246638 );
nor ( n247909 , n247907 , n247908 );
or ( n247910 , n246642 , n246778 );
not ( n247911 , n247910 );
nor ( n247912 , n246782 , n246911 );
nor ( n247913 , n247911 , n247912 );
nand ( n247914 , n247909 , n247913 );
not ( n247915 , n247035 );
not ( n247916 , n247149 );
and ( n247917 , n247915 , n247916 );
nor ( n247918 , n247031 , n246915 );
nor ( n247919 , n247917 , n247918 );
or ( n247920 , n247363 , n247445 );
not ( n247921 , n247920 );
nor ( n247922 , n247359 , n247258 );
nor ( n247923 , n247153 , n247254 );
nor ( n247924 , n247921 , n247922 , n247923 );
nand ( n247925 , n247919 , n247924 );
nor ( n247926 , n247914 , n247925 );
nand ( n247927 , n247906 , n247926 );
nor ( n247928 , n247899 , n247927 );
or ( n247929 , n247530 , n247449 );
nor ( n247930 , n247593 , n247534 );
not ( n247931 , n247930 );
nand ( n247932 , n247929 , n247931 );
or ( n247933 , n247659 , n247707 );
or ( n247934 , n247597 , n247655 );
or ( n247935 , n247711 , n247758 );
nand ( n247936 , n247933 , n247934 , n247935 );
nor ( n247937 , n247932 , n247936 );
and ( n247938 , n247928 , n247937 );
not ( n247939 , n247938 );
or ( n247940 , n238563 , n238160 );
buf ( n247941 , n238567 );
buf ( n247942 , n238955 );
nor ( n247943 , n247941 , n247942 );
not ( n247944 , n247943 );
not ( n247945 , n239343 );
not ( n247946 , n239722 );
nand ( n247947 , n247945 , n247946 );
not ( n247948 , n238959 );
not ( n247949 , n239339 );
nand ( n247950 , n247948 , n247949 );
buf ( n247951 , n247950 );
nand ( n247952 , n247940 , n247944 , n247947 , n247951 );
nor ( n247953 , n240800 , n241131 );
nor ( n247954 , n241465 , n241135 );
nor ( n247955 , n247953 , n247954 );
nor ( n247956 , n241776 , n241469 );
nor ( n247957 , n241780 , n242091 );
nor ( n247958 , n247956 , n247957 );
and ( n247959 , n247955 , n247958 );
not ( n247960 , n240796 );
not ( n247961 , n240453 );
nand ( n247962 , n247960 , n247961 );
not ( n247963 , n240086 );
not ( n247964 , n239726 );
nand ( n247965 , n247963 , n247964 );
not ( n247966 , n240090 );
not ( n247967 , n240449 );
nand ( n247968 , n247966 , n247967 );
and ( n247969 , n247962 , n247965 , n247968 );
nand ( n247970 , n247959 , n247969 );
nor ( n247971 , n247952 , n247970 );
buf ( n247972 , n242691 );
buf ( n247973 , n242393 );
nor ( n247974 , n247972 , n247973 );
not ( n247975 , n247974 );
not ( n247976 , n242695 );
not ( n247977 , n242979 );
nand ( n247978 , n247976 , n247977 );
buf ( n247979 , n247978 );
or ( n247980 , n242389 , n242095 );
not ( n247981 , n243259 );
not ( n247982 , n242983 );
nand ( n247983 , n247981 , n247982 );
and ( n247984 , n247975 , n247979 , n247980 , n247983 );
nor ( n247985 , n244302 , n244055 );
nor ( n247986 , n244536 , n244306 );
nor ( n247987 , n247985 , n247986 );
nor ( n247988 , n244766 , n244540 );
nor ( n247989 , n244770 , n244981 );
nor ( n247990 , n247988 , n247989 );
nand ( n247991 , n247987 , n247990 );
not ( n247992 , n243803 );
not ( n247993 , n243536 );
nand ( n247994 , n247992 , n247993 );
not ( n247995 , n243263 );
not ( n247996 , n243532 );
nand ( n247997 , n247995 , n247996 );
not ( n247998 , n244051 );
not ( n247999 , n243807 );
nand ( n248000 , n247998 , n247999 );
nand ( n248001 , n247994 , n247997 , n248000 );
nor ( n248002 , n247991 , n248001 );
nand ( n248003 , n247984 , n248002 );
not ( n248004 , n248003 );
and ( n248005 , n247971 , n248004 );
not ( n248006 , n248005 );
not ( n248007 , n237339 );
not ( n248008 , n236928 );
nand ( n248009 , n248007 , n248008 );
not ( n248010 , n237343 );
not ( n248011 , n237756 );
nand ( n248012 , n248010 , n248011 );
not ( n248013 , n236499 );
not ( n248014 , n236924 );
nand ( n248015 , n248013 , n248014 );
and ( n248016 , n248009 , n248012 , n248015 );
buf ( n248017 , n234199 );
buf ( n248018 , n233713 );
nor ( n248019 , n248017 , n248018 );
nor ( n248020 , n233709 , n233230 );
nor ( n248021 , n248019 , n248020 );
not ( n248022 , n235139 );
not ( n248023 , n234680 );
and ( n248024 , n248022 , n248023 );
not ( n248025 , n234676 );
not ( n248026 , n234203 );
nand ( n248027 , n248025 , n248026 );
not ( n248028 , n248027 );
nor ( n248029 , n248024 , n248028 );
nand ( n248030 , n248021 , n248029 );
not ( n248031 , n248030 );
nor ( n248032 , n236048 , n235593 );
nor ( n248033 , n236052 , n236495 );
nor ( n248034 , n235589 , n235143 );
nor ( n248035 , n248032 , n248033 , n248034 );
or ( n248036 , n238156 , n237760 );
and ( n248037 , n248016 , n248031 , n248035 , n248036 );
not ( n248038 , n248037 );
nor ( n248039 , n230104 , n230636 );
nor ( n248040 , n231198 , n230640 );
nor ( n248041 , n248039 , n248040 );
buf ( n248042 , n231714 );
not ( n248043 , n248042 );
not ( n248044 , n231202 );
nand ( n248045 , n248043 , n248044 );
or ( n248046 , n232220 , n231718 );
nand ( n248047 , n248041 , n248045 , n248046 );
or ( n248048 , n232727 , n232224 );
or ( n248049 , n233226 , n232731 );
nand ( n248050 , n248048 , n248049 );
nor ( n248051 , n248047 , n248050 );
not ( n248052 , n248051 );
or ( n248053 , n229063 , n229556 );
not ( n248054 , n248053 );
nor ( n248055 , n229059 , n228553 );
not ( n248056 , n248055 );
not ( n248057 , n248056 );
not ( n248058 , n228549 );
not ( n248059 , n228055 );
nand ( n248060 , n248058 , n248059 );
not ( n248061 , n248060 );
nor ( n248062 , n228051 , n227551 );
nand ( n248063 , n227547 , n227090 );
or ( n248064 , n248062 , n248063 );
nand ( n248065 , n228051 , n227551 );
nand ( n248066 , n248064 , n248065 );
not ( n248067 , n248066 );
or ( n248068 , n248061 , n248067 );
nand ( n248069 , n228549 , n228055 );
nand ( n248070 , n248068 , n248069 );
not ( n248071 , n248070 );
or ( n248072 , n248057 , n248071 );
nand ( n248073 , n229059 , n228553 );
nand ( n248074 , n248072 , n248073 );
not ( n248075 , n248074 );
or ( n248076 , n248054 , n248075 );
nand ( n248077 , n229063 , n229556 );
nand ( n248078 , n248076 , n248077 );
nor ( n248079 , n230100 , n229560 );
not ( n248080 , n248079 );
nand ( n248081 , n248078 , n248080 );
nor ( n248082 , n225244 , n224778 );
not ( n248083 , n248082 );
or ( n248084 , n225248 , n225672 );
or ( n248085 , n226130 , n225676 );
nand ( n248086 , n248083 , n248084 , n248085 );
or ( n248087 , n227086 , n226584 );
or ( n248088 , n226580 , n226134 );
nand ( n248089 , n248087 , n248088 );
nor ( n248090 , n248086 , n248089 );
not ( n248091 , n248090 );
nor ( n248092 , n223467 , n223884 );
nor ( n248093 , n223463 , n223040 );
nor ( n248094 , n248092 , n248093 );
not ( n248095 , n224774 );
not ( n248096 , n224344 );
nand ( n248097 , n248095 , n248096 );
or ( n248098 , n224340 , n223888 );
and ( n248099 , n248094 , n248097 , n248098 );
not ( n248100 , n248099 );
nor ( n248101 , n222648 , n222229 );
nor ( n248102 , n222652 , n223036 );
nor ( n248103 , n222225 , n221834 );
nor ( n248104 , n248101 , n248102 , n248103 );
not ( n248105 , n248104 );
nor ( n248106 , n221830 , n221437 );
nor ( n248107 , n221085 , n221433 );
nor ( n248108 , n221081 , n220693 );
nor ( n248109 , n248106 , n248107 , n248108 );
not ( n248110 , n248109 );
not ( n248111 , n220689 );
not ( n248112 , n220336 );
and ( n248113 , n248111 , n248112 );
not ( n248114 , n220332 );
not ( n248115 , n219964 );
and ( n248116 , n248114 , n248115 );
nor ( n248117 , n248113 , n248116 );
not ( n248118 , n248117 );
nor ( n248119 , n218940 , n218613 );
nor ( n248120 , n218609 , n218320 );
nor ( n248121 , n218316 , n218014 );
nor ( n248122 , n248119 , n248120 , n248121 );
not ( n248123 , n248122 );
nor ( n248124 , n218010 , n217735 );
nor ( n248125 , n217731 , n217427 );
nor ( n248126 , n248124 , n248125 );
not ( n248127 , n248126 );
nor ( n248128 , n217423 , n217169 );
nor ( n248129 , n217165 , n216877 );
nor ( n248130 , n248128 , n248129 );
not ( n248131 , n248130 );
nor ( n248132 , n216873 , n216642 );
nor ( n248133 , n216638 , n216357 );
nor ( n248134 , n248132 , n248133 );
not ( n248135 , n248134 );
not ( n248136 , n215679 );
not ( n248137 , n215466 );
and ( n248138 , n248136 , n248137 );
nor ( n248139 , n215462 , n215264 );
nor ( n248140 , n248138 , n248139 );
not ( n248141 , n248140 );
nor ( n248142 , n215260 , n215048 );
nor ( n248143 , n215044 , n214866 );
nor ( n248144 , n248142 , n248143 );
not ( n248145 , n248144 );
or ( n248146 , n214862 , n214671 );
not ( n248147 , n248146 );
nor ( n248148 , n214667 , n214514 );
not ( n248149 , n248148 );
not ( n248150 , n248149 );
nor ( n248151 , n214510 , n214343 );
not ( n248152 , n248151 );
not ( n248153 , n248152 );
nor ( n248154 , n214339 , n214216 );
nor ( n248155 , n214212 , n214053 );
nor ( n248156 , n248154 , n248155 );
not ( n248157 , n248156 );
or ( n248158 , n214049 , n213936 );
not ( n248159 , n248158 );
or ( n248160 , n213932 , n213797 );
not ( n248161 , n248160 );
or ( n248162 , n213793 , n213682 );
not ( n248163 , n248162 );
or ( n248164 , n213678 , n213569 );
not ( n248165 , n248164 );
nor ( n248166 , n213483 , n213398 );
or ( n248167 , n213394 , n213334 );
xor ( n248168 , n213180 , n213239 );
xor ( n248169 , n213090 , n213097 );
not ( n248170 , n211314 );
and ( n248171 , n213087 , n213144 );
not ( n248172 , n213087 );
and ( n248173 , n248172 , n213421 );
or ( n248174 , n248171 , n248173 );
not ( n248175 , n248174 );
or ( n248176 , n248170 , n248175 );
and ( n248177 , n213087 , n30666 );
not ( n248178 , n213087 );
and ( n248179 , n248178 , n213062 );
or ( n248180 , n248177 , n248179 );
or ( n248181 , n248180 , n213172 );
nand ( n248182 , n248176 , n248181 );
xor ( n248183 , n248169 , n248182 );
nor ( n248184 , n213057 , n213104 );
xnor ( n248185 , n168522 , n37684 );
not ( n248186 , n248185 );
not ( n248187 , n213171 );
and ( n248188 , n248186 , n248187 );
and ( n248189 , n213086 , n209375 );
nor ( n248190 , n248189 , n213084 );
nor ( n248191 , n248190 , n213172 );
nor ( n248192 , n248188 , n248191 );
nor ( n248193 , n213084 , n213171 );
not ( n248194 , n248193 );
nand ( n248195 , n248194 , n213087 );
nor ( n248196 , n248192 , n248195 );
xor ( n248197 , n248184 , n248196 );
or ( n248198 , n248180 , n213171 );
or ( n248199 , n248185 , n213172 );
nand ( n248200 , n248198 , n248199 );
and ( n248201 , n248197 , n248200 );
or ( n248202 , n248201 , C0 );
and ( n248203 , n248183 , n248202 );
and ( n248204 , n248169 , n248182 );
or ( n248205 , n248203 , n248204 );
not ( n248206 , n248205 );
not ( n248207 , n213099 );
and ( n248208 , n213170 , n211314 );
not ( n248209 , n248174 );
nor ( n248210 , n248209 , n213172 );
nor ( n248211 , n248208 , n248210 );
nand ( n248212 , n248207 , n248211 );
not ( n248213 , n248212 );
or ( n248214 , n248206 , n248213 );
not ( n248215 , n248207 );
not ( n248216 , n248211 );
nand ( n248217 , n248215 , n248216 );
nand ( n248218 , n248214 , n248217 );
xor ( n248219 , n213103 , n248218 );
and ( n248220 , n248219 , n213176 );
and ( n248221 , n213103 , n248218 );
or ( n248222 , n248220 , n248221 );
and ( n248223 , n248168 , n248222 );
and ( n248224 , n213180 , n213239 );
or ( n248225 , n248223 , n248224 );
not ( n248226 , n248225 );
or ( n248227 , n213330 , n213243 );
not ( n248228 , n248227 );
or ( n248229 , n248226 , n248228 );
nand ( n248230 , n213243 , n213330 );
nand ( n248231 , n248229 , n248230 );
and ( n248232 , n248167 , n248231 );
and ( n248233 , n213394 , n213334 );
nor ( n248234 , n248232 , n248233 );
or ( n248235 , n248166 , n248234 );
nand ( n248236 , n213483 , n213398 );
nand ( n248237 , n248235 , n248236 );
not ( n248238 , n248237 );
or ( n248239 , n213565 , n213487 );
not ( n248240 , n248239 );
or ( n248241 , n248238 , n248240 );
nand ( n248242 , n213565 , n213487 );
nand ( n248243 , n248241 , n248242 );
not ( n248244 , n248243 );
or ( n248245 , n248165 , n248244 );
nand ( n248246 , n213678 , n213569 );
nand ( n248247 , n248245 , n248246 );
not ( n248248 , n248247 );
or ( n248249 , n248163 , n248248 );
nand ( n248250 , n213793 , n213682 );
nand ( n248251 , n248249 , n248250 );
not ( n248252 , n248251 );
or ( n248253 , n248161 , n248252 );
nand ( n248254 , n213932 , n213797 );
nand ( n248255 , n248253 , n248254 );
not ( n248256 , n248255 );
or ( n248257 , n248159 , n248256 );
nand ( n248258 , n214049 , n213936 );
nand ( n248259 , n248257 , n248258 );
not ( n248260 , n248259 );
or ( n248261 , n248157 , n248260 );
nand ( n248262 , n214212 , n214053 );
not ( n248263 , n248262 );
nand ( n248264 , n214339 , n214216 );
not ( n248265 , n248264 );
or ( n248266 , n248263 , n248265 );
not ( n248267 , n248154 );
nand ( n248268 , n248266 , n248267 );
nand ( n248269 , n248261 , n248268 );
not ( n248270 , n248269 );
or ( n248271 , n248153 , n248270 );
nand ( n248272 , n214510 , n214343 );
nand ( n248273 , n248271 , n248272 );
not ( n248274 , n248273 );
or ( n248275 , n248150 , n248274 );
nand ( n248276 , n214667 , n214514 );
nand ( n248277 , n248275 , n248276 );
not ( n248278 , n248277 );
or ( n248279 , n248147 , n248278 );
nand ( n248280 , n214862 , n214671 );
nand ( n248281 , n248279 , n248280 );
not ( n248282 , n248281 );
or ( n248283 , n248145 , n248282 );
not ( n248284 , n248142 );
and ( n248285 , n215044 , n214866 );
and ( n248286 , n248284 , n248285 );
nand ( n248287 , n215260 , n215048 );
not ( n248288 , n248287 );
nor ( n248289 , n248286 , n248288 );
nand ( n248290 , n248283 , n248289 );
not ( n248291 , n248290 );
or ( n248292 , n248141 , n248291 );
or ( n248293 , n215679 , n215466 );
and ( n248294 , n215462 , n215264 );
and ( n248295 , n248293 , n248294 );
and ( n248296 , n215679 , n215466 );
nor ( n248297 , n248295 , n248296 );
nand ( n248298 , n248292 , n248297 );
nor ( n248299 , n216101 , n215860 );
nor ( n248300 , n215856 , n215683 );
nor ( n248301 , n248299 , n248300 );
nor ( n248302 , n216353 , n216105 );
not ( n248303 , n248302 );
nand ( n248304 , n248298 , n248301 , n248303 );
nand ( n248305 , n216101 , n215860 );
nand ( n248306 , n215856 , n215683 );
and ( n248307 , n248305 , n248306 );
nor ( n248308 , n248307 , n248299 );
nand ( n248309 , n248303 , n248308 );
nand ( n248310 , n216105 , n216353 );
nand ( n248311 , n248304 , n248309 , n248310 );
not ( n248312 , n248311 );
or ( n248313 , n248135 , n248312 );
not ( n248314 , n248132 );
nand ( n248315 , n216638 , n216357 );
not ( n248316 , n248315 );
and ( n248317 , n248314 , n248316 );
nand ( n248318 , n216873 , n216642 );
not ( n248319 , n248318 );
nor ( n248320 , n248317 , n248319 );
nand ( n248321 , n248313 , n248320 );
not ( n248322 , n248321 );
or ( n248323 , n248131 , n248322 );
not ( n248324 , n248128 );
nand ( n248325 , n217165 , n216877 );
not ( n248326 , n248325 );
and ( n248327 , n248324 , n248326 );
and ( n248328 , n217423 , n217169 );
nor ( n248329 , n248327 , n248328 );
nand ( n248330 , n248323 , n248329 );
not ( n248331 , n248330 );
or ( n248332 , n248127 , n248331 );
not ( n248333 , n248124 );
nand ( n248334 , n217731 , n217427 );
not ( n248335 , n248334 );
and ( n248336 , n248333 , n248335 );
nand ( n248337 , n218010 , n217735 );
not ( n248338 , n248337 );
nor ( n248339 , n248336 , n248338 );
nand ( n248340 , n248332 , n248339 );
not ( n248341 , n248340 );
or ( n248342 , n248123 , n248341 );
nand ( n248343 , n218316 , n218014 );
nor ( n248344 , n248120 , n248343 );
not ( n248345 , n218613 );
not ( n248346 , n218940 );
or ( n248347 , n248345 , n248346 );
nand ( n248348 , n218609 , n218320 );
nand ( n248349 , n248347 , n248348 );
or ( n248350 , n248344 , n248349 );
or ( n248351 , n218940 , n218613 );
nand ( n248352 , n248350 , n248351 );
nand ( n248353 , n248342 , n248352 );
not ( n248354 , n248353 );
nor ( n248355 , n219626 , n219270 );
nor ( n248356 , n219266 , n218944 );
nor ( n248357 , n248355 , n248356 );
not ( n248358 , n219960 );
not ( n248359 , n219630 );
nand ( n248360 , n248358 , n248359 );
nand ( n248361 , n248357 , n248360 );
not ( n248362 , n248361 );
not ( n248363 , n248362 );
or ( n248364 , n248354 , n248363 );
nand ( n248365 , n219266 , n218944 );
or ( n248366 , n248355 , n248365 );
nand ( n248367 , n219626 , n219270 );
nand ( n248368 , n248366 , n248367 );
not ( n248369 , n219960 );
nand ( n248370 , n248369 , n248359 );
and ( n248371 , n248368 , n248370 );
and ( n248372 , n219960 , n219630 );
nor ( n248373 , n248371 , n248372 );
nand ( n248374 , n248364 , n248373 );
not ( n248375 , n248374 );
or ( n248376 , n248118 , n248375 );
nor ( n248377 , n220689 , n220336 );
not ( n248378 , n248377 );
nand ( n248379 , n220332 , n219964 );
not ( n248380 , n248379 );
and ( n248381 , n248378 , n248380 );
and ( n248382 , n220689 , n220336 );
nor ( n248383 , n248381 , n248382 );
nand ( n248384 , n248376 , n248383 );
not ( n248385 , n248384 );
or ( n248386 , n248110 , n248385 );
nor ( n248387 , n221433 , n221085 );
nand ( n248388 , n221081 , n220693 );
or ( n248389 , n248387 , n248388 );
nand ( n248390 , n221433 , n221085 );
nand ( n248391 , n248389 , n248390 );
or ( n248392 , n221830 , n221437 );
and ( n248393 , n248391 , n248392 );
and ( n248394 , n221830 , n221437 );
nor ( n248395 , n248393 , n248394 );
nand ( n248396 , n248386 , n248395 );
not ( n248397 , n248396 );
or ( n248398 , n248105 , n248397 );
nor ( n248399 , n222648 , n222229 );
nand ( n248400 , n222225 , n221834 );
or ( n248401 , n248399 , n248400 );
nand ( n248402 , n222229 , n222648 );
nand ( n248403 , n248401 , n248402 );
or ( n248404 , n222652 , n223036 );
and ( n248405 , n248403 , n248404 );
nand ( n248406 , n222652 , n223036 );
not ( n248407 , n248406 );
nor ( n248408 , n248405 , n248407 );
nand ( n248409 , n248398 , n248408 );
not ( n248410 , n248409 );
or ( n248411 , n248100 , n248410 );
nand ( n248412 , n224340 , n223888 );
not ( n248413 , n248412 );
and ( n248414 , n224774 , n224344 );
nor ( n248415 , n248413 , n248414 );
not ( n248416 , n248415 );
nand ( n248417 , n223463 , n223040 );
or ( n248418 , n248092 , n248417 );
nand ( n248419 , n223884 , n223467 );
nand ( n248420 , n248418 , n248419 );
nand ( n248421 , n248098 , n248420 );
not ( n248422 , n248421 );
or ( n248423 , n248416 , n248422 );
not ( n248424 , n224774 );
nand ( n248425 , n248424 , n248096 );
nand ( n248426 , n248423 , n248425 );
nand ( n248427 , n248411 , n248426 );
not ( n248428 , n248427 );
or ( n248429 , n248091 , n248428 );
nand ( n248430 , n227086 , n226584 );
not ( n248431 , n248430 );
not ( n248432 , n248431 );
not ( n248433 , n248432 );
nor ( n248434 , n227086 , n226584 );
not ( n248435 , n248434 );
or ( n248436 , n248433 , n248435 );
not ( n248437 , n226130 );
not ( n248438 , n225676 );
nand ( n248439 , n248437 , n248438 );
not ( n248440 , n248439 );
nor ( n248441 , n225672 , n225248 );
nand ( n248442 , n224778 , n225244 );
or ( n248443 , n248441 , n248442 );
nand ( n248444 , n225248 , n225672 );
nand ( n248445 , n248443 , n248444 );
not ( n248446 , n248445 );
or ( n248447 , n248440 , n248446 );
nand ( n248448 , n226130 , n225676 );
nand ( n248449 , n248447 , n248448 );
or ( n248450 , n226580 , n226134 );
nand ( n248451 , n248449 , n248450 );
nand ( n248452 , n226580 , n226134 );
nand ( n248453 , n248451 , n248432 , n248452 );
nand ( n248454 , n248436 , n248453 );
nand ( n248455 , n248429 , n248454 );
nor ( n248456 , n229059 , n228553 );
not ( n248457 , n248456 );
buf ( n248458 , n227547 );
buf ( n248459 , n227090 );
nor ( n248460 , n248458 , n248459 );
buf ( n248461 , n248062 );
nor ( n248462 , n248460 , n248461 );
not ( n248463 , n228549 );
nand ( n248464 , n248463 , n248059 );
nand ( n248465 , n248457 , n248462 , n248464 );
not ( n248466 , n248079 );
nand ( n248467 , n248466 , n248053 );
nor ( n248468 , n248465 , n248467 );
nand ( n248469 , n248455 , n248468 );
nand ( n248470 , n230100 , n229560 );
nand ( n248471 , n248081 , n248469 , n248470 );
not ( n248472 , n248471 );
or ( n248473 , n248052 , n248472 );
buf ( n248474 , n232727 );
not ( n248475 , n248474 );
not ( n248476 , n232224 );
and ( n248477 , n248475 , n248476 );
buf ( n248478 , n232731 );
nor ( n248479 , n248478 , n233226 );
nor ( n248480 , n248477 , n248479 );
nand ( n248481 , n233226 , n248478 );
not ( n248482 , n248481 );
or ( n248483 , n248480 , n248482 );
not ( n248484 , n231718 );
not ( n248485 , n248484 );
not ( n248486 , n232220 );
not ( n248487 , n248486 );
or ( n248488 , n248485 , n248487 );
not ( n248489 , n231714 );
nand ( n248490 , n248489 , n248044 );
not ( n248491 , n248490 );
nor ( n248492 , n231198 , n230640 );
nand ( n248493 , n230636 , n230104 );
or ( n248494 , n248492 , n248493 );
nand ( n248495 , n231198 , n230640 );
nand ( n248496 , n248494 , n248495 );
not ( n248497 , n248496 );
or ( n248498 , n248491 , n248497 );
nand ( n248499 , n248042 , n231202 );
nand ( n248500 , n248498 , n248499 );
nand ( n248501 , n248488 , n248500 );
nand ( n248502 , n248474 , n232224 );
nand ( n248503 , n232220 , n231718 );
nand ( n248504 , n248501 , n248502 , n248481 , n248503 );
nand ( n248505 , n248483 , n248504 );
nand ( n248506 , n248473 , n248505 );
not ( n248507 , n248506 );
or ( n248508 , n248038 , n248507 );
not ( n248509 , n248035 );
not ( n248510 , n235139 );
not ( n248511 , n234680 );
nand ( n248512 , n248510 , n248511 );
not ( n248513 , n248512 );
not ( n248514 , n234676 );
nand ( n248515 , n248514 , n248026 );
not ( n248516 , n248515 );
nor ( n248517 , n234199 , n233713 );
nand ( n248518 , n233709 , n233230 );
or ( n248519 , n248517 , n248518 );
nand ( n248520 , n234199 , n233713 );
nand ( n248521 , n248519 , n248520 );
not ( n248522 , n248521 );
or ( n248523 , n248516 , n248522 );
buf ( n248524 , n234676 );
nand ( n248525 , n248524 , n234203 );
nand ( n248526 , n248523 , n248525 );
not ( n248527 , n248526 );
or ( n248528 , n248513 , n248527 );
or ( n248529 , n248510 , n248511 );
nand ( n248530 , n248528 , n248529 );
not ( n248531 , n248530 );
or ( n248532 , n248509 , n248531 );
nor ( n248533 , n235593 , n236048 );
nand ( n248534 , n235589 , n235143 );
or ( n248535 , n248533 , n248534 );
nand ( n248536 , n236048 , n235593 );
nand ( n248537 , n248535 , n248536 );
or ( n248538 , n236052 , n236495 );
and ( n248539 , n248537 , n248538 );
nand ( n248540 , n236495 , n236052 );
not ( n248541 , n248540 );
nor ( n248542 , n248539 , n248541 );
nand ( n248543 , n248532 , n248542 );
nand ( n248544 , n248013 , n248014 );
and ( n248545 , n248009 , n248012 , n248036 , n248544 );
and ( n248546 , n248543 , n248545 );
not ( n248547 , n248011 );
nand ( n248548 , n248547 , n237343 );
not ( n248549 , n248548 );
nand ( n248550 , n248549 , n248036 );
nor ( n248551 , n248013 , n248014 );
not ( n248552 , n248551 );
not ( n248553 , n248009 );
or ( n248554 , n248552 , n248553 );
or ( n248555 , n248007 , n248008 );
nand ( n248556 , n248554 , n248555 );
nand ( n248557 , n248036 , n248556 , n248012 );
nand ( n248558 , n238156 , n237760 );
nand ( n248559 , n248550 , n248557 , n248558 );
nor ( n248560 , n248546 , n248559 );
nand ( n248561 , n248508 , n248560 );
not ( n248562 , n248561 );
or ( n248563 , n248006 , n248562 );
not ( n248564 , n247959 );
and ( n248565 , n247962 , n247965 , n247968 );
not ( n248566 , n248565 );
not ( n248567 , n247947 );
not ( n248568 , n247950 );
nor ( n248569 , n238567 , n238955 );
nand ( n248570 , n238563 , n238160 );
or ( n248571 , n248569 , n248570 );
nand ( n248572 , n238567 , n238955 );
nand ( n248573 , n248571 , n248572 );
not ( n248574 , n248573 );
or ( n248575 , n248568 , n248574 );
not ( n248576 , n247949 );
nand ( n248577 , n248576 , n238959 );
nand ( n248578 , n248575 , n248577 );
not ( n248579 , n248578 );
or ( n248580 , n248567 , n248579 );
not ( n248581 , n247946 );
nand ( n248582 , n248581 , n239343 );
nand ( n248583 , n248580 , n248582 );
not ( n248584 , n248583 );
or ( n248585 , n248566 , n248584 );
nand ( n248586 , n240086 , n239726 );
nor ( n248587 , n240449 , n240090 );
or ( n248588 , n248586 , n248587 );
nand ( n248589 , n240449 , n240090 );
nand ( n248590 , n248588 , n248589 );
nand ( n248591 , n247960 , n247961 );
and ( n248592 , n248590 , n248591 );
nor ( n248593 , n247960 , n247961 );
nor ( n248594 , n248592 , n248593 );
nand ( n248595 , n248585 , n248594 );
not ( n248596 , n248595 );
or ( n248597 , n248564 , n248596 );
not ( n248598 , n247956 );
not ( n248599 , n248598 );
nand ( n248600 , n240800 , n241131 );
or ( n248601 , n248600 , n247954 );
nand ( n248602 , n241465 , n241135 );
nand ( n248603 , n248601 , n248602 );
not ( n248604 , n248603 );
or ( n248605 , n248599 , n248604 );
nand ( n248606 , n241776 , n241469 );
nand ( n248607 , n248605 , n248606 );
not ( n248608 , n247957 );
and ( n248609 , n248607 , n248608 );
and ( n248610 , n241780 , n242091 );
nor ( n248611 , n248609 , n248610 );
nand ( n248612 , n248597 , n248611 );
and ( n248613 , n248612 , n248004 );
not ( n248614 , n247991 );
not ( n248615 , n248614 );
not ( n248616 , n248001 );
not ( n248617 , n248616 );
not ( n248618 , n247983 );
not ( n248619 , n247978 );
nor ( n248620 , n242691 , n242393 );
nand ( n248621 , n242389 , n242095 );
or ( n248622 , n248620 , n248621 );
nand ( n248623 , n242691 , n242393 );
nand ( n248624 , n248622 , n248623 );
not ( n248625 , n248624 );
or ( n248626 , n248619 , n248625 );
not ( n248627 , n247977 );
nand ( n248628 , n248627 , n242695 );
nand ( n248629 , n248626 , n248628 );
not ( n248630 , n248629 );
or ( n248631 , n248618 , n248630 );
nand ( n248632 , n243259 , n242983 );
nand ( n248633 , n248631 , n248632 );
not ( n248634 , n248633 );
or ( n248635 , n248617 , n248634 );
nor ( n248636 , n243803 , n243536 );
nand ( n248637 , n243263 , n243532 );
or ( n248638 , n248636 , n248637 );
nand ( n248639 , n243803 , n243536 );
nand ( n248640 , n248638 , n248639 );
buf ( n248641 , n248000 );
and ( n248642 , n248640 , n248641 );
nor ( n248643 , n247998 , n247999 );
nor ( n248644 , n248642 , n248643 );
nand ( n248645 , n248635 , n248644 );
not ( n248646 , n248645 );
or ( n248647 , n248615 , n248646 );
not ( n248648 , n247988 );
not ( n248649 , n248648 );
nor ( n248650 , n244536 , n244306 );
nand ( n248651 , n244302 , n244055 );
or ( n248652 , n248650 , n248651 );
nand ( n248653 , n244306 , n244536 );
nand ( n248654 , n248652 , n248653 );
not ( n248655 , n248654 );
or ( n248656 , n248649 , n248655 );
nand ( n248657 , n244766 , n244540 );
nand ( n248658 , n248656 , n248657 );
not ( n248659 , n247989 );
buf ( n248660 , n248659 );
and ( n248661 , n248658 , n248660 );
and ( n248662 , n244770 , n244981 );
nor ( n248663 , n248661 , n248662 );
nand ( n248664 , n248647 , n248663 );
nor ( n248665 , n248613 , n248664 );
nand ( n248666 , n248563 , n248665 );
not ( n248667 , n248666 );
or ( n248668 , n247939 , n248667 );
not ( n248669 , n247937 );
not ( n248670 , n247926 );
not ( n248671 , n247905 );
not ( n248672 , n247897 );
not ( n248673 , n247895 );
nand ( n248674 , n245197 , n244985 );
or ( n248675 , n247891 , n248674 );
nand ( n248676 , n245402 , n245201 );
nand ( n248677 , n248675 , n248676 );
not ( n248678 , n248677 );
or ( n248679 , n248673 , n248678 );
nand ( n248680 , n245603 , n245406 );
nand ( n248681 , n248679 , n248680 );
not ( n248682 , n248681 );
or ( n248683 , n248672 , n248682 );
nand ( n248684 , n245607 , n245785 );
nand ( n248685 , n248683 , n248684 );
not ( n248686 , n248685 );
or ( n248687 , n248671 , n248686 );
not ( n248688 , n247902 );
nand ( n248689 , n245789 , n245965 );
or ( n248690 , n248689 , n247900 );
nand ( n248691 , n245969 , n246135 );
nand ( n248692 , n248690 , n248691 );
not ( n248693 , n248692 );
or ( n248694 , n248688 , n248693 );
nand ( n248695 , n246139 , n246301 );
nand ( n248696 , n248694 , n248695 );
not ( n248697 , n248696 );
nand ( n248698 , n248687 , n248697 );
not ( n248699 , n248698 );
or ( n248700 , n248670 , n248699 );
not ( n248701 , n247919 );
not ( n248702 , n247912 );
not ( n248703 , n248702 );
not ( n248704 , n247910 );
nand ( n248705 , n246486 , n246305 );
or ( n248706 , n247908 , n248705 );
nand ( n248707 , n246490 , n246638 );
nand ( n248708 , n248706 , n248707 );
not ( n248709 , n248708 );
or ( n248710 , n248704 , n248709 );
nand ( n248711 , n246642 , n246778 );
nand ( n248712 , n248710 , n248711 );
not ( n248713 , n248712 );
or ( n248714 , n248703 , n248713 );
nand ( n248715 , n246782 , n246911 );
nand ( n248716 , n248714 , n248715 );
not ( n248717 , n248716 );
or ( n248718 , n248701 , n248717 );
or ( n248719 , n247149 , n247035 );
and ( n248720 , n246915 , n247031 );
and ( n248721 , n248719 , n248720 );
nand ( n248722 , n247149 , n247035 );
not ( n248723 , n248722 );
nor ( n248724 , n248721 , n248723 );
nand ( n248725 , n248718 , n248724 );
and ( n248726 , n248725 , n247924 );
not ( n248727 , n247920 );
nand ( n248728 , n247153 , n247254 );
or ( n248729 , n248728 , n247922 );
nand ( n248730 , n247359 , n247258 );
nand ( n248731 , n248729 , n248730 );
not ( n248732 , n248731 );
or ( n248733 , n248727 , n248732 );
nand ( n248734 , n247363 , n247445 );
nand ( n248735 , n248733 , n248734 );
nor ( n248736 , n248726 , n248735 );
nand ( n248737 , n248700 , n248736 );
not ( n248738 , n248737 );
or ( n248739 , n248669 , n248738 );
nand ( n248740 , n247530 , n247449 );
or ( n248741 , n248740 , n247930 );
nand ( n248742 , n247593 , n247534 );
nand ( n248743 , n248741 , n248742 );
not ( n248744 , n247936 );
and ( n248745 , n248743 , n248744 );
not ( n248746 , n247935 );
nor ( n248747 , n247659 , n247707 );
nand ( n248748 , n247597 , n247655 );
or ( n248749 , n248747 , n248748 );
nand ( n248750 , n247659 , n247707 );
nand ( n248751 , n248749 , n248750 );
not ( n248752 , n248751 );
or ( n248753 , n248746 , n248752 );
nand ( n248754 , n247711 , n247758 );
nand ( n248755 , n248753 , n248754 );
nor ( n248756 , n248745 , n248755 );
nand ( n248757 , n248739 , n248756 );
buf ( n248758 , n248757 );
not ( n248759 , n248758 );
nand ( n248760 , n248668 , n248759 );
not ( n248761 , n248760 );
or ( n248762 , n247889 , n248761 );
nand ( n248763 , n247762 , n247793 );
nand ( n248764 , n248762 , n248763 );
nor ( n248765 , n247797 , n247829 );
not ( n248766 , n248765 );
nand ( n248767 , n247797 , n247829 );
nand ( n248768 , n248766 , n248767 );
not ( n248769 , n248768 );
and ( n248770 , n248764 , n248769 );
not ( n248771 , n248764 );
and ( n248772 , n248771 , n248768 );
nor ( n248773 , n248770 , n248772 );
not ( n248774 , n247896 );
not ( n248775 , n247892 );
not ( n248776 , n248666 );
or ( n248777 , n248775 , n248776 );
not ( n248778 , n248677 );
nand ( n248779 , n248777 , n248778 );
not ( n248780 , n248779 );
or ( n248781 , n248774 , n248780 );
nand ( n248782 , n248781 , n248680 );
nand ( n248783 , n247897 , n248684 );
not ( n248784 , n248783 );
and ( n248785 , n248782 , n248784 );
not ( n248786 , n248782 );
and ( n248787 , n248786 , n248783 );
nor ( n248788 , n248785 , n248787 );
not ( n248789 , n248598 );
buf ( n248790 , n247969 );
buf ( n248791 , n247955 );
and ( n248792 , n248790 , n248791 );
not ( n248793 , n248792 );
not ( n248794 , n247952 );
not ( n248795 , n248794 );
not ( n248796 , n248561 );
or ( n248797 , n248795 , n248796 );
buf ( n248798 , n248583 );
not ( n248799 , n248798 );
nand ( n248800 , n248797 , n248799 );
not ( n248801 , n248800 );
or ( n248802 , n248793 , n248801 );
buf ( n248803 , n248594 );
not ( n248804 , n248803 );
and ( n248805 , n248804 , n248791 );
buf ( n248806 , n248603 );
nor ( n248807 , n248805 , n248806 );
nand ( n248808 , n248802 , n248807 );
not ( n248809 , n248808 );
or ( n248810 , n248789 , n248809 );
nand ( n248811 , n248810 , n248606 );
not ( n248812 , n248610 );
nand ( n248813 , n248812 , n248608 );
not ( n248814 , n248813 );
and ( n248815 , n248811 , n248814 );
not ( n248816 , n248811 );
and ( n248817 , n248816 , n248813 );
nor ( n248818 , n248815 , n248817 );
not ( n248819 , n247929 );
buf ( n248820 , n248004 );
not ( n248821 , n247898 );
nor ( n248822 , n248821 , n247927 );
nand ( n248823 , n248820 , n248822 );
not ( n248824 , n248823 );
not ( n248825 , n248824 );
buf ( n248826 , n247971 );
not ( n248827 , n248826 );
not ( n248828 , n248037 );
not ( n248829 , n248506 );
or ( n248830 , n248828 , n248829 );
and ( n248831 , n248543 , n248545 );
nor ( n248832 , n248831 , n248559 );
nand ( n248833 , n248830 , n248832 );
not ( n248834 , n248833 );
or ( n248835 , n248827 , n248834 );
not ( n248836 , n248612 );
nand ( n248837 , n248835 , n248836 );
not ( n248838 , n248837 );
or ( n248839 , n248825 , n248838 );
not ( n248840 , n248822 );
not ( n248841 , n248664 );
or ( n248842 , n248840 , n248841 );
not ( n248843 , n248737 );
nand ( n248844 , n248842 , n248843 );
not ( n248845 , n248844 );
nand ( n248846 , n248839 , n248845 );
not ( n248847 , n248846 );
or ( n248848 , n248819 , n248847 );
nand ( n248849 , n248848 , n248740 );
nand ( n248850 , n247931 , n248742 );
not ( n248851 , n248850 );
and ( n248852 , n248849 , n248851 );
not ( n248853 , n248849 );
and ( n248854 , n248853 , n248850 );
nor ( n248855 , n248852 , n248854 );
not ( n248856 , n247914 );
and ( n248857 , n247906 , n248856 );
not ( n248858 , n248857 );
nor ( n248859 , n248858 , n247918 );
not ( n248860 , n248859 );
buf ( n248861 , n248833 );
buf ( n248862 , n247898 );
nand ( n248863 , n248005 , n248862 );
not ( n248864 , n248863 );
nand ( n248865 , n248861 , n248864 );
and ( n248866 , n248004 , n247898 );
and ( n248867 , n248866 , n248612 );
not ( n248868 , n248614 );
not ( n248869 , n248645 );
or ( n248870 , n248868 , n248869 );
nand ( n248871 , n248870 , n248663 );
nand ( n248872 , n248871 , n247898 );
buf ( n248873 , n248685 );
not ( n248874 , n248873 );
nand ( n248875 , n248872 , n248874 );
nor ( n248876 , n248867 , n248875 );
nand ( n248877 , n248865 , n248876 );
not ( n248878 , n248877 );
or ( n248879 , n248860 , n248878 );
not ( n248880 , n248856 );
not ( n248881 , n248696 );
or ( n248882 , n248880 , n248881 );
not ( n248883 , n248716 );
nand ( n248884 , n248882 , n248883 );
not ( n248885 , n247918 );
and ( n248886 , n248884 , n248885 );
nor ( n248887 , n248886 , n248720 );
nand ( n248888 , n248879 , n248887 );
nand ( n248889 , n248719 , n248722 );
not ( n248890 , n248889 );
and ( n248891 , n248888 , n248890 );
not ( n248892 , n248888 );
and ( n248893 , n248892 , n248889 );
nor ( n248894 , n248891 , n248893 );
not ( n248895 , n247904 );
not ( n248896 , n248895 );
not ( n248897 , n248877 );
or ( n248898 , n248896 , n248897 );
nand ( n248899 , n248898 , n248689 );
nand ( n248900 , n247901 , n248691 );
not ( n248901 , n248900 );
and ( n248902 , n248899 , n248901 );
not ( n248903 , n248899 );
and ( n248904 , n248903 , n248900 );
nor ( n248905 , n248902 , n248904 );
nand ( n248906 , n247906 , n247909 );
nor ( n248907 , n248906 , n247911 );
not ( n248908 , n248907 );
not ( n248909 , n248877 );
or ( n248910 , n248908 , n248909 );
not ( n248911 , n247909 );
not ( n248912 , n248696 );
or ( n248913 , n248911 , n248912 );
not ( n248914 , n248708 );
nand ( n248915 , n248913 , n248914 );
or ( n248916 , n246642 , n246778 );
and ( n248917 , n248915 , n248916 );
not ( n248918 , n248711 );
nor ( n248919 , n248917 , n248918 );
nand ( n248920 , n248910 , n248919 );
nand ( n248921 , n248702 , n248715 );
not ( n248922 , n248921 );
and ( n248923 , n248920 , n248922 );
not ( n248924 , n248920 );
and ( n248925 , n248924 , n248921 );
nor ( n248926 , n248923 , n248925 );
not ( n248927 , n247906 );
not ( n248928 , n248877 );
or ( n248929 , n248927 , n248928 );
nand ( n248930 , n248929 , n248697 );
not ( n248931 , n247907 );
nand ( n248932 , n248931 , n248705 );
not ( n248933 , n248932 );
and ( n248934 , n248930 , n248933 );
not ( n248935 , n248930 );
and ( n248936 , n248935 , n248932 );
nor ( n248937 , n248934 , n248936 );
not ( n248938 , n247987 );
and ( n248939 , n247984 , n248616 );
nand ( n248940 , n248861 , n248826 , n248939 );
not ( n248941 , n248836 );
and ( n248942 , n248941 , n248939 );
buf ( n248943 , n248645 );
nor ( n248944 , n248942 , n248943 );
nand ( n248945 , n248940 , n248944 );
not ( n248946 , n248945 );
or ( n248947 , n248938 , n248946 );
not ( n248948 , n248654 );
nand ( n248949 , n248947 , n248948 );
nand ( n248950 , n248648 , n248657 );
not ( n248951 , n248950 );
and ( n248952 , n248949 , n248951 );
not ( n248953 , n248949 );
and ( n248954 , n248953 , n248950 );
nor ( n248955 , n248952 , n248954 );
not ( n248956 , n247985 );
not ( n248957 , n248956 );
not ( n248958 , n248945 );
or ( n248959 , n248957 , n248958 );
nand ( n248960 , n248959 , n248651 );
not ( n248961 , n248650 );
nand ( n248962 , n248961 , n248653 );
not ( n248963 , n248962 );
and ( n248964 , n248960 , n248963 );
not ( n248965 , n248960 );
and ( n248966 , n248965 , n248962 );
nor ( n248967 , n248964 , n248966 );
not ( n248968 , n248794 );
not ( n248969 , n248561 );
or ( n248970 , n248968 , n248969 );
not ( n248971 , n248798 );
nand ( n248972 , n248970 , n248971 );
nand ( n248973 , n248972 , n248790 );
buf ( n248974 , n247953 );
or ( n248975 , n248973 , n248974 );
not ( n248976 , n248974 );
and ( n248977 , n248804 , n248976 );
not ( n248978 , n248600 );
nor ( n248979 , n248977 , n248978 );
nand ( n248980 , n248975 , n248979 );
or ( n248981 , n241465 , n241135 );
nand ( n248982 , n248981 , n248602 );
not ( n248983 , n248982 );
and ( n248984 , n248980 , n248983 );
not ( n248985 , n248980 );
and ( n248986 , n248985 , n248982 );
nor ( n248987 , n248984 , n248986 );
not ( n248988 , n247965 );
nor ( n248989 , n248988 , n248587 );
not ( n248990 , n248989 );
not ( n248991 , n248972 );
or ( n248992 , n248990 , n248991 );
not ( n248993 , n248590 );
nand ( n248994 , n248992 , n248993 );
not ( n248995 , n248593 );
nand ( n248996 , n248995 , n248591 );
not ( n248997 , n248996 );
and ( n248998 , n248994 , n248997 );
not ( n248999 , n248994 );
and ( n249000 , n248999 , n248996 );
nor ( n249001 , n248998 , n249000 );
not ( n249002 , n247888 );
nor ( n249003 , n249002 , n248765 );
nand ( n249004 , n247937 , n249003 );
nor ( n249005 , n248823 , n249004 );
not ( n249006 , n249005 );
not ( n249007 , n248837 );
or ( n249008 , n249006 , n249007 );
not ( n249009 , n249004 );
and ( n249010 , n249009 , n248844 );
not ( n249011 , n248756 );
and ( n249012 , n249011 , n247888 );
not ( n249013 , n248763 );
nor ( n249014 , n249012 , n249013 );
or ( n249015 , n249014 , n248765 );
nand ( n249016 , n249015 , n248767 );
nor ( n249017 , n249010 , n249016 );
nand ( n249018 , n249008 , n249017 );
nor ( n249019 , n247833 , n247853 );
not ( n249020 , n249019 );
nand ( n249021 , n247833 , n247853 );
nand ( n249022 , n249020 , n249021 );
not ( n249023 , n249022 );
and ( n249024 , n249018 , n249023 );
not ( n249025 , n249018 );
and ( n249026 , n249025 , n249022 );
nor ( n249027 , n249024 , n249026 );
nor ( n249028 , n247923 , n247922 );
nand ( n249029 , n247919 , n249028 );
nor ( n249030 , n248858 , n249029 );
not ( n249031 , n249030 );
not ( n249032 , n248877 );
or ( n249033 , n249031 , n249032 );
not ( n249034 , n249029 );
and ( n249035 , n248884 , n249034 );
not ( n249036 , n248724 );
not ( n249037 , n247923 );
and ( n249038 , n249036 , n249037 );
not ( n249039 , n248728 );
nor ( n249040 , n249038 , n249039 );
or ( n249041 , n249040 , n247922 );
nand ( n249042 , n249041 , n248730 );
nor ( n249043 , n249035 , n249042 );
nand ( n249044 , n249033 , n249043 );
nand ( n249045 , n247920 , n248734 );
not ( n249046 , n249045 );
and ( n249047 , n249044 , n249046 );
not ( n249048 , n249044 );
and ( n249049 , n249048 , n249045 );
nor ( n249050 , n249047 , n249049 );
and ( n249051 , n247975 , n247983 , n247979 , n247980 );
nand ( n249052 , n249051 , n247997 );
not ( n249053 , n249052 );
not ( n249054 , n249053 );
buf ( n249055 , n248837 );
not ( n249056 , n249055 );
or ( n249057 , n249054 , n249056 );
not ( n249058 , n247997 );
not ( n249059 , n248633 );
or ( n249060 , n249058 , n249059 );
nand ( n249061 , n249060 , n248637 );
not ( n249062 , n249061 );
nand ( n249063 , n249057 , n249062 );
nand ( n249064 , n247994 , n248639 );
not ( n249065 , n249064 );
and ( n249066 , n249063 , n249065 );
not ( n249067 , n249063 );
and ( n249068 , n249067 , n249064 );
nor ( n249069 , n249066 , n249068 );
nor ( n249070 , n249052 , n248636 );
not ( n249071 , n249070 );
not ( n249072 , n249055 );
or ( n249073 , n249071 , n249072 );
nand ( n249074 , n249061 , n247994 );
and ( n249075 , n249074 , n248639 );
nand ( n249076 , n249073 , n249075 );
not ( n249077 , n248643 );
nand ( n249078 , n249077 , n248000 );
not ( n249079 , n249078 );
and ( n249080 , n249076 , n249079 );
not ( n249081 , n249076 );
and ( n249082 , n249081 , n249078 );
nor ( n249083 , n249080 , n249082 );
not ( n249084 , n247890 );
not ( n249085 , n249084 );
buf ( n249086 , n248666 );
not ( n249087 , n249086 );
or ( n249088 , n249085 , n249087 );
nand ( n249089 , n249088 , n248674 );
not ( n249090 , n247891 );
nand ( n249091 , n249090 , n248676 );
not ( n249092 , n249091 );
and ( n249093 , n249089 , n249092 );
not ( n249094 , n249089 );
and ( n249095 , n249094 , n249091 );
nor ( n249096 , n249093 , n249095 );
not ( n249097 , n248862 );
nand ( n249098 , n248895 , n247901 );
nor ( n249099 , n249097 , n249098 );
not ( n249100 , n249099 );
not ( n249101 , n249086 );
or ( n249102 , n249100 , n249101 );
not ( n249103 , n248895 );
not ( n249104 , n248873 );
or ( n249105 , n249103 , n249104 );
nand ( n249106 , n249105 , n248689 );
and ( n249107 , n249106 , n247901 );
not ( n249108 , n248691 );
nor ( n249109 , n249107 , n249108 );
nand ( n249110 , n249102 , n249109 );
nand ( n249111 , n247902 , n248695 );
not ( n249112 , n249111 );
and ( n249113 , n249110 , n249112 );
not ( n249114 , n249110 );
and ( n249115 , n249114 , n249111 );
nor ( n249116 , n249113 , n249115 );
nor ( n249117 , n249097 , n248906 );
not ( n249118 , n249117 );
not ( n249119 , n249086 );
or ( n249120 , n249118 , n249119 );
buf ( n249121 , n248698 );
and ( n249122 , n249121 , n247909 );
buf ( n249123 , n248708 );
nor ( n249124 , n249122 , n249123 );
nand ( n249125 , n249120 , n249124 );
nand ( n249126 , n248916 , n248711 );
not ( n249127 , n249126 );
and ( n249128 , n249125 , n249127 );
not ( n249129 , n249125 );
and ( n249130 , n249129 , n249126 );
nor ( n249131 , n249128 , n249130 );
nand ( n249132 , n247906 , n248931 );
nor ( n249133 , n249097 , n249132 );
not ( n249134 , n249133 );
not ( n249135 , n249086 );
or ( n249136 , n249134 , n249135 );
and ( n249137 , n249121 , n248931 );
not ( n249138 , n248705 );
nor ( n249139 , n249137 , n249138 );
nand ( n249140 , n249136 , n249139 );
not ( n249141 , n247908 );
nand ( n249142 , n249141 , n248707 );
not ( n249143 , n249142 );
and ( n249144 , n249140 , n249143 );
not ( n249145 , n249140 );
and ( n249146 , n249145 , n249142 );
nor ( n249147 , n249144 , n249146 );
nand ( n249148 , n247919 , n249037 );
nor ( n249149 , n247914 , n249148 );
nand ( n249150 , n247906 , n249149 );
nor ( n249151 , n249097 , n249150 );
not ( n249152 , n249151 );
not ( n249153 , n249086 );
or ( n249154 , n249152 , n249153 );
and ( n249155 , n249121 , n249149 );
not ( n249156 , n249037 );
not ( n249157 , n248725 );
or ( n249158 , n249156 , n249157 );
nand ( n249159 , n249158 , n248728 );
nor ( n249160 , n249155 , n249159 );
nand ( n249161 , n249154 , n249160 );
not ( n249162 , n247922 );
nand ( n249163 , n249162 , n248730 );
not ( n249164 , n249163 );
and ( n249165 , n249161 , n249164 );
not ( n249166 , n249161 );
and ( n249167 , n249166 , n249163 );
nor ( n249168 , n249165 , n249167 );
nand ( n249169 , n248857 , n248862 );
not ( n249170 , n249169 );
not ( n249171 , n249170 );
not ( n249172 , n249086 );
or ( n249173 , n249171 , n249172 );
and ( n249174 , n248873 , n248857 );
nor ( n249175 , n249174 , n248884 );
nand ( n249176 , n249173 , n249175 );
nor ( n249177 , n248720 , n247918 );
and ( n249178 , n249176 , n249177 );
not ( n249179 , n249176 );
not ( n249180 , n249177 );
and ( n249181 , n249179 , n249180 );
nor ( n249182 , n249178 , n249181 );
not ( n249183 , n248822 );
not ( n249184 , n249086 );
or ( n249185 , n249183 , n249184 );
nand ( n249186 , n249185 , n248843 );
nand ( n249187 , n247929 , n248740 );
not ( n249188 , n249187 );
and ( n249189 , n249186 , n249188 );
not ( n249190 , n249186 );
and ( n249191 , n249190 , n249187 );
nor ( n249192 , n249189 , n249191 );
not ( n249193 , n247979 );
not ( n249194 , n247980 );
nor ( n249195 , n249193 , n247974 , n249194 );
not ( n249196 , n249195 );
not ( n249197 , n249055 );
or ( n249198 , n249196 , n249197 );
not ( n249199 , n247978 );
buf ( n249200 , n248624 );
not ( n249201 , n249200 );
or ( n249202 , n249199 , n249201 );
nand ( n249203 , n249202 , n248628 );
not ( n249204 , n249203 );
nand ( n249205 , n249198 , n249204 );
nand ( n249206 , n247983 , n248632 );
not ( n249207 , n249206 );
and ( n249208 , n249205 , n249207 );
not ( n249209 , n249205 );
and ( n249210 , n249209 , n249206 );
nor ( n249211 , n249208 , n249210 );
nor ( n249212 , n247974 , n249194 );
not ( n249213 , n249212 );
not ( n249214 , n249055 );
or ( n249215 , n249213 , n249214 );
not ( n249216 , n249200 );
nand ( n249217 , n249215 , n249216 );
nand ( n249218 , n247979 , n248628 );
not ( n249219 , n249218 );
and ( n249220 , n249217 , n249219 );
not ( n249221 , n249217 );
and ( n249222 , n249221 , n249218 );
nor ( n249223 , n249220 , n249222 );
not ( n249224 , n247980 );
not ( n249225 , n249055 );
or ( n249226 , n249224 , n249225 );
buf ( n249227 , n248621 );
nand ( n249228 , n249226 , n249227 );
nand ( n249229 , n247975 , n248623 );
not ( n249230 , n249229 );
and ( n249231 , n249228 , n249230 );
not ( n249232 , n249228 );
and ( n249233 , n249232 , n249229 );
nor ( n249234 , n249231 , n249233 );
nand ( n249235 , n248598 , n248606 );
not ( n249236 , n249235 );
and ( n249237 , n248808 , n249236 );
not ( n249238 , n248808 );
and ( n249239 , n249238 , n249235 );
nor ( n249240 , n249237 , n249239 );
not ( n249241 , n248790 );
not ( n249242 , n248800 );
or ( n249243 , n249241 , n249242 );
nand ( n249244 , n249243 , n248803 );
nand ( n249245 , n248976 , n248600 );
not ( n249246 , n249245 );
and ( n249247 , n249244 , n249246 );
not ( n249248 , n249244 );
and ( n249249 , n249248 , n249245 );
nor ( n249250 , n249247 , n249249 );
not ( n249251 , n247965 );
not ( n249252 , n248800 );
or ( n249253 , n249251 , n249252 );
nand ( n249254 , n249253 , n248586 );
nand ( n249255 , n247968 , n248589 );
not ( n249256 , n249255 );
and ( n249257 , n249254 , n249256 );
not ( n249258 , n249254 );
and ( n249259 , n249258 , n249255 );
nor ( n249260 , n249257 , n249259 );
not ( n249261 , n247951 );
not ( n249262 , n247940 );
nor ( n249263 , n249262 , n247943 );
not ( n249264 , n249263 );
not ( n249265 , n248561 );
or ( n249266 , n249264 , n249265 );
buf ( n249267 , n248573 );
not ( n249268 , n249267 );
nand ( n249269 , n249266 , n249268 );
not ( n249270 , n249269 );
or ( n249271 , n249261 , n249270 );
buf ( n249272 , n248577 );
nand ( n249273 , n249271 , n249272 );
nand ( n249274 , n247947 , n248582 );
not ( n249275 , n249274 );
and ( n249276 , n249273 , n249275 );
not ( n249277 , n249273 );
and ( n249278 , n249277 , n249274 );
nor ( n249279 , n249276 , n249278 );
not ( n249280 , n248544 );
buf ( n249281 , n248035 );
not ( n249282 , n249281 );
not ( n249283 , n248031 );
not ( n249284 , n248506 );
or ( n249285 , n249283 , n249284 );
buf ( n249286 , n248530 );
not ( n249287 , n249286 );
nand ( n249288 , n249285 , n249287 );
not ( n249289 , n249288 );
or ( n249290 , n249282 , n249289 );
and ( n249291 , n248537 , n248538 );
nor ( n249292 , n249291 , n248541 );
not ( n249293 , n249292 );
not ( n249294 , n249293 );
nand ( n249295 , n249290 , n249294 );
not ( n249296 , n249295 );
or ( n249297 , n249280 , n249296 );
not ( n249298 , n248014 );
nand ( n249299 , n249298 , n236499 );
nand ( n249300 , n249297 , n249299 );
nand ( n249301 , n248009 , n248555 );
not ( n249302 , n249301 );
and ( n249303 , n249300 , n249302 );
not ( n249304 , n249300 );
and ( n249305 , n249304 , n249301 );
nor ( n249306 , n249303 , n249305 );
nor ( n249307 , n248765 , n249019 );
not ( n249308 , n247857 );
not ( n249309 , n247873 );
nand ( n249310 , n249308 , n249309 );
and ( n249311 , n249307 , n249310 );
nand ( n249312 , n247938 , n249311 , n247888 );
not ( n249313 , n249312 );
not ( n249314 , n249313 );
not ( n249315 , n249086 );
or ( n249316 , n249314 , n249315 );
not ( n249317 , n249311 );
not ( n249318 , n247888 );
not ( n249319 , n248757 );
or ( n249320 , n249318 , n249319 );
nand ( n249321 , n249320 , n248763 );
not ( n249322 , n249321 );
or ( n249323 , n249317 , n249322 );
or ( n249324 , n248767 , n249019 );
nand ( n249325 , n249324 , n249021 );
and ( n249326 , n249325 , n249310 );
nor ( n249327 , n249308 , n249309 );
nor ( n249328 , n249326 , n249327 );
nand ( n249329 , n249323 , n249328 );
not ( n249330 , n249329 );
nand ( n249331 , n249316 , n249330 );
nor ( n249332 , n247877 , n247883 );
and ( n249333 , n247877 , n247883 );
nor ( n249334 , n249332 , n249333 );
and ( n249335 , n249331 , n249334 );
not ( n249336 , n249331 );
not ( n249337 , n249334 );
and ( n249338 , n249336 , n249337 );
nor ( n249339 , n249335 , n249338 );
not ( n249340 , n247938 );
nand ( n249341 , n247888 , n249307 );
nor ( n249342 , n249340 , n249341 );
not ( n249343 , n249342 );
not ( n249344 , n249086 );
or ( n249345 , n249343 , n249344 );
not ( n249346 , n249341 );
and ( n249347 , n248758 , n249346 );
not ( n249348 , n249020 );
or ( n249349 , n248763 , n248765 );
nand ( n249350 , n249349 , n248767 );
not ( n249351 , n249350 );
or ( n249352 , n249348 , n249351 );
nand ( n249353 , n249352 , n249021 );
nor ( n249354 , n249347 , n249353 );
nand ( n249355 , n249345 , n249354 );
not ( n249356 , n249327 );
nand ( n249357 , n249356 , n249310 );
not ( n249358 , n249357 );
and ( n249359 , n249355 , n249358 );
not ( n249360 , n249355 );
and ( n249361 , n249360 , n249357 );
nor ( n249362 , n249359 , n249361 );
not ( n249363 , n247934 );
nor ( n249364 , n249363 , n247932 );
and ( n249365 , n247928 , n249364 );
not ( n249366 , n249365 );
not ( n249367 , n249086 );
or ( n249368 , n249366 , n249367 );
not ( n249369 , n247932 );
not ( n249370 , n249369 );
not ( n249371 , n248737 );
or ( n249372 , n249370 , n249371 );
not ( n249373 , n248743 );
nand ( n249374 , n249372 , n249373 );
and ( n249375 , n249374 , n247934 );
not ( n249376 , n248748 );
nor ( n249377 , n249375 , n249376 );
nand ( n249378 , n249368 , n249377 );
nand ( n249379 , n247933 , n248750 );
not ( n249380 , n249379 );
and ( n249381 , n249378 , n249380 );
not ( n249382 , n249378 );
and ( n249383 , n249382 , n249379 );
nor ( n249384 , n249381 , n249383 );
not ( n249385 , n248027 );
buf ( n249386 , n248021 );
not ( n249387 , n249386 );
buf ( n249388 , n248506 );
not ( n249389 , n249388 );
or ( n249390 , n249387 , n249389 );
buf ( n249391 , n248521 );
not ( n249392 , n249391 );
nand ( n249393 , n249390 , n249392 );
not ( n249394 , n249393 );
or ( n249395 , n249385 , n249394 );
buf ( n249396 , n248525 );
nand ( n249397 , n249395 , n249396 );
nand ( n249398 , n248512 , n248529 );
not ( n249399 , n249398 );
and ( n249400 , n249397 , n249399 );
not ( n249401 , n249397 );
and ( n249402 , n249401 , n249398 );
nor ( n249403 , n249400 , n249402 );
nand ( n249404 , n248544 , n249299 );
not ( n249405 , n249404 );
and ( n249406 , n249295 , n249405 );
not ( n249407 , n249295 );
and ( n249408 , n249407 , n249404 );
nor ( n249409 , n249406 , n249408 );
and ( n249410 , n248016 , n249281 );
not ( n249411 , n249410 );
buf ( n249412 , n249288 );
not ( n249413 , n249412 );
or ( n249414 , n249411 , n249413 );
and ( n249415 , n248544 , n248009 );
not ( n249416 , n249415 );
not ( n249417 , n249293 );
or ( n249418 , n249416 , n249417 );
not ( n249419 , n248556 );
nand ( n249420 , n249418 , n249419 );
and ( n249421 , n249420 , n248012 );
nor ( n249422 , n249421 , n248549 );
nand ( n249423 , n249414 , n249422 );
nand ( n249424 , n248036 , n248558 );
not ( n249425 , n249424 );
and ( n249426 , n249423 , n249425 );
not ( n249427 , n249423 );
and ( n249428 , n249427 , n249424 );
nor ( n249429 , n249426 , n249428 );
not ( n249430 , n247940 );
buf ( n249431 , n248861 );
not ( n249432 , n249431 );
or ( n249433 , n249430 , n249432 );
buf ( n249434 , n248570 );
buf ( n249435 , n249434 );
nand ( n249436 , n249433 , n249435 );
nand ( n249437 , n247944 , n248572 );
not ( n249438 , n249437 );
and ( n249439 , n249436 , n249438 );
not ( n249440 , n249436 );
and ( n249441 , n249440 , n249437 );
nor ( n249442 , n249439 , n249441 );
nand ( n249443 , n247965 , n248586 );
not ( n249444 , n249443 );
and ( n249445 , n248972 , n249444 );
not ( n249446 , n248972 );
and ( n249447 , n249446 , n249443 );
nor ( n249448 , n249445 , n249447 );
nand ( n249449 , n247980 , n249227 );
not ( n249450 , n249449 );
and ( n249451 , n249055 , n249450 );
not ( n249452 , n249055 );
and ( n249453 , n249452 , n249449 );
nor ( n249454 , n249451 , n249453 );
not ( n249455 , n248045 );
not ( n249456 , n248041 );
buf ( n249457 , n248469 );
buf ( n249458 , n248081 );
nand ( n249459 , n249457 , n249458 , n248470 );
buf ( n249460 , n249459 );
not ( n249461 , n249460 );
or ( n249462 , n249456 , n249461 );
buf ( n249463 , n248496 );
not ( n249464 , n249463 );
nand ( n249465 , n249462 , n249464 );
not ( n249466 , n249465 );
or ( n249467 , n249455 , n249466 );
nand ( n249468 , n249467 , n248499 );
nand ( n249469 , n248503 , n248046 );
not ( n249470 , n249469 );
and ( n249471 , n249468 , n249470 );
not ( n249472 , n249468 );
and ( n249473 , n249472 , n249469 );
nor ( n249474 , n249471 , n249473 );
nand ( n249475 , n247940 , n249435 );
not ( n249476 , n249475 );
and ( n249477 , n249431 , n249476 );
not ( n249478 , n249431 );
and ( n249479 , n249478 , n249475 );
nor ( n249480 , n249477 , n249479 );
not ( n249481 , n248034 );
nand ( n249482 , n249481 , n248534 );
not ( n249483 , n249482 );
and ( n249484 , n249412 , n249483 );
not ( n249485 , n249412 );
and ( n249486 , n249485 , n249482 );
nor ( n249487 , n249484 , n249486 );
or ( n249488 , n248474 , n232224 );
not ( n249489 , n249488 );
buf ( n249490 , n248047 );
not ( n249491 , n249490 );
not ( n249492 , n249491 );
not ( n249493 , n249460 );
or ( n249494 , n249492 , n249493 );
and ( n249495 , n248501 , n248503 );
nand ( n249496 , n249494 , n249495 );
not ( n249497 , n249496 );
or ( n249498 , n249489 , n249497 );
nand ( n249499 , n249498 , n248502 );
or ( n249500 , n248482 , n248479 );
not ( n249501 , n249500 );
and ( n249502 , n249499 , n249501 );
not ( n249503 , n249499 );
and ( n249504 , n249503 , n249500 );
nor ( n249505 , n249502 , n249504 );
not ( n249506 , n248020 );
not ( n249507 , n249506 );
not ( n249508 , n249388 );
or ( n249509 , n249507 , n249508 );
buf ( n249510 , n248518 );
nand ( n249511 , n249509 , n249510 );
not ( n249512 , n248019 );
nand ( n249513 , n249512 , n248520 );
not ( n249514 , n249513 );
and ( n249515 , n249511 , n249514 );
not ( n249516 , n249511 );
and ( n249517 , n249516 , n249513 );
nor ( n249518 , n249515 , n249517 );
nand ( n249519 , n249506 , n249510 );
not ( n249520 , n249519 );
and ( n249521 , n249388 , n249520 );
not ( n249522 , n249388 );
and ( n249523 , n249522 , n249519 );
nor ( n249524 , n249521 , n249523 );
nand ( n249525 , n249488 , n248502 );
not ( n249526 , n249525 );
and ( n249527 , n249496 , n249526 );
not ( n249528 , n249496 );
and ( n249529 , n249528 , n249525 );
nor ( n249530 , n249527 , n249529 );
nand ( n249531 , n248045 , n248499 );
not ( n249532 , n249531 );
and ( n249533 , n249465 , n249532 );
not ( n249534 , n249465 );
and ( n249535 , n249534 , n249531 );
nor ( n249536 , n249533 , n249535 );
not ( n249537 , n248039 );
not ( n249538 , n249537 );
not ( n249539 , n249460 );
or ( n249540 , n249538 , n249539 );
buf ( n249541 , n248493 );
nand ( n249542 , n249540 , n249541 );
not ( n249543 , n248040 );
nand ( n249544 , n249543 , n248495 );
not ( n249545 , n249544 );
and ( n249546 , n249542 , n249545 );
not ( n249547 , n249542 );
and ( n249548 , n249547 , n249544 );
nor ( n249549 , n249546 , n249548 );
not ( n249550 , n248053 );
buf ( n249551 , n248074 );
buf ( n249552 , n249551 );
not ( n249553 , n249552 );
not ( n249554 , n248465 );
buf ( n249555 , n248455 );
nand ( n249556 , n249554 , n249555 );
nand ( n249557 , n249553 , n249556 );
not ( n249558 , n249557 );
or ( n249559 , n249550 , n249558 );
nand ( n249560 , n249559 , n248077 );
nand ( n249561 , n248080 , n248470 );
not ( n249562 , n249561 );
and ( n249563 , n249560 , n249562 );
not ( n249564 , n249560 );
and ( n249565 , n249564 , n249561 );
nor ( n249566 , n249563 , n249565 );
not ( n249567 , n248464 );
not ( n249568 , n248462 );
not ( n249569 , n249555 );
or ( n249570 , n249568 , n249569 );
buf ( n249571 , n248066 );
not ( n249572 , n249571 );
nand ( n249573 , n249570 , n249572 );
not ( n249574 , n249573 );
or ( n249575 , n249567 , n249574 );
nand ( n249576 , n249575 , n248069 );
not ( n249577 , n248456 );
nand ( n249578 , n249577 , n248073 );
not ( n249579 , n249578 );
and ( n249580 , n249576 , n249579 );
not ( n249581 , n249576 );
and ( n249582 , n249581 , n249578 );
nor ( n249583 , n249580 , n249582 );
nand ( n249584 , n248053 , n248077 );
not ( n249585 , n249584 );
and ( n249586 , n249557 , n249585 );
not ( n249587 , n249557 );
and ( n249588 , n249587 , n249584 );
nor ( n249589 , n249586 , n249588 );
not ( n249590 , n248460 );
not ( n249591 , n249590 );
not ( n249592 , n249555 );
or ( n249593 , n249591 , n249592 );
buf ( n249594 , n248063 );
nand ( n249595 , n249593 , n249594 );
not ( n249596 , n248461 );
buf ( n249597 , n248065 );
nand ( n249598 , n249596 , n249597 );
not ( n249599 , n249598 );
and ( n249600 , n249595 , n249599 );
not ( n249601 , n249595 );
and ( n249602 , n249601 , n249598 );
nor ( n249603 , n249600 , n249602 );
buf ( n249604 , n248427 );
not ( n249605 , n248086 );
and ( n249606 , n249604 , n249605 );
nor ( n249607 , n249606 , n248449 );
not ( n249608 , n248088 );
or ( n249609 , n249607 , n249608 );
nand ( n249610 , n249609 , n248452 );
not ( n249611 , n248434 );
buf ( n249612 , n248430 );
nand ( n249613 , n249611 , n249612 );
not ( n249614 , n249613 );
and ( n249615 , n249610 , n249614 );
not ( n249616 , n249610 );
and ( n249617 , n249616 , n249613 );
nor ( n249618 , n249615 , n249617 );
not ( n249619 , n248082 );
nand ( n249620 , n249619 , n249604 );
not ( n249621 , n248084 );
or ( n249622 , n249620 , n249621 );
not ( n249623 , n248445 );
nand ( n249624 , n249622 , n249623 );
nand ( n249625 , n248085 , n248448 );
not ( n249626 , n249625 );
and ( n249627 , n249624 , n249626 );
not ( n249628 , n249624 );
and ( n249629 , n249628 , n249625 );
nor ( n249630 , n249627 , n249629 );
not ( n249631 , n249607 );
nand ( n249632 , n248452 , n248450 );
not ( n249633 , n249632 );
and ( n249634 , n249631 , n249633 );
not ( n249635 , n249631 );
and ( n249636 , n249635 , n249632 );
nor ( n249637 , n249634 , n249636 );
buf ( n249638 , n248442 );
nand ( n249639 , n249638 , n249620 );
nand ( n249640 , n248084 , n248444 );
not ( n249641 , n249640 );
and ( n249642 , n249639 , n249641 );
not ( n249643 , n249639 );
and ( n249644 , n249643 , n249640 );
nor ( n249645 , n249642 , n249644 );
buf ( n249646 , n248409 );
not ( n249647 , n249646 );
not ( n249648 , n248094 );
or ( n249649 , n249647 , n249648 );
buf ( n249650 , n248420 );
not ( n249651 , n249650 );
nand ( n249652 , n249649 , n249651 );
buf ( n249653 , n248412 );
nand ( n249654 , n248098 , n249653 );
not ( n249655 , n249654 );
and ( n249656 , n249652 , n249655 );
not ( n249657 , n249652 );
and ( n249658 , n249657 , n249654 );
nor ( n249659 , n249656 , n249658 );
buf ( n249660 , n248093 );
not ( n249661 , n249660 );
not ( n249662 , n249661 );
not ( n249663 , n249646 );
or ( n249664 , n249662 , n249663 );
buf ( n249665 , n248417 );
nand ( n249666 , n249664 , n249665 );
not ( n249667 , n248092 );
nand ( n249668 , n249667 , n248419 );
not ( n249669 , n249668 );
and ( n249670 , n249666 , n249669 );
not ( n249671 , n249666 );
and ( n249672 , n249671 , n249668 );
nor ( n249673 , n249670 , n249672 );
buf ( n249674 , n248384 );
not ( n249675 , n248108 );
nand ( n249676 , n249674 , n249675 );
or ( n249677 , n249676 , n248107 );
not ( n249678 , n248391 );
nand ( n249679 , n249677 , n249678 );
not ( n249680 , n248394 );
nand ( n249681 , n249680 , n248392 );
not ( n249682 , n249681 );
and ( n249683 , n249679 , n249682 );
not ( n249684 , n249679 );
and ( n249685 , n249684 , n249681 );
nor ( n249686 , n249683 , n249685 );
not ( n249687 , n248103 );
not ( n249688 , n249687 );
buf ( n249689 , n248396 );
buf ( n249690 , n249689 );
not ( n249691 , n249690 );
or ( n249692 , n249688 , n249691 );
nand ( n249693 , n249692 , n248400 );
not ( n249694 , n248356 );
not ( n249695 , n249694 );
not ( n249696 , n248122 );
not ( n249697 , n248340 );
or ( n249698 , n249696 , n249697 );
nand ( n249699 , n249698 , n248352 );
buf ( n249700 , n249699 );
not ( n249701 , n249700 );
or ( n249702 , n249695 , n249701 );
nand ( n249703 , n249702 , n248365 );
buf ( n249704 , n248340 );
not ( n249705 , n248121 );
nand ( n249706 , n249704 , n249705 );
nand ( n249707 , n248343 , n249706 );
not ( n249708 , n248125 );
not ( n249709 , n249708 );
not ( n249710 , n248330 );
or ( n249711 , n249709 , n249710 );
nand ( n249712 , n249711 , n248334 );
buf ( n249713 , n248298 );
nand ( n249714 , n249713 , n248301 );
nand ( n249715 , n249594 , n249590 );
not ( n249716 , n249715 );
nand ( n249717 , n248027 , n249396 );
nand ( n249718 , n249619 , n249638 );
not ( n249719 , n248143 );
not ( n249720 , n249719 );
not ( n249721 , n248281 );
or ( n249722 , n249720 , n249721 );
not ( n249723 , n248285 );
nand ( n249724 , n249722 , n249723 );
not ( n249725 , n247987 );
not ( n249726 , n248644 );
not ( n249727 , n249726 );
or ( n249728 , n249725 , n249727 );
nand ( n249729 , n249728 , n248948 );
and ( n249730 , n249729 , n248648 );
not ( n249731 , n248657 );
nor ( n249732 , n249730 , n249731 );
nor ( n249733 , n248101 , n248103 );
not ( n249734 , n248533 );
buf ( n249735 , n248536 );
nand ( n249736 , n249734 , n249735 );
nand ( n249737 , n249661 , n249665 );
nand ( n249738 , n249687 , n248400 );
nand ( n249739 , n249675 , n248388 );
not ( n249740 , n248368 );
not ( n249741 , n248148 );
nand ( n249742 , n249741 , n248276 );
not ( n249743 , n249742 );
buf ( n249744 , n248273 );
not ( n249745 , n249744 );
or ( n249746 , n249743 , n249745 );
or ( n249747 , n249744 , n249742 );
nand ( n249748 , n249746 , n249747 );
nand ( n249749 , n249694 , n248365 );
not ( n249750 , n248120 );
nand ( n249751 , n249750 , n248348 );
nand ( n249752 , n247997 , n248637 );
not ( n249753 , n249752 );
nor ( n249754 , n249312 , n249332 );
nand ( n249755 , n248333 , n248337 );
nand ( n249756 , n248956 , n248651 );
buf ( n249757 , n248259 );
not ( n249758 , n248155 );
and ( n249759 , n249757 , n249758 );
not ( n249760 , n248262 );
nor ( n249761 , n249759 , n249760 );
not ( n249762 , n249761 );
and ( n249763 , n248267 , n248264 );
not ( n249764 , n249763 );
or ( n249765 , n249762 , n249764 );
or ( n249766 , n249763 , n249761 );
nand ( n249767 , n249765 , n249766 );
not ( n249768 , n248884 );
nand ( n249769 , n249708 , n248334 );
not ( n249770 , n248662 );
nand ( n249771 , n249770 , n248659 );
not ( n249772 , n249771 );
nand ( n249773 , n249758 , n248262 );
not ( n249774 , n249773 );
not ( n249775 , n249757 );
or ( n249776 , n249774 , n249775 );
or ( n249777 , n249757 , n249773 );
nand ( n249778 , n249776 , n249777 );
not ( n249779 , n248129 );
nand ( n249780 , n249779 , n248325 );
not ( n249781 , n248133 );
nand ( n249782 , n249781 , n248315 );
nand ( n249783 , n248314 , n248318 );
nand ( n249784 , n248303 , n248310 );
not ( n249785 , n248255 );
not ( n249786 , n249785 );
and ( n249787 , n248158 , n248258 );
not ( n249788 , n249787 );
or ( n249789 , n249786 , n249788 );
or ( n249790 , n249785 , n249787 );
nand ( n249791 , n249789 , n249790 );
not ( n249792 , n248674 );
nor ( n249793 , n249792 , n247890 );
not ( n249794 , n248300 );
nand ( n249795 , n249794 , n248306 );
not ( n249796 , n248293 );
nor ( n249797 , n249796 , n248296 );
nand ( n249798 , n247896 , n248680 );
nand ( n249799 , n249719 , n249723 );
nand ( n249800 , n248284 , n248287 );
nand ( n249801 , n248146 , n248280 );
and ( n249802 , n248743 , n247934 );
nor ( n249803 , n249802 , n249376 );
or ( n249804 , n249803 , n248747 );
nand ( n249805 , n249804 , n248750 );
not ( n249806 , n248247 );
not ( n249807 , n249806 );
and ( n249808 , n248162 , n248250 );
not ( n249809 , n249808 );
or ( n249810 , n249807 , n249809 );
or ( n249811 , n249806 , n249808 );
nand ( n249812 , n249810 , n249811 );
nand ( n249813 , n249364 , n247933 );
not ( n249814 , n249813 );
nand ( n249815 , n249037 , n248728 );
not ( n249816 , n249815 );
nand ( n249817 , n248164 , n248246 );
not ( n249818 , n249817 );
not ( n249819 , n248243 );
or ( n249820 , n249818 , n249819 );
or ( n249821 , n248243 , n249817 );
nand ( n249822 , n249820 , n249821 );
not ( n249823 , n248237 );
not ( n249824 , n249823 );
and ( n249825 , n248239 , n248242 );
not ( n249826 , n249825 );
or ( n249827 , n249824 , n249826 );
or ( n249828 , n249825 , n249823 );
nand ( n249829 , n249827 , n249828 );
nand ( n249830 , n248160 , n248254 );
not ( n249831 , n248166 );
nand ( n249832 , n249831 , n248236 );
not ( n249833 , n249832 );
not ( n249834 , n248234 );
not ( n249835 , n249834 );
or ( n249836 , n249833 , n249835 );
or ( n249837 , n249834 , n249832 );
nand ( n249838 , n249836 , n249837 );
nand ( n249839 , n247888 , n248763 );
not ( n249840 , n248231 );
not ( n249841 , n249840 );
not ( n249842 , n248167 );
nor ( n249843 , n249842 , n248233 );
not ( n249844 , n249843 );
or ( n249845 , n249841 , n249844 );
or ( n249846 , n249840 , n249843 );
nand ( n249847 , n249845 , n249846 );
nand ( n249848 , n248227 , n248230 );
not ( n249849 , n249848 );
not ( n249850 , n248225 );
or ( n249851 , n249849 , n249850 );
or ( n249852 , n248225 , n249848 );
nand ( n249853 , n249851 , n249852 );
xor ( n249854 , n213180 , n213239 );
xor ( n249855 , n249854 , n248222 );
xor ( n249856 , n213103 , n248218 );
xor ( n249857 , n249856 , n213176 );
not ( n249858 , n249332 );
not ( n249859 , n248205 );
nand ( n249860 , n248212 , n248217 );
not ( n249861 , n249860 );
or ( n249862 , n249859 , n249861 );
or ( n249863 , n248205 , n249860 );
nand ( n249864 , n249862 , n249863 );
xor ( n249865 , n248169 , n248182 );
xor ( n249866 , n249865 , n248202 );
xor ( n249867 , n248184 , n248196 );
xor ( n249868 , n249867 , n248200 );
and ( n249869 , n248192 , n248195 );
nor ( n249870 , n249869 , n248196 );
not ( n249871 , n247881 );
not ( n249872 , n247879 );
buf ( n249873 , n248098 );
not ( n249874 , n249873 );
not ( n249875 , n249652 );
or ( n249876 , n249874 , n249875 );
nand ( n249877 , n249876 , n249653 );
not ( n249878 , n248425 );
nor ( n249879 , n249878 , n248414 );
xor ( n249880 , n249877 , n249879 );
not ( n249881 , n248101 );
nand ( n249882 , n249881 , n248402 );
xnor ( n249883 , n249693 , n249882 );
xnor ( n249884 , n249690 , n249738 );
nand ( n249885 , n247951 , n248577 );
xnor ( n249886 , n249269 , n249885 );
xnor ( n249887 , n249674 , n249739 );
xnor ( n249888 , n248277 , n249801 );
not ( n249889 , n248355 );
nand ( n249890 , n249889 , n248367 );
xnor ( n249891 , n249703 , n249890 );
xnor ( n249892 , n249700 , n249749 );
xnor ( n249893 , n249707 , n249751 );
nand ( n249894 , n249705 , n248343 );
xnor ( n249895 , n249704 , n249894 );
xnor ( n249896 , n249712 , n249755 );
xnor ( n249897 , n248330 , n249769 );
not ( n249898 , n249779 );
not ( n249899 , n248321 );
or ( n249900 , n249898 , n249899 );
nand ( n249901 , n249900 , n248325 );
nor ( n249902 , n248328 , n248128 );
xor ( n249903 , n249901 , n249902 );
not ( n249904 , n249781 );
buf ( n249905 , n248311 );
not ( n249906 , n249905 );
or ( n249907 , n249904 , n249906 );
nand ( n249908 , n249907 , n248315 );
xnor ( n249909 , n249908 , n249783 );
not ( n249910 , n248308 );
nand ( n249911 , n249910 , n249714 );
xnor ( n249912 , n249911 , n249784 );
xnor ( n249913 , n249713 , n249795 );
not ( n249914 , n248139 );
not ( n249915 , n249914 );
not ( n249916 , n248290 );
or ( n249917 , n249915 , n249916 );
not ( n249918 , n248294 );
nand ( n249919 , n249917 , n249918 );
xor ( n249920 , n249919 , n249797 );
xnor ( n249921 , n248779 , n249798 );
nand ( n249922 , n249918 , n249914 );
xnor ( n249923 , n248290 , n249922 );
xnor ( n249924 , n248281 , n249799 );
xnor ( n249925 , n249724 , n249800 );
not ( n249926 , n247666 );
nor ( n249927 , n249926 , n209973 );
and ( n249928 , n239270 , n247666 );
nor ( n249929 , n249928 , n249872 );
xor ( n249930 , n249929 , n249927 );
xor ( n249931 , n249930 , n249871 );
xor ( n249932 , n210193 , n210359 );
and ( n249933 , n210224 , n210226 , n210221 );
nor ( n249934 , n249933 , n209441 );
not ( n249935 , n249934 );
xor ( n249936 , n249935 , n210374 );
xnor ( n249937 , n248945 , n249756 );
xor ( n249938 , n249086 , n249793 );
not ( n249939 , n249481 );
not ( n249940 , n249288 );
or ( n249941 , n249939 , n249940 );
nand ( n249942 , n249941 , n248534 );
xnor ( n249943 , n249942 , n249736 );
xnor ( n249944 , n249393 , n249717 );
xnor ( n249945 , n248251 , n249830 );
not ( n249946 , n248664 );
not ( n249947 , n249311 );
not ( n249948 , n249321 );
or ( n249949 , n249947 , n249948 );
nand ( n249950 , n249949 , n249328 );
and ( n249951 , n249950 , n249858 );
nor ( n249952 , n249951 , n249333 );
nor ( n249953 , n248377 , n248382 );
not ( n249954 , n247919 );
nor ( n249955 , n249954 , n249169 );
and ( n249956 , n249955 , n248820 );
not ( n249957 , n249956 );
not ( n249958 , n249055 );
or ( n249959 , n249957 , n249958 );
nor ( n249960 , n248857 , n249036 );
nand ( n249961 , n249768 , n249960 );
not ( n249962 , n249036 );
nand ( n249963 , n249962 , n249768 , n248872 , n248874 );
or ( n249964 , n249036 , n247919 );
nand ( n249965 , n249961 , n249963 , n249964 );
nand ( n249966 , n249959 , n249965 );
and ( n249967 , n249966 , n249816 );
not ( n249968 , n249966 );
and ( n249969 , n249968 , n249815 );
nor ( n249970 , n249967 , n249969 );
not ( n249971 , n249754 );
not ( n249972 , n249086 );
or ( n249973 , n249971 , n249972 );
nand ( n249974 , n249973 , n249952 );
not ( n249975 , n247887 );
not ( n249976 , n249931 );
or ( n249977 , n249975 , n249976 );
or ( n249978 , n249931 , n247887 );
nand ( n249979 , n249977 , n249978 );
not ( n249980 , n249979 );
and ( n249981 , n249974 , n249980 );
not ( n249982 , n249974 );
and ( n249983 , n249982 , n249979 );
nor ( n249984 , n249981 , n249983 );
not ( n249985 , n248759 );
nor ( n249986 , n249985 , n249839 );
not ( n249987 , n249986 );
not ( n249988 , n249946 );
nand ( n249989 , n248820 , n248837 );
not ( n249990 , n249989 );
or ( n249991 , n249988 , n249990 );
nand ( n249992 , n249991 , n247938 );
not ( n249993 , n249992 );
or ( n249994 , n249987 , n249993 );
and ( n249995 , n248759 , n249946 );
not ( n249996 , n249995 );
not ( n249997 , n249989 );
or ( n249998 , n249996 , n249997 );
not ( n249999 , n247938 );
and ( n250000 , n249999 , n248759 );
not ( n250001 , n249839 );
nor ( n250002 , n250000 , n250001 );
nand ( n250003 , n249998 , n250002 );
nand ( n250004 , n249994 , n250003 );
not ( n250005 , n249051 );
not ( n250006 , n248837 );
or ( n250007 , n250005 , n250006 );
buf ( n250008 , n248633 );
not ( n250009 , n250008 );
nand ( n250010 , n250007 , n250009 );
and ( n250011 , n250010 , n249753 );
not ( n250012 , n250010 );
and ( n250013 , n250012 , n249752 );
nor ( n250014 , n250011 , n250013 );
not ( n250015 , n249782 );
not ( n250016 , n249905 );
or ( n250017 , n250015 , n250016 );
or ( n250018 , n249782 , n249905 );
nand ( n250019 , n250017 , n250018 );
or ( n250020 , n248120 , n248343 );
nand ( n250021 , n250020 , n248348 );
and ( n250022 , n249690 , n249733 );
or ( n250023 , n248400 , n248399 );
nand ( n250024 , n250023 , n248402 );
nor ( n250025 , n250022 , n250024 );
and ( n250026 , n249555 , n249716 );
not ( n250027 , n249555 );
and ( n250028 , n250027 , n249715 );
nor ( n250029 , n250026 , n250028 );
not ( n250030 , n249718 );
not ( n250031 , n249604 );
or ( n250032 , n250030 , n250031 );
or ( n250033 , n249718 , n249604 );
nand ( n250034 , n250032 , n250033 );
not ( n250035 , n249737 );
not ( n250036 , n249646 );
or ( n250037 , n250035 , n250036 );
or ( n250038 , n249737 , n249646 );
nand ( n250039 , n250037 , n250038 );
not ( n250040 , n249369 );
not ( n250041 , n248846 );
or ( n250042 , n250040 , n250041 );
buf ( n250043 , n249373 );
nand ( n250044 , n250042 , n250043 );
nand ( n250045 , n247934 , n248748 );
not ( n250046 , n250045 );
and ( n250047 , n250044 , n250046 );
not ( n250048 , n250044 );
and ( n250049 , n250048 , n250045 );
nor ( n250050 , n250047 , n250049 );
nand ( n250051 , n218613 , n218940 );
nand ( n250052 , n248114 , n248115 );
buf ( n250053 , n248379 );
not ( n250054 , n248362 );
not ( n250055 , n248353 );
or ( n250056 , n250054 , n250055 );
buf ( n250057 , n248373 );
nand ( n250058 , n250056 , n250057 );
nand ( n250059 , n250052 , n250058 );
nand ( n250060 , n250053 , n250059 );
xor ( n250061 , n250060 , n249953 );
and ( n250062 , n248844 , n249814 );
nor ( n250063 , n250062 , n249805 );
not ( n250064 , n249813 );
nand ( n250065 , n250064 , n248837 , n248824 );
nand ( n250066 , n248464 , n248069 );
not ( n250067 , n250066 );
not ( n250068 , n249573 );
or ( n250069 , n250067 , n250068 );
or ( n250070 , n250066 , n249573 );
nand ( n250071 , n250069 , n250070 );
nand ( n250072 , n209591 , n209770 );
and ( n250073 , n250072 , n209712 );
not ( n250074 , n250072 );
and ( n250075 , n250074 , n209711 );
nor ( n250076 , n250073 , n250075 );
nand ( n250077 , n250065 , n250063 );
nand ( n250078 , n247935 , n248754 );
not ( n250079 , n250078 );
and ( n250080 , n250077 , n250079 );
not ( n250081 , n250077 );
and ( n250082 , n250081 , n250078 );
nor ( n250083 , n250080 , n250082 );
nand ( n250084 , n249537 , n249541 );
not ( n250085 , n250084 );
and ( n250086 , n249460 , n250085 );
not ( n250087 , n249460 );
and ( n250088 , n250087 , n250084 );
nor ( n250089 , n250086 , n250088 );
nand ( n250090 , n249704 , n249705 , n249750 );
not ( n250091 , n212462 );
not ( n250092 , n211459 );
or ( n250093 , n250091 , n250092 );
nand ( n250094 , n250093 , n211507 );
not ( n250095 , n250094 );
nand ( n250096 , n211428 , n211517 );
not ( n250097 , n250096 );
or ( n250098 , n250095 , n250097 );
or ( n250099 , n250096 , n250094 );
nand ( n250100 , n250098 , n250099 );
not ( n250101 , n248151 );
nand ( n250102 , n250101 , n248272 );
not ( n250103 , n250102 );
buf ( n250104 , n248269 );
not ( n250105 , n250104 );
or ( n250106 , n250103 , n250105 );
or ( n250107 , n250104 , n250102 );
nand ( n250108 , n250106 , n250107 );
not ( n250109 , n250025 );
and ( n250110 , n248404 , n248406 );
not ( n250111 , n250110 );
or ( n250112 , n250109 , n250111 );
or ( n250113 , n250110 , n250025 );
nand ( n250114 , n250112 , n250113 );
nand ( n250115 , n210999 , n210995 );
not ( n250116 , n250115 );
not ( n250117 , n212199 );
or ( n250118 , n250116 , n250117 );
or ( n250119 , n250115 , n212199 );
nand ( n250120 , n250118 , n250119 );
not ( n250121 , n248372 );
buf ( n250122 , n248370 );
nand ( n250123 , n250121 , n250122 );
not ( n250124 , n250123 );
not ( n250125 , n249700 );
not ( n250126 , n248357 );
or ( n250127 , n250125 , n250126 );
nand ( n250128 , n250127 , n249740 );
not ( n250129 , n250128 );
or ( n250130 , n250124 , n250129 );
or ( n250131 , n250123 , n250128 );
nand ( n250132 , n250130 , n250131 );
buf ( n250133 , n248351 );
nand ( n250134 , n250133 , n250051 );
not ( n250135 , n250134 );
not ( n250136 , n250021 );
nand ( n250137 , n250136 , n250090 );
not ( n250138 , n250137 );
or ( n250139 , n250135 , n250138 );
or ( n250140 , n250134 , n250137 );
nand ( n250141 , n250139 , n250140 );
nand ( n250142 , n40316 , n209518 );
not ( n250143 , n250142 );
nand ( n250144 , n209513 , n210062 );
not ( n250145 , n250144 );
or ( n250146 , n250143 , n250145 );
or ( n250147 , n250142 , n250144 );
nand ( n250148 , n250146 , n250147 );
nand ( n250149 , n250053 , n250052 );
not ( n250150 , n250149 );
and ( n250151 , n250058 , n250150 );
not ( n250152 , n250058 );
and ( n250153 , n250152 , n250149 );
nor ( n250154 , n250151 , n250153 );
not ( n250155 , n212048 );
nand ( n250156 , n250155 , n212070 );
not ( n250157 , n250156 );
nand ( n250158 , n212044 , n212065 );
not ( n250159 , n250158 );
or ( n250160 , n250157 , n250159 );
or ( n250161 , n250156 , n250158 );
nand ( n250162 , n250160 , n250161 );
nand ( n250163 , n211812 , n211890 );
not ( n250164 , n250163 );
not ( n250165 , n211820 );
not ( n250166 , n212381 );
or ( n250167 , n250165 , n250166 );
nand ( n250168 , n250167 , n212784 );
not ( n250169 , n250168 );
or ( n250170 , n250164 , n250169 );
or ( n250171 , n250163 , n250168 );
nand ( n250172 , n250170 , n250171 );
not ( n250173 , n248107 );
nand ( n250174 , n250173 , n248390 );
not ( n250175 , n250174 );
nand ( n250176 , n248388 , n249676 );
not ( n250177 , n250176 );
or ( n250178 , n250175 , n250177 );
or ( n250179 , n250174 , n250176 );
nand ( n250180 , n250178 , n250179 );
not ( n250181 , n41568 );
nand ( n250182 , n250181 , n209448 );
not ( n250183 , n250182 );
not ( n250184 , n209442 );
not ( n250185 , n249935 );
or ( n250186 , n250184 , n250185 );
nand ( n250187 , n250186 , n209444 );
not ( n250188 , n250187 );
or ( n250189 , n250183 , n250188 );
or ( n250190 , n250182 , n250187 );
nand ( n250191 , n250189 , n250190 );
not ( n250192 , n211689 );
nand ( n250193 , n250192 , n211720 );
not ( n250194 , n250193 );
nand ( n250195 , n212351 , n211714 );
not ( n250196 , n250195 );
or ( n250197 , n250194 , n250196 );
or ( n250198 , n250193 , n250195 );
nand ( n250199 , n250197 , n250198 );
nand ( n250200 , n210226 , n209438 );
not ( n250201 , n250200 );
not ( n250202 , n210224 );
or ( n250203 , n250201 , n250202 );
or ( n250204 , n250200 , n210224 );
nand ( n250205 , n250203 , n250204 );
or ( n250206 , n210877 , n212032 );
not ( n250207 , n250206 );
not ( n250208 , n211998 );
not ( n250209 , n212256 );
or ( n250210 , n250208 , n250209 );
nand ( n250211 , n250210 , n212021 );
not ( n250212 , n250211 );
or ( n250213 , n250207 , n250212 );
or ( n250214 , n250206 , n250211 );
nand ( n250215 , n250213 , n250214 );
not ( n250216 , n210780 );
not ( n250217 , n212088 );
or ( n250218 , n250216 , n250217 );
nand ( n250219 , n250218 , n212095 );
nor ( n250220 , n210786 , n212104 );
and ( n250221 , n250219 , n250220 );
not ( n250222 , n250219 );
not ( n250223 , n250220 );
and ( n250224 , n250222 , n250223 );
nor ( n250225 , n250221 , n250224 );
not ( n250226 , n248299 );
nand ( n250227 , n250226 , n248305 );
not ( n250228 , n250227 );
not ( n250229 , n249794 );
not ( n250230 , n249713 );
or ( n250231 , n250229 , n250230 );
nand ( n250232 , n250231 , n248306 );
not ( n250233 , n250232 );
or ( n250234 , n250228 , n250233 );
or ( n250235 , n250227 , n250232 );
nand ( n250236 , n250234 , n250235 );
not ( n250237 , n209383 );
nand ( n250238 , n209363 , n209386 );
not ( n250239 , n250238 );
or ( n250240 , n250237 , n250239 );
or ( n250241 , n209383 , n250238 );
nand ( n250242 , n250240 , n250241 );
not ( n250243 , n249734 );
not ( n250244 , n249942 );
or ( n250245 , n250243 , n250244 );
nand ( n250246 , n250245 , n249735 );
nand ( n250247 , n248538 , n248540 );
not ( n250248 , n250247 );
and ( n250249 , n250246 , n250248 );
not ( n250250 , n250246 );
and ( n250251 , n250250 , n250247 );
nor ( n250252 , n250249 , n250251 );
buf ( n250253 , n212897 );
buf ( n250254 , n212119 );
xor ( n250255 , n250253 , n250254 );
buf ( n250256 , n250255 );
not ( n250257 , n249415 );
not ( n250258 , n249295 );
or ( n250259 , n250257 , n250258 );
nand ( n250260 , n250259 , n249419 );
nand ( n250261 , n248548 , n248012 );
not ( n250262 , n250261 );
and ( n250263 , n250260 , n250262 );
not ( n250264 , n250260 );
and ( n250265 , n250264 , n250261 );
nor ( n250266 , n250263 , n250265 );
nand ( n250267 , n248895 , n248689 );
not ( n250268 , n250267 );
and ( n250269 , n248877 , n250268 );
not ( n250270 , n248877 );
and ( n250271 , n250270 , n250267 );
nor ( n250272 , n250269 , n250271 );
xor ( n250273 , n199344 , n213750 );
not ( n250274 , n210158 );
and ( n250275 , n209479 , n209482 );
not ( n250276 , n250275 );
or ( n250277 , n250274 , n250276 );
or ( n250278 , n250275 , n210158 );
nand ( n250279 , n250277 , n250278 );
xnor ( n250280 , n248321 , n249780 );
buf ( n250281 , n209348 );
buf ( n250282 , n211314 );
xor ( n250283 , n250281 , n250282 );
buf ( n250284 , n250283 );
xnor ( n250285 , n212165 , n212763 );
and ( n250286 , n248616 , n247987 , n248648 );
not ( n250287 , n249771 );
nand ( n250288 , n250287 , n249732 );
or ( n250289 , n250288 , n250010 );
not ( n250290 , n250286 );
nor ( n250291 , n250290 , n249772 );
nand ( n250292 , n250291 , n250010 );
not ( n250293 , n249732 );
not ( n250294 , n249772 );
and ( n250295 , n250293 , n250294 );
nor ( n250296 , n250286 , n249771 );
and ( n250297 , n249732 , n250296 );
nor ( n250298 , n250295 , n250297 );
nand ( n250299 , n250289 , n250292 , n250298 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
