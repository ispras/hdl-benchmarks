module logical_not_1_3(a, b);
  input a;
  output [2:0] b;
  assign b = !a;
endmodule
