module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n108233 , n681 , n682 , n683 , 
 n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , 
 n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , 
 n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , 
 n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , 
 n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , 
 n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , 
 n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , 
 n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , 
 n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , 
 n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , 
 n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , 
 n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , 
 n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , 
 n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , 
 n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , 
 n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , 
 n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , 
 n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , 
 n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , 
 n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , 
 n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , 
 n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , 
 n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , 
 n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , 
 n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , 
 n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , 
 n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , 
 n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , 
 n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , 
 n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , 
 n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , 
 n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , 
 n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , 
 n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , 
 n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , 
 n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , 
 n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , 
 n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , 
 n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , 
 n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , 
 n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , 
 n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , 
 n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , 
 n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , 
 n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , 
 n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , 
 n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , 
 n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , 
 n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , 
 n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , 
 n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , 
 n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , 
 n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , 
 n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , 
 n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , 
 n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , 
 n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , 
 n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , 
 n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , 
 n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , 
 n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , 
 n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , 
 n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , 
 n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , 
 n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , 
 n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , 
 n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , 
 n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , 
 n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , 
 n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , 
 n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , 
 n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , 
 n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , 
 n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , 
 n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , 
 n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , 
 n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , 
 n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , 
 n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , 
 n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , 
 n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , 
 n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , 
 n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , 
 n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , 
 n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , 
 n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , 
 n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , 
 n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , 
 n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , 
 n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , 
 n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , 
 n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , 
 n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , 
 n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , 
 n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , 
 n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , 
 n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , 
 n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , 
 n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , 
 n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , 
 n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , 
 n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , 
 n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , 
 n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , 
 n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , 
 n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , 
 n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , 
 n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , 
 n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , 
 n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , 
 n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , 
 n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , 
 n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , 
 n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , 
 n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , 
 n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , 
 n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , 
 n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , 
 n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , 
 n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , 
 n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , 
 n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , 
 n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , 
 n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , 
 n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , 
 n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , 
 n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , 
 n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , 
 n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , 
 n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , 
 n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , 
 n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , 
 n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , 
 n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , 
 n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , 
 n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , 
 n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , 
 n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , 
 n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , 
 n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , 
 n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , 
 n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , 
 n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , 
 n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , 
 n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , 
 n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , 
 n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , 
 n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , 
 n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , 
 n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , 
 n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , 
 n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , 
 n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , 
 n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , 
 n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , 
 n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , 
 n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , 
 n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , 
 n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , 
 n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , 
 n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , 
 n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , 
 n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , 
 n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , 
 n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , 
 n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , 
 n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , 
 n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , 
 n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , 
 n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , 
 n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , 
 n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , 
 n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , 
 n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , 
 n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , 
 n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , 
 n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , 
 n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , 
 n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , 
 n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , 
 n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , 
 n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , 
 n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , 
 n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , 
 n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , 
 n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , 
 n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , 
 n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , 
 n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , 
 n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , 
 n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , 
 n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , 
 n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , 
 n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , 
 n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , 
 n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , 
 n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , 
 n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , 
 n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , 
 n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , 
 n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , 
 n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , 
 n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , 
 n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , 
 n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , 
 n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , 
 n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , 
 n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , 
 n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , 
 n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , 
 n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , 
 n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , 
 n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , 
 n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , 
 n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , 
 n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , 
 n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , 
 n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , 
 n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , 
 n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , 
 n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , 
 n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , 
 n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , 
 n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , 
 n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , 
 n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , 
 n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , 
 n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , 
 n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , 
 n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , 
 n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , 
 n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , 
 n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , 
 n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , 
 n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , 
 n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , 
 n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , 
 n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , 
 n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , 
 n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , 
 n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , 
 n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , 
 n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , 
 n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , 
 n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , 
 n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , 
 n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , 
 n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , 
 n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , 
 n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , 
 n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , 
 n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , 
 n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , 
 n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , 
 n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , 
 n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , 
 n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , 
 n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , 
 n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , 
 n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , 
 n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , 
 n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , 
 n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , 
 n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , 
 n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , 
 n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , 
 n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , 
 n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , 
 n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , 
 n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , 
 n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , 
 n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , 
 n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , 
 n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , 
 n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , 
 n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , 
 n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , 
 n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , 
 n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , 
 n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , 
 n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , 
 n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , 
 n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , 
 n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , 
 n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , 
 n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , 
 n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , 
 n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , 
 n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , 
 n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , 
 n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , 
 n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , 
 n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , 
 n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , 
 n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , 
 n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , 
 n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , 
 n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , 
 n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , 
 n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , 
 n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , 
 n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , 
 n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , 
 n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , 
 n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , 
 n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , 
 n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , 
 n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , 
 n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , 
 n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , 
 n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , 
 n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , 
 n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , 
 n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , 
 n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , 
 n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , 
 n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , 
 n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , 
 n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , 
 n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , 
 n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , 
 n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , 
 n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , 
 n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , 
 n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , 
 n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , 
 n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , 
 n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , 
 n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , 
 n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , 
 n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , 
 n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , 
 n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , 
 n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , 
 n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , 
 n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , 
 n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , 
 n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , 
 n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , 
 n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , 
 n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , 
 n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , 
 n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , 
 n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , 
 n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , 
 n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , 
 n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , 
 n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , 
 n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , 
 n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , 
 n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , 
 n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , 
 n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , 
 n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , 
 n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , 
 n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , 
 n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , 
 n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n111813 , n111814 , n4262 , n4263 , 
 n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , 
 n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , 
 n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , 
 n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , 
 n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , 
 n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , 
 n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , 
 n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , 
 n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , 
 n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , 
 n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , 
 n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , 
 n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , 
 n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , 
 n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , 
 n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , 
 n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , 
 n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , 
 n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , 
 n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , 
 n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , 
 n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , 
 n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , 
 n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , 
 n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , 
 n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , 
 n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , 
 n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , 
 n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , 
 n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , 
 n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , 
 n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , 
 n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , 
 n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , 
 n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , 
 n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , 
 n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , 
 n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , 
 n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , 
 n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , 
 n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , 
 n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , 
 n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , 
 n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , 
 n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , 
 n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , 
 n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , 
 n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , 
 n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , 
 n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , 
 n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , 
 n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , 
 n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , 
 n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , 
 n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , 
 n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , 
 n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , 
 n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , 
 n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , 
 n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , 
 n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , 
 n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , 
 n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , 
 n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , 
 n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , 
 n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , 
 n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , 
 n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , 
 n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , 
 n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , 
 n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , 
 n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , 
 n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , 
 n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , 
 n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , 
 n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , 
 n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , 
 n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , 
 n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , 
 n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , 
 n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , 
 n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , 
 n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , 
 n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , 
 n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , 
 n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , 
 n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , 
 n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , 
 n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , 
 n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , 
 n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , 
 n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , 
 n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , 
 n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , 
 n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , 
 n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , 
 n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , 
 n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , 
 n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , 
 n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , 
 n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , 
 n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , 
 n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , 
 n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , 
 n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , 
 n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , 
 n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , 
 n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , 
 n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , 
 n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , 
 n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , 
 n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , 
 n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , 
 n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , 
 n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , 
 n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , 
 n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , 
 n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , 
 n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , 
 n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , 
 n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , 
 n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , 
 n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , 
 n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , 
 n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , 
 n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , 
 n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , 
 n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , 
 n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , 
 n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , 
 n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , 
 n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , 
 n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , 
 n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , 
 n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , 
 n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , 
 n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , 
 n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , 
 n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , 
 n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , 
 n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , 
 n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , 
 n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , 
 n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , 
 n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , 
 n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , 
 n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , 
 n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , 
 n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , 
 n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , 
 n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , 
 n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , 
 n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , 
 n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , 
 n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , 
 n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , 
 n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , 
 n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , 
 n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , 
 n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , 
 n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , 
 n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , 
 n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , 
 n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , 
 n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , 
 n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , 
 n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , 
 n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , 
 n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , 
 n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , 
 n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , 
 n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , 
 n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , 
 n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , 
 n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , 
 n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , 
 n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , 
 n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , 
 n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , 
 n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , 
 n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , 
 n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , 
 n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , 
 n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , 
 n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , 
 n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , 
 n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , 
 n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , 
 n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , 
 n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , 
 n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , 
 n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , 
 n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , 
 n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , 
 n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , 
 n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , 
 n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , 
 n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , 
 n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , 
 n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , 
 n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , 
 n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , 
 n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , 
 n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , 
 n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , 
 n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , 
 n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , 
 n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , 
 n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , 
 n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , 
 n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , 
 n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , 
 n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , 
 n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , 
 n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , 
 n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , 
 n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , 
 n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , 
 n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , 
 n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , 
 n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , 
 n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , 
 n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , 
 n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , 
 n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , 
 n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , 
 n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , 
 n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , 
 n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , 
 n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , 
 n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , 
 n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6583 , n6584 , 
 n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , 
 n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , 
 n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , 
 n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , 
 n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , 
 n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , 
 n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , 
 n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , 
 n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , 
 n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , 
 n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , 
 n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , 
 n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , 
 n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , 
 n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , 
 n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , 
 n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , 
 n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , 
 n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , 
 n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , 
 n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , 
 n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , 
 n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , 
 n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , 
 n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , 
 n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , 
 n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , 
 n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , 
 n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , 
 n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , 
 n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , 
 n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , 
 n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , 
 n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , 
 n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , 
 n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , 
 n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , 
 n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , 
 n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , 
 n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , 
 n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , 
 n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , 
 n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , 
 n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , 
 n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , 
 n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , 
 n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , 
 n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , 
 n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , 
 n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , 
 n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , 
 n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , 
 n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , 
 n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , 
 n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , 
 n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , 
 n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , 
 n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , 
 n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , 
 n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , 
 n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , 
 n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , 
 n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , 
 n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , 
 n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , 
 n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , 
 n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , 
 n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , 
 n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , 
 n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , 
 n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , 
 n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , 
 n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , 
 n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , 
 n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , 
 n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , 
 n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , 
 n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , 
 n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , 
 n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , 
 n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , 
 n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , 
 n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , 
 n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , 
 n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , 
 n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , 
 n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , 
 n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , 
 n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , 
 n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , 
 n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , 
 n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , 
 n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , 
 n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , 
 n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , 
 n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , 
 n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , 
 n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , 
 n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , 
 n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , 
 n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , 
 n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , 
 n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , 
 n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , 
 n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , 
 n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , 
 n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , 
 n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , 
 n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , 
 n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , 
 n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , 
 n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , 
 n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , 
 n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , 
 n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , 
 n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , 
 n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , 
 n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , 
 n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , 
 n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , 
 n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , 
 n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , 
 n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , 
 n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , 
 n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , 
 n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , 
 n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , 
 n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , 
 n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , 
 n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , 
 n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , 
 n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , 
 n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , 
 n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , 
 n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , 
 n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , 
 n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , 
 n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , 
 n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , 
 n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , 
 n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , 
 n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , 
 n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , 
 n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , 
 n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , 
 n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , 
 n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , 
 n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , 
 n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , 
 n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , 
 n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , 
 n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , 
 n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , 
 n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , 
 n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , 
 n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , 
 n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , 
 n8555 , n8556 , n8557 , n8558 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , 
 n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , 
 n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , 
 n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , 
 n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , 
 n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , 
 n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , 
 n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , 
 n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , 
 n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , 
 n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , 
 n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , 
 n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , 
 n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , 
 n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , 
 n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , 
 n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , 
 n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , 
 n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , 
 n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , 
 n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , 
 n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , 
 n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , 
 n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , 
 n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , 
 n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , 
 n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , 
 n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , 
 n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , 
 n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , 
 n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , 
 n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , 
 n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , 
 n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , 
 n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , 
 n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , 
 n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , 
 n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , 
 n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , 
 n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , 
 n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , 
 n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , 
 n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , 
 n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , 
 n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , 
 n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , 
 n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , 
 n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , 
 n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , 
 n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , 
 n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , 
 n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , 
 n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , 
 n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , 
 n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , 
 n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , 
 n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , 
 n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , 
 n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , 
 n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , 
 n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , 
 n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , 
 n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , 
 n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , 
 n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , 
 n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , 
 n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , 
 n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , 
 n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n116794 , n9243 , n9244 , 
 n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , 
 n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , 
 n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , 
 n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , 
 n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , 
 n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , 
 n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , 
 n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , 
 n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , 
 n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , 
 n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , 
 n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , 
 n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , 
 n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , 
 n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , 
 n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , 
 n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , 
 n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , 
 n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , 
 n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , 
 n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , 
 n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , 
 n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , 
 n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , 
 n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , 
 n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , 
 n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , 
 n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , 
 n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , 
 n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , 
 n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , 
 n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , 
 n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , 
 n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , 
 n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , 
 n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , 
 n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , 
 n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , 
 n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , 
 n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , 
 n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , 
 n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , 
 n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , 
 n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , 
 n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , 
 n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , 
 n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , 
 n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , 
 n9725 , n9726 , n9727 , n9728 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , 
 n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , 
 n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , 
 n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , 
 n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
 n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
 n9786 , n9787 , n9788 , n9789 , n9790 , n9792 , n9793 , n9794 , n9795 , n9796 , 
 n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , 
 n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , 
 n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , 
 n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , 
 n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , 
 n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , 
 n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , 
 n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , 
 n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , 
 n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , 
 n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , 
 n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , 
 n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , 
 n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , 
 n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , 
 n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , 
 n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , 
 n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , 
 n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , 
 n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , 
 n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , 
 n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , 
 n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , 
 n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , 
 n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , 
 n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , 
 n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , 
 n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , 
 n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , 
 n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
 n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , 
 n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , 
 n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , 
 n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , 
 n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
 n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , 
 n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , 
 n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , 
 n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , 
 n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , 
 n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , 
 n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , 
 n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , 
 n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , 
 n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , 
 n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , 
 n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , 
 n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , 
 n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , 
 n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , 
 n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , 
 n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , 
 n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , 
 n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , 
 n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , 
 n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , 
 n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , 
 n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , 
 n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , 
 n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , 
 n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , 
 n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , 
 n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , 
 n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , 
 n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , 
 n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , 
 n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , 
 n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , 
 n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , 
 n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , 
 n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , 
 n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , 
 n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , 
 n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , 
 n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , 
 n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , 
 n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , 
 n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , 
 n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , 
 n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , 
 n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , 
 n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , 
 n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , 
 n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , 
 n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , 
 n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , 
 n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , 
 n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , 
 n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , 
 n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , 
 n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , 
 n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , 
 n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , 
 n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , 
 n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , 
 n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , 
 n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , 
 n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , 
 n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , 
 n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , 
 n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , 
 n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , 
 n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , 
 n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , 
 n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , 
 n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , 
 n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , 
 n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , 
 n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , 
 n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , 
 n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , 
 n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , 
 n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , 
 n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , 
 n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , 
 n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , 
 n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , 
 n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , 
 n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , 
 n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , 
 n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , 
 n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , 
 n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , 
 n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , 
 n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , 
 n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , 
 n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , 
 n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , 
 n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , 
 n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , 
 n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , 
 n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , 
 n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , 
 n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , 
 n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , 
 n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , 
 n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , 
 n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , 
 n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , 
 n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , 
 n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , 
 n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , 
 n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , 
 n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , 
 n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , 
 n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , 
 n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , 
 n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , 
 n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , 
 n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , 
 n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , 
 n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , 
 n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , 
 n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , 
 n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , 
 n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , 
 n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , 
 n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , 
 n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , 
 n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , 
 n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , 
 n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , 
 n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , 
 n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , 
 n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , 
 n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , 
 n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
 n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , 
 n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , 
 n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , 
 n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , 
 n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , 
 n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , 
 n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , 
 n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , 
 n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , 
 n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , 
 n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , 
 n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , 
 n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , 
 n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , 
 n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , 
 n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , 
 n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , 
 n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , 
 n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , 
 n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , 
 n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , 
 n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , 
 n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , 
 n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , 
 n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , 
 n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , 
 n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , 
 n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , 
 n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , 
 n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , 
 n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , 
 n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , 
 n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , 
 n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , 
 n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , 
 n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , 
 n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , 
 n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , 
 n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , 
 n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , 
 n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , 
 n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , 
 n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , 
 n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , 
 n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , 
 n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , 
 n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , 
 n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , 
 n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , 
 n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , 
 n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , 
 n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , 
 n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , 
 n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , 
 n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , 
 n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , 
 n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , 
 n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , 
 n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , 
 n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , 
 n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , 
 n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , 
 n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , 
 n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , 
 n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , 
 n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , 
 n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , 
 n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , 
 n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , 
 n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , 
 n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , 
 n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , 
 n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , 
 n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , 
 n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , 
 n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , 
 n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , 
 n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , 
 n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , 
 n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , 
 n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , 
 n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , 
 n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , 
 n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , 
 n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , 
 n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , 
 n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , 
 n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , 
 n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , 
 n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , 
 n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , 
 n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , 
 n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , 
 n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , 
 n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , 
 n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , 
 n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , 
 n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , 
 n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , 
 n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , 
 n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , 
 n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , 
 n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , 
 n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , 
 n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , 
 n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , 
 n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , 
 n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , 
 n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , 
 n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , 
 n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , 
 n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , 
 n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , 
 n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , 
 n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , 
 n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , 
 n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , 
 n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , 
 n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , 
 n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , 
 n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , 
 n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , 
 n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , 
 n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , 
 n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , 
 n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , 
 n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , 
 n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , 
 n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , 
 n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , 
 n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , 
 n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , 
 n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , 
 n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , 
 n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , 
 n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , 
 n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , 
 n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , 
 n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , 
 n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , 
 n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , 
 n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , 
 n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , 
 n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , 
 n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , 
 n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , 
 n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , 
 n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , 
 n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , 
 n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , 
 n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , 
 n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , 
 n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , 
 n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , 
 n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , 
 n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , 
 n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , 
 n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , 
 n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , 
 n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , 
 n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , 
 n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , 
 n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , 
 n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , 
 n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , 
 n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , 
 n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , 
 n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , 
 n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , 
 n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , 
 n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , 
 n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , 
 n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , 
 n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , 
 n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , 
 n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , 
 n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , 
 n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , 
 n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , 
 n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , 
 n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , 
 n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , 
 n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , 
 n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , 
 n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , 
 n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , 
 n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , 
 n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , 
 n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , 
 n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , 
 n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , 
 n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , 
 n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , 
 n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , 
 n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , 
 n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , 
 n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
 n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
 n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , 
 n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , 
 n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , 
 n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , 
 n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , 
 n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , 
 n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , 
 n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , 
 n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , 
 n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , 
 n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , 
 n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , 
 n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , 
 n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , 
 n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , 
 n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , 
 n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , 
 n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , 
 n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , 
 n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , 
 n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , 
 n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , 
 n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , 
 n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , 
 n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , 
 n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , 
 n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , 
 n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , 
 n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , 
 n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , 
 n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , 
 n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , 
 n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , 
 n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , 
 n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , 
 n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , 
 n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , 
 n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , 
 n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , 
 n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , 
 n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , 
 n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , 
 n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , 
 n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , 
 n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , 
 n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , 
 n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , 
 n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , 
 n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , 
 n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , 
 n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , 
 n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , 
 n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
 n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
 n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
 n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
 n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , 
 n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
 n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
 n121587 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , 
 n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , 
 n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , 
 n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , 
 n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , 
 n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , 
 n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , 
 n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , 
 n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , 
 n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , 
 n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , 
 n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , 
 n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , 
 n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , 
 n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , 
 n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , 
 n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , 
 n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , 
 n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , 
 n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , 
 n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , 
 n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , 
 n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , 
 n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , 
 n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , 
 n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , 
 n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , 
 n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , 
 n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , 
 n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , 
 n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , 
 n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , 
 n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , 
 n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , 
 n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , 
 n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , 
 n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , 
 n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , 
 n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , 
 n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , 
 n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , 
 n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , 
 n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , 
 n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , 
 n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , 
 n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , 
 n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , 
 n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , 
 n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , 
 n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , 
 n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , 
 n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , 
 n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , 
 n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , 
 n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , 
 n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , 
 n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , 
 n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , 
 n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , 
 n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , 
 n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , 
 n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , 
 n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , 
 n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , 
 n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , 
 n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , 
 n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , 
 n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , 
 n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , 
 n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , 
 n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , 
 n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , 
 n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , 
 n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , 
 n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , 
 n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , 
 n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , 
 n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , 
 n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , 
 n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , 
 n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , 
 n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , 
 n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , 
 n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , 
 n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , 
 n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , 
 n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , 
 n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , 
 n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , 
 n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , 
 n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , 
 n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , 
 n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , 
 n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , 
 n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , 
 n14986 , n14987 , n14988 , n14989 , n14990 , n122542 , n14991 , n14992 , n14993 , n14994 , 
 n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , 
 n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , 
 n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , 
 n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , 
 n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , 
 n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , 
 n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , 
 n122617 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , 
 n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , 
 n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , 
 n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , 
 n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , 
 n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , 
 n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , 
 n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , 
 n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , 
 n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , 
 n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , 
 n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , 
 n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , 
 n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , 
 n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , 
 n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , 
 n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , 
 n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , 
 n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , 
 n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , 
 n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , 
 n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , 
 n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , 
 n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , 
 n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , 
 n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , 
 n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , 
 n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , 
 n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , 
 n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , 
 n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , 
 n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , 
 n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , 
 n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , 
 n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , 
 n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , 
 n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , 
 n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , 
 n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , 
 n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , 
 n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , 
 n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , 
 n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , 
 n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , 
 n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , 
 n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , 
 n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , 
 n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , 
 n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , 
 n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , 
 n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , 
 n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , 
 n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , 
 n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , 
 n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , 
 n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , 
 n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , 
 n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , 
 n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , 
 n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , 
 n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , 
 n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , 
 n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , 
 n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , 
 n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , 
 n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , 
 n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , 
 n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , 
 n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , 
 n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , 
 n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , 
 n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , 
 n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , 
 n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , 
 n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , 
 n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , 
 n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , 
 n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , 
 n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , 
 n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , 
 n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , 
 n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , 
 n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , 
 n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , 
 n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , 
 n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , 
 n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , 
 n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , 
 n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , 
 n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , 
 n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , 
 n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , 
 n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , 
 n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , 
 n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , 
 n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , 
 n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , 
 n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , 
 n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , 
 n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , 
 n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , 
 n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , 
 n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , 
 n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , 
 n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , 
 n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , 
 n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , 
 n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , 
 n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , 
 n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , 
 n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , 
 n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , 
 n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , 
 n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , 
 n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , 
 n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , 
 n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , 
 n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , 
 n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , 
 n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , 
 n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , 
 n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , 
 n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , 
 n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , 
 n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , 
 n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , 
 n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , 
 n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , 
 n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , 
 n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , 
 n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , 
 n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , 
 n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , 
 n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , 
 n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , 
 n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , 
 n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , 
 n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , 
 n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , 
 n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , 
 n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , 
 n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , 
 n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , 
 n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , 
 n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , 
 n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , 
 n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , 
 n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , 
 n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , 
 n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , 
 n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , 
 n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , 
 n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , 
 n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , 
 n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , 
 n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , 
 n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , 
 n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , 
 n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , 
 n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , 
 n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , 
 n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , 
 n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , 
 n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , 
 n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , 
 n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , 
 n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , 
 n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , 
 n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , 
 n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , 
 n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , 
 n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , 
 n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , 
 n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , 
 n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , 
 n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , 
 n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , 
 n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , 
 n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , 
 n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , 
 n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , 
 n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , 
 n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , 
 n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , 
 n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , 
 n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , 
 n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , 
 n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , 
 n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , 
 n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , 
 n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , 
 n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , 
 n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , 
 n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , 
 n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , 
 n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , 
 n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , 
 n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , 
 n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , 
 n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , 
 n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , 
 n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , 
 n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , 
 n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , 
 n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , 
 n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , 
 n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , 
 n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , 
 n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , 
 n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , 
 n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , 
 n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , 
 n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , 
 n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , 
 n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , 
 n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , 
 n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , 
 n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , 
 n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , 
 n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , 
 n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , 
 n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , 
 n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , 
 n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , 
 n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , 
 n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , 
 n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , 
 n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , 
 n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , 
 n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , 
 n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , 
 n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , 
 n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , 
 n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , 
 n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , 
 n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , 
 n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , 
 n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , 
 n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , 
 n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , 
 n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , 
 n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , 
 n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , 
 n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , 
 n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , 
 n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , 
 n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , 
 n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , 
 n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , 
 n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , 
 n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , 
 n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , 
 n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , 
 n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , 
 n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , 
 n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , 
 n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , 
 n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , 
 n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , 
 n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , 
 n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , 
 n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , 
 n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , 
 n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , 
 n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , 
 n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , 
 n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , 
 n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , 
 n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , 
 n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , 
 n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , 
 n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , 
 n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , 
 n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , 
 n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , 
 n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , 
 n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , 
 n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , 
 n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , 
 n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , 
 n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , 
 n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , 
 n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , 
 n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , 
 n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , 
 n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , 
 n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , 
 n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , 
 n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , 
 n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , 
 n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , 
 n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , 
 n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , 
 n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , 
 n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , 
 n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , 
 n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , 
 n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , 
 n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , 
 n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , 
 n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , 
 n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , 
 n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , 
 n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , 
 n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , 
 n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , 
 n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , 
 n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , 
 n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , 
 n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , 
 n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , 
 n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , 
 n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , 
 n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , 
 n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , 
 n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , 
 n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , 
 n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , 
 n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , 
 n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , 
 n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , 
 n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , 
 n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , 
 n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , 
 n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , 
 n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , 
 n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , 
 n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , 
 n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , 
 n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , 
 n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , 
 n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , 
 n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , 
 n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , 
 n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , 
 n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , 
 n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , 
 n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , 
 n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , 
 n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , 
 n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , 
 n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , 
 n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , 
 n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , 
 n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , 
 n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , 
 n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , 
 n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , 
 n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , 
 n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , 
 n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , 
 n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , 
 n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , 
 n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , 
 n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , 
 n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , 
 n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , 
 n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , 
 n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , 
 n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , 
 n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , 
 n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , 
 n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , 
 n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , 
 n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , 
 n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , 
 n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , 
 n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , 
 n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , 
 n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , 
 n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , 
 n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , 
 n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , 
 n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , 
 n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , 
 n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , 
 n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , 
 n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , 
 n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , 
 n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , 
 n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , 
 n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , 
 n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , 
 n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , 
 n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , 
 n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , 
 n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , 
 n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , 
 n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , 
 n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , 
 n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , 
 n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , 
 n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , 
 n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , 
 n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , 
 n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , 
 n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , 
 n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , 
 n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , 
 n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , 
 n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , 
 n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , 
 n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , 
 n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , 
 n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , 
 n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , 
 n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , 
 n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , 
 n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , 
 n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , 
 n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , 
 n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , 
 n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , 
 n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , 
 n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , 
 n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , 
 n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , 
 n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , 
 n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , 
 n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , 
 n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , 
 n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , 
 n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , 
 n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , 
 n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , 
 n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , 
 n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , 
 n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , 
 n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , 
 n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , 
 n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , 
 n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , 
 n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , 
 n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , 
 n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , 
 n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , 
 n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , 
 n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , 
 n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , 
 n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , 
 n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , 
 n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , 
 n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , 
 n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , 
 n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , 
 n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , 
 n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , 
 n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , 
 n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , 
 n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , 
 n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , 
 n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , 
 n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , 
 n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , 
 n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , 
 n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , 
 n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , 
 n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , 
 n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , 
 n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , 
 n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , 
 n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , 
 n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , 
 n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , 
 n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , 
 n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , 
 n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , 
 n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , 
 n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , 
 n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , 
 n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , 
 n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , 
 n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , 
 n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , 
 n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , 
 n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , 
 n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , 
 n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , 
 n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , 
 n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , 
 n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , 
 n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , 
 n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , 
 n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , 
 n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , 
 n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , 
 n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , 
 n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , 
 n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , 
 n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , 
 n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , 
 n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , 
 n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , 
 n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , 
 n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , 
 n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , 
 n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , 
 n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , 
 n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , 
 n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , 
 n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , 
 n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , 
 n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , 
 n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , 
 n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , 
 n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , 
 n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , 
 n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , 
 n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , 
 n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , 
 n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , 
 n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , 
 n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , 
 n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , 
 n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , 
 n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , 
 n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , 
 n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , 
 n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , 
 n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , 
 n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , 
 n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , 
 n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , 
 n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , 
 n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , 
 n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , 
 n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , 
 n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , 
 n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , 
 n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , 
 n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , 
 n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , 
 n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , 
 n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , 
 n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , 
 n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , 
 n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , 
 n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , 
 n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , 
 n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , 
 n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , 
 n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , 
 n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , 
 n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , 
 n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , 
 n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , 
 n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , 
 n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , 
 n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , 
 n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , 
 n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , 
 n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , 
 n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , 
 n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , 
 n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , 
 n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , 
 n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , 
 n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , 
 n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , 
 n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , 
 n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , 
 n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , 
 n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , 
 n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , 
 n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , 
 n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , 
 n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , 
 n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , 
 n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , 
 n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , 
 n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , 
 n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , 
 n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , 
 n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , 
 n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , 
 n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , 
 n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , 
 n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , 
 n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , 
 n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , 
 n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , 
 n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , 
 n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , 
 n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , 
 n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , 
 n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , 
 n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , 
 n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , 
 n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , 
 n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , 
 n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , 
 n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , 
 n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , 
 n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , 
 n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , 
 n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , 
 n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , 
 n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , 
 n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , 
 n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , 
 n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , 
 n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , 
 n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , 
 n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , 
 n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , 
 n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , 
 n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , 
 n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , 
 n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , 
 n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , 
 n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , 
 n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , 
 n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , 
 n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , 
 n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , 
 n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , 
 n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , 
 n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , 
 n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , 
 n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , 
 n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , 
 n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , 
 n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , 
 n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , 
 n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , 
 n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , 
 n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , 
 n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , 
 n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , 
 n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , 
 n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , 
 n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , 
 n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , 
 n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , 
 n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , 
 n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , 
 n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , 
 n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , 
 n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , 
 n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , 
 n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , 
 n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , 
 n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , 
 n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , 
 n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , 
 n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , 
 n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , 
 n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , 
 n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , 
 n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , 
 n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , 
 n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , 
 n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , 
 n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , 
 n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , 
 n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , 
 n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , 
 n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , 
 n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , 
 n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , 
 n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , 
 n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , 
 n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , 
 n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , 
 n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , 
 n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , 
 n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , 
 n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , 
 n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , 
 n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , 
 n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , 
 n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , 
 n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , 
 n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , 
 n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , 
 n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , 
 n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , 
 n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , 
 n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , 
 n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , 
 n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , 
 n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , 
 n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , 
 n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , 
 n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , 
 n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , 
 n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , 
 n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , 
 n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , 
 n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , 
 n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , 
 n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , 
 n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , 
 n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , 
 n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , 
 n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , 
 n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , 
 n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , 
 n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , 
 n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , 
 n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , 
 n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , 
 n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , 
 n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , 
 n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , 
 n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , 
 n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , 
 n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , 
 n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , 
 n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , 
 n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , 
 n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , 
 n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , 
 n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , 
 n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , 
 n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , 
 n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , 
 n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , 
 n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , 
 n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , 
 n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , 
 n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , 
 n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , 
 n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , 
 n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , 
 n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , 
 n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , 
 n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , 
 n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , 
 n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , 
 n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , 
 n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , 
 n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , 
 n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , 
 n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , 
 n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , 
 n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , 
 n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , 
 n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , 
 n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , 
 n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , 
 n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , 
 n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , 
 n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , 
 n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , 
 n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , 
 n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , 
 n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , 
 n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , 
 n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , 
 n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , 
 n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , 
 n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , 
 n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , 
 n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , 
 n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , 
 n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , 
 n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , 
 n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , 
 n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , 
 n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , 
 n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , 
 n22684 , n22685 , n22686 , n130240 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , 
 n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , 
 n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , 
 n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , 
 n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , 
 n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , 
 n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , 
 n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , 
 n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , 
 n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , 
 n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , 
 n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , 
 n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , 
 n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , 
 n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , 
 n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , 
 n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , 
 n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , 
 n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , 
 n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , 
 n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , 
 n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , 
 n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , 
 n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , 
 n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , 
 n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , 
 n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , 
 n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , 
 n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , 
 n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , 
 n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , 
 n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , 
 n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , 
 n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , 
 n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , 
 n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , 
 n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , 
 n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , 
 n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , 
 n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , 
 n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , 
 n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , 
 n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , 
 n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , 
 n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , 
 n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , 
 n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , 
 n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , 
 n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , 
 n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , 
 n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , 
 n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , 
 n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , 
 n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , 
 n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , 
 n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , 
 n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , 
 n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , 
 n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , 
 n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , 
 n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , 
 n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , 
 n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , 
 n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , 
 n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , 
 n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , 
 n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , 
 n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , 
 n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , 
 n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , 
 n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , 
 n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , 
 n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , 
 n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , 
 n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , 
 n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , 
 n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , 
 n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , 
 n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , 
 n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , 
 n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , 
 n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , 
 n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , 
 n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , 
 n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , 
 n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , 
 n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , 
 n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , 
 n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , 
 n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , 
 n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , 
 n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , 
 n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , 
 n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , 
 n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , 
 n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , 
 n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , 
 n23653 , n131208 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , 
 n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , 
 n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , 
 n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , 
 n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , 
 n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , 
 n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , 
 n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , 
 n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , 
 n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , 
 n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , 
 n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , 
 n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , 
 n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , 
 n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , 
 n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , 
 n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , 
 n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , 
 n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , 
 n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , 
 n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , 
 n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , 
 n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , 
 n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , 
 n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , 
 n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , 
 n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , 
 n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , 
 n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , 
 n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , 
 n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , 
 n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , 
 n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , 
 n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , 
 n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , 
 n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , 
 n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , 
 n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , 
 n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , 
 n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , 
 n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , 
 n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , 
 n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , 
 n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , 
 n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , 
 n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , 
 n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , 
 n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , 
 n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , 
 n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , 
 n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , 
 n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , 
 n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , 
 n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , 
 n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , 
 n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , 
 n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , 
 n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , 
 n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , 
 n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , 
 n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , 
 n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , 
 n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , 
 n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , 
 n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , 
 n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , 
 n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , 
 n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , 
 n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , 
 n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , 
 n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , 
 n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , 
 n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , 
 n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , 
 n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , 
 n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , 
 n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , 
 n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , 
 n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , 
 n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , 
 n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , 
 n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , 
 n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , 
 n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , 
 n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , 
 n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , 
 n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , 
 n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , 
 n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , 
 n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , 
 n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , 
 n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , 
 n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , 
 n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , 
 n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , 
 n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , 
 n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , 
 n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , 
 n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , 
 n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , 
 n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24660 , n24661 , n24662 , 
 n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , 
 n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , 
 n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , 
 n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , 
 n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , 
 n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , 
 n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , 
 n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , 
 n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , 
 n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , 
 n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , 
 n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , 
 n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , 
 n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , 
 n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , 
 n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , 
 n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , 
 n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , 
 n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , 
 n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , 
 n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , 
 n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , 
 n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , 
 n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , 
 n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , 
 n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , 
 n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , 
 n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , 
 n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , 
 n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , 
 n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , 
 n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , 
 n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , 
 n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , 
 n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , 
 n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , 
 n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , 
 n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , 
 n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , 
 n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , 
 n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , 
 n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , 
 n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , 
 n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , 
 n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , 
 n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , 
 n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , 
 n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , 
 n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , 
 n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , 
 n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , 
 n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , 
 n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , 
 n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , 
 n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , 
 n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , 
 n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , 
 n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , 
 n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , 
 n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , 
 n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , 
 n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , 
 n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , 
 n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , 
 n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , 
 n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , 
 n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , 
 n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , 
 n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , 
 n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , 
 n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , 
 n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , 
 n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , 
 n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , 
 n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , 
 n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , 
 n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , 
 n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , 
 n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , 
 n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , 
 n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , 
 n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , 
 n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , 
 n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , 
 n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , 
 n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , 
 n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , 
 n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25543 , 
 n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , 
 n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , 
 n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , 
 n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , 
 n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , 
 n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , 
 n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , 
 n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , 
 n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , 
 n25634 , n25635 , n25636 , n25637 , n25638 , n25640 , n25641 , n25642 , n25643 , n25644 , 
 n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , 
 n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , 
 n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , 
 n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , 
 n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , 
 n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , 
 n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , 
 n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , 
 n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , 
 n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , 
 n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , 
 n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , 
 n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , 
 n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , 
 n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , 
 n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , 
 n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , 
 n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , 
 n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , 
 n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , 
 n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , 
 n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , 
 n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , 
 n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , 
 n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , 
 n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , 
 n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , 
 n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , 
 n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , 
 n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , 
 n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , 
 n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , 
 n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , 
 n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , 
 n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , 
 n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , 
 n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , 
 n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , 
 n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , 
 n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , 
 n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , 
 n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , 
 n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , 
 n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , 
 n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , 
 n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , 
 n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , 
 n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , 
 n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , 
 n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , 
 n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , 
 n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , 
 n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , 
 n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , 
 n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , 
 n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , 
 n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , 
 n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , 
 n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , 
 n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , 
 n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , 
 n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , 
 n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , 
 n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , 
 n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , 
 n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , 
 n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , 
 n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , 
 n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , 
 n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , 
 n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , 
 n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , 
 n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , 
 n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , 
 n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , 
 n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , 
 n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , 
 n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , 
 n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , 
 n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , 
 n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , 
 n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , 
 n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , 
 n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , 
 n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , 
 n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , 
 n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , 
 n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , 
 n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , 
 n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , 
 n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , 
 n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , 
 n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , 
 n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , 
 n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , 
 n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , 
 n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , 
 n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , 
 n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , 
 n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , 
 n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , 
 n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , 
 n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , 
 n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , 
 n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , 
 n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , 
 n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , 
 n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , 
 n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , 
 n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , 
 n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , 
 n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , 
 n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , 
 n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , 
 n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , 
 n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , 
 n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , 
 n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , 
 n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , 
 n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , 
 n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , 
 n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , 
 n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , 
 n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , 
 n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , 
 n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , 
 n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , 
 n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , 
 n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , 
 n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , 
 n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , 
 n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , 
 n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , 
 n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , 
 n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , 
 n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , 
 n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , 
 n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , 
 n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , 
 n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , 
 n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , 
 n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , 
 n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , 
 n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , 
 n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , 
 n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , 
 n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , 
 n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , 
 n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , 
 n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , 
 n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , 
 n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , 
 n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , 
 n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , 
 n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , 
 n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , 
 n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , 
 n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , 
 n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , 
 n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , 
 n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , 
 n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , 
 n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , 
 n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , 
 n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , 
 n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , 
 n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , 
 n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , 
 n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , 
 n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , 
 n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , 
 n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , 
 n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , 
 n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , 
 n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , 
 n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , 
 n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , 
 n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , 
 n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , 
 n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , 
 n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27454 , n27455 , 
 n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , 
 n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , 
 n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , 
 n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , 
 n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , 
 n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , 
 n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , 
 n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , 
 n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , 
 n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27554 , n27555 , n27556 , 
 n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , 
 n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , 
 n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , 
 n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , 
 n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , 
 n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , 
 n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , 
 n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , 
 n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , 
 n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , 
 n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , 
 n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , 
 n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , 
 n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , 
 n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , 
 n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , 
 n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , 
 n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , 
 n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , 
 n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , 
 n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , 
 n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , 
 n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , 
 n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , 
 n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , 
 n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , 
 n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , 
 n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , 
 n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , 
 n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , 
 n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , 
 n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , 
 n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , 
 n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , 
 n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , 
 n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , 
 n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , 
 n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , 
 n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , 
 n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , 
 n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , 
 n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , 
 n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , 
 n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , 
 n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , 
 n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , 
 n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , 
 n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , 
 n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , 
 n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , 
 n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , 
 n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , 
 n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , 
 n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , 
 n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , 
 n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , 
 n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , 
 n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , 
 n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , 
 n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , 
 n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , 
 n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , 
 n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , 
 n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , 
 n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , 
 n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , 
 n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , 
 n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , 
 n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , 
 n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , 
 n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , 
 n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , 
 n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , 
 n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , 
 n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , 
 n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , 
 n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , 
 n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , 
 n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , 
 n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , 
 n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , 
 n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28375 , n28376 , C0n , 
 C0 , C1n , C1 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , n27914 );
buf ( n570 , n27919 );
buf ( n571 , n27836 );
buf ( n572 , n27858 );
buf ( n573 , n27764 );
buf ( n574 , n27251 );
buf ( n575 , n26152 );
buf ( n576 , n26079 );
buf ( n577 , n26003 );
buf ( n578 , n19166 );
buf ( n579 , n19175 );
buf ( n580 , n18047 );
buf ( n581 , n17721 );
buf ( n582 , n17810 );
buf ( n583 , n17782 );
buf ( n584 , n17752 );
buf ( n585 , n17851 );
buf ( n586 , n17871 );
buf ( n587 , n17912 );
buf ( n588 , n17685 );
buf ( n589 , n18238 );
buf ( n590 , n18226 );
buf ( n591 , n13996 );
buf ( n592 , n18258 );
buf ( n593 , n14029 );
buf ( n594 , n18323 );
buf ( n595 , n18446 );
buf ( n596 , n18481 );
buf ( n597 , n18516 );
buf ( n598 , n9909 );
buf ( n599 , n9920 );
buf ( n600 , n18572 );
buf ( n601 , n9937 );
buf ( n602 , n18634 );
buf ( n603 , n18668 );
buf ( n604 , n9953 );
buf ( n605 , n9971 );
buf ( n606 , n9987 );
buf ( n607 , n10008 );
buf ( n608 , n10028 );
buf ( n609 , n18788 );
buf ( n610 , n18806 );
buf ( n611 , n14012 );
buf ( n612 , n26634 );
buf ( n613 , n28357 );
buf ( n614 , n28356 );
buf ( n615 , n28308 );
buf ( n616 , n28355 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , n27399 );
buf ( n634 , n28317 );
buf ( n635 , n28376 );
buf ( n636 , n28247 );
buf ( n637 , n28144 );
buf ( n638 , n28090 );
buf ( n639 , n28132 );
buf ( n640 , n28167 );
buf ( n641 , n28211 );
buf ( n642 , n28121 );
buf ( n643 , n27302 );
buf ( n644 , n26407 );
buf ( n645 , n26455 );
buf ( n646 , n25890 );
buf ( n647 , n28368 );
buf ( n648 , n28181 );
buf ( n649 , n26558 );
buf ( n650 , n26597 );
buf ( n651 , n26614 );
buf ( n652 , n28278 );
buf ( n653 , n28257 );
buf ( n654 , n25922 );
buf ( n655 , n28230 );
buf ( n656 , n25939 );
buf ( n657 , n25953 );
buf ( n658 , n25961 );
buf ( n659 , n25981 );
buf ( n660 , n26419 );
buf ( n661 , n26432 );
buf ( n662 , n26447 );
buf ( n663 , n26469 );
buf ( n664 , n26480 );
buf ( n665 , n26497 );
buf ( n666 , n26505 );
buf ( n667 , n26526 );
buf ( n668 , n28327 );
buf ( n669 , n28337 );
buf ( n670 , n28342 );
buf ( n671 , n28322 );
buf ( n672 , n26567 );
buf ( n673 , n28332 );
buf ( n674 , n26622 );
buf ( n675 , n27317 );
buf ( n676 , n28354 );
buf ( n677 , n28373 );
buf ( n678 , n28347 );
buf ( n679 , n28295 );
buf ( n680 , n28292 );
not ( n108233 , n456 );
nand ( n681 , n108233 , n470 );
nand ( n682 , n486 , n456 );
nand ( n683 , n681 , n682 );
buf ( n684 , n683 );
buf ( n685 , n684 );
and ( n686 , n456 , n485 );
not ( n687 , n456 );
and ( n688 , n687 , n469 );
nor ( n689 , n686 , n688 );
not ( n690 , n689 );
buf ( n691 , n690 );
and ( n692 , n456 , n480 );
not ( n693 , n456 );
and ( n694 , n693 , n464 );
nor ( n695 , n692 , n694 );
not ( n696 , n695 );
buf ( n697 , n696 );
and ( n698 , n456 , n484 );
not ( n699 , n456 );
and ( n700 , n699 , n468 );
nor ( n701 , n698 , n700 );
not ( n702 , n701 );
buf ( n703 , n702 );
and ( n704 , n544 , n545 );
not ( n705 , n544 );
not ( n706 , n545 );
and ( n707 , n705 , n706 );
nor ( n708 , n704 , n707 );
not ( n709 , n708 );
and ( n710 , n543 , n544 );
nor ( n711 , n543 , n544 );
nor ( n712 , n710 , n711 );
nand ( n713 , n709 , n712 );
not ( n714 , n713 );
not ( n715 , n714 );
not ( n716 , n455 );
not ( n717 , n716 );
not ( n718 , n494 );
not ( n719 , n495 );
not ( n720 , n719 );
or ( n721 , n718 , n720 );
not ( n722 , n494 );
nand ( n723 , n722 , n495 );
nand ( n724 , n721 , n723 );
not ( n725 , n724 );
not ( n726 , n493 );
not ( n727 , n456 );
nand ( n728 , n727 , n471 );
nand ( n729 , n456 , n487 );
nand ( n730 , n728 , n729 );
not ( n731 , n730 );
not ( n732 , n731 );
or ( n733 , n726 , n732 );
and ( n734 , n456 , n487 );
not ( n735 , n456 );
and ( n736 , n735 , n471 );
nor ( n737 , n734 , n736 );
not ( n738 , n737 );
not ( n739 , n493 );
nand ( n740 , n738 , n739 );
nand ( n741 , n733 , n740 );
not ( n742 , n741 );
or ( n743 , n725 , n742 );
not ( n744 , n493 );
not ( n745 , n488 );
and ( n746 , n456 , n745 );
not ( n747 , n456 );
not ( n748 , n472 );
and ( n749 , n747 , n748 );
nor ( n750 , n746 , n749 );
buf ( n751 , n750 );
not ( n752 , n751 );
not ( n753 , n752 );
or ( n754 , n744 , n753 );
buf ( n755 , n751 );
nand ( n756 , n755 , n739 );
nand ( n757 , n754 , n756 );
xor ( n758 , n494 , n495 );
xnor ( n759 , n493 , n494 );
nor ( n760 , n758 , n759 );
nand ( n761 , n757 , n760 );
nand ( n762 , n743 , n761 );
not ( n763 , n499 );
nor ( n764 , n500 , n501 );
not ( n765 , n764 );
or ( n766 , n763 , n765 );
not ( n767 , n499 );
nand ( n768 , n767 , n501 , n500 );
nand ( n769 , n766 , n768 );
buf ( n770 , n769 );
not ( n771 , n770 );
not ( n772 , n499 );
and ( n773 , n456 , n482 );
not ( n774 , n456 );
and ( n775 , n774 , n466 );
nor ( n776 , n773 , n775 );
not ( n777 , n776 );
buf ( n778 , n777 );
not ( n779 , n778 );
not ( n780 , n779 );
or ( n781 , n772 , n780 );
not ( n782 , n499 );
nand ( n783 , n778 , n782 );
nand ( n784 , n781 , n783 );
not ( n785 , n784 );
or ( n786 , n771 , n785 );
not ( n787 , n499 );
and ( n788 , n456 , n481 );
not ( n789 , n456 );
and ( n790 , n789 , n465 );
nor ( n791 , n788 , n790 );
not ( n792 , n791 );
or ( n793 , n787 , n792 );
and ( n794 , n456 , n481 );
not ( n795 , n456 );
and ( n796 , n795 , n465 );
nor ( n797 , n794 , n796 );
not ( n798 , n797 );
nand ( n799 , n798 , n782 );
nand ( n800 , n793 , n799 );
not ( n801 , n501 );
not ( n802 , n801 );
not ( n803 , n500 );
or ( n804 , n802 , n803 );
not ( n805 , n500 );
nand ( n806 , n805 , n501 );
nand ( n807 , n804 , n806 );
nand ( n808 , n800 , n807 );
nand ( n809 , n786 , n808 );
xor ( n810 , n762 , n809 );
buf ( n811 , n751 );
nor ( n812 , n811 , n494 );
not ( n813 , n495 );
or ( n814 , n812 , n813 );
and ( n815 , n755 , n494 );
nor ( n816 , n815 , n739 );
nand ( n817 , n814 , n816 );
not ( n818 , n503 );
not ( n819 , n502 );
nand ( n820 , n818 , n819 );
not ( n821 , n820 );
nand ( n822 , n503 , n502 );
not ( n823 , n822 );
or ( n824 , n821 , n823 );
not ( n825 , n502 );
or ( n826 , n825 , n501 );
not ( n827 , n502 );
nand ( n828 , n501 , n827 );
nand ( n829 , n826 , n828 );
nand ( n830 , n824 , n829 );
not ( n831 , n830 );
not ( n832 , n831 );
not ( n833 , n501 );
and ( n834 , n696 , n833 );
not ( n835 , n696 );
and ( n836 , n835 , n501 );
or ( n837 , n834 , n836 );
not ( n838 , n837 );
or ( n839 , n832 , n838 );
not ( n840 , n501 );
and ( n841 , n456 , n479 );
not ( n842 , n456 );
and ( n843 , n842 , n463 );
nor ( n844 , n841 , n843 );
not ( n845 , n844 );
or ( n846 , n840 , n845 );
and ( n847 , n456 , n479 );
not ( n848 , n456 );
and ( n849 , n848 , n463 );
nor ( n850 , n847 , n849 );
not ( n851 , n850 );
nand ( n852 , n851 , n833 );
nand ( n853 , n846 , n852 );
and ( n854 , n503 , n827 );
not ( n855 , n503 );
and ( n856 , n855 , n502 );
nor ( n857 , n854 , n856 );
not ( n858 , n857 );
nand ( n859 , n853 , n858 );
nand ( n860 , n839 , n859 );
not ( n861 , n860 );
xor ( n862 , n817 , n861 );
xor ( n863 , n810 , n862 );
and ( n864 , n751 , n758 );
not ( n865 , n831 );
not ( n866 , n501 );
and ( n867 , n456 , n481 );
not ( n868 , n456 );
and ( n869 , n868 , n465 );
nor ( n870 , n867 , n869 );
not ( n871 , n870 );
or ( n872 , n866 , n871 );
not ( n873 , n791 );
nand ( n874 , n873 , n833 );
nand ( n875 , n872 , n874 );
not ( n876 , n875 );
or ( n877 , n865 , n876 );
not ( n878 , n503 );
or ( n879 , n878 , n502 );
not ( n880 , n503 );
nand ( n881 , n880 , n502 );
nand ( n882 , n879 , n881 );
nand ( n883 , n837 , n882 );
nand ( n884 , n877 , n883 );
xor ( n885 , n864 , n884 );
not ( n886 , n497 );
nor ( n887 , n498 , n499 );
not ( n888 , n887 );
or ( n889 , n886 , n888 );
not ( n890 , n497 );
nand ( n891 , n890 , n498 , n499 );
nand ( n892 , n889 , n891 );
buf ( n893 , n892 );
not ( n894 , n893 );
not ( n895 , n497 );
not ( n896 , n690 );
not ( n897 , n896 );
or ( n898 , n895 , n897 );
not ( n899 , n690 );
not ( n900 , n899 );
not ( n901 , n497 );
nand ( n902 , n900 , n901 );
nand ( n903 , n898 , n902 );
not ( n904 , n903 );
or ( n905 , n894 , n904 );
not ( n906 , n497 );
not ( n907 , n701 );
or ( n908 , n906 , n907 );
nand ( n909 , n702 , n901 );
nand ( n910 , n908 , n909 );
xor ( n911 , n498 , n499 );
buf ( n912 , n911 );
nand ( n913 , n910 , n912 );
nand ( n914 , n905 , n913 );
and ( n915 , n885 , n914 );
and ( n916 , n864 , n884 );
or ( n917 , n915 , n916 );
xor ( n918 , n496 , n497 );
not ( n919 , n918 );
not ( n920 , n495 );
not ( n921 , n684 );
not ( n922 , n921 );
or ( n923 , n920 , n922 );
nand ( n924 , n684 , n813 );
nand ( n925 , n923 , n924 );
not ( n926 , n925 );
or ( n927 , n919 , n926 );
not ( n928 , n495 );
not ( n929 , n730 );
not ( n930 , n929 );
or ( n931 , n928 , n930 );
nand ( n932 , n738 , n813 );
nand ( n933 , n931 , n932 );
not ( n934 , n495 );
nand ( n935 , n496 , n497 );
not ( n936 , n935 );
and ( n937 , n934 , n936 );
nor ( n938 , n496 , n497 );
and ( n939 , n938 , n495 );
nor ( n940 , n937 , n939 );
not ( n941 , n940 );
nand ( n942 , n933 , n941 );
nand ( n943 , n927 , n942 );
not ( n944 , n504 );
nand ( n945 , n944 , n503 );
not ( n946 , n945 );
not ( n947 , n946 );
not ( n948 , n503 );
not ( n949 , n844 );
or ( n950 , n948 , n949 );
buf ( n951 , n851 );
nand ( n952 , n951 , n878 );
nand ( n953 , n950 , n952 );
not ( n954 , n953 );
or ( n955 , n947 , n954 );
not ( n956 , n503 );
and ( n957 , n456 , n478 );
not ( n958 , n456 );
and ( n959 , n958 , n462 );
nor ( n960 , n957 , n959 );
not ( n961 , n960 );
or ( n962 , n956 , n961 );
and ( n963 , n456 , n478 );
not ( n964 , n456 );
and ( n965 , n964 , n462 );
nor ( n966 , n963 , n965 );
not ( n967 , n966 );
nand ( n968 , n967 , n878 );
nand ( n969 , n962 , n968 );
nand ( n970 , n969 , n504 );
nand ( n971 , n955 , n970 );
xor ( n972 , n943 , n971 );
not ( n973 , n807 );
not ( n974 , n784 );
or ( n975 , n973 , n974 );
not ( n976 , n782 );
not ( n977 , n483 );
and ( n978 , n456 , n977 );
not ( n979 , n456 );
not ( n980 , n467 );
and ( n981 , n979 , n980 );
nor ( n982 , n978 , n981 );
not ( n983 , n982 );
or ( n984 , n976 , n983 );
and ( n985 , n456 , n483 );
not ( n986 , n456 );
and ( n987 , n986 , n467 );
nor ( n988 , n985 , n987 );
not ( n989 , n988 );
not ( n990 , n989 );
nand ( n991 , n990 , n499 );
nand ( n992 , n984 , n991 );
not ( n993 , n769 );
not ( n994 , n993 );
nand ( n995 , n992 , n994 );
nand ( n996 , n975 , n995 );
and ( n997 , n972 , n996 );
and ( n998 , n943 , n971 );
or ( n999 , n997 , n998 );
xor ( n1000 , n917 , n999 );
not ( n1001 , n893 );
not ( n1002 , n910 );
or ( n1003 , n1001 , n1002 );
and ( n1004 , n456 , n483 );
not ( n1005 , n456 );
and ( n1006 , n1005 , n467 );
or ( n1007 , n1004 , n1006 );
or ( n1008 , n1007 , n901 );
not ( n1009 , n497 );
nand ( n1010 , n1007 , n1009 );
nand ( n1011 , n1008 , n1010 );
nand ( n1012 , n1011 , n911 );
nand ( n1013 , n1003 , n1012 );
not ( n1014 , n941 );
not ( n1015 , n925 );
or ( n1016 , n1014 , n1015 );
not ( n1017 , n899 );
not ( n1018 , n495 );
or ( n1019 , n1017 , n1018 );
and ( n1020 , n456 , n485 );
not ( n1021 , n456 );
and ( n1022 , n1021 , n469 );
or ( n1023 , n1020 , n1022 );
nand ( n1024 , n1023 , n813 );
nand ( n1025 , n1019 , n1024 );
buf ( n1026 , n918 );
nand ( n1027 , n1025 , n1026 );
nand ( n1028 , n1016 , n1027 );
xor ( n1029 , n1013 , n1028 );
nand ( n1030 , n969 , n946 );
not ( n1031 , n878 );
and ( n1032 , n456 , n477 );
not ( n1033 , n456 );
and ( n1034 , n1033 , n461 );
nor ( n1035 , n1032 , n1034 );
not ( n1036 , n1035 );
buf ( n1037 , n1036 );
not ( n1038 , n1037 );
or ( n1039 , n1031 , n1038 );
and ( n1040 , n456 , n477 );
not ( n1041 , n456 );
and ( n1042 , n1041 , n461 );
nor ( n1043 , n1040 , n1042 );
nand ( n1044 , n503 , n1043 );
nand ( n1045 , n1039 , n1044 );
nand ( n1046 , n1045 , n504 );
nand ( n1047 , n1030 , n1046 );
xor ( n1048 , n1029 , n1047 );
xor ( n1049 , n1000 , n1048 );
xor ( n1050 , n863 , n1049 );
not ( n1051 , n938 );
and ( n1052 , n755 , n1051 );
nand ( n1053 , n496 , n497 );
nand ( n1054 , n1053 , n495 );
nor ( n1055 , n1052 , n1054 );
not ( n1056 , n882 );
not ( n1057 , n875 );
or ( n1058 , n1056 , n1057 );
not ( n1059 , n501 );
and ( n1060 , n456 , n482 );
not ( n1061 , n456 );
and ( n1062 , n1061 , n466 );
nor ( n1063 , n1060 , n1062 );
not ( n1064 , n1063 );
not ( n1065 , n1064 );
not ( n1066 , n1065 );
or ( n1067 , n1059 , n1066 );
nand ( n1068 , n1064 , n833 );
nand ( n1069 , n1067 , n1068 );
nand ( n1070 , n1069 , n831 );
nand ( n1071 , n1058 , n1070 );
and ( n1072 , n1055 , n1071 );
not ( n1073 , n893 );
not ( n1074 , n684 );
not ( n1075 , n901 );
or ( n1076 , n1074 , n1075 );
not ( n1077 , n456 );
nand ( n1078 , n1077 , n470 );
nand ( n1079 , n456 , n486 );
nand ( n1080 , n1078 , n1079 , n497 );
nand ( n1081 , n1076 , n1080 );
not ( n1082 , n1081 );
or ( n1083 , n1073 , n1082 );
nand ( n1084 , n903 , n912 );
nand ( n1085 , n1083 , n1084 );
not ( n1086 , n940 );
not ( n1087 , n1086 );
not ( n1088 , n751 );
and ( n1089 , n813 , n1088 );
not ( n1090 , n813 );
and ( n1091 , n1090 , n751 );
nor ( n1092 , n1089 , n1091 );
not ( n1093 , n1092 );
or ( n1094 , n1087 , n1093 );
nand ( n1095 , n933 , n1026 );
nand ( n1096 , n1094 , n1095 );
xor ( n1097 , n1085 , n1096 );
not ( n1098 , n504 );
not ( n1099 , n953 );
or ( n1100 , n1098 , n1099 );
not ( n1101 , n503 );
not ( n1102 , n695 );
or ( n1103 , n1101 , n1102 );
nand ( n1104 , n696 , n878 );
nand ( n1105 , n1103 , n1104 );
nand ( n1106 , n1105 , n946 );
nand ( n1107 , n1100 , n1106 );
and ( n1108 , n1097 , n1107 );
and ( n1109 , n1085 , n1096 );
or ( n1110 , n1108 , n1109 );
xor ( n1111 , n1072 , n1110 );
xor ( n1112 , n864 , n884 );
xor ( n1113 , n1112 , n914 );
and ( n1114 , n1111 , n1113 );
and ( n1115 , n1072 , n1110 );
or ( n1116 , n1114 , n1115 );
xor ( n1117 , n1050 , n1116 );
not ( n1118 , n1117 );
xor ( n1119 , n943 , n971 );
xor ( n1120 , n1119 , n996 );
not ( n1121 , n992 );
xor ( n1122 , n500 , n501 );
not ( n1123 , n1122 );
or ( n1124 , n1121 , n1123 );
not ( n1125 , n782 );
and ( n1126 , n456 , n484 );
not ( n1127 , n456 );
and ( n1128 , n1127 , n468 );
nor ( n1129 , n1126 , n1128 );
not ( n1130 , n1129 );
not ( n1131 , n1130 );
or ( n1132 , n1125 , n1131 );
nand ( n1133 , n1129 , n499 );
nand ( n1134 , n1132 , n1133 );
nand ( n1135 , n770 , n1134 );
nand ( n1136 , n1124 , n1135 );
xor ( n1137 , n1055 , n1071 );
xor ( n1138 , n1136 , n1137 );
and ( n1139 , n751 , n918 );
not ( n1140 , n504 );
not ( n1141 , n1105 );
or ( n1142 , n1140 , n1141 );
not ( n1143 , n503 );
not ( n1144 , n797 );
or ( n1145 , n1143 , n1144 );
nand ( n1146 , n873 , n878 );
nand ( n1147 , n1145 , n1146 );
nand ( n1148 , n1147 , n946 );
nand ( n1149 , n1142 , n1148 );
xor ( n1150 , n1139 , n1149 );
not ( n1151 , n912 );
not ( n1152 , n1081 );
or ( n1153 , n1151 , n1152 );
not ( n1154 , n497 );
not ( n1155 , n731 );
or ( n1156 , n1154 , n1155 );
nand ( n1157 , n738 , n901 );
nand ( n1158 , n1156 , n1157 );
nand ( n1159 , n1158 , n893 );
nand ( n1160 , n1153 , n1159 );
and ( n1161 , n1150 , n1160 );
and ( n1162 , n1139 , n1149 );
or ( n1163 , n1161 , n1162 );
and ( n1164 , n1138 , n1163 );
and ( n1165 , n1136 , n1137 );
or ( n1166 , n1164 , n1165 );
xor ( n1167 , n1120 , n1166 );
xor ( n1168 , n1072 , n1110 );
xor ( n1169 , n1168 , n1113 );
and ( n1170 , n1167 , n1169 );
and ( n1171 , n1120 , n1166 );
or ( n1172 , n1170 , n1171 );
not ( n1173 , n1172 );
nand ( n1174 , n1118 , n1173 );
nand ( n1175 , n1172 , n1117 );
nand ( n1176 , n1174 , n1175 );
xor ( n1177 , n1120 , n1166 );
xor ( n1178 , n1177 , n1169 );
not ( n1179 , n1178 );
xor ( n1180 , n1085 , n1096 );
xor ( n1181 , n1180 , n1107 );
not ( n1182 , n822 );
not ( n1183 , n820 );
or ( n1184 , n1182 , n1183 );
nor ( n1185 , n825 , n501 );
nor ( n1186 , n801 , n502 );
or ( n1187 , n1185 , n1186 );
nand ( n1188 , n1184 , n1187 );
not ( n1189 , n1188 );
not ( n1190 , n1189 );
nand ( n1191 , n989 , n833 );
and ( n1192 , n456 , n483 );
not ( n1193 , n456 );
and ( n1194 , n1193 , n467 );
nor ( n1195 , n1192 , n1194 );
nand ( n1196 , n1195 , n501 );
nand ( n1197 , n1191 , n1196 );
not ( n1198 , n1197 );
or ( n1199 , n1190 , n1198 );
nand ( n1200 , n1069 , n882 );
nand ( n1201 , n1199 , n1200 );
not ( n1202 , n770 );
not ( n1203 , n499 );
not ( n1204 , n900 );
not ( n1205 , n1204 );
or ( n1206 , n1203 , n1205 );
not ( n1207 , n896 );
nand ( n1208 , n1207 , n782 );
nand ( n1209 , n1206 , n1208 );
not ( n1210 , n1209 );
or ( n1211 , n1202 , n1210 );
nand ( n1212 , n1134 , n1122 );
nand ( n1213 , n1211 , n1212 );
xor ( n1214 , n1201 , n1213 );
buf ( n1215 , n751 );
nor ( n1216 , n498 , n499 );
not ( n1217 , n1216 );
and ( n1218 , n1215 , n1217 );
nand ( n1219 , n498 , n499 );
nand ( n1220 , n1219 , n497 );
nor ( n1221 , n1218 , n1220 );
not ( n1222 , n946 );
not ( n1223 , n1064 );
not ( n1224 , n878 );
or ( n1225 , n1223 , n1224 );
nand ( n1226 , n503 , n1063 );
nand ( n1227 , n1225 , n1226 );
not ( n1228 , n1227 );
or ( n1229 , n1222 , n1228 );
nand ( n1230 , n1147 , n504 );
nand ( n1231 , n1229 , n1230 );
and ( n1232 , n1221 , n1231 );
and ( n1233 , n1214 , n1232 );
and ( n1234 , n1201 , n1213 );
or ( n1235 , n1233 , n1234 );
xor ( n1236 , n1181 , n1235 );
xor ( n1237 , n1136 , n1137 );
xor ( n1238 , n1237 , n1163 );
and ( n1239 , n1236 , n1238 );
and ( n1240 , n1181 , n1235 );
or ( n1241 , n1239 , n1240 );
not ( n1242 , n1241 );
nand ( n1243 , n1179 , n1242 );
not ( n1244 , n1243 );
xor ( n1245 , n1181 , n1235 );
xor ( n1246 , n1245 , n1238 );
not ( n1247 , n912 );
not ( n1248 , n1158 );
or ( n1249 , n1247 , n1248 );
not ( n1250 , n751 );
and ( n1251 , n1216 , n497 );
and ( n1252 , n1250 , n1251 );
nor ( n1253 , n1219 , n497 );
and ( n1254 , n751 , n1253 );
nor ( n1255 , n1252 , n1254 );
nand ( n1256 , n1249 , n1255 );
not ( n1257 , n702 );
not ( n1258 , n833 );
or ( n1259 , n1257 , n1258 );
and ( n1260 , n456 , n484 );
not ( n1261 , n456 );
and ( n1262 , n1261 , n468 );
nor ( n1263 , n1260 , n1262 );
nand ( n1264 , n1263 , n501 );
nand ( n1265 , n1259 , n1264 );
not ( n1266 , n1265 );
not ( n1267 , n1189 );
or ( n1268 , n1266 , n1267 );
not ( n1269 , n1196 );
not ( n1270 , n1191 );
or ( n1271 , n1269 , n1270 );
nand ( n1272 , n1271 , n858 );
nand ( n1273 , n1268 , n1272 );
xor ( n1274 , n1256 , n1273 );
not ( n1275 , n807 );
not ( n1276 , n1209 );
or ( n1277 , n1275 , n1276 );
not ( n1278 , n499 );
not ( n1279 , n684 );
not ( n1280 , n1279 );
or ( n1281 , n1278 , n1280 );
nand ( n1282 , n684 , n782 );
nand ( n1283 , n1281 , n1282 );
nand ( n1284 , n1283 , n770 );
nand ( n1285 , n1277 , n1284 );
and ( n1286 , n1274 , n1285 );
and ( n1287 , n1256 , n1273 );
or ( n1288 , n1286 , n1287 );
xor ( n1289 , n1139 , n1149 );
xor ( n1290 , n1289 , n1160 );
xor ( n1291 , n1288 , n1290 );
xor ( n1292 , n1201 , n1213 );
xor ( n1293 , n1292 , n1232 );
and ( n1294 , n1291 , n1293 );
and ( n1295 , n1288 , n1290 );
or ( n1296 , n1294 , n1295 );
nor ( n1297 , n1246 , n1296 );
xor ( n1298 , n1288 , n1290 );
xor ( n1299 , n1298 , n1293 );
xor ( n1300 , n1221 , n1231 );
and ( n1301 , n751 , n911 );
not ( n1302 , n946 );
not ( n1303 , n503 );
not ( n1304 , n1195 );
or ( n1305 , n1303 , n1304 );
and ( n1306 , n456 , n483 );
not ( n1307 , n456 );
and ( n1308 , n1307 , n467 );
or ( n1309 , n1306 , n1308 );
nand ( n1310 , n1309 , n878 );
nand ( n1311 , n1305 , n1310 );
not ( n1312 , n1311 );
or ( n1313 , n1302 , n1312 );
nand ( n1314 , n1227 , n504 );
nand ( n1315 , n1313 , n1314 );
xor ( n1316 , n1301 , n1315 );
not ( n1317 , n858 );
not ( n1318 , n1265 );
or ( n1319 , n1317 , n1318 );
not ( n1320 , n501 );
and ( n1321 , n456 , n485 );
not ( n1322 , n456 );
and ( n1323 , n1322 , n469 );
nor ( n1324 , n1321 , n1323 );
not ( n1325 , n1324 );
or ( n1326 , n1320 , n1325 );
nand ( n1327 , n900 , n833 );
nand ( n1328 , n1326 , n1327 );
nand ( n1329 , n1328 , n831 );
nand ( n1330 , n1319 , n1329 );
and ( n1331 , n1316 , n1330 );
and ( n1332 , n1301 , n1315 );
or ( n1333 , n1331 , n1332 );
xor ( n1334 , n1300 , n1333 );
xor ( n1335 , n1256 , n1273 );
xor ( n1336 , n1335 , n1285 );
and ( n1337 , n1334 , n1336 );
and ( n1338 , n1300 , n1333 );
or ( n1339 , n1337 , n1338 );
nor ( n1340 , n1299 , n1339 );
nor ( n1341 , n1297 , n1340 );
not ( n1342 , n1341 );
not ( n1343 , n858 );
not ( n1344 , n1328 );
or ( n1345 , n1343 , n1344 );
not ( n1346 , n501 );
not ( n1347 , n1279 );
or ( n1348 , n1346 , n1347 );
nand ( n1349 , n684 , n833 );
nand ( n1350 , n1348 , n1349 );
nand ( n1351 , n1350 , n831 );
nand ( n1352 , n1345 , n1351 );
not ( n1353 , n807 );
not ( n1354 , n499 );
not ( n1355 , n731 );
or ( n1356 , n1354 , n1355 );
nand ( n1357 , n738 , n782 );
nand ( n1358 , n1356 , n1357 );
not ( n1359 , n1358 );
or ( n1360 , n1353 , n1359 );
not ( n1361 , n499 );
nand ( n1362 , n1361 , n751 );
not ( n1363 , n1362 );
not ( n1364 , n782 );
nand ( n1365 , n1364 , n1250 );
not ( n1366 , n1365 );
or ( n1367 , n1363 , n1366 );
nand ( n1368 , n1367 , n770 );
nand ( n1369 , n1360 , n1368 );
xor ( n1370 , n1352 , n1369 );
not ( n1371 , n764 );
and ( n1372 , n811 , n1371 );
not ( n1373 , n500 );
not ( n1374 , n501 );
or ( n1375 , n1373 , n1374 );
nand ( n1376 , n1375 , n499 );
nor ( n1377 , n1372 , n1376 );
not ( n1378 , n946 );
and ( n1379 , n702 , n878 );
not ( n1380 , n702 );
and ( n1381 , n1380 , n503 );
or ( n1382 , n1379 , n1381 );
not ( n1383 , n1382 );
or ( n1384 , n1378 , n1383 );
nand ( n1385 , n1311 , n504 );
nand ( n1386 , n1384 , n1385 );
xor ( n1387 , n1377 , n1386 );
and ( n1388 , n1370 , n1387 );
and ( n1389 , n1352 , n1369 );
or ( n1390 , n1388 , n1389 );
not ( n1391 , n807 );
not ( n1392 , n1283 );
or ( n1393 , n1391 , n1392 );
nand ( n1394 , n1358 , n994 );
nand ( n1395 , n1393 , n1394 );
and ( n1396 , n1377 , n1386 );
xor ( n1397 , n1395 , n1396 );
xor ( n1398 , n1301 , n1315 );
xor ( n1399 , n1398 , n1330 );
xor ( n1400 , n1397 , n1399 );
nand ( n1401 , n1390 , n1400 );
not ( n1402 , n946 );
not ( n1403 , n503 );
not ( n1404 , n921 );
or ( n1405 , n1403 , n1404 );
nand ( n1406 , n684 , n878 );
nand ( n1407 , n1405 , n1406 );
not ( n1408 , n1407 );
or ( n1409 , n1402 , n1408 );
not ( n1410 , n690 );
not ( n1411 , n878 );
or ( n1412 , n1410 , n1411 );
nand ( n1413 , n1324 , n503 );
nand ( n1414 , n1412 , n1413 );
nand ( n1415 , n1414 , n504 );
nand ( n1416 , n1409 , n1415 );
not ( n1417 , n811 );
nand ( n1418 , n1417 , n819 );
and ( n1419 , n1418 , n503 );
not ( n1420 , n502 );
not ( n1421 , n751 );
or ( n1422 , n1420 , n1421 );
nand ( n1423 , n1422 , n501 );
nor ( n1424 , n1419 , n1423 );
xor ( n1425 , n1416 , n1424 );
not ( n1426 , n831 );
and ( n1427 , n833 , n755 );
not ( n1428 , n833 );
and ( n1429 , n1428 , n1088 );
or ( n1430 , n1427 , n1429 );
not ( n1431 , n1430 );
or ( n1432 , n1426 , n1431 );
not ( n1433 , n501 );
not ( n1434 , n929 );
or ( n1435 , n1433 , n1434 );
nand ( n1436 , n738 , n833 );
nand ( n1437 , n1435 , n1436 );
nand ( n1438 , n1437 , n858 );
nand ( n1439 , n1432 , n1438 );
or ( n1440 , n1425 , n1439 );
nand ( n1441 , n503 , n504 );
nor ( n1442 , n811 , n1441 );
not ( n1443 , n1442 );
and ( n1444 , n731 , n503 );
not ( n1445 , n731 );
and ( n1446 , n1445 , n878 );
or ( n1447 , n1444 , n1446 );
not ( n1448 , n1447 );
or ( n1449 , n1443 , n1448 );
nand ( n1450 , n811 , n858 );
nand ( n1451 , n1449 , n1450 );
and ( n1452 , n503 , n755 );
not ( n1453 , n503 );
and ( n1454 , n1453 , n752 );
nor ( n1455 , n1452 , n1454 );
and ( n1456 , n1455 , n946 );
or ( n1457 , n1451 , n1456 );
not ( n1458 , n946 );
not ( n1459 , n1447 );
or ( n1460 , n1458 , n1459 );
nand ( n1461 , n1407 , n504 );
nand ( n1462 , n1460 , n1461 );
nand ( n1463 , n1457 , n1462 );
nand ( n1466 , n1463 , C1 );
nand ( n1467 , n1440 , n1466 );
nand ( n1468 , n1439 , n1425 );
nand ( n1469 , n1467 , n1468 );
not ( n1470 , n1469 );
and ( n1471 , n1215 , n807 );
not ( n1472 , n501 );
not ( n1473 , n1279 );
or ( n1474 , n1472 , n1473 );
nand ( n1475 , n1474 , n1349 );
not ( n1476 , n1475 );
not ( n1477 , n882 );
or ( n1478 , n1476 , n1477 );
nand ( n1479 , n1437 , n831 );
nand ( n1480 , n1478 , n1479 );
xor ( n1481 , n1471 , n1480 );
not ( n1482 , n504 );
not ( n1483 , n1382 );
or ( n1484 , n1482 , n1483 );
nand ( n1485 , n1414 , n946 );
nand ( n1486 , n1484 , n1485 );
xor ( n1487 , n1481 , n1486 );
and ( n1488 , n1416 , n1424 );
nor ( n1489 , n1487 , n1488 );
or ( n1490 , n1470 , n1489 );
nand ( n1491 , n1487 , n1488 );
nand ( n1492 , n1490 , n1491 );
xor ( n1493 , n1352 , n1369 );
xor ( n1494 , n1493 , n1387 );
not ( n1495 , n1494 );
xor ( n1496 , n1471 , n1480 );
and ( n1497 , n1496 , n1486 );
and ( n1498 , n1471 , n1480 );
or ( n1499 , n1497 , n1498 );
not ( n1500 , n1499 );
nand ( n1501 , n1495 , n1500 );
nand ( n1502 , n1492 , n1501 );
nand ( n1503 , n1494 , n1499 );
nand ( n1504 , n1401 , n1502 , n1503 );
xor ( n1505 , n1300 , n1333 );
xor ( n1506 , n1505 , n1336 );
xor ( n1507 , n1395 , n1396 );
and ( n1508 , n1507 , n1399 );
and ( n1509 , n1395 , n1396 );
or ( n1510 , n1508 , n1509 );
nor ( n1511 , n1506 , n1510 );
nor ( n1512 , n1400 , n1390 );
nor ( n1513 , n1511 , n1512 );
nand ( n1514 , n1504 , n1513 );
buf ( n1515 , n1506 );
nand ( n1516 , n1515 , n1510 );
nand ( n1517 , n1299 , n1339 );
nand ( n1518 , n1514 , n1516 , n1517 );
not ( n1519 , n1518 );
or ( n1520 , n1342 , n1519 );
buf ( n1521 , n1246 );
nand ( n1522 , n1521 , n1296 );
nand ( n1523 , n1520 , n1522 );
not ( n1524 , n1523 );
or ( n1525 , n1244 , n1524 );
buf ( n1526 , n1178 );
nand ( n1527 , n1526 , n1241 );
nand ( n1528 , n1525 , n1527 );
buf ( n1529 , n1528 );
not ( n1530 , n1529 );
and ( n1531 , n1176 , n1530 );
not ( n1532 , n1176 );
and ( n1533 , n1532 , n1529 );
nor ( n1534 , n1531 , n1533 );
not ( n1535 , n1534 );
or ( n1536 , n717 , n1535 );
xor ( n1537 , n514 , n501 );
not ( n1538 , n1537 );
xor ( n1539 , n502 , n503 );
not ( n1540 , n1539 );
and ( n1541 , n502 , n501 );
not ( n1542 , n502 );
not ( n1543 , n501 );
and ( n1544 , n1542 , n1543 );
nor ( n1545 , n1541 , n1544 );
and ( n1546 , n1540 , n1545 );
not ( n1547 , n1546 );
or ( n1548 , n1538 , n1547 );
buf ( n1549 , n1539 );
xor ( n1550 , n513 , n501 );
nand ( n1551 , n1549 , n1550 );
nand ( n1552 , n1548 , n1551 );
not ( n1553 , n1552 );
not ( n1554 , n495 );
not ( n1555 , n1554 );
nand ( n1556 , n520 , n496 );
or ( n1557 , n520 , n496 );
nand ( n1558 , n1557 , n497 );
nand ( n1559 , n1555 , n1556 , n1558 );
nor ( n1560 , n1553 , n1559 );
xor ( n1561 , n494 , n495 );
and ( n1562 , n1561 , n520 );
xor ( n1563 , n498 , n499 );
xor ( n1564 , n517 , n497 );
xor ( n1565 , n498 , n497 );
nand ( n1566 , n1564 , n1565 );
or ( n1567 , n1563 , n1566 );
xor ( n1568 , n516 , n497 );
nand ( n1569 , n1563 , n1568 );
nand ( n1570 , n1567 , n1569 );
xor ( n1571 , n1562 , n1570 );
not ( n1572 , n1550 );
nand ( n1573 , n1540 , n1545 );
not ( n1574 , n1573 );
not ( n1575 , n1574 );
or ( n1576 , n1572 , n1575 );
xor ( n1577 , n512 , n501 );
nand ( n1578 , n1549 , n1577 );
nand ( n1579 , n1576 , n1578 );
xor ( n1580 , n1571 , n1579 );
xor ( n1581 , n1560 , n1580 );
xor ( n1582 , n520 , n495 );
not ( n1583 , n1582 );
xor ( n1584 , n495 , n496 );
and ( n1585 , n496 , n497 );
not ( n1586 , n496 );
not ( n1587 , n497 );
and ( n1588 , n1586 , n1587 );
nor ( n1589 , n1585 , n1588 );
not ( n1590 , n1589 );
nand ( n1591 , n1584 , n1590 );
not ( n1592 , n1591 );
not ( n1593 , n1592 );
or ( n1594 , n1583 , n1593 );
xor ( n1595 , n496 , n497 );
xor ( n1596 , n519 , n495 );
nand ( n1597 , n1595 , n1596 );
nand ( n1598 , n1594 , n1597 );
not ( n1599 , n1598 );
not ( n1600 , n504 );
nand ( n1601 , n1600 , n503 );
not ( n1602 , n1601 );
not ( n1603 , n1602 );
xor ( n1604 , n512 , n503 );
not ( n1605 , n1604 );
or ( n1606 , n1603 , n1605 );
xor ( n1607 , n511 , n503 );
nand ( n1608 , n1607 , n504 );
nand ( n1609 , n1606 , n1608 );
not ( n1610 , n1609 );
or ( n1611 , n1599 , n1610 );
nor ( n1612 , n1598 , n1609 );
not ( n1613 , n1563 );
xor ( n1614 , n518 , n497 );
nand ( n1615 , n1613 , n1565 , n1614 );
xor ( n1616 , n498 , n499 );
nand ( n1617 , n1616 , n1564 );
and ( n1618 , n1615 , n1617 );
or ( n1619 , n1612 , n1618 );
nand ( n1620 , n1611 , n1619 );
xor ( n1621 , n1581 , n1620 );
not ( n1622 , n1621 );
xor ( n1623 , n516 , n499 );
not ( n1624 , n1623 );
and ( n1625 , n501 , n805 );
not ( n1626 , n501 );
and ( n1627 , n1626 , n500 );
nor ( n1628 , n1625 , n1627 );
xor ( n1629 , n500 , n499 );
and ( n1630 , n1628 , n1629 );
not ( n1631 , n1630 );
or ( n1632 , n1624 , n1631 );
xor ( n1633 , n500 , n501 );
buf ( n1634 , n1633 );
xor ( n1635 , n515 , n499 );
nand ( n1636 , n1634 , n1635 );
nand ( n1637 , n1632 , n1636 );
not ( n1638 , n1637 );
xor ( n1639 , n1559 , n1552 );
nand ( n1640 , n1638 , n1639 );
not ( n1641 , n1640 );
and ( n1642 , n1595 , n520 );
xor ( n1643 , n513 , n503 );
not ( n1644 , n1643 );
not ( n1645 , n1602 );
or ( n1646 , n1644 , n1645 );
nand ( n1647 , n1604 , n504 );
nand ( n1648 , n1646 , n1647 );
xor ( n1649 , n1642 , n1648 );
and ( n1650 , n497 , n519 );
not ( n1651 , n497 );
not ( n1652 , n519 );
and ( n1653 , n1651 , n1652 );
nor ( n1654 , n1650 , n1653 );
not ( n1655 , n1654 );
not ( n1656 , n499 );
nand ( n1657 , n1656 , n498 );
not ( n1658 , n498 );
nand ( n1659 , n1658 , n499 );
and ( n1660 , n1657 , n1565 , n1659 );
not ( n1661 , n1660 );
or ( n1662 , n1655 , n1661 );
and ( n1663 , n498 , n499 );
not ( n1664 , n498 );
not ( n1665 , n499 );
and ( n1666 , n1664 , n1665 );
nor ( n1667 , n1663 , n1666 );
nand ( n1668 , n1667 , n1614 );
nand ( n1669 , n1662 , n1668 );
and ( n1670 , n1649 , n1669 );
and ( n1671 , n1642 , n1648 );
or ( n1672 , n1670 , n1671 );
not ( n1673 , n1672 );
or ( n1674 , n1641 , n1673 );
not ( n1675 , n1639 );
nand ( n1676 , n1675 , n1637 );
nand ( n1677 , n1674 , n1676 );
not ( n1678 , n1677 );
not ( n1679 , n1607 );
buf ( n1680 , n1602 );
not ( n1681 , n1680 );
or ( n1682 , n1679 , n1681 );
xor ( n1683 , n510 , n503 );
nand ( n1684 , n1683 , n504 );
nand ( n1685 , n1682 , n1684 );
not ( n1686 , n1596 );
not ( n1687 , n1591 );
not ( n1688 , n1687 );
or ( n1689 , n1686 , n1688 );
xor ( n1690 , n518 , n495 );
nand ( n1691 , n1595 , n1690 );
nand ( n1692 , n1689 , n1691 );
xor ( n1693 , n1685 , n1692 );
not ( n1694 , n1629 );
not ( n1695 , n1694 );
nand ( n1696 , n1635 , n1695 );
or ( n1697 , n1634 , n1696 );
xor ( n1698 , n499 , n514 );
nand ( n1699 , n1634 , n1698 );
nand ( n1700 , n1697 , n1699 );
buf ( n1701 , n1700 );
xor ( n1702 , n1693 , n1701 );
not ( n1703 , n1702 );
not ( n1704 , n1703 );
and ( n1705 , n1678 , n1704 );
and ( n1706 , n1677 , n1703 );
nor ( n1707 , n1705 , n1706 );
not ( n1708 , n1707 );
and ( n1709 , n1622 , n1708 );
and ( n1710 , n1621 , n1707 );
nor ( n1711 , n1709 , n1710 );
xor ( n1712 , n1637 , n1639 );
xor ( n1713 , n1712 , n1672 );
not ( n1714 , n1713 );
xor ( n1715 , n517 , n499 );
and ( n1716 , n1715 , n1695 );
not ( n1717 , n1716 );
not ( n1718 , n1634 );
not ( n1719 , n1718 );
or ( n1720 , n1717 , n1719 );
nand ( n1721 , n1634 , n1623 );
nand ( n1722 , n1720 , n1721 );
not ( n1723 , n1722 );
not ( n1724 , n1723 );
not ( n1725 , n1724 );
nand ( n1726 , n520 , n498 );
or ( n1727 , n520 , n498 );
nand ( n1728 , n1727 , n499 );
nand ( n1729 , n1726 , n1728 , n497 );
not ( n1730 , n1729 );
and ( n1731 , n514 , n503 );
not ( n1732 , n514 );
not ( n1733 , n503 );
and ( n1734 , n1732 , n1733 );
nor ( n1735 , n1731 , n1734 );
not ( n1736 , n1735 );
not ( n1737 , n1602 );
or ( n1738 , n1736 , n1737 );
nand ( n1739 , n1643 , n504 );
nand ( n1740 , n1738 , n1739 );
nand ( n1741 , n1730 , n1740 );
not ( n1742 , n1741 );
not ( n1743 , n1742 );
or ( n1744 , n1725 , n1743 );
not ( n1745 , n1723 );
not ( n1746 , n1741 );
or ( n1747 , n1745 , n1746 );
xor ( n1748 , n515 , n501 );
not ( n1749 , n1748 );
not ( n1750 , n1573 );
not ( n1751 , n1750 );
or ( n1752 , n1749 , n1751 );
nand ( n1753 , n1549 , n1537 );
nand ( n1754 , n1752 , n1753 );
nand ( n1755 , n1747 , n1754 );
nand ( n1756 , n1744 , n1755 );
not ( n1757 , n1756 );
and ( n1758 , n1618 , n1609 );
not ( n1759 , n1618 );
not ( n1760 , n1609 );
and ( n1761 , n1759 , n1760 );
nor ( n1762 , n1758 , n1761 );
and ( n1763 , n1762 , n1598 );
not ( n1764 , n1762 );
not ( n1765 , n1598 );
and ( n1766 , n1764 , n1765 );
nor ( n1767 , n1763 , n1766 );
nand ( n1768 , n1757 , n1767 );
and ( n1769 , n1714 , n1768 );
not ( n1770 , n1756 );
nor ( n1771 , n1770 , n1767 );
nor ( n1772 , n1769 , n1771 );
nand ( n1773 , n1711 , n1772 );
not ( n1774 , n1773 );
not ( n1775 , n1729 );
not ( n1776 , n1740 );
or ( n1777 , n1775 , n1776 );
or ( n1778 , n1740 , n1729 );
nand ( n1779 , n1777 , n1778 );
and ( n1780 , n1616 , n520 );
xor ( n1781 , n515 , n503 );
not ( n1782 , n1781 );
not ( n1783 , n1602 );
or ( n1784 , n1782 , n1783 );
nand ( n1785 , n1735 , n504 );
nand ( n1786 , n1784 , n1785 );
xor ( n1787 , n1780 , n1786 );
xor ( n1788 , n517 , n501 );
not ( n1789 , n1788 );
not ( n1790 , n1574 );
or ( n1791 , n1789 , n1790 );
xor ( n1792 , n516 , n501 );
nand ( n1793 , n1549 , n1792 );
nand ( n1794 , n1791 , n1793 );
and ( n1795 , n1787 , n1794 );
and ( n1796 , n1780 , n1786 );
or ( n1797 , n1795 , n1796 );
xor ( n1798 , n1779 , n1797 );
not ( n1799 , n1616 );
not ( n1800 , n1654 );
or ( n1801 , n1799 , n1800 );
xor ( n1802 , n497 , n520 );
nand ( n1803 , n1565 , n1799 , n1802 );
nand ( n1804 , n1801 , n1803 );
xor ( n1805 , n501 , n500 );
and ( n1806 , n518 , n499 );
not ( n1807 , n518 );
not ( n1808 , n499 );
and ( n1809 , n1807 , n1808 );
nor ( n1810 , n1806 , n1809 );
nand ( n1811 , n1629 , n1810 );
or ( n1812 , n1805 , n1811 );
nand ( n1813 , n1633 , n1715 );
nand ( n1814 , n1812 , n1813 );
xor ( n1815 , n1804 , n1814 );
not ( n1816 , n1792 );
not ( n1817 , n1546 );
or ( n1818 , n1816 , n1817 );
nand ( n1819 , n1549 , n1748 );
nand ( n1820 , n1818 , n1819 );
xor ( n1821 , n1815 , n1820 );
xor ( n1822 , n1798 , n1821 );
not ( n1823 , n1822 );
xor ( n1824 , n519 , n499 );
not ( n1825 , n1824 );
not ( n1826 , n1630 );
or ( n1827 , n1825 , n1826 );
nand ( n1828 , n1634 , n1810 );
nand ( n1829 , n1827 , n1828 );
or ( n1830 , n520 , n500 );
nand ( n1831 , n1830 , n501 );
nand ( n1832 , n520 , n500 );
and ( n1833 , n1831 , n1832 , n499 );
and ( n1834 , n503 , n516 );
not ( n1835 , n503 );
not ( n1836 , n516 );
and ( n1837 , n1835 , n1836 );
nor ( n1838 , n1834 , n1837 );
not ( n1839 , n1838 );
not ( n1840 , n1602 );
or ( n1841 , n1839 , n1840 );
nand ( n1842 , n1781 , n504 );
nand ( n1843 , n1841 , n1842 );
and ( n1844 , n1833 , n1843 );
xor ( n1845 , n1829 , n1844 );
xor ( n1846 , n1780 , n1786 );
xor ( n1847 , n1846 , n1794 );
and ( n1848 , n1845 , n1847 );
and ( n1849 , n1829 , n1844 );
or ( n1850 , n1848 , n1849 );
not ( n1851 , n1850 );
nand ( n1852 , n1823 , n1851 );
not ( n1853 , n1852 );
nand ( n1854 , n1822 , n1850 );
xor ( n1855 , n1829 , n1844 );
xor ( n1856 , n1855 , n1847 );
and ( n1857 , n1634 , n1824 );
not ( n1858 , n1634 );
xor ( n1859 , n520 , n499 );
and ( n1860 , n1695 , n1859 );
and ( n1861 , n1858 , n1860 );
or ( n1862 , n1857 , n1861 );
xor ( n1863 , n518 , n501 );
not ( n1864 , n1863 );
not ( n1865 , n1750 );
or ( n1866 , n1864 , n1865 );
buf ( n1867 , n1549 );
nand ( n1868 , n1867 , n1788 );
nand ( n1869 , n1866 , n1868 );
xor ( n1870 , n1862 , n1869 );
xor ( n1871 , n1833 , n1843 );
and ( n1872 , n1870 , n1871 );
and ( n1873 , n1862 , n1869 );
or ( n1874 , n1872 , n1873 );
nand ( n1875 , n1856 , n1874 );
nand ( n1876 , n1854 , n1875 );
not ( n1877 , n1876 );
or ( n1878 , n1853 , n1877 );
and ( n1879 , n1633 , n520 );
and ( n1880 , n503 , n517 );
not ( n1881 , n503 );
not ( n1882 , n517 );
and ( n1883 , n1881 , n1882 );
nor ( n1884 , n1880 , n1883 );
nand ( n1885 , n1884 , n1600 , n503 );
nand ( n1886 , n1838 , n504 );
nand ( n1887 , n1885 , n1886 );
xor ( n1888 , n1879 , n1887 );
not ( n1889 , n1549 );
xor ( n1890 , n519 , n501 );
nand ( n1891 , n1889 , n1890 , n1545 );
nand ( n1892 , n1549 , n1863 );
nand ( n1893 , n1891 , n1892 );
and ( n1894 , n1888 , n1893 );
and ( n1895 , n1879 , n1887 );
or ( n1896 , n1894 , n1895 );
xor ( n1897 , n1862 , n1869 );
xor ( n1898 , n1897 , n1871 );
xor ( n1899 , n1896 , n1898 );
or ( n1900 , n520 , n502 );
nand ( n1901 , n1900 , n503 );
nand ( n1902 , n520 , n502 );
and ( n1903 , n1901 , n1902 , n501 );
xor ( n1904 , n518 , n503 );
not ( n1905 , n1904 );
not ( n1906 , n1602 );
or ( n1907 , n1905 , n1906 );
nand ( n1908 , n1884 , n504 );
nand ( n1909 , n1907 , n1908 );
and ( n1910 , n1903 , n1909 );
xor ( n1911 , n1879 , n1887 );
xor ( n1912 , n1911 , n1893 );
xor ( n1913 , n1910 , n1912 );
xor ( n1914 , n1903 , n1909 );
xor ( n1915 , n520 , n501 );
not ( n1916 , n1915 );
not ( n1917 , n1750 );
or ( n1918 , n1916 , n1917 );
nand ( n1919 , n1867 , n1890 );
nand ( n1920 , n1918 , n1919 );
nor ( n1921 , n1914 , n1920 );
xor ( n1922 , n520 , n503 );
nand ( n1923 , n1680 , n1922 );
not ( n1924 , n1923 );
xor ( n1925 , n519 , n503 );
not ( n1926 , n1925 );
nor ( n1927 , n520 , n1441 );
not ( n1928 , n1927 );
or ( n1929 , n1926 , n1928 );
nand ( n1930 , n1549 , n520 );
nand ( n1931 , n1929 , n1930 );
not ( n1932 , n1931 );
not ( n1933 , n1932 );
or ( n1934 , n1924 , n1933 );
not ( n1935 , n1925 );
not ( n1936 , n1680 );
or ( n1937 , n1935 , n1936 );
nand ( n1938 , n1904 , n504 );
nand ( n1939 , n1937 , n1938 );
nand ( n1940 , n1934 , n1939 );
nand ( n1941 , n1940 , C1 );
not ( n1942 , n1941 );
or ( n1943 , n1921 , n1942 );
nand ( n1944 , n1914 , n1920 );
nand ( n1945 , n1943 , n1944 );
and ( n1946 , n1913 , n1945 );
and ( n1947 , n1910 , n1912 );
or ( n1948 , n1946 , n1947 );
and ( n1949 , n1899 , n1948 );
and ( n1950 , n1896 , n1898 );
or ( n1951 , n1949 , n1950 );
or ( n1952 , n1856 , n1874 );
nand ( n1953 , n1951 , n1852 , n1952 );
nand ( n1954 , n1878 , n1953 );
not ( n1955 , n1767 );
not ( n1956 , n1955 );
not ( n1957 , n1756 );
or ( n1958 , n1956 , n1957 );
not ( n1959 , n1756 );
nand ( n1960 , n1959 , n1767 );
nand ( n1961 , n1958 , n1960 );
and ( n1962 , n1961 , n1713 );
not ( n1963 , n1961 );
and ( n1964 , n1963 , n1714 );
nor ( n1965 , n1962 , n1964 );
not ( n1966 , n1965 );
xor ( n1967 , n1642 , n1648 );
xor ( n1968 , n1967 , n1669 );
xor ( n1969 , n1804 , n1814 );
and ( n1970 , n1969 , n1820 );
and ( n1971 , n1804 , n1814 );
or ( n1972 , n1970 , n1971 );
xor ( n1973 , n1968 , n1972 );
xor ( n1974 , n1722 , n1754 );
xnor ( n1975 , n1974 , n1741 );
and ( n1976 , n1973 , n1975 );
and ( n1977 , n1968 , n1972 );
or ( n1978 , n1976 , n1977 );
not ( n1979 , n1978 );
nand ( n1980 , n1966 , n1979 );
xor ( n1981 , n1968 , n1972 );
xor ( n1982 , n1981 , n1975 );
not ( n1983 , n1982 );
xor ( n1984 , n1779 , n1797 );
and ( n1985 , n1984 , n1821 );
and ( n1986 , n1779 , n1797 );
or ( n1987 , n1985 , n1986 );
not ( n1988 , n1987 );
nand ( n1989 , n1983 , n1988 );
nand ( n1990 , n1954 , n1980 , n1989 );
nand ( n1991 , n1965 , n1978 );
nand ( n1992 , n1982 , n1987 );
nand ( n1993 , n1991 , n1992 );
nand ( n1994 , n1980 , n1993 );
nand ( n1995 , n1990 , n1994 );
not ( n1996 , n1995 );
or ( n1997 , n1774 , n1996 );
not ( n1998 , n1711 );
not ( n1999 , n1772 );
nand ( n2000 , n1998 , n1999 );
nand ( n2001 , n1997 , n2000 );
not ( n2002 , n2001 );
or ( n2003 , n520 , n494 );
nand ( n2004 , n2003 , n495 );
nand ( n2005 , n520 , n494 );
nand ( n2006 , n2004 , n2005 , n493 );
not ( n2007 , n2006 );
not ( n2008 , n1577 );
not ( n2009 , n1750 );
or ( n2010 , n2008 , n2009 );
xor ( n2011 , n511 , n501 );
nand ( n2012 , n1867 , n2011 );
nand ( n2013 , n2010 , n2012 );
not ( n2014 , n2013 );
or ( n2015 , n2007 , n2014 );
or ( n2016 , n2013 , n2006 );
nand ( n2017 , n2015 , n2016 );
xor ( n2018 , n520 , n493 );
not ( n2019 , n2018 );
and ( n2020 , n494 , n493 );
not ( n2021 , n494 );
not ( n2022 , n493 );
and ( n2023 , n2021 , n2022 );
nor ( n2024 , n2020 , n2023 );
xor ( n2025 , n494 , n495 );
not ( n2026 , n2025 );
nand ( n2027 , n2024 , n2026 );
not ( n2028 , n2027 );
not ( n2029 , n2028 );
or ( n2030 , n2019 , n2029 );
xor ( n2031 , n494 , n495 );
xor ( n2032 , n519 , n493 );
nand ( n2033 , n2031 , n2032 );
nand ( n2034 , n2030 , n2033 );
not ( n2035 , n2034 );
not ( n2036 , n2035 );
not ( n2037 , n1698 );
not ( n2038 , n1630 );
or ( n2039 , n2037 , n2038 );
xor ( n2040 , n513 , n499 );
nand ( n2041 , n1634 , n2040 );
nand ( n2042 , n2039 , n2041 );
not ( n2043 , n2042 );
or ( n2044 , n2036 , n2043 );
or ( n2045 , n2042 , n2035 );
nand ( n2046 , n2044 , n2045 );
xor ( n2047 , n2017 , n2046 );
not ( n2048 , n1700 );
not ( n2049 , n1685 );
or ( n2050 , n2048 , n2049 );
or ( n2051 , n1685 , n1700 );
nand ( n2052 , n2051 , n1692 );
nand ( n2053 , n2050 , n2052 );
xor ( n2054 , n1562 , n1570 );
and ( n2055 , n2054 , n1579 );
and ( n2056 , n1562 , n1570 );
or ( n2057 , n2055 , n2056 );
and ( n2058 , n2053 , n2057 );
not ( n2059 , n2053 );
not ( n2060 , n2057 );
and ( n2061 , n2059 , n2060 );
or ( n2062 , n2058 , n2061 );
not ( n2063 , n1683 );
not ( n2064 , n1680 );
or ( n2065 , n2063 , n2064 );
and ( n2066 , n509 , n503 );
not ( n2067 , n509 );
not ( n2068 , n503 );
and ( n2069 , n2067 , n2068 );
nor ( n2070 , n2066 , n2069 );
nand ( n2071 , n2070 , n504 );
nand ( n2072 , n2065 , n2071 );
not ( n2073 , n1690 );
not ( n2074 , n1687 );
or ( n2075 , n2073 , n2074 );
xor ( n2076 , n517 , n495 );
nand ( n2077 , n1595 , n2076 );
nand ( n2078 , n2075 , n2077 );
xor ( n2079 , n2072 , n2078 );
not ( n2080 , n1568 );
or ( n2081 , n1665 , n498 );
nand ( n2082 , n2081 , n1657 , n1565 );
not ( n2083 , n2082 );
not ( n2084 , n2083 );
or ( n2085 , n2080 , n2084 );
xor ( n2086 , n498 , n499 );
xor ( n2087 , n497 , n515 );
nand ( n2088 , n2086 , n2087 );
nand ( n2089 , n2085 , n2088 );
xor ( n2090 , n2079 , n2089 );
not ( n2091 , n2090 );
and ( n2092 , n2062 , n2091 );
not ( n2093 , n2062 );
and ( n2094 , n2093 , n2090 );
nor ( n2095 , n2092 , n2094 );
xor ( n2096 , n2047 , n2095 );
xor ( n2097 , n1560 , n1580 );
and ( n2098 , n2097 , n1620 );
and ( n2099 , n1560 , n1580 );
or ( n2100 , n2098 , n2099 );
xor ( n2101 , n2096 , n2100 );
not ( n2102 , n1702 );
not ( n2103 , n1621 );
or ( n2104 , n2102 , n2103 );
not ( n2105 , n1703 );
not ( n2106 , n1621 );
not ( n2107 , n2106 );
or ( n2108 , n2105 , n2107 );
nand ( n2109 , n2108 , n1677 );
nand ( n2110 , n2104 , n2109 );
nand ( n2111 , n2101 , n2110 );
nor ( n2112 , n2101 , n2110 );
not ( n2113 , n2112 );
nand ( n2114 , n2111 , n2113 );
and ( n2115 , n2002 , n2114 );
not ( n2116 , n2002 );
not ( n2117 , n2114 );
and ( n2118 , n2116 , n2117 );
nor ( n2119 , n2115 , n2118 );
nand ( n2120 , n2119 , n455 );
nand ( n2121 , n1536 , n2120 );
buf ( n2122 , n2121 );
not ( n2123 , n543 );
nand ( n2124 , n2122 , n2123 );
not ( n2125 , n2122 );
nand ( n2126 , n2125 , n543 );
nand ( n2127 , n2124 , n2126 );
not ( n2128 , n2127 );
or ( n2129 , n715 , n2128 );
not ( n2130 , n716 );
not ( n2131 , n1174 );
not ( n2132 , n1528 );
or ( n2133 , n2131 , n2132 );
buf ( n2134 , n1175 );
nand ( n2135 , n2133 , n2134 );
not ( n2136 , n770 );
not ( n2137 , n800 );
or ( n2138 , n2136 , n2137 );
not ( n2139 , n499 );
not ( n2140 , n695 );
or ( n2141 , n2139 , n2140 );
nand ( n2142 , n696 , n782 );
nand ( n2143 , n2141 , n2142 );
nand ( n2144 , n2143 , n1122 );
nand ( n2145 , n2138 , n2144 );
nor ( n2146 , n861 , n817 );
xor ( n2147 , n2145 , n2146 );
xor ( n2148 , n1013 , n1028 );
and ( n2149 , n2148 , n1047 );
and ( n2150 , n1013 , n1028 );
or ( n2151 , n2149 , n2150 );
xor ( n2152 , n2147 , n2151 );
xor ( n2153 , n917 , n999 );
and ( n2154 , n2153 , n1048 );
and ( n2155 , n917 , n999 );
or ( n2156 , n2154 , n2155 );
xor ( n2157 , n2152 , n2156 );
not ( n2158 , n702 );
not ( n2159 , n813 );
or ( n2160 , n2158 , n2159 );
not ( n2161 , n495 );
or ( n2162 , n1130 , n2161 );
nand ( n2163 , n2160 , n2162 );
not ( n2164 , n2163 );
not ( n2165 , n1026 );
or ( n2166 , n2164 , n2165 );
nand ( n2167 , n1025 , n941 );
nand ( n2168 , n2166 , n2167 );
not ( n2169 , n946 );
not ( n2170 , n1045 );
or ( n2171 , n2169 , n2170 );
not ( n2172 , n503 );
and ( n2173 , n456 , n476 );
not ( n2174 , n456 );
and ( n2175 , n2174 , n460 );
nor ( n2176 , n2173 , n2175 );
not ( n2177 , n2176 );
not ( n2178 , n2177 );
not ( n2179 , n2178 );
or ( n2180 , n2172 , n2179 );
nand ( n2181 , n878 , n2177 );
nand ( n2182 , n2180 , n2181 );
nand ( n2183 , n2182 , n504 );
nand ( n2184 , n2171 , n2183 );
xor ( n2185 , n2168 , n2184 );
not ( n2186 , n760 );
not ( n2187 , n741 );
or ( n2188 , n2186 , n2187 );
nand ( n2189 , n684 , n739 );
not ( n2190 , n2189 );
not ( n2191 , n739 );
nand ( n2192 , n2191 , n1078 , n1079 );
not ( n2193 , n2192 );
or ( n2194 , n2190 , n2193 );
not ( n2195 , n758 );
not ( n2196 , n2195 );
nand ( n2197 , n2194 , n2196 );
nand ( n2198 , n2188 , n2197 );
xor ( n2199 , n2185 , n2198 );
xnor ( n2200 , n492 , n493 );
nor ( n2201 , n1088 , n2200 );
not ( n2202 , n1189 );
not ( n2203 , n853 );
or ( n2204 , n2202 , n2203 );
not ( n2205 , n501 );
not ( n2206 , n966 );
or ( n2207 , n2205 , n2206 );
and ( n2208 , n456 , n478 );
not ( n2209 , n456 );
and ( n2210 , n2209 , n462 );
or ( n2211 , n2208 , n2210 );
nand ( n2212 , n2211 , n833 );
nand ( n2213 , n2207 , n2212 );
nand ( n2214 , n2213 , n882 );
nand ( n2215 , n2204 , n2214 );
xor ( n2216 , n2201 , n2215 );
not ( n2217 , n912 );
not ( n2218 , n497 );
not ( n2219 , n1065 );
or ( n2220 , n2218 , n2219 );
nand ( n2221 , n1064 , n901 );
nand ( n2222 , n2220 , n2221 );
not ( n2223 , n2222 );
or ( n2224 , n2217 , n2223 );
nand ( n2225 , n893 , n1011 );
nand ( n2226 , n2224 , n2225 );
xor ( n2227 , n2216 , n2226 );
xor ( n2228 , n2199 , n2227 );
xor ( n2229 , n762 , n809 );
and ( n2230 , n2229 , n862 );
and ( n2231 , n762 , n809 );
or ( n2232 , n2230 , n2231 );
xor ( n2233 , n2228 , n2232 );
xor ( n2234 , n2157 , n2233 );
xor ( n2235 , n863 , n1049 );
and ( n2236 , n2235 , n1116 );
and ( n2237 , n863 , n1049 );
or ( n2238 , n2236 , n2237 );
nor ( n2239 , n2234 , n2238 );
not ( n2240 , n2239 );
buf ( n2241 , n2234 );
buf ( n2242 , n2238 );
nand ( n2243 , n2241 , n2242 );
nand ( n2244 , n2240 , n2243 );
not ( n2245 , n2244 );
and ( n2246 , n2135 , n2245 );
not ( n2247 , n2135 );
and ( n2248 , n2247 , n2244 );
nor ( n2249 , n2246 , n2248 );
not ( n2250 , n2249 );
or ( n2251 , n2130 , n2250 );
nand ( n2252 , n2001 , n2113 );
nand ( n2253 , n2252 , n2111 );
not ( n2254 , n2060 );
not ( n2255 , n2053 );
not ( n2256 , n2255 );
or ( n2257 , n2254 , n2256 );
nand ( n2258 , n2257 , n2090 );
not ( n2259 , n2255 );
nand ( n2260 , n2259 , n2057 );
nand ( n2261 , n2258 , n2260 );
not ( n2262 , n2040 );
not ( n2263 , n1630 );
or ( n2264 , n2262 , n2263 );
xor ( n2265 , n512 , n499 );
nand ( n2266 , n1634 , n2265 );
nand ( n2267 , n2264 , n2266 );
not ( n2268 , n2013 );
nor ( n2269 , n2268 , n2006 );
xor ( n2270 , n2267 , n2269 );
xor ( n2271 , n2072 , n2078 );
and ( n2272 , n2271 , n2089 );
and ( n2273 , n2072 , n2078 );
or ( n2274 , n2272 , n2273 );
xor ( n2275 , n2270 , n2274 );
xor ( n2276 , n2261 , n2275 );
xor ( n2277 , n492 , n493 );
not ( n2278 , n2277 );
not ( n2279 , n2278 );
and ( n2280 , n2279 , n520 );
xor ( n2281 , n514 , n497 );
and ( n2282 , n1563 , n2281 );
not ( n2283 , n1563 );
and ( n2284 , n1565 , n2087 );
and ( n2285 , n2283 , n2284 );
or ( n2286 , n2282 , n2285 );
xor ( n2287 , n2280 , n2286 );
not ( n2288 , n2011 );
not ( n2289 , n1574 );
or ( n2290 , n2288 , n2289 );
xor ( n2291 , n510 , n501 );
nand ( n2292 , n1549 , n2291 );
nand ( n2293 , n2290 , n2292 );
xor ( n2294 , n2287 , n2293 );
buf ( n2295 , n1589 );
not ( n2296 , n2295 );
and ( n2297 , n516 , n495 );
not ( n2298 , n516 );
and ( n2299 , n2298 , n719 );
nor ( n2300 , n2297 , n2299 );
not ( n2301 , n2300 );
not ( n2302 , n2301 );
or ( n2303 , n2296 , n2302 );
not ( n2304 , n1584 );
not ( n2305 , n2076 );
or ( n2306 , n2304 , n2305 );
not ( n2307 , n2295 );
nand ( n2308 , n2306 , n2307 );
nand ( n2309 , n2303 , n2308 );
not ( n2310 , n2070 );
not ( n2311 , n1602 );
or ( n2312 , n2310 , n2311 );
not ( n2313 , n508 );
not ( n2314 , n1733 );
or ( n2315 , n2313 , n2314 );
not ( n2316 , n508 );
nand ( n2317 , n2316 , n503 );
nand ( n2318 , n2315 , n2317 );
nand ( n2319 , n2318 , n504 );
nand ( n2320 , n2312 , n2319 );
xor ( n2321 , n2309 , n2320 );
not ( n2322 , n2032 );
not ( n2323 , n2028 );
or ( n2324 , n2322 , n2323 );
xor ( n2325 , n518 , n493 );
nand ( n2326 , n2031 , n2325 );
nand ( n2327 , n2324 , n2326 );
xor ( n2328 , n2321 , n2327 );
not ( n2329 , n2328 );
xor ( n2330 , n2294 , n2329 );
not ( n2331 , n2042 );
nand ( n2332 , n2331 , n2035 );
not ( n2333 , n2332 );
not ( n2334 , n2017 );
or ( n2335 , n2333 , n2334 );
nand ( n2336 , n2042 , n2034 );
nand ( n2337 , n2335 , n2336 );
xor ( n2338 , n2330 , n2337 );
xor ( n2339 , n2276 , n2338 );
xor ( n2340 , n2047 , n2095 );
and ( n2341 , n2340 , n2100 );
and ( n2342 , n2047 , n2095 );
or ( n2343 , n2341 , n2342 );
nand ( n2344 , n2339 , n2343 );
nor ( n2345 , n2339 , n2343 );
not ( n2346 , n2345 );
nand ( n2347 , n2344 , n2346 );
not ( n2348 , n2347 );
and ( n2349 , n2253 , n2348 );
not ( n2350 , n2253 );
and ( n2351 , n2350 , n2347 );
nor ( n2352 , n2349 , n2351 );
nand ( n2353 , n2352 , n455 );
nand ( n2354 , n2251 , n2353 );
buf ( n2355 , n2354 );
not ( n2356 , n2355 );
and ( n2357 , n2356 , n543 );
not ( n2358 , n2356 );
and ( n2359 , n2358 , n2123 );
or ( n2360 , n2357 , n2359 );
buf ( n2361 , n708 );
buf ( n2362 , n2361 );
nand ( n2363 , n2360 , n2362 );
nand ( n2364 , n2129 , n2363 );
not ( n2365 , n546 );
not ( n2366 , n2365 );
not ( n2367 , n547 );
and ( n2368 , n2366 , n2367 );
not ( n2369 , n547 );
nor ( n2370 , n2369 , n546 );
nor ( n2371 , n2368 , n2370 );
and ( n2372 , n546 , n545 );
nor ( n2373 , n545 , n546 );
nor ( n2374 , n2372 , n2373 );
and ( n2375 , n2371 , n2374 );
buf ( n2376 , n2375 );
not ( n2377 , n2376 );
not ( n2378 , n545 );
not ( n2379 , n455 );
xor ( n2380 , n2261 , n2275 );
and ( n2381 , n2380 , n2338 );
and ( n2382 , n2261 , n2275 );
or ( n2383 , n2381 , n2382 );
not ( n2384 , n2383 );
not ( n2385 , n504 );
xor ( n2386 , n507 , n503 );
not ( n2387 , n2386 );
or ( n2388 , n2385 , n2387 );
nand ( n2389 , n2318 , n1602 );
nand ( n2390 , n2388 , n2389 );
or ( n2391 , n520 , n492 );
nand ( n2392 , n2391 , n493 );
nand ( n2393 , n520 , n492 );
nand ( n2394 , n2392 , n2393 , n491 );
not ( n2395 , n2394 );
and ( n2396 , n2390 , n2395 );
not ( n2397 , n2390 );
and ( n2398 , n2397 , n2394 );
nor ( n2399 , n2396 , n2398 );
not ( n2400 , n2309 );
not ( n2401 , n2320 );
not ( n2402 , n2401 );
or ( n2403 , n2400 , n2402 );
nand ( n2404 , n2403 , n2327 );
not ( n2405 , n2309 );
nand ( n2406 , n2405 , n2320 );
nand ( n2407 , n2404 , n2406 );
xor ( n2408 , n2399 , n2407 );
xor ( n2409 , n2280 , n2286 );
and ( n2410 , n2409 , n2293 );
and ( n2411 , n2280 , n2286 );
or ( n2412 , n2410 , n2411 );
xor ( n2413 , n2408 , n2412 );
not ( n2414 , n2294 );
nand ( n2415 , n2414 , n2328 );
not ( n2416 , n2415 );
not ( n2417 , n2337 );
or ( n2418 , n2416 , n2417 );
nand ( n2419 , n2329 , n2294 );
nand ( n2420 , n2418 , n2419 );
and ( n2421 , n2413 , n2420 );
not ( n2422 , n2413 );
not ( n2423 , n2420 );
and ( n2424 , n2422 , n2423 );
nor ( n2425 , n2421 , n2424 );
not ( n2426 , n2291 );
not ( n2427 , n1574 );
or ( n2428 , n2426 , n2427 );
xor ( n2429 , n509 , n501 );
nand ( n2430 , n1549 , n2429 );
nand ( n2431 , n2428 , n2430 );
not ( n2432 , n2281 );
not ( n2433 , n1660 );
or ( n2434 , n2432 , n2433 );
xor ( n2435 , n513 , n497 );
nand ( n2436 , n1667 , n2435 );
nand ( n2437 , n2434 , n2436 );
xor ( n2438 , n2431 , n2437 );
not ( n2439 , n2300 );
not ( n2440 , n1592 );
or ( n2441 , n2439 , n2440 );
xor ( n2442 , n515 , n495 );
nand ( n2443 , n1595 , n2442 );
nand ( n2444 , n2441 , n2443 );
xnor ( n2445 , n2438 , n2444 );
xor ( n2446 , n520 , n491 );
not ( n2447 , n2446 );
not ( n2448 , n2277 );
and ( n2449 , n491 , n492 );
not ( n2450 , n491 );
not ( n2451 , n492 );
and ( n2452 , n2450 , n2451 );
nor ( n2453 , n2449 , n2452 );
nand ( n2454 , n2448 , n2453 );
not ( n2455 , n2454 );
not ( n2456 , n2455 );
or ( n2457 , n2447 , n2456 );
xor ( n2458 , n519 , n491 );
nand ( n2459 , n2458 , n2279 );
nand ( n2460 , n2457 , n2459 );
not ( n2461 , n1694 );
nand ( n2462 , n2461 , n2265 );
or ( n2463 , n1633 , n2462 );
and ( n2464 , n499 , n511 );
not ( n2465 , n499 );
not ( n2466 , n511 );
and ( n2467 , n2465 , n2466 );
nor ( n2468 , n2464 , n2467 );
nand ( n2469 , n2468 , n1633 );
nand ( n2470 , n2463 , n2469 );
not ( n2471 , n2470 );
xor ( n2472 , n2460 , n2471 );
not ( n2473 , n2031 );
not ( n2474 , n2473 );
not ( n2475 , n493 );
not ( n2476 , n722 );
or ( n2477 , n2475 , n2476 );
nand ( n2478 , n2022 , n494 );
nand ( n2479 , n2477 , n2478 );
and ( n2480 , n2479 , n2325 );
not ( n2481 , n2480 );
or ( n2482 , n2474 , n2481 );
xor ( n2483 , n517 , n493 );
nand ( n2484 , n2031 , n2483 );
nand ( n2485 , n2482 , n2484 );
xor ( n2486 , n2472 , n2485 );
not ( n2487 , n2486 );
and ( n2488 , n2445 , n2487 );
not ( n2489 , n2445 );
and ( n2490 , n2489 , n2486 );
nor ( n2491 , n2488 , n2490 );
xor ( n2492 , n2267 , n2269 );
and ( n2493 , n2492 , n2274 );
and ( n2494 , n2267 , n2269 );
or ( n2495 , n2493 , n2494 );
not ( n2496 , n2495 );
and ( n2497 , n2491 , n2496 );
not ( n2498 , n2491 );
and ( n2499 , n2498 , n2495 );
nor ( n2500 , n2497 , n2499 );
and ( n2501 , n2425 , n2500 );
not ( n2502 , n2425 );
not ( n2503 , n2500 );
and ( n2504 , n2502 , n2503 );
nor ( n2505 , n2501 , n2504 );
not ( n2506 , n2505 );
nand ( n2507 , n2384 , n2506 );
not ( n2508 , n2507 );
not ( n2509 , n2508 );
nand ( n2510 , n2505 , n2383 );
nand ( n2511 , n2509 , n2510 );
nor ( n2512 , n2345 , n2112 );
nand ( n2513 , n2001 , n2512 );
not ( n2514 , n2513 );
not ( n2515 , n2514 );
not ( n2516 , n2111 );
not ( n2517 , n2516 );
not ( n2518 , n2346 );
or ( n2519 , n2517 , n2518 );
nand ( n2520 , n2519 , n2344 );
not ( n2521 , n2520 );
nand ( n2522 , n2515 , n2521 );
not ( n2523 , n2522 );
and ( n2524 , n2511 , n2523 );
not ( n2525 , n2511 );
and ( n2526 , n2525 , n2522 );
nor ( n2527 , n2524 , n2526 );
not ( n2528 , n2527 );
or ( n2529 , n2379 , n2528 );
not ( n2530 , n2240 );
not ( n2531 , n2135 );
or ( n2532 , n2530 , n2531 );
nand ( n2533 , n2532 , n2243 );
or ( n2534 , n2451 , n739 );
nand ( n2535 , n2534 , n491 );
or ( n2536 , n2535 , n811 );
not ( n2537 , n492 );
nand ( n2538 , n2537 , n739 , n491 );
nand ( n2539 , n2536 , n2538 );
not ( n2540 , n946 );
not ( n2541 , n2182 );
or ( n2542 , n2540 , n2541 );
and ( n2543 , n456 , n475 );
not ( n2544 , n456 );
and ( n2545 , n2544 , n459 );
nor ( n2546 , n2543 , n2545 );
not ( n2547 , n2546 );
or ( n2548 , n2547 , n878 );
nand ( n2549 , n2547 , n878 );
nand ( n2550 , n2548 , n2549 );
nand ( n2551 , n2550 , n504 );
nand ( n2552 , n2542 , n2551 );
xor ( n2553 , n2539 , n2552 );
xor ( n2554 , n2201 , n2215 );
and ( n2555 , n2554 , n2226 );
and ( n2556 , n2201 , n2215 );
or ( n2557 , n2555 , n2556 );
xor ( n2558 , n2553 , n2557 );
xor ( n2559 , n2168 , n2184 );
and ( n2560 , n2559 , n2198 );
and ( n2561 , n2168 , n2184 );
or ( n2562 , n2560 , n2561 );
xor ( n2563 , n2558 , n2562 );
xor ( n2564 , n2199 , n2227 );
and ( n2565 , n2564 , n2232 );
and ( n2566 , n2199 , n2227 );
or ( n2567 , n2565 , n2566 );
xor ( n2568 , n2563 , n2567 );
not ( n2569 , n769 );
not ( n2570 , n2143 );
or ( n2571 , n2569 , n2570 );
not ( n2572 , n499 );
and ( n2573 , n456 , n479 );
not ( n2574 , n456 );
and ( n2575 , n2574 , n463 );
nor ( n2576 , n2573 , n2575 );
not ( n2577 , n2576 );
or ( n2578 , n2572 , n2577 );
nand ( n2579 , n851 , n782 );
nand ( n2580 , n2578 , n2579 );
nand ( n2581 , n2580 , n807 );
nand ( n2582 , n2571 , n2581 );
not ( n2583 , n2196 );
not ( n2584 , n493 );
not ( n2585 , n896 );
or ( n2586 , n2584 , n2585 );
not ( n2587 , n1324 );
nand ( n2588 , n2587 , n739 );
nand ( n2589 , n2586 , n2588 );
not ( n2590 , n2589 );
or ( n2591 , n2583 , n2590 );
not ( n2592 , n493 );
nor ( n2593 , n2592 , n495 , n494 );
not ( n2594 , n2593 );
not ( n2595 , n1279 );
or ( n2596 , n2594 , n2595 );
not ( n2597 , n495 );
not ( n2598 , n493 );
nand ( n2599 , n2598 , n494 );
nor ( n2600 , n2597 , n2599 );
nand ( n2601 , n684 , n2600 );
nand ( n2602 , n2596 , n2601 );
not ( n2603 , n2602 );
nand ( n2604 , n2591 , n2603 );
xor ( n2605 , n2582 , n2604 );
not ( n2606 , n2200 );
not ( n2607 , n2606 );
not ( n2608 , n491 );
not ( n2609 , n730 );
not ( n2610 , n2609 );
or ( n2611 , n2608 , n2610 );
not ( n2612 , n731 );
not ( n2613 , n491 );
nand ( n2614 , n2612 , n2613 );
nand ( n2615 , n2611 , n2614 );
not ( n2616 , n2615 );
or ( n2617 , n2607 , n2616 );
not ( n2618 , n491 );
not ( n2619 , n752 );
or ( n2620 , n2618 , n2619 );
nand ( n2621 , n755 , n2613 );
nand ( n2622 , n2620 , n2621 );
xor ( n2623 , n491 , n492 );
and ( n2624 , n2200 , n2623 );
nand ( n2625 , n2622 , n2624 );
nand ( n2626 , n2617 , n2625 );
xor ( n2627 , n2605 , n2626 );
not ( n2628 , n882 );
not ( n2629 , n501 );
and ( n2630 , n456 , n477 );
not ( n2631 , n456 );
and ( n2632 , n2631 , n461 );
nor ( n2633 , n2630 , n2632 );
not ( n2634 , n2633 );
or ( n2635 , n2629 , n2634 );
nand ( n2636 , n1036 , n833 );
nand ( n2637 , n2635 , n2636 );
not ( n2638 , n2637 );
or ( n2639 , n2628 , n2638 );
nand ( n2640 , n1189 , n2213 );
nand ( n2641 , n2639 , n2640 );
not ( n2642 , n893 );
not ( n2643 , n2222 );
or ( n2644 , n2642 , n2643 );
not ( n2645 , n497 );
not ( n2646 , n797 );
or ( n2647 , n2645 , n2646 );
or ( n2648 , n456 , n465 );
not ( n2649 , n481 );
nand ( n2650 , n2649 , n456 );
nand ( n2651 , n2648 , n2650 , n901 );
nand ( n2652 , n2647 , n2651 );
nand ( n2653 , n2652 , n912 );
nand ( n2654 , n2644 , n2653 );
xor ( n2655 , n2641 , n2654 );
not ( n2656 , n1026 );
not ( n2657 , n495 );
not ( n2658 , n989 );
not ( n2659 , n2658 );
or ( n2660 , n2657 , n2659 );
nand ( n2661 , n982 , n813 );
nand ( n2662 , n2660 , n2661 );
not ( n2663 , n2662 );
or ( n2664 , n2656 , n2663 );
nand ( n2665 , n2163 , n1086 );
nand ( n2666 , n2664 , n2665 );
xor ( n2667 , n2655 , n2666 );
xor ( n2668 , n2627 , n2667 );
xor ( n2669 , n2145 , n2146 );
and ( n2670 , n2669 , n2151 );
and ( n2671 , n2145 , n2146 );
or ( n2672 , n2670 , n2671 );
xor ( n2673 , n2668 , n2672 );
xor ( n2674 , n2568 , n2673 );
xor ( n2675 , n2152 , n2156 );
and ( n2676 , n2675 , n2233 );
and ( n2677 , n2152 , n2156 );
or ( n2678 , n2676 , n2677 );
nor ( n2679 , n2674 , n2678 );
not ( n2680 , n2679 );
nand ( n2681 , n2674 , n2678 );
buf ( n2682 , n2681 );
nand ( n2683 , n2680 , n2682 , n716 );
nor ( n2684 , n2533 , n2683 );
buf ( n2685 , n2240 );
and ( n2686 , n2135 , n2685 );
not ( n2687 , n2243 );
nor ( n2688 , n2686 , n2687 );
not ( n2689 , n2682 );
or ( n2690 , n2674 , n2678 );
not ( n2691 , n2690 );
or ( n2692 , n2689 , n2691 );
nand ( n2693 , n2692 , n716 );
nor ( n2694 , n2688 , n2693 );
nor ( n2695 , n2684 , n2694 );
nand ( n2696 , n2529 , n2695 );
buf ( n2697 , n2696 );
not ( n2698 , n2697 );
not ( n2699 , n2698 );
or ( n2700 , n2378 , n2699 );
not ( n2701 , n2697 );
not ( n2702 , n2701 );
nand ( n2703 , n2702 , n706 );
nand ( n2704 , n2700 , n2703 );
not ( n2705 , n2704 );
or ( n2706 , n2377 , n2705 );
not ( n2707 , n2346 );
nor ( n2708 , n2707 , n2508 );
not ( n2709 , n2708 );
not ( n2710 , n2252 );
not ( n2711 , n2710 );
or ( n2712 , n2709 , n2711 );
and ( n2713 , n2708 , n2516 );
or ( n2714 , n2508 , n2344 );
nand ( n2715 , n2714 , n2510 );
nor ( n2716 , n2713 , n2715 );
nand ( n2717 , n2712 , n2716 );
or ( n2718 , n2444 , n2431 );
nand ( n2719 , n2718 , n2437 );
nand ( n2720 , n2431 , n2444 );
nand ( n2721 , n2719 , n2720 );
not ( n2722 , n2485 );
not ( n2723 , n2470 );
or ( n2724 , n2722 , n2723 );
or ( n2725 , n2470 , n2485 );
nand ( n2726 , n2725 , n2460 );
nand ( n2727 , n2724 , n2726 );
and ( n2728 , n2721 , n2727 );
not ( n2729 , n2721 );
not ( n2730 , n2727 );
and ( n2731 , n2729 , n2730 );
nor ( n2732 , n2728 , n2731 );
xor ( n2733 , n490 , n491 );
nand ( n2734 , n2733 , n520 );
not ( n2735 , n2734 );
not ( n2736 , n1602 );
not ( n2737 , n2386 );
or ( n2738 , n2736 , n2737 );
and ( n2739 , n503 , n506 );
not ( n2740 , n503 );
not ( n2741 , n506 );
and ( n2742 , n2740 , n2741 );
nor ( n2743 , n2739 , n2742 );
nand ( n2744 , n2743 , n504 );
nand ( n2745 , n2738 , n2744 );
not ( n2746 , n2745 );
not ( n2747 , n2746 );
or ( n2748 , n2735 , n2747 );
not ( n2749 , n2734 );
nand ( n2750 , n2749 , n2745 );
nand ( n2751 , n2748 , n2750 );
not ( n2752 , n2429 );
not ( n2753 , n1750 );
or ( n2754 , n2752 , n2753 );
xor ( n2755 , n508 , n501 );
nand ( n2756 , n1867 , n2755 );
nand ( n2757 , n2754 , n2756 );
xor ( n2758 , n2751 , n2757 );
and ( n2759 , n2732 , n2758 );
not ( n2760 , n2732 );
not ( n2761 , n2758 );
and ( n2762 , n2760 , n2761 );
nor ( n2763 , n2759 , n2762 );
buf ( n2764 , n2277 );
xor ( n2765 , n518 , n491 );
not ( n2766 , n2765 );
and ( n2767 , n2764 , n2766 );
not ( n2768 , n2764 );
nand ( n2769 , n2458 , n2453 );
and ( n2770 , n2768 , n2769 );
nor ( n2771 , n2767 , n2770 );
not ( n2772 , n1561 );
nand ( n2773 , n2479 , n2483 );
and ( n2774 , n2772 , n2773 );
not ( n2775 , n2772 );
xor ( n2776 , n516 , n493 );
not ( n2777 , n2776 );
and ( n2778 , n2775 , n2777 );
nor ( n2779 , n2774 , n2778 );
and ( n2780 , n2771 , n2779 );
not ( n2781 , n2771 );
not ( n2782 , n2779 );
and ( n2783 , n2781 , n2782 );
nor ( n2784 , n2780 , n2783 );
nand ( n2785 , n2395 , n2390 );
and ( n2786 , n2784 , n2785 );
not ( n2787 , n2784 );
not ( n2788 , n2785 );
and ( n2789 , n2787 , n2788 );
nor ( n2790 , n2786 , n2789 );
and ( n2791 , n510 , n499 );
not ( n2792 , n510 );
and ( n2793 , n2792 , n1808 );
nor ( n2794 , n2791 , n2793 );
not ( n2795 , n2794 );
not ( n2796 , n1633 );
or ( n2797 , n2795 , n2796 );
nand ( n2798 , n1629 , n2468 , n1628 );
nand ( n2799 , n2797 , n2798 );
not ( n2800 , n2799 );
not ( n2801 , n1616 );
xor ( n2802 , n512 , n497 );
not ( n2803 , n2802 );
or ( n2804 , n2801 , n2803 );
not ( n2805 , n1667 );
nand ( n2806 , n2805 , n1565 , n2435 );
nand ( n2807 , n2804 , n2806 );
not ( n2808 , n2807 );
xor ( n2809 , n2800 , n2808 );
not ( n2810 , n2442 );
not ( n2811 , n1687 );
or ( n2812 , n2810 , n2811 );
xor ( n2813 , n514 , n495 );
nand ( n2814 , n1595 , n2813 );
nand ( n2815 , n2812 , n2814 );
xor ( n2816 , n2809 , n2815 );
xor ( n2817 , n2790 , n2816 );
xor ( n2818 , n2399 , n2407 );
and ( n2819 , n2818 , n2412 );
and ( n2820 , n2399 , n2407 );
or ( n2821 , n2819 , n2820 );
xor ( n2822 , n2817 , n2821 );
xor ( n2823 , n2763 , n2822 );
nand ( n2824 , n2445 , n2486 );
not ( n2825 , n2824 );
not ( n2826 , n2495 );
or ( n2827 , n2825 , n2826 );
not ( n2828 , n2445 );
nand ( n2829 , n2828 , n2487 );
nand ( n2830 , n2827 , n2829 );
xnor ( n2831 , n2823 , n2830 );
not ( n2832 , n2831 );
not ( n2833 , n2413 );
nand ( n2834 , n2833 , n2423 );
not ( n2835 , n2834 );
not ( n2836 , n2500 );
or ( n2837 , n2835 , n2836 );
not ( n2838 , n2423 );
nand ( n2839 , n2838 , n2413 );
nand ( n2840 , n2837 , n2839 );
nand ( n2841 , n2832 , n2840 );
not ( n2842 , n2832 );
not ( n2843 , n2840 );
nand ( n2844 , n2842 , n2843 );
nand ( n2845 , n2841 , n2844 );
not ( n2846 , n2845 );
and ( n2847 , n2717 , n2846 );
not ( n2848 , n2717 );
and ( n2849 , n2848 , n2845 );
nor ( n2850 , n2847 , n2849 );
or ( n2851 , n2850 , n716 );
nand ( n2852 , n2238 , n2234 );
nand ( n2853 , n2681 , n2852 , n1175 );
not ( n2854 , n2853 );
and ( n2855 , n2681 , n2239 );
nor ( n2856 , n2855 , n2679 );
not ( n2857 , n2856 );
or ( n2858 , n2854 , n2857 );
not ( n2859 , n2234 );
not ( n2860 , n2238 );
and ( n2861 , n2859 , n2860 );
nor ( n2862 , n1117 , n1172 );
nor ( n2863 , n2861 , n2862 );
not ( n2864 , n1243 );
not ( n2865 , n1523 );
or ( n2866 , n2864 , n2865 );
nand ( n2867 , n2866 , n1527 );
nand ( n2868 , n2863 , n2690 , n2867 );
nand ( n2869 , n2858 , n2868 );
not ( n2870 , n2869 );
not ( n2871 , n2870 );
xor ( n2872 , n2563 , n2567 );
and ( n2873 , n2872 , n2673 );
and ( n2874 , n2563 , n2567 );
or ( n2875 , n2873 , n2874 );
not ( n2876 , n2875 );
xor ( n2877 , n2641 , n2654 );
and ( n2878 , n2877 , n2666 );
and ( n2879 , n2641 , n2654 );
or ( n2880 , n2878 , n2879 );
xor ( n2881 , n2582 , n2604 );
and ( n2882 , n2881 , n2626 );
and ( n2883 , n2582 , n2604 );
or ( n2884 , n2882 , n2883 );
xor ( n2885 , n2880 , n2884 );
not ( n2886 , n490 );
not ( n2887 , n491 );
not ( n2888 , n2887 );
or ( n2889 , n2886 , n2888 );
not ( n2890 , n490 );
nand ( n2891 , n2890 , n491 );
nand ( n2892 , n2889 , n2891 );
and ( n2893 , n751 , n2892 );
not ( n2894 , n946 );
not ( n2895 , n2550 );
or ( n2896 , n2894 , n2895 );
not ( n2897 , n503 );
and ( n2898 , n456 , n474 );
not ( n2899 , n456 );
and ( n2900 , n2899 , n458 );
nor ( n2901 , n2898 , n2900 );
not ( n2902 , n2901 );
or ( n2903 , n2897 , n2902 );
or ( n2904 , n2901 , n503 );
nand ( n2905 , n2903 , n2904 );
nand ( n2906 , n2905 , n504 );
nand ( n2907 , n2896 , n2906 );
xor ( n2908 , n2893 , n2907 );
not ( n2909 , n858 );
and ( n2910 , n456 , n476 );
not ( n2911 , n456 );
and ( n2912 , n2911 , n460 );
nor ( n2913 , n2910 , n2912 );
not ( n2914 , n501 );
and ( n2915 , n2913 , n2914 );
not ( n2916 , n2913 );
and ( n2917 , n2916 , n501 );
nor ( n2918 , n2915 , n2917 );
not ( n2919 , n2918 );
or ( n2920 , n2909 , n2919 );
nand ( n2921 , n831 , n2637 );
nand ( n2922 , n2920 , n2921 );
xor ( n2923 , n2908 , n2922 );
xor ( n2924 , n2885 , n2923 );
not ( n2925 , n912 );
not ( n2926 , n497 );
not ( n2927 , n695 );
or ( n2928 , n2926 , n2927 );
nand ( n2929 , n696 , n901 );
nand ( n2930 , n2928 , n2929 );
not ( n2931 , n2930 );
or ( n2932 , n2925 , n2931 );
nand ( n2933 , n893 , n2652 );
nand ( n2934 , n2932 , n2933 );
not ( n2935 , n1086 );
not ( n2936 , n2662 );
or ( n2937 , n2935 , n2936 );
not ( n2938 , n495 );
not ( n2939 , n776 );
or ( n2940 , n2938 , n2939 );
nand ( n2941 , n777 , n813 );
nand ( n2942 , n2940 , n2941 );
nand ( n2943 , n2942 , n1026 );
nand ( n2944 , n2937 , n2943 );
xor ( n2945 , n2934 , n2944 );
not ( n2946 , n807 );
not ( n2947 , n499 );
not ( n2948 , n960 );
not ( n2949 , n2948 );
not ( n2950 , n2949 );
or ( n2951 , n2947 , n2950 );
nand ( n2952 , n2948 , n782 );
nand ( n2953 , n2951 , n2952 );
not ( n2954 , n2953 );
or ( n2955 , n2946 , n2954 );
nand ( n2956 , n994 , n2580 );
nand ( n2957 , n2955 , n2956 );
xor ( n2958 , n2945 , n2957 );
not ( n2959 , n2195 );
not ( n2960 , n2959 );
nand ( n2961 , n702 , n739 );
nand ( n2962 , n1263 , n493 );
nand ( n2963 , n2961 , n2962 );
not ( n2964 , n2963 );
or ( n2965 , n2960 , n2964 );
nor ( n2966 , n724 , n759 );
buf ( n2967 , n2966 );
nand ( n2968 , n2589 , n2967 );
nand ( n2969 , n2965 , n2968 );
not ( n2970 , n2606 );
not ( n2971 , n491 );
not ( n2972 , n684 );
not ( n2973 , n2972 );
or ( n2974 , n2971 , n2973 );
not ( n2975 , n2972 );
nand ( n2976 , n2975 , n2613 );
nand ( n2977 , n2974 , n2976 );
not ( n2978 , n2977 );
or ( n2979 , n2970 , n2978 );
nand ( n2980 , n2615 , n2624 );
nand ( n2981 , n2979 , n2980 );
xor ( n2982 , n2969 , n2981 );
and ( n2983 , n2539 , n2552 );
xor ( n2984 , n2982 , n2983 );
xor ( n2985 , n2958 , n2984 );
xor ( n2986 , n2553 , n2557 );
and ( n2987 , n2986 , n2562 );
and ( n2988 , n2553 , n2557 );
or ( n2989 , n2987 , n2988 );
xor ( n2990 , n2985 , n2989 );
xor ( n2991 , n2924 , n2990 );
xor ( n2992 , n2627 , n2667 );
and ( n2993 , n2992 , n2672 );
and ( n2994 , n2627 , n2667 );
or ( n2995 , n2993 , n2994 );
xor ( n2996 , n2991 , n2995 );
not ( n2997 , n2996 );
not ( n2998 , n2997 );
not ( n2999 , n2998 );
or ( n3000 , n2876 , n2999 );
not ( n3001 , n2875 );
nand ( n3002 , n2997 , n3001 );
nand ( n3003 , n3000 , n3002 );
nand ( n3004 , n3003 , n716 );
not ( n3005 , n3004 );
or ( n3006 , n2871 , n3005 );
or ( n3007 , n3003 , n455 );
nand ( n3008 , n3007 , n2869 );
nand ( n3009 , n3006 , n3008 );
nand ( n3010 , n2851 , n3009 );
not ( n3011 , n3010 );
not ( n3012 , n3011 );
and ( n3013 , n3012 , n545 );
not ( n3014 , n3012 );
and ( n3015 , n3014 , n706 );
or ( n3016 , n3013 , n3015 );
not ( n3017 , n2371 );
nand ( n3018 , n3016 , n3017 );
nand ( n3019 , n2706 , n3018 );
xor ( n3020 , n2364 , n3019 );
not ( n3021 , n540 );
or ( n3022 , n3021 , n541 );
not ( n3023 , n541 );
or ( n3024 , n3023 , n540 );
nand ( n3025 , n3022 , n3024 );
buf ( n3026 , n3025 );
not ( n3027 , n3026 );
not ( n3028 , n539 );
not ( n3029 , n1952 );
buf ( n3030 , n1951 );
not ( n3031 , n3030 );
or ( n3032 , n3029 , n3031 );
nand ( n3033 , n3032 , n1875 );
nand ( n3034 , n1852 , n1854 );
not ( n3035 , n3034 );
and ( n3036 , n3033 , n3035 );
not ( n3037 , n3033 );
and ( n3038 , n3037 , n3034 );
nor ( n3039 , n3036 , n3038 );
and ( n3040 , n3039 , n455 );
not ( n3041 , n1510 );
not ( n3042 , n1515 );
or ( n3043 , n3041 , n3042 );
not ( n3044 , n1511 );
nand ( n3045 , n3043 , n3044 );
not ( n3046 , n3045 );
not ( n3047 , n1512 );
not ( n3048 , n3047 );
not ( n3049 , n1501 );
not ( n3050 , n1492 );
or ( n3051 , n3049 , n3050 );
nand ( n3052 , n3051 , n1503 );
not ( n3053 , n3052 );
or ( n3054 , n3048 , n3053 );
nand ( n3055 , n1400 , n1390 );
nand ( n3056 , n3054 , n3055 );
not ( n3057 , n3056 );
not ( n3058 , n455 );
nand ( n3059 , n3046 , n3057 , n3058 );
nand ( n3060 , n3056 , n3045 , n3058 );
nand ( n3061 , n3059 , n3060 );
nor ( n3062 , n3040 , n3061 );
not ( n3063 , n3062 );
not ( n3064 , n3063 );
not ( n3065 , n3064 );
or ( n3066 , n3028 , n3065 );
not ( n3067 , n3063 );
not ( n3068 , n3067 );
not ( n3069 , n539 );
nand ( n3070 , n3068 , n3069 );
nand ( n3071 , n3066 , n3070 );
not ( n3072 , n3071 );
or ( n3073 , n3027 , n3072 );
not ( n3074 , n539 );
not ( n3075 , n3030 );
nand ( n3076 , n1875 , n1952 );
not ( n3077 , n3076 );
or ( n3078 , n3075 , n3077 );
or ( n3079 , n3076 , n3030 );
nand ( n3080 , n3078 , n3079 );
and ( n3081 , n455 , n3080 );
not ( n3082 , n455 );
not ( n3083 , n3052 );
nand ( n3084 , n3047 , n3055 );
and ( n3085 , n3083 , n3084 );
not ( n3086 , n3083 );
not ( n3087 , n3084 );
and ( n3088 , n3086 , n3087 );
nor ( n3089 , n3085 , n3088 );
and ( n3090 , n3082 , n3089 );
nor ( n3091 , n3081 , n3090 );
not ( n3092 , n3091 );
not ( n3093 , n3092 );
not ( n3094 , n3093 );
or ( n3095 , n3074 , n3094 );
not ( n3096 , n3093 );
nand ( n3097 , n3096 , n3069 );
nand ( n3098 , n3095 , n3097 );
and ( n3099 , n539 , n540 );
nor ( n3100 , n539 , n540 );
nor ( n3101 , n3099 , n3025 , n3100 );
not ( n3102 , n3101 );
not ( n3103 , n3102 );
nand ( n3104 , n3098 , n3103 );
nand ( n3105 , n3073 , n3104 );
not ( n3106 , n455 );
not ( n3107 , n1921 );
nand ( n3108 , n3107 , n1944 );
and ( n3109 , n3108 , n1942 );
not ( n3110 , n3108 );
and ( n3111 , n3110 , n1941 );
nor ( n3112 , n3109 , n3111 );
not ( n3113 , n3112 );
or ( n3114 , n3106 , n3113 );
not ( n3115 , n455 );
not ( n3116 , n1439 );
not ( n3117 , n1425 );
nand ( n3118 , n3116 , n3117 );
nand ( n3119 , n3118 , n1468 );
buf ( n3120 , n1466 );
not ( n3121 , n3120 );
and ( n3122 , n3119 , n3121 );
not ( n3123 , n3119 );
and ( n3124 , n3123 , n3120 );
nor ( n3125 , n3122 , n3124 );
nand ( n3126 , n3115 , n3125 );
nand ( n3127 , n3114 , n3126 );
buf ( n3128 , n3127 );
and ( n3129 , n3128 , n537 );
not ( n3130 , n538 );
or ( n3131 , n3130 , n539 );
or ( n3132 , n3069 , n538 );
nand ( n3133 , n3131 , n3132 );
buf ( n3134 , n3133 );
not ( n3135 , n3134 );
xor ( n3136 , n1896 , n1898 );
xor ( n3137 , n3136 , n1948 );
and ( n3138 , n455 , n3137 );
not ( n3139 , n455 );
or ( n3140 , n1494 , n1499 );
nand ( n3141 , n3140 , n1503 );
buf ( n3142 , n1492 );
not ( n3143 , n3142 );
and ( n3144 , n3141 , n3143 );
not ( n3145 , n3141 );
and ( n3146 , n3145 , n3142 );
nor ( n3147 , n3144 , n3146 );
and ( n3148 , n3139 , n3147 );
or ( n3149 , n3138 , n3148 );
xor ( n3150 , n537 , n3149 );
not ( n3151 , n3150 );
or ( n3152 , n3135 , n3151 );
not ( n3153 , n537 );
buf ( n3154 , n1470 );
not ( n3155 , n3154 );
not ( n3156 , n3155 );
not ( n3157 , n1488 );
not ( n3158 , n3157 );
not ( n3159 , n1487 );
not ( n3160 , n3159 );
or ( n3161 , n3158 , n3160 );
nand ( n3162 , n3161 , n1491 );
nor ( n3163 , n3162 , n455 );
not ( n3164 , n3163 );
or ( n3165 , n3156 , n3164 );
not ( n3166 , n455 );
and ( n3167 , n3162 , n3166 , n3154 );
xor ( n3168 , n1910 , n1912 );
xor ( n3169 , n3168 , n1945 );
nor ( n3170 , n3169 , n3166 );
nor ( n3171 , n3167 , n3170 );
nand ( n3172 , n3165 , n3171 );
buf ( n3173 , n3172 );
not ( n3174 , n3173 );
or ( n3175 , n3153 , n3174 );
not ( n3176 , n3173 );
not ( n3177 , n537 );
nand ( n3178 , n3176 , n3177 );
nand ( n3179 , n3175 , n3178 );
and ( n3180 , n3177 , n3130 );
and ( n3181 , n537 , n538 );
nor ( n3182 , n3180 , n3181 , n3133 );
nand ( n3183 , n3179 , n3182 );
nand ( n3184 , n3152 , n3183 );
xor ( n3185 , n3129 , n3184 );
buf ( n3186 , n3133 );
not ( n3187 , n3186 );
not ( n3188 , n3179 );
or ( n3189 , n3187 , n3188 );
not ( n3190 , n3127 );
nand ( n3191 , n3190 , n537 );
nand ( n3192 , n3177 , n3128 );
and ( n3193 , n3191 , n3192 );
not ( n3194 , n3182 );
nor ( n3195 , n3193 , n3194 );
not ( n3196 , n3195 );
nand ( n3197 , n3189 , n3196 );
not ( n3198 , n3197 );
not ( n3199 , n3190 );
and ( n3200 , n3199 , n538 );
nor ( n3201 , n3200 , n3177 );
not ( n3202 , n3130 );
not ( n3203 , n3128 );
not ( n3204 , n3203 );
or ( n3205 , n3202 , n3204 );
nand ( n3206 , n3205 , n539 );
nand ( n3207 , n3201 , n3206 );
nor ( n3208 , n3198 , n3207 );
xor ( n3209 , n3185 , n3208 );
xor ( n3210 , n3105 , n3209 );
or ( n3211 , n2123 , n542 );
not ( n3212 , n543 );
nand ( n3213 , n3212 , n542 );
nand ( n3214 , n3211 , n3213 );
not ( n3215 , n3214 );
not ( n3216 , n541 );
not ( n3217 , n1989 );
buf ( n3218 , n1954 );
not ( n3219 , n3218 );
or ( n3220 , n3217 , n3219 );
buf ( n3221 , n1991 );
buf ( n3222 , n1980 );
and ( n3223 , n3221 , n3222 );
not ( n3224 , n1992 );
nor ( n3225 , n3223 , n3224 );
nand ( n3226 , n3220 , n3225 );
nand ( n3227 , n3221 , n3222 , n1989 , n3218 );
and ( n3228 , n3222 , n3224 , n3221 );
not ( n3229 , n455 );
nor ( n3230 , n3228 , n3229 );
nand ( n3231 , n3226 , n3227 , n3230 );
nor ( n3232 , n1521 , n1296 );
not ( n3233 , n1522 );
nor ( n3234 , n3232 , n3233 );
not ( n3235 , n3234 );
and ( n3236 , n1516 , n1517 );
buf ( n3237 , n1514 );
and ( n3238 , n3236 , n3237 );
not ( n3239 , n1340 );
not ( n3240 , n3239 );
nor ( n3241 , n3238 , n3240 );
nand ( n3242 , n3235 , n3241 , n716 );
not ( n3243 , n455 );
not ( n3244 , n3232 );
not ( n3245 , n3241 );
not ( n3246 , n3233 );
nand ( n3247 , n3243 , n3244 , n3245 , n3246 );
nand ( n3248 , n3231 , n3242 , n3247 );
buf ( n3249 , n3248 );
not ( n3250 , n3249 );
not ( n3251 , n3250 );
or ( n3252 , n3216 , n3251 );
nand ( n3253 , n3249 , n3023 );
nand ( n3254 , n3252 , n3253 );
not ( n3255 , n3254 );
or ( n3256 , n3215 , n3255 );
not ( n3257 , n541 );
nand ( n3258 , n1992 , n1989 );
not ( n3259 , n3258 );
not ( n3260 , n3218 );
or ( n3261 , n3259 , n3260 );
or ( n3262 , n3258 , n3218 );
nand ( n3263 , n3261 , n3262 );
not ( n3264 , n3263 );
not ( n3265 , n455 );
or ( n3266 , n3264 , n3265 );
nand ( n3267 , n1515 , n1510 );
nand ( n3268 , n3237 , n3267 );
buf ( n3269 , n1299 );
nand ( n3270 , n3269 , n1339 );
nand ( n3271 , n3239 , n3270 );
and ( n3272 , n3271 , n716 );
and ( n3273 , n3268 , n3272 );
not ( n3274 , n3268 );
nor ( n3275 , n455 , n3271 );
and ( n3276 , n3274 , n3275 );
nor ( n3277 , n3273 , n3276 );
nand ( n3278 , n3266 , n3277 );
buf ( n3279 , n3278 );
not ( n3280 , n3279 );
not ( n3281 , n3280 );
or ( n3282 , n3257 , n3281 );
nand ( n3283 , n3279 , n3023 );
nand ( n3284 , n3282 , n3283 );
and ( n3285 , n541 , n542 );
nor ( n3286 , n541 , n542 );
nor ( n3287 , n3285 , n3214 , n3286 );
buf ( n3288 , n3287 );
nand ( n3289 , n3284 , n3288 );
nand ( n3290 , n3256 , n3289 );
and ( n3291 , n3210 , n3290 );
and ( n3292 , n3105 , n3209 );
or ( n3293 , n3291 , n3292 );
xor ( n3294 , n3020 , n3293 );
not ( n3295 , n548 );
and ( n3296 , n2369 , n3295 );
and ( n3297 , n547 , n548 );
xor ( n3298 , n548 , n549 );
nor ( n3299 , n3296 , n3297 , n3298 );
buf ( n3300 , n3299 );
not ( n3301 , n3300 );
not ( n3302 , n547 );
not ( n3303 , n2843 );
not ( n3304 , n2831 );
or ( n3305 , n3303 , n3304 );
not ( n3306 , n2510 );
nand ( n3307 , n3305 , n3306 );
nand ( n3308 , n3307 , n2841 );
not ( n3309 , n3308 );
or ( n3310 , n2514 , n2520 );
not ( n3311 , n2843 );
not ( n3312 , n2831 );
or ( n3313 , n3311 , n3312 );
nand ( n3314 , n3313 , n2507 );
not ( n3315 , n3314 );
nand ( n3316 , n3310 , n3315 );
nand ( n3317 , n3309 , n3316 );
not ( n3318 , n2830 );
not ( n3319 , n3318 );
not ( n3320 , n2763 );
or ( n3321 , n3319 , n3320 );
not ( n3322 , n2822 );
nand ( n3323 , n3321 , n3322 );
or ( n3324 , n3318 , n2763 );
nand ( n3325 , n3323 , n3324 );
not ( n3326 , n2799 );
not ( n3327 , n2807 );
or ( n3328 , n3326 , n3327 );
or ( n3329 , n2807 , n2799 );
nand ( n3330 , n3329 , n2815 );
nand ( n3331 , n3328 , n3330 );
not ( n3332 , n2776 );
not ( n3333 , n2028 );
or ( n3334 , n3332 , n3333 );
xor ( n3335 , n515 , n493 );
nand ( n3336 , n2031 , n3335 );
nand ( n3337 , n3334 , n3336 );
not ( n3338 , n2794 );
and ( n3339 , n1628 , n1629 );
not ( n3340 , n3339 );
or ( n3341 , n3338 , n3340 );
xor ( n3342 , n509 , n499 );
nand ( n3343 , n1634 , n3342 );
nand ( n3344 , n3341 , n3343 );
xor ( n3345 , n3337 , n3344 );
not ( n3346 , n2813 );
not ( n3347 , n1687 );
or ( n3348 , n3346 , n3347 );
xor ( n3349 , n513 , n495 );
nand ( n3350 , n1595 , n3349 );
nand ( n3351 , n3348 , n3350 );
xor ( n3352 , n3345 , n3351 );
xor ( n3353 , n3331 , n3352 );
not ( n3354 , n2802 );
not ( n3355 , n1660 );
or ( n3356 , n3354 , n3355 );
not ( n3357 , n2805 );
xor ( n3358 , n511 , n497 );
nand ( n3359 , n3357 , n3358 );
nand ( n3360 , n3356 , n3359 );
not ( n3361 , n2755 );
not ( n3362 , n1546 );
or ( n3363 , n3361 , n3362 );
xor ( n3364 , n507 , n501 );
nand ( n3365 , n1549 , n3364 );
nand ( n3366 , n3363 , n3365 );
xor ( n3367 , n3360 , n3366 );
xor ( n3368 , n490 , n491 );
xor ( n3369 , n519 , n489 );
and ( n3370 , n3368 , n3369 );
not ( n3371 , n3368 );
xor ( n3372 , n520 , n489 );
not ( n3373 , n3372 );
and ( n3374 , n489 , n490 );
not ( n3375 , n489 );
and ( n3376 , n3375 , n2890 );
nor ( n3377 , n3374 , n3376 );
not ( n3378 , n3377 );
nor ( n3379 , n3373 , n3378 );
and ( n3380 , n3371 , n3379 );
or ( n3381 , n3370 , n3380 );
xnor ( n3382 , n3367 , n3381 );
xnor ( n3383 , n3353 , n3382 );
not ( n3384 , n3383 );
not ( n3385 , n2771 );
not ( n3386 , n3385 );
not ( n3387 , n2785 );
or ( n3388 , n3386 , n3387 );
nand ( n3389 , n3388 , n2779 );
nand ( n3390 , n2771 , n2788 );
nand ( n3391 , n3389 , n3390 );
not ( n3392 , n2734 );
not ( n3393 , n2746 );
or ( n3394 , n3392 , n3393 );
nand ( n3395 , n3394 , n2757 );
nand ( n3396 , n3395 , n2750 );
not ( n3397 , n3396 );
not ( n3398 , n2743 );
not ( n3399 , n1602 );
or ( n3400 , n3398 , n3399 );
xor ( n3401 , n503 , n505 );
nand ( n3402 , n3401 , n504 );
nand ( n3403 , n3400 , n3402 );
not ( n3404 , n3403 );
nand ( n3405 , n520 , n490 );
or ( n3406 , n520 , n490 );
nand ( n3407 , n3406 , n491 );
nand ( n3408 , n3405 , n489 , n3407 );
not ( n3409 , n3408 );
and ( n3410 , n3404 , n3409 );
and ( n3411 , n3403 , n3408 );
nor ( n3412 , n3410 , n3411 );
not ( n3413 , n3412 );
not ( n3414 , n2765 );
not ( n3415 , n2455 );
or ( n3416 , n3414 , n3415 );
xor ( n3417 , n517 , n491 );
nand ( n3418 , n2764 , n3417 );
nand ( n3419 , n3416 , n3418 );
not ( n3420 , n3419 );
and ( n3421 , n3413 , n3420 );
and ( n3422 , n3412 , n3419 );
nor ( n3423 , n3421 , n3422 );
not ( n3424 , n3423 );
or ( n3425 , n3397 , n3424 );
or ( n3426 , n3396 , n3423 );
nand ( n3427 , n3425 , n3426 );
xor ( n3428 , n3391 , n3427 );
not ( n3429 , n2761 );
not ( n3430 , n2727 );
or ( n3431 , n3429 , n3430 );
not ( n3432 , n2730 );
not ( n3433 , n2758 );
or ( n3434 , n3432 , n3433 );
nand ( n3435 , n3434 , n2721 );
nand ( n3436 , n3431 , n3435 );
xor ( n3437 , n3428 , n3436 );
not ( n3438 , n3437 );
not ( n3439 , n3438 );
or ( n3440 , n3384 , n3439 );
not ( n3441 , n3383 );
nand ( n3442 , n3441 , n3437 );
nand ( n3443 , n3440 , n3442 );
not ( n3444 , n2790 );
or ( n3445 , n2821 , n3444 );
nand ( n3446 , n3445 , n2816 );
nand ( n3447 , n2821 , n3444 );
and ( n3448 , n3446 , n3447 );
not ( n3449 , n3448 );
and ( n3450 , n3443 , n3449 );
not ( n3451 , n3443 );
and ( n3452 , n3451 , n3448 );
nor ( n3453 , n3450 , n3452 );
nand ( n3454 , n3325 , n3453 );
not ( n3455 , n3453 );
not ( n3456 , n3325 );
nand ( n3457 , n3455 , n3456 );
nand ( n3458 , n3454 , n3457 );
xnor ( n3459 , n3317 , n3458 );
and ( n3460 , n455 , n3459 );
not ( n3461 , n455 );
not ( n3462 , n3002 );
not ( n3463 , n2853 );
not ( n3464 , n2856 );
or ( n3465 , n3463 , n3464 );
nand ( n3466 , n3465 , n2868 );
not ( n3467 , n3466 );
or ( n3468 , n3462 , n3467 );
nand ( n3469 , n2875 , n2998 );
nand ( n3470 , n3468 , n3469 );
xor ( n3471 , n2934 , n2944 );
and ( n3472 , n3471 , n2957 );
and ( n3473 , n2934 , n2944 );
or ( n3474 , n3472 , n3473 );
not ( n3475 , n1086 );
not ( n3476 , n2942 );
or ( n3477 , n3475 , n3476 );
and ( n3478 , n870 , n495 );
not ( n3479 , n870 );
and ( n3480 , n3479 , n813 );
or ( n3481 , n3478 , n3480 );
nand ( n3482 , n3481 , n918 );
nand ( n3483 , n3477 , n3482 );
not ( n3484 , n770 );
not ( n3485 , n2953 );
or ( n3486 , n3484 , n3485 );
not ( n3487 , n499 );
not ( n3488 , n1043 );
or ( n3489 , n3487 , n3488 );
nand ( n3490 , n1036 , n782 );
nand ( n3491 , n3489 , n3490 );
nand ( n3492 , n3491 , n1122 );
nand ( n3493 , n3486 , n3492 );
xor ( n3494 , n3483 , n3493 );
not ( n3495 , n2967 );
not ( n3496 , n2963 );
or ( n3497 , n3495 , n3496 );
not ( n3498 , n2658 );
nand ( n3499 , n3498 , n739 );
not ( n3500 , n3499 );
not ( n3501 , n982 );
nand ( n3502 , n3501 , n493 );
not ( n3503 , n3502 );
or ( n3504 , n3500 , n3503 );
nand ( n3505 , n3504 , n2959 );
nand ( n3506 , n3497 , n3505 );
xor ( n3507 , n3494 , n3506 );
xor ( n3508 , n3474 , n3507 );
not ( n3509 , n1189 );
not ( n3510 , n2918 );
or ( n3511 , n3509 , n3510 );
not ( n3512 , n833 );
not ( n3513 , n2547 );
or ( n3514 , n3512 , n3513 );
or ( n3515 , n2547 , n801 );
nand ( n3516 , n3514 , n3515 );
nand ( n3517 , n858 , n3516 );
nand ( n3518 , n3511 , n3517 );
nand ( n3519 , n490 , n491 );
or ( n3520 , n3519 , n489 );
nor ( n3521 , n490 , n491 );
nand ( n3522 , n3521 , n489 );
nand ( n3523 , n3520 , n3522 );
not ( n3524 , n3523 );
not ( n3525 , n489 );
not ( n3526 , n1250 );
or ( n3527 , n3525 , n3526 );
not ( n3528 , n489 );
nand ( n3529 , n3528 , n751 );
nand ( n3530 , n3527 , n3529 );
not ( n3531 , n3530 );
or ( n3532 , n3524 , n3531 );
nand ( n3533 , n728 , n729 , n489 );
not ( n3534 , n489 );
nand ( n3535 , n3534 , n738 );
nand ( n3536 , n3533 , n3535 );
nand ( n3537 , n3536 , n2892 );
nand ( n3538 , n3532 , n3537 );
xor ( n3539 , n3518 , n3538 );
not ( n3540 , n2930 );
not ( n3541 , n893 );
or ( n3542 , n3540 , n3541 );
not ( n3543 , n901 );
not ( n3544 , n951 );
or ( n3545 , n3543 , n3544 );
nand ( n3546 , n844 , n497 );
nand ( n3547 , n3545 , n3546 );
nand ( n3548 , n3547 , n912 );
nand ( n3549 , n3542 , n3548 );
xor ( n3550 , n3539 , n3549 );
xor ( n3551 , n3508 , n3550 );
xor ( n3552 , n2958 , n2984 );
and ( n3553 , n3552 , n2989 );
and ( n3554 , n2958 , n2984 );
or ( n3555 , n3553 , n3554 );
xor ( n3556 , n3551 , n3555 );
xor ( n3557 , n2969 , n2981 );
and ( n3558 , n3557 , n2983 );
and ( n3559 , n2969 , n2981 );
or ( n3560 , n3558 , n3559 );
not ( n3561 , n2606 );
and ( n3562 , n456 , n485 );
not ( n3563 , n456 );
and ( n3564 , n3563 , n469 );
nor ( n3565 , n3562 , n3564 );
and ( n3566 , n3565 , n491 );
not ( n3567 , n3565 );
and ( n3568 , n3567 , n2613 );
or ( n3569 , n3566 , n3568 );
not ( n3570 , n3569 );
or ( n3571 , n3561 , n3570 );
nand ( n3572 , n2200 , n2623 );
not ( n3573 , n3572 );
nand ( n3574 , n2977 , n3573 );
nand ( n3575 , n3571 , n3574 );
not ( n3576 , n3521 );
not ( n3577 , n3576 );
not ( n3578 , n1215 );
or ( n3579 , n3577 , n3578 );
and ( n3580 , n3519 , n489 );
nand ( n3581 , n3579 , n3580 );
not ( n3582 , n3581 );
not ( n3583 , n946 );
not ( n3584 , n2905 );
or ( n3585 , n3583 , n3584 );
not ( n3586 , n473 );
and ( n3587 , n456 , n3586 );
not ( n3588 , n456 );
not ( n3589 , n457 );
and ( n3590 , n3588 , n3589 );
nor ( n3591 , n3587 , n3590 );
not ( n3592 , n3591 );
and ( n3593 , n3592 , n2068 );
not ( n3594 , n3592 );
and ( n3595 , n3594 , n503 );
nor ( n3596 , n3593 , n3595 );
nand ( n3597 , n3596 , n504 );
nand ( n3598 , n3585 , n3597 );
xor ( n3599 , n3582 , n3598 );
xor ( n3600 , n3575 , n3599 );
xor ( n3601 , n2893 , n2907 );
and ( n3602 , n3601 , n2922 );
and ( n3603 , n2893 , n2907 );
or ( n3604 , n3602 , n3603 );
xor ( n3605 , n3600 , n3604 );
xor ( n3606 , n3560 , n3605 );
xor ( n3607 , n2880 , n2884 );
and ( n3608 , n3607 , n2923 );
and ( n3609 , n2880 , n2884 );
or ( n3610 , n3608 , n3609 );
xor ( n3611 , n3606 , n3610 );
xor ( n3612 , n3556 , n3611 );
buf ( n3613 , n3612 );
xor ( n3614 , n2924 , n2990 );
and ( n3615 , n3614 , n2995 );
and ( n3616 , n2924 , n2990 );
or ( n3617 , n3615 , n3616 );
and ( n3618 , n3613 , n3617 );
not ( n3619 , n3613 );
not ( n3620 , n3617 );
and ( n3621 , n3619 , n3620 );
or ( n3622 , n3618 , n3621 );
not ( n3623 , n3622 );
and ( n3624 , n3470 , n3623 );
not ( n3625 , n3470 );
and ( n3626 , n3625 , n3622 );
nor ( n3627 , n3624 , n3626 );
and ( n3628 , n3461 , n3627 );
nor ( n3629 , n3460 , n3628 );
not ( n3630 , n3629 );
buf ( n3631 , n3630 );
not ( n3632 , n3631 );
not ( n3633 , n3632 );
or ( n3634 , n3302 , n3633 );
nand ( n3635 , n3631 , n2369 );
nand ( n3636 , n3634 , n3635 );
not ( n3637 , n3636 );
or ( n3638 , n3301 , n3637 );
not ( n3639 , n547 );
not ( n3640 , n455 );
nor ( n3641 , n3325 , n3453 );
nor ( n3642 , n3641 , n3314 );
not ( n3643 , n3642 );
not ( n3644 , n2522 );
or ( n3645 , n3643 , n3644 );
and ( n3646 , n3308 , n3457 );
not ( n3647 , n3454 );
nor ( n3648 , n3646 , n3647 );
nand ( n3649 , n3645 , n3648 );
not ( n3650 , n3419 );
nand ( n3651 , n3650 , n3412 );
not ( n3652 , n3651 );
not ( n3653 , n3396 );
or ( n3654 , n3652 , n3653 );
not ( n3655 , n3412 );
nand ( n3656 , n3655 , n3419 );
nand ( n3657 , n3654 , n3656 );
not ( n3658 , n3657 );
not ( n3659 , n3408 );
and ( n3660 , n3659 , n3403 );
or ( n3661 , n3366 , n3381 );
nand ( n3662 , n3661 , n3360 );
nand ( n3663 , n3366 , n3381 );
nand ( n3664 , n3662 , n3663 );
xor ( n3665 , n3660 , n3664 );
not ( n3666 , n3351 );
not ( n3667 , n3344 );
or ( n3668 , n3666 , n3667 );
or ( n3669 , n3344 , n3351 );
nand ( n3670 , n3669 , n3337 );
nand ( n3671 , n3668 , n3670 );
xnor ( n3672 , n3665 , n3671 );
xor ( n3673 , n3658 , n3672 );
not ( n3674 , n3352 );
not ( n3675 , n3331 );
nand ( n3676 , n3675 , n3382 );
not ( n3677 , n3676 );
or ( n3678 , n3674 , n3677 );
not ( n3679 , n3382 );
nand ( n3680 , n3679 , n3331 );
nand ( n3681 , n3678 , n3680 );
xnor ( n3682 , n3673 , n3681 );
not ( n3683 , n3401 );
not ( n3684 , n1602 );
or ( n3685 , n3683 , n3684 );
nand ( n3686 , n3685 , n1441 );
not ( n3687 , n3686 );
nand ( n3688 , n520 , n489 );
not ( n3689 , n3688 );
and ( n3690 , n3687 , n3689 );
and ( n3691 , n3686 , n3688 );
nor ( n3692 , n3690 , n3691 );
not ( n3693 , n3364 );
not ( n3694 , n1574 );
or ( n3695 , n3693 , n3694 );
xor ( n3696 , n506 , n501 );
nand ( n3697 , n1867 , n3696 );
nand ( n3698 , n3695 , n3697 );
buf ( n3699 , n3698 );
xor ( n3700 , n3692 , n3699 );
not ( n3701 , n3700 );
not ( n3702 , n3342 );
not ( n3703 , n3339 );
or ( n3704 , n3702 , n3703 );
xor ( n3705 , n508 , n499 );
nand ( n3706 , n1634 , n3705 );
nand ( n3707 , n3704 , n3706 );
not ( n3708 , n3417 );
not ( n3709 , n2455 );
or ( n3710 , n3708 , n3709 );
not ( n3711 , n2277 );
not ( n3712 , n3711 );
xor ( n3713 , n516 , n491 );
nand ( n3714 , n3712 , n3713 );
nand ( n3715 , n3710 , n3714 );
xor ( n3716 , n3707 , n3715 );
not ( n3717 , n3335 );
not ( n3718 , n2028 );
or ( n3719 , n3717 , n3718 );
xor ( n3720 , n493 , n514 );
nand ( n3721 , n2031 , n3720 );
nand ( n3722 , n3719 , n3721 );
not ( n3723 , n3722 );
and ( n3724 , n3716 , n3723 );
not ( n3725 , n3716 );
not ( n3726 , n3723 );
and ( n3727 , n3725 , n3726 );
nor ( n3728 , n3724 , n3727 );
not ( n3729 , n3728 );
or ( n3730 , n3701 , n3729 );
or ( n3731 , n3700 , n3728 );
nand ( n3732 , n3730 , n3731 );
not ( n3733 , n3369 );
nor ( n3734 , n3378 , n3368 );
not ( n3735 , n3734 );
or ( n3736 , n3733 , n3735 );
xor ( n3737 , n489 , n518 );
nand ( n3738 , n2733 , n3737 );
nand ( n3739 , n3736 , n3738 );
not ( n3740 , n3349 );
not ( n3741 , n1687 );
or ( n3742 , n3740 , n3741 );
xor ( n3743 , n512 , n495 );
nand ( n3744 , n1595 , n3743 );
nand ( n3745 , n3742 , n3744 );
xor ( n3746 , n3739 , n3745 );
not ( n3747 , n3358 );
not ( n3748 , n2083 );
or ( n3749 , n3747 , n3748 );
xor ( n3750 , n510 , n497 );
nand ( n3751 , n2086 , n3750 );
nand ( n3752 , n3749 , n3751 );
xnor ( n3753 , n3746 , n3752 );
not ( n3754 , n3753 );
and ( n3755 , n3732 , n3754 );
not ( n3756 , n3732 );
and ( n3757 , n3756 , n3753 );
nor ( n3758 , n3755 , n3757 );
not ( n3759 , n3758 );
xor ( n3760 , n3391 , n3427 );
and ( n3761 , n3760 , n3436 );
and ( n3762 , n3391 , n3427 );
or ( n3763 , n3761 , n3762 );
not ( n3764 , n3763 );
or ( n3765 , n3759 , n3764 );
or ( n3766 , n3763 , n3758 );
nand ( n3767 , n3765 , n3766 );
not ( n3768 , n3767 );
and ( n3769 , n3682 , n3768 );
not ( n3770 , n3682 );
and ( n3771 , n3770 , n3767 );
nor ( n3772 , n3769 , n3771 );
not ( n3773 , n3449 );
not ( n3774 , n3383 );
or ( n3775 , n3773 , n3774 );
not ( n3776 , n3441 );
not ( n3777 , n3448 );
or ( n3778 , n3776 , n3777 );
buf ( n3779 , n3437 );
nand ( n3780 , n3778 , n3779 );
nand ( n3781 , n3775 , n3780 );
nand ( n3782 , n3772 , n3781 );
not ( n3783 , n3772 );
not ( n3784 , n3781 );
nand ( n3785 , n3783 , n3784 );
nand ( n3786 , n3782 , n3785 );
xnor ( n3787 , n3649 , n3786 );
not ( n3788 , n3787 );
or ( n3789 , n3640 , n3788 );
not ( n3790 , n3617 );
not ( n3791 , n3612 );
and ( n3792 , n3790 , n3791 );
and ( n3793 , n2997 , n3001 );
nor ( n3794 , n3792 , n3793 );
not ( n3795 , n3794 );
not ( n3796 , n3466 );
or ( n3797 , n3795 , n3796 );
nand ( n3798 , n2996 , n2875 );
not ( n3799 , n3798 );
nand ( n3800 , n3617 , n3612 );
not ( n3801 , n3800 );
or ( n3802 , n3799 , n3801 );
not ( n3803 , n3612 );
nand ( n3804 , n3803 , n3620 );
nand ( n3805 , n3802 , n3804 );
buf ( n3806 , n3805 );
nand ( n3807 , n3797 , n3806 );
not ( n3808 , n807 );
and ( n3809 , n2177 , n782 );
not ( n3810 , n2177 );
and ( n3811 , n3810 , n499 );
or ( n3812 , n3809 , n3811 );
not ( n3813 , n3812 );
or ( n3814 , n3808 , n3813 );
nand ( n3815 , n769 , n3491 );
nand ( n3816 , n3814 , n3815 );
not ( n3817 , n2196 );
not ( n3818 , n493 );
not ( n3819 , n776 );
or ( n3820 , n3818 , n3819 );
nand ( n3821 , n739 , n1064 );
nand ( n3822 , n3820 , n3821 );
not ( n3823 , n3822 );
or ( n3824 , n3817 , n3823 );
not ( n3825 , n2599 );
nand ( n3826 , n3825 , n495 );
and ( n3827 , n989 , n3826 );
not ( n3828 , n989 );
not ( n3829 , n2593 );
and ( n3830 , n3828 , n3829 );
or ( n3831 , n3827 , n3830 );
nand ( n3832 , n3824 , n3831 );
xor ( n3833 , n3816 , n3832 );
not ( n3834 , n2624 );
not ( n3835 , n3569 );
or ( n3836 , n3834 , n3835 );
not ( n3837 , n2200 );
or ( n3838 , n1130 , n2887 );
nand ( n3839 , n1130 , n2613 );
nand ( n3840 , n3838 , n3839 );
nand ( n3841 , n3837 , n3840 );
nand ( n3842 , n3836 , n3841 );
xor ( n3843 , n3833 , n3842 );
and ( n3844 , n1215 , n489 );
not ( n3845 , n946 );
not ( n3846 , n3596 );
or ( n3847 , n3845 , n3846 );
nand ( n3848 , n3847 , n1441 );
xor ( n3849 , n3844 , n3848 );
not ( n3850 , n831 );
not ( n3851 , n3516 );
or ( n3852 , n3850 , n3851 );
not ( n3853 , n501 );
and ( n3854 , n456 , n474 );
not ( n3855 , n456 );
and ( n3856 , n3855 , n458 );
nor ( n3857 , n3854 , n3856 );
not ( n3858 , n3857 );
not ( n3859 , n3858 );
not ( n3860 , n3859 );
or ( n3861 , n3853 , n3860 );
nand ( n3862 , n3858 , n833 );
nand ( n3863 , n3861 , n3862 );
nand ( n3864 , n3863 , n858 );
nand ( n3865 , n3852 , n3864 );
xor ( n3866 , n3849 , n3865 );
xor ( n3867 , n3843 , n3866 );
not ( n3868 , n3523 );
not ( n3869 , n3536 );
or ( n3870 , n3868 , n3869 );
xor ( n3871 , n489 , n684 );
nand ( n3872 , n2892 , n3871 );
nand ( n3873 , n3870 , n3872 );
not ( n3874 , n893 );
not ( n3875 , n3547 );
or ( n3876 , n3874 , n3875 );
not ( n3877 , n497 );
not ( n3878 , n966 );
or ( n3879 , n3877 , n3878 );
nand ( n3880 , n2948 , n901 );
nand ( n3881 , n3879 , n3880 );
nand ( n3882 , n912 , n3881 );
nand ( n3883 , n3876 , n3882 );
xor ( n3884 , n3873 , n3883 );
not ( n3885 , n1086 );
not ( n3886 , n3481 );
or ( n3887 , n3885 , n3886 );
not ( n3888 , n495 );
and ( n3889 , n456 , n480 );
not ( n3890 , n456 );
and ( n3891 , n3890 , n464 );
nor ( n3892 , n3889 , n3891 );
not ( n3893 , n3892 );
or ( n3894 , n3888 , n3893 );
nand ( n3895 , n696 , n813 );
nand ( n3896 , n3894 , n3895 );
nand ( n3897 , n3896 , n1026 );
nand ( n3898 , n3887 , n3897 );
xor ( n3899 , n3884 , n3898 );
xor ( n3900 , n3867 , n3899 );
xor ( n3901 , n3560 , n3605 );
and ( n3902 , n3901 , n3610 );
and ( n3903 , n3560 , n3605 );
or ( n3904 , n3902 , n3903 );
xor ( n3905 , n3900 , n3904 );
xor ( n3906 , n3575 , n3599 );
and ( n3907 , n3906 , n3604 );
and ( n3908 , n3575 , n3599 );
or ( n3909 , n3907 , n3908 );
and ( n3910 , n3598 , n3582 );
xor ( n3911 , n3518 , n3538 );
and ( n3912 , n3911 , n3549 );
and ( n3913 , n3518 , n3538 );
or ( n3914 , n3912 , n3913 );
xor ( n3915 , n3910 , n3914 );
xor ( n3916 , n3483 , n3493 );
and ( n3917 , n3916 , n3506 );
and ( n3918 , n3483 , n3493 );
or ( n3919 , n3917 , n3918 );
xor ( n3920 , n3915 , n3919 );
xor ( n3921 , n3909 , n3920 );
xor ( n3922 , n3474 , n3507 );
and ( n3923 , n3922 , n3550 );
and ( n3924 , n3474 , n3507 );
or ( n3925 , n3923 , n3924 );
xor ( n3926 , n3921 , n3925 );
xor ( n3927 , n3905 , n3926 );
xor ( n3928 , n3551 , n3555 );
and ( n3929 , n3928 , n3611 );
and ( n3930 , n3551 , n3555 );
or ( n3931 , n3929 , n3930 );
or ( n3932 , n3927 , n3931 );
nand ( n3933 , n3927 , n3931 );
nand ( n3934 , n3932 , n3933 );
not ( n3935 , n3934 );
and ( n3936 , n3807 , n3935 );
not ( n3937 , n3807 );
and ( n3938 , n3937 , n3934 );
nor ( n3939 , n3936 , n3938 );
not ( n3940 , n455 );
nand ( n3941 , n3939 , n3940 );
nand ( n3942 , n3789 , n3941 );
not ( n3943 , n3942 );
not ( n3944 , n3943 );
or ( n3945 , n3639 , n3944 );
not ( n3946 , n3943 );
nand ( n3947 , n3946 , n2369 );
nand ( n3948 , n3945 , n3947 );
nand ( n3949 , n3948 , n3298 );
nand ( n3950 , n3638 , n3949 );
xor ( n3951 , n3129 , n3184 );
and ( n3952 , n3951 , n3208 );
and ( n3953 , n3129 , n3184 );
or ( n3954 , n3952 , n3953 );
buf ( n3955 , n3214 );
not ( n3956 , n3955 );
not ( n3957 , n1242 );
not ( n3958 , n1526 );
or ( n3959 , n3957 , n3958 );
or ( n3960 , n1526 , n1242 );
nand ( n3961 , n3959 , n3960 );
buf ( n3962 , n1523 );
and ( n3963 , n3961 , n3962 );
nor ( n3964 , n3963 , n455 );
not ( n3965 , n3964 );
not ( n3966 , n3962 );
not ( n3967 , n3961 );
nand ( n3968 , n3966 , n3967 );
not ( n3969 , n3968 );
or ( n3970 , n3965 , n3969 );
nand ( n3971 , n2000 , n1773 );
and ( n3972 , n3971 , n455 );
buf ( n3973 , n1995 );
buf ( n3974 , n3973 );
and ( n3975 , n3972 , n3974 );
not ( n3976 , n455 );
nor ( n3977 , n3976 , n3971 , n3973 );
nor ( n3978 , n3975 , n3977 );
nand ( n3979 , n3970 , n3978 );
buf ( n3980 , n3979 );
buf ( n3981 , n3980 );
and ( n3982 , n3981 , n3023 );
not ( n3983 , n3981 );
and ( n3984 , n3983 , n541 );
or ( n3985 , n3982 , n3984 );
not ( n3986 , n3985 );
or ( n3987 , n3956 , n3986 );
nand ( n3988 , n3254 , n3288 );
nand ( n3989 , n3987 , n3988 );
xor ( n3990 , n3954 , n3989 );
nor ( n3991 , n3173 , n3177 );
not ( n3992 , n3134 );
xor ( n3993 , n537 , n3096 );
not ( n3994 , n3993 );
or ( n3995 , n3992 , n3994 );
nand ( n3996 , n3150 , n3182 );
nand ( n3997 , n3995 , n3996 );
xor ( n3998 , n3991 , n3997 );
not ( n3999 , n3026 );
not ( n4000 , n539 );
not ( n4001 , n3279 );
not ( n4002 , n4001 );
or ( n4003 , n4000 , n4002 );
nand ( n4004 , n3279 , n3069 );
nand ( n4005 , n4003 , n4004 );
not ( n4006 , n4005 );
or ( n4007 , n3999 , n4006 );
nand ( n4008 , n3071 , n3103 );
nand ( n4009 , n4007 , n4008 );
xor ( n4010 , n3998 , n4009 );
xor ( n4011 , n3990 , n4010 );
xor ( n4012 , n3950 , n4011 );
not ( n4013 , n549 );
not ( n4014 , n550 );
and ( n4015 , n4013 , n4014 );
and ( n4016 , n549 , n550 );
or ( n4017 , n4014 , n551 );
not ( n4018 , n551 );
or ( n4019 , n4018 , n550 );
nand ( n4020 , n4017 , n4019 );
nor ( n4021 , n4015 , n4016 , n4020 );
buf ( n4022 , n4021 );
not ( n4023 , n4022 );
not ( n4024 , n549 );
not ( n4025 , n716 );
nand ( n4026 , n3466 , n3932 , n3794 );
nor ( n4027 , n3927 , n3931 );
nor ( n4028 , n3805 , n4027 );
not ( n4029 , n3933 );
nor ( n4030 , n4028 , n4029 );
nand ( n4031 , n4026 , n4030 );
not ( n4032 , n912 );
not ( n4033 , n901 );
not ( n4034 , n1036 );
or ( n4035 , n4033 , n4034 );
nand ( n4036 , n2633 , n497 );
nand ( n4037 , n4035 , n4036 );
not ( n4038 , n4037 );
or ( n4039 , n4032 , n4038 );
nand ( n4040 , n3881 , n893 );
nand ( n4041 , n4039 , n4040 );
not ( n4042 , n2892 );
not ( n4043 , n489 );
not ( n4044 , n1204 );
or ( n4045 , n4043 , n4044 );
not ( n4046 , n489 );
nand ( n4047 , n900 , n4046 );
nand ( n4048 , n4045 , n4047 );
not ( n4049 , n4048 );
or ( n4050 , n4042 , n4049 );
not ( n4051 , n489 );
not ( n4052 , n3521 );
or ( n4053 , n4051 , n4052 );
not ( n4054 , n3519 );
nand ( n4055 , n4054 , n4046 );
nand ( n4056 , n4053 , n4055 );
nand ( n4057 , n3871 , n4056 );
nand ( n4058 , n4050 , n4057 );
xor ( n4059 , n4041 , n4058 );
not ( n4060 , n489 );
nor ( n4061 , n4060 , n2609 );
xor ( n4062 , n4059 , n4061 );
not ( n4063 , n1026 );
and ( n4064 , n844 , n495 );
not ( n4065 , n844 );
and ( n4066 , n4065 , n813 );
or ( n4067 , n4064 , n4066 );
not ( n4068 , n4067 );
or ( n4069 , n4063 , n4068 );
nand ( n4070 , n941 , n3896 );
nand ( n4071 , n4069 , n4070 );
not ( n4072 , n831 );
not ( n4073 , n3863 );
or ( n4074 , n4072 , n4073 );
not ( n4075 , n501 );
not ( n4076 , n3592 );
not ( n4077 , n4076 );
not ( n4078 , n4077 );
or ( n4079 , n4075 , n4078 );
nand ( n4080 , n4076 , n833 );
nand ( n4081 , n4079 , n4080 );
nand ( n4082 , n4081 , n858 );
nand ( n4083 , n4074 , n4082 );
xor ( n4084 , n4071 , n4083 );
not ( n4085 , n807 );
not ( n4086 , n499 );
and ( n4087 , n456 , n475 );
not ( n4088 , n456 );
and ( n4089 , n4088 , n459 );
nor ( n4090 , n4087 , n4089 );
not ( n4091 , n4090 );
or ( n4092 , n4086 , n4091 );
not ( n4093 , n4090 );
nand ( n4094 , n4093 , n782 );
nand ( n4095 , n4092 , n4094 );
not ( n4096 , n4095 );
or ( n4097 , n4085 , n4096 );
nand ( n4098 , n770 , n3812 );
nand ( n4099 , n4097 , n4098 );
xor ( n4100 , n4084 , n4099 );
xor ( n4101 , n4062 , n4100 );
not ( n4102 , n2959 );
not ( n4103 , n493 );
not ( n4104 , n791 );
or ( n4105 , n4103 , n4104 );
nand ( n4106 , n798 , n739 );
nand ( n4107 , n4105 , n4106 );
not ( n4108 , n4107 );
or ( n4109 , n4102 , n4108 );
nand ( n4110 , n3822 , n2967 );
nand ( n4111 , n4109 , n4110 );
not ( n4112 , n2606 );
not ( n4113 , n491 );
not ( n4114 , n2658 );
or ( n4115 , n4113 , n4114 );
nand ( n4116 , n982 , n2613 );
nand ( n4117 , n4115 , n4116 );
not ( n4118 , n4117 );
or ( n4119 , n4112 , n4118 );
nand ( n4120 , n3840 , n3573 );
nand ( n4121 , n4119 , n4120 );
xor ( n4122 , n4111 , n4121 );
nand ( n4123 , n945 , n1441 );
xor ( n4124 , n4122 , n4123 );
xor ( n4125 , n4101 , n4124 );
xor ( n4126 , n3909 , n3920 );
and ( n4127 , n4126 , n3925 );
and ( n4128 , n3909 , n3920 );
or ( n4129 , n4127 , n4128 );
xor ( n4130 , n4125 , n4129 );
xor ( n4131 , n3910 , n3914 );
and ( n4132 , n4131 , n3919 );
and ( n4133 , n3910 , n3914 );
or ( n4134 , n4132 , n4133 );
xor ( n4135 , n3816 , n3832 );
and ( n4136 , n4135 , n3842 );
and ( n4137 , n3816 , n3832 );
or ( n4138 , n4136 , n4137 );
xor ( n4139 , n3873 , n3883 );
and ( n4140 , n4139 , n3898 );
and ( n4141 , n3873 , n3883 );
or ( n4142 , n4140 , n4141 );
xor ( n4143 , n4138 , n4142 );
xor ( n4144 , n3844 , n3848 );
and ( n4145 , n4144 , n3865 );
and ( n4146 , n3844 , n3848 );
or ( n4147 , n4145 , n4146 );
xor ( n4148 , n4143 , n4147 );
xor ( n4149 , n4134 , n4148 );
xor ( n4150 , n3843 , n3866 );
and ( n4151 , n4150 , n3899 );
and ( n4152 , n3843 , n3866 );
or ( n4153 , n4151 , n4152 );
xor ( n4154 , n4149 , n4153 );
xor ( n4155 , n4130 , n4154 );
buf ( n4156 , n4155 );
not ( n4157 , n4156 );
xor ( n4158 , n3900 , n3904 );
and ( n4159 , n4158 , n3926 );
and ( n4160 , n3900 , n3904 );
or ( n4161 , n4159 , n4160 );
not ( n4162 , n4161 );
nand ( n4163 , n4157 , n4162 );
nand ( n4164 , n4156 , n4161 );
nand ( n4165 , n4163 , n4164 );
not ( n4166 , n4165 );
and ( n4167 , n4031 , n4166 );
not ( n4168 , n4031 );
and ( n4169 , n4168 , n4165 );
nor ( n4170 , n4167 , n4169 );
not ( n4171 , n4170 );
or ( n4172 , n4025 , n4171 );
nand ( n4173 , n3457 , n3785 );
not ( n4174 , n4173 );
not ( n4175 , n4174 );
not ( n4176 , n3317 );
or ( n4177 , n4175 , n4176 );
not ( n4178 , n3782 );
not ( n4179 , n3454 );
or ( n4180 , n4178 , n4179 );
nand ( n4181 , n4180 , n3785 );
buf ( n4182 , n4181 );
nand ( n4183 , n4177 , n4182 );
not ( n4184 , n3657 );
not ( n4185 , n3672 );
not ( n4186 , n4185 );
or ( n4187 , n4184 , n4186 );
not ( n4188 , n3658 );
not ( n4189 , n3672 );
or ( n4190 , n4188 , n4189 );
nand ( n4191 , n4190 , n3681 );
nand ( n4192 , n4187 , n4191 );
not ( n4193 , n4192 );
not ( n4194 , n3660 );
not ( n4195 , n3671 );
or ( n4196 , n4194 , n4195 );
or ( n4197 , n3671 , n3660 );
nand ( n4198 , n4197 , n3664 );
nand ( n4199 , n4196 , n4198 );
not ( n4200 , n503 );
not ( n4201 , n1602 );
or ( n4202 , n4200 , n4201 );
nand ( n4203 , n4202 , n1441 );
not ( n4204 , n4203 );
nand ( n4205 , n519 , n489 );
and ( n4206 , n4204 , n4205 );
not ( n4207 , n4204 );
not ( n4208 , n4205 );
and ( n4209 , n4207 , n4208 );
nor ( n4210 , n4206 , n4209 );
not ( n4211 , n3737 );
not ( n4212 , n3734 );
or ( n4213 , n4211 , n4212 );
xor ( n4214 , n489 , n517 );
nand ( n4215 , n2733 , n4214 );
nand ( n4216 , n4213 , n4215 );
xor ( n4217 , n4210 , n4216 );
not ( n4218 , n4217 );
not ( n4219 , n3696 );
not ( n4220 , n1574 );
or ( n4221 , n4219 , n4220 );
xor ( n4222 , n505 , n501 );
nand ( n4223 , n1867 , n4222 );
nand ( n4224 , n4221 , n4223 );
not ( n4225 , n3743 );
not ( n4226 , n1687 );
or ( n4227 , n4225 , n4226 );
xor ( n4228 , n511 , n495 );
nand ( n4229 , n1595 , n4228 );
nand ( n4230 , n4227 , n4229 );
xor ( n4231 , n4224 , n4230 );
not ( n4232 , n3705 );
not ( n4233 , n1630 );
or ( n4234 , n4232 , n4233 );
xor ( n4235 , n499 , n507 );
nand ( n4236 , n1634 , n4235 );
nand ( n4237 , n4234 , n4236 );
xor ( n4238 , n4231 , n4237 );
not ( n4239 , n4238 );
or ( n4240 , n4218 , n4239 );
or ( n4241 , n4238 , n4217 );
nand ( n4242 , n4240 , n4241 );
xnor ( n4243 , n4199 , n4242 );
not ( n4244 , n4243 );
and ( n4245 , n4193 , n4244 );
and ( n4246 , n4192 , n4243 );
nor ( n4247 , n4245 , n4246 );
not ( n4248 , n3700 );
nand ( n4249 , n3754 , n4248 );
not ( n4250 , n3700 );
not ( n4251 , n3753 );
or ( n4252 , n4250 , n4251 );
and ( n4253 , n3716 , n3723 );
not ( n4254 , n3716 );
and ( n4255 , n4254 , n3726 );
or ( n4256 , n4253 , n4255 );
nand ( n4257 , n4252 , n4256 );
nand ( n4258 , n4249 , n4257 );
not ( n4259 , n4258 );
not ( n4260 , n2025 );
and ( n4261 , n493 , n722 );
not ( n111813 , n493 );
and ( n111814 , n111813 , n494 );
or ( n4262 , n4261 , n111814 );
nand ( n4263 , n4260 , n4262 , n3720 );
xor ( n4264 , n513 , n493 );
nand ( n4265 , n2031 , n4264 );
nand ( n4266 , n4263 , n4265 );
not ( n4267 , n4266 );
not ( n4268 , n3713 );
not ( n4269 , n2455 );
or ( n4270 , n4268 , n4269 );
xor ( n4271 , n515 , n491 );
nand ( n4272 , n2764 , n4271 );
nand ( n4273 , n4270 , n4272 );
not ( n4274 , n4273 );
and ( n4275 , n4267 , n4274 );
not ( n4276 , n4267 );
and ( n4277 , n4276 , n4273 );
or ( n4278 , n4275 , n4277 );
not ( n4279 , n3750 );
not ( n4280 , n2083 );
or ( n4281 , n4279 , n4280 );
xor ( n4282 , n497 , n509 );
nand ( n4283 , n2086 , n4282 );
nand ( n4284 , n4281 , n4283 );
not ( n4285 , n4284 );
xor ( n4286 , n4278 , n4285 );
not ( n4287 , n3688 );
or ( n4288 , n3686 , n4287 );
nand ( n4289 , n4288 , n3698 );
nand ( n4290 , n3686 , n4287 );
nand ( n4291 , n4289 , n4290 );
not ( n4292 , n3722 );
not ( n4293 , n3707 );
or ( n4294 , n4292 , n4293 );
or ( n4295 , n3722 , n3707 );
nand ( n4296 , n4295 , n3715 );
nand ( n4297 , n4294 , n4296 );
xor ( n4298 , n4291 , n4297 );
or ( n4299 , n3745 , n3739 );
nand ( n4300 , n4299 , n3752 );
nand ( n4301 , n3739 , n3745 );
nand ( n4302 , n4300 , n4301 );
xor ( n4303 , n4298 , n4302 );
buf ( n4304 , n4303 );
xnor ( n4305 , n4286 , n4304 );
not ( n4306 , n4305 );
or ( n4307 , n4259 , n4306 );
not ( n4308 , n4286 );
not ( n4309 , n4303 );
or ( n4310 , n4308 , n4309 );
nand ( n4311 , n4310 , n4249 );
not ( n4312 , n4311 );
not ( n4313 , n4286 );
not ( n4314 , n4303 );
nand ( n4315 , n4313 , n4314 );
nand ( n4316 , n4312 , n4315 , n4257 );
nand ( n4317 , n4307 , n4316 );
xor ( n4318 , n4247 , n4317 );
not ( n4319 , n3758 );
not ( n4320 , n3763 );
not ( n4321 , n4320 );
or ( n4322 , n4319 , n4321 );
not ( n4323 , n3682 );
nand ( n4324 , n4322 , n4323 );
not ( n4325 , n3758 );
nand ( n4326 , n4325 , n3763 );
nand ( n4327 , n4324 , n4326 );
nor ( n4328 , n4318 , n4327 );
not ( n4329 , n4328 );
nand ( n4330 , n4318 , n4327 );
nand ( n4331 , n4329 , n4330 );
not ( n4332 , n4331 );
and ( n4333 , n4183 , n4332 );
not ( n4334 , n4183 );
and ( n4335 , n4334 , n4331 );
nor ( n4336 , n4333 , n4335 );
nand ( n4337 , n4336 , n455 );
nand ( n4338 , n4172 , n4337 );
not ( n4339 , n4338 );
not ( n4340 , n4339 );
or ( n4341 , n4024 , n4340 );
not ( n4342 , n4339 );
nand ( n4343 , n4342 , n4013 );
nand ( n4344 , n4341 , n4343 );
not ( n4345 , n4344 );
or ( n4346 , n4023 , n4345 );
nor ( n4347 , n4173 , n4328 );
not ( n4348 , n4347 );
not ( n4349 , n3317 );
or ( n4350 , n4348 , n4349 );
or ( n4351 , n4181 , n4328 );
nand ( n4352 , n4351 , n4330 );
not ( n4353 , n4352 );
nand ( n4354 , n4350 , n4353 );
not ( n4355 , n4354 );
not ( n4356 , n4286 );
not ( n4357 , n4314 );
or ( n4358 , n4356 , n4357 );
nand ( n4359 , n4358 , n4258 );
not ( n4360 , n4286 );
nand ( n4361 , n4360 , n4303 );
nand ( n4362 , n4359 , n4361 );
not ( n4363 , n4228 );
not ( n4364 , n1687 );
or ( n4365 , n4363 , n4364 );
xor ( n4366 , n510 , n495 );
nand ( n4367 , n1595 , n4366 );
nand ( n4368 , n4365 , n4367 );
not ( n4369 , n1805 );
xor ( n4370 , n506 , n499 );
not ( n4371 , n4370 );
or ( n4372 , n4369 , n4371 );
not ( n4373 , n1805 );
and ( n4374 , n1629 , n4235 );
nand ( n4375 , n4373 , n4374 );
nand ( n4376 , n4372 , n4375 );
nand ( n4377 , n518 , n489 );
and ( n4378 , n4376 , n4377 );
not ( n4379 , n4376 );
not ( n4380 , n4377 );
and ( n4381 , n4379 , n4380 );
nor ( n4382 , n4378 , n4381 );
xnor ( n4383 , n4368 , n4382 );
xor ( n4384 , n4291 , n4297 );
and ( n4385 , n4384 , n4302 );
and ( n4386 , n4291 , n4297 );
or ( n4387 , n4385 , n4386 );
xor ( n4388 , n4383 , n4387 );
not ( n4389 , n4214 );
not ( n4390 , n3734 );
or ( n4391 , n4389 , n4390 );
xor ( n4392 , n516 , n489 );
nand ( n4393 , n2733 , n4392 );
nand ( n4394 , n4391 , n4393 );
not ( n4395 , n4222 );
not ( n4396 , n1750 );
or ( n4397 , n4395 , n4396 );
nand ( n4398 , n1867 , n501 );
nand ( n4399 , n4397 , n4398 );
not ( n4400 , n4399 );
xor ( n4401 , n4394 , n4400 );
xor ( n4402 , n4401 , n4284 );
not ( n4403 , n4402 );
xor ( n4404 , n4388 , n4403 );
not ( n4405 , n4404 );
and ( n4406 , n4362 , n4405 );
not ( n4407 , n4362 );
and ( n4408 , n4407 , n4404 );
nor ( n4409 , n4406 , n4408 );
not ( n4410 , n4274 );
not ( n4411 , n4267 );
or ( n4412 , n4410 , n4411 );
nand ( n4413 , n4412 , n4285 );
nand ( n4414 , n4266 , n4273 );
nand ( n4415 , n4413 , n4414 );
not ( n4416 , n4415 );
not ( n4417 , n4204 );
not ( n4418 , n4208 );
or ( n4419 , n4417 , n4418 );
not ( n4420 , n4205 );
not ( n4421 , n4203 );
or ( n4422 , n4420 , n4421 );
nand ( n4423 , n4422 , n4216 );
nand ( n4424 , n4419 , n4423 );
not ( n4425 , n4230 );
not ( n4426 , n4237 );
or ( n4427 , n4425 , n4426 );
nor ( n4428 , n4237 , n4230 );
not ( n4429 , n4224 );
or ( n4430 , n4428 , n4429 );
nand ( n4431 , n4427 , n4430 );
xor ( n4432 , n4424 , n4431 );
xor ( n4433 , n514 , n491 );
not ( n4434 , n4433 );
not ( n4435 , n2277 );
or ( n4436 , n4434 , n4435 );
nand ( n4437 , n2278 , n4271 , n2453 );
nand ( n4438 , n4436 , n4437 );
not ( n4439 , n2479 );
not ( n4440 , n4264 );
or ( n4441 , n4439 , n4440 );
nand ( n4442 , n4441 , n2772 );
xor ( n4443 , n493 , n512 );
not ( n4444 , n4443 );
nand ( n4445 , n4444 , n1561 );
nand ( n4446 , n4442 , n4445 );
not ( n4447 , n4446 );
xor ( n4448 , n4438 , n4447 );
not ( n4449 , n4282 );
not ( n4450 , n1660 );
or ( n4451 , n4449 , n4450 );
xor ( n4452 , n497 , n508 );
nand ( n4453 , n1563 , n4452 );
nand ( n4454 , n4451 , n4453 );
xor ( n4455 , n4448 , n4454 );
xnor ( n4456 , n4432 , n4455 );
xor ( n4457 , n4416 , n4456 );
not ( n4458 , n4238 );
nand ( n4459 , n4458 , n4217 );
not ( n4460 , n4459 );
not ( n4461 , n4199 );
or ( n4462 , n4460 , n4461 );
not ( n4463 , n4217 );
nand ( n4464 , n4463 , n4238 );
nand ( n4465 , n4462 , n4464 );
xnor ( n4466 , n4457 , n4465 );
not ( n4467 , n4466 );
and ( n4468 , n4409 , n4467 );
not ( n4469 , n4409 );
and ( n4470 , n4469 , n4466 );
or ( n4471 , n4468 , n4470 );
buf ( n4472 , n4243 );
not ( n4473 , n4472 );
not ( n4474 , n4258 );
not ( n4475 , n4305 );
or ( n4476 , n4474 , n4475 );
nand ( n4477 , n4476 , n4316 );
not ( n4478 , n4477 );
and ( n4479 , n4473 , n4478 );
nand ( n4480 , n4477 , n4472 );
buf ( n4481 , n4192 );
and ( n4482 , n4480 , n4481 );
nor ( n4483 , n4479 , n4482 );
nor ( n4484 , n4471 , n4483 );
not ( n4485 , n4484 );
nand ( n4486 , n4483 , n4471 );
nand ( n4487 , n4485 , n4486 );
not ( n4488 , n4487 );
nand ( n4489 , n4355 , n4488 );
not ( n4490 , n4489 );
nand ( n4491 , n4354 , n4487 );
not ( n4492 , n4491 );
or ( n4493 , n4490 , n4492 );
nand ( n4494 , n4493 , n455 );
not ( n4495 , n4164 );
not ( n4496 , n4030 );
not ( n4497 , n4026 );
or ( n4498 , n4496 , n4497 );
nand ( n4499 , n4498 , n4163 );
not ( n4500 , n4499 );
or ( n4501 , n4495 , n4500 );
not ( n4502 , n769 );
not ( n4503 , n4095 );
or ( n4504 , n4502 , n4503 );
not ( n4505 , n499 );
not ( n4506 , n3859 );
or ( n4507 , n4505 , n4506 );
nand ( n4508 , n3858 , n782 );
nand ( n4509 , n4507 , n4508 );
nand ( n4510 , n4509 , n1122 );
nand ( n4511 , n4504 , n4510 );
and ( n4512 , n2975 , n489 );
xor ( n4513 , n4511 , n4512 );
not ( n4514 , n1026 );
not ( n4515 , n495 );
not ( n4516 , n2949 );
or ( n4517 , n4515 , n4516 );
not ( n4518 , n960 );
nand ( n4519 , n4518 , n813 );
nand ( n4520 , n4517 , n4519 );
not ( n4521 , n4520 );
or ( n4522 , n4514 , n4521 );
nand ( n4523 , n4067 , n1086 );
nand ( n4524 , n4522 , n4523 );
xor ( n4525 , n4513 , n4524 );
xor ( n4526 , n4111 , n4121 );
and ( n4527 , n4526 , n4123 );
and ( n4528 , n4111 , n4121 );
or ( n4529 , n4527 , n4528 );
xor ( n4530 , n4525 , n4529 );
xor ( n4531 , n4138 , n4142 );
and ( n4532 , n4531 , n4147 );
and ( n4533 , n4138 , n4142 );
or ( n4534 , n4532 , n4533 );
xor ( n4535 , n4530 , n4534 );
xor ( n4536 , n4134 , n4148 );
and ( n4537 , n4536 , n4153 );
and ( n4538 , n4134 , n4148 );
or ( n4539 , n4537 , n4538 );
xor ( n4540 , n4535 , n4539 );
not ( n4541 , n489 );
not ( n4542 , n1263 );
or ( n4543 , n4541 , n4542 );
or ( n4544 , n1263 , n489 );
nand ( n4545 , n4543 , n4544 );
not ( n4546 , n4545 );
buf ( n4547 , n2892 );
not ( n4548 , n4547 );
or ( n4549 , n4546 , n4548 );
not ( n4550 , n4046 );
not ( n4551 , n4054 );
or ( n4552 , n4550 , n4551 );
nand ( n4553 , n4552 , n3522 );
nand ( n4554 , n4048 , n4553 );
nand ( n4555 , n4549 , n4554 );
not ( n4556 , n4081 );
not ( n4557 , n831 );
or ( n4558 , n4556 , n4557 );
nand ( n4559 , n858 , n501 );
nand ( n4560 , n4558 , n4559 );
not ( n4561 , n4560 );
xor ( n4562 , n4555 , n4561 );
not ( n4563 , n4123 );
xor ( n4564 , n4562 , n4563 );
xor ( n4565 , n4041 , n4058 );
and ( n4566 , n4565 , n4061 );
and ( n4567 , n4041 , n4058 );
or ( n4568 , n4566 , n4567 );
xor ( n4569 , n4071 , n4083 );
and ( n4570 , n4569 , n4099 );
and ( n4571 , n4071 , n4083 );
or ( n4572 , n4570 , n4571 );
xor ( n4573 , n4568 , n4572 );
not ( n4574 , n724 );
not ( n4575 , n493 );
not ( n4576 , n3892 );
or ( n4577 , n4575 , n4576 );
nor ( n4578 , n456 , n464 );
not ( n4579 , n4578 );
not ( n4580 , n480 );
nand ( n4581 , n4580 , n456 );
nand ( n4582 , n4579 , n4581 , n739 );
nand ( n4583 , n4577 , n4582 );
not ( n4584 , n4583 );
or ( n4585 , n4574 , n4584 );
nand ( n4586 , n4107 , n760 );
nand ( n4587 , n4585 , n4586 );
not ( n4588 , n912 );
not ( n4589 , n497 );
not ( n4590 , n2178 );
or ( n4591 , n4589 , n4590 );
nand ( n4592 , n2177 , n901 );
nand ( n4593 , n4591 , n4592 );
not ( n4594 , n4593 );
or ( n4595 , n4588 , n4594 );
nand ( n4596 , n4037 , n893 );
nand ( n4597 , n4595 , n4596 );
xor ( n4598 , n4587 , n4597 );
not ( n4599 , n3573 );
not ( n4600 , n4117 );
or ( n4601 , n4599 , n4600 );
not ( n4602 , n491 );
not ( n4603 , n779 );
or ( n4604 , n4602 , n4603 );
nand ( n4605 , n778 , n2613 );
nand ( n4606 , n4604 , n4605 );
nand ( n4607 , n4606 , n2606 );
nand ( n4608 , n4601 , n4607 );
xor ( n4609 , n4598 , n4608 );
xor ( n4610 , n4573 , n4609 );
xor ( n4611 , n4564 , n4610 );
xor ( n4612 , n4062 , n4100 );
and ( n4613 , n4612 , n4124 );
and ( n4614 , n4062 , n4100 );
or ( n4615 , n4613 , n4614 );
xor ( n4616 , n4611 , n4615 );
xor ( n4617 , n4540 , n4616 );
not ( n4618 , n4617 );
xor ( n4619 , n4125 , n4129 );
and ( n4620 , n4619 , n4154 );
and ( n4621 , n4125 , n4129 );
or ( n4622 , n4620 , n4621 );
not ( n4623 , n4622 );
nand ( n4624 , n4618 , n4623 );
buf ( n4625 , n4624 );
nand ( n4626 , n4617 , n4622 );
and ( n4627 , n4625 , n4626 );
nor ( n4628 , n4627 , n455 );
nand ( n4629 , n4501 , n4628 );
not ( n4630 , n455 );
nand ( n4631 , n4630 , n4626 );
not ( n4632 , n4631 );
nand ( n4633 , n4632 , n4499 , n4164 , n4625 );
nand ( n4634 , n4494 , n4629 , n4633 );
not ( n4635 , n4634 );
and ( n4636 , n4013 , n4635 );
not ( n4637 , n4013 );
buf ( n4638 , n4634 );
and ( n4639 , n4637 , n4638 );
nor ( n4640 , n4636 , n4639 );
nand ( n4641 , n4640 , n4020 );
nand ( n4642 , n4346 , n4641 );
xor ( n4643 , n4012 , n4642 );
xor ( n4644 , n3294 , n4643 );
not ( n4645 , n4020 );
not ( n4646 , n4344 );
or ( n4647 , n4645 , n4646 );
not ( n4648 , n549 );
not ( n4649 , n455 );
not ( n4650 , n3787 );
or ( n4651 , n4649 , n4650 );
nand ( n4652 , n4651 , n3941 );
not ( n4653 , n4652 );
not ( n4654 , n4653 );
or ( n4655 , n4648 , n4654 );
nand ( n4656 , n4652 , n4013 );
nand ( n4657 , n4655 , n4656 );
nand ( n4658 , n4657 , n4022 );
nand ( n4659 , n4647 , n4658 );
not ( n4660 , n3186 );
not ( n4661 , n3179 );
or ( n4662 , n4660 , n4661 );
not ( n4663 , n3195 );
nand ( n4664 , n4662 , n4663 );
xnor ( n4665 , n4664 , n3207 );
not ( n4666 , n3026 );
not ( n4667 , n3098 );
or ( n4668 , n4666 , n4667 );
not ( n4669 , n539 );
not ( n4670 , n3149 );
not ( n4671 , n4670 );
or ( n4672 , n4669 , n4671 );
nand ( n4673 , n3149 , n3069 );
nand ( n4674 , n4672 , n4673 );
nand ( n4675 , n4674 , n3103 );
nand ( n4676 , n4668 , n4675 );
xor ( n4677 , n4665 , n4676 );
and ( n4678 , n3128 , n3186 );
not ( n4679 , n3026 );
not ( n4680 , n4674 );
or ( n4681 , n4679 , n4680 );
not ( n4682 , n3069 );
not ( n4683 , n3176 );
or ( n4684 , n4682 , n4683 );
nand ( n4685 , n539 , n3173 );
nand ( n4686 , n4684 , n4685 );
nand ( n4687 , n4686 , n3101 );
nand ( n4688 , n4681 , n4687 );
xor ( n4689 , n4678 , n4688 );
not ( n4690 , n3021 );
not ( n4691 , n3190 );
or ( n4692 , n4690 , n4691 );
nand ( n4693 , n4692 , n541 );
and ( n4694 , n3128 , n540 );
nor ( n4695 , n4694 , n3069 );
and ( n4696 , n4693 , n4695 );
and ( n4697 , n3069 , n3026 );
nand ( n4698 , n3176 , n4697 );
nor ( n4699 , n3102 , n539 );
and ( n4700 , n3128 , n4699 );
and ( n4701 , n3101 , n539 );
not ( n4702 , n4701 );
not ( n4703 , n3127 );
not ( n4704 , n4703 );
nor ( n4705 , n4702 , n4704 );
nor ( n4706 , n4700 , n4705 );
nand ( n4707 , n3173 , n3026 , n539 );
nand ( n4708 , n4698 , n4706 , n4707 );
and ( n4709 , n4696 , n4708 );
and ( n4710 , n4689 , n4709 );
and ( n4711 , n4678 , n4688 );
or ( n4712 , n4710 , n4711 );
and ( n4713 , n4677 , n4712 );
and ( n4714 , n4665 , n4676 );
or ( n4715 , n4713 , n4714 );
not ( n4716 , n2362 );
not ( n4717 , n2127 );
or ( n4718 , n4716 , n4717 );
not ( n4719 , n543 );
not ( n4720 , n3980 );
not ( n4721 , n4720 );
or ( n4722 , n4719 , n4721 );
nand ( n4723 , n3980 , n2123 );
nand ( n4724 , n4722 , n4723 );
nand ( n4725 , n4724 , n714 );
nand ( n4726 , n4718 , n4725 );
xor ( n4727 , n4715 , n4726 );
not ( n4728 , n3017 );
not ( n4729 , n2704 );
or ( n4730 , n4728 , n4729 );
not ( n4731 , n545 );
not ( n4732 , n2355 );
not ( n4733 , n4732 );
or ( n4734 , n4731 , n4733 );
nand ( n4735 , n2355 , n706 );
nand ( n4736 , n4734 , n4735 );
nand ( n4737 , n4736 , n2376 );
nand ( n4738 , n4730 , n4737 );
xor ( n4739 , n4727 , n4738 );
xor ( n4740 , n4659 , n4739 );
xor ( n4741 , n4665 , n4676 );
xor ( n4742 , n4741 , n4712 );
not ( n4743 , n3214 );
not ( n4744 , n541 );
not ( n4745 , n3067 );
or ( n4746 , n4744 , n4745 );
nand ( n4747 , n3068 , n3023 );
nand ( n4748 , n4746 , n4747 );
not ( n4749 , n4748 );
or ( n4750 , n4743 , n4749 );
not ( n4751 , n541 );
not ( n4752 , n3093 );
or ( n4753 , n4751 , n4752 );
nand ( n4754 , n3092 , n3023 );
nand ( n4755 , n4753 , n4754 );
nand ( n4756 , n4755 , n3288 );
nand ( n4757 , n4750 , n4756 );
xor ( n4758 , n4678 , n4688 );
xor ( n4759 , n4758 , n4709 );
xor ( n4760 , n4757 , n4759 );
not ( n4761 , n2361 );
not ( n4762 , n543 );
not ( n4763 , n3250 );
or ( n4764 , n4762 , n4763 );
nand ( n4765 , n3249 , n2123 );
nand ( n4766 , n4764 , n4765 );
not ( n4767 , n4766 );
or ( n4768 , n4761 , n4767 );
not ( n4769 , n543 );
not ( n4770 , n4001 );
or ( n4771 , n4769 , n4770 );
nand ( n4772 , n3279 , n2123 );
nand ( n4773 , n4771 , n4772 );
nand ( n4774 , n4773 , n714 );
nand ( n4775 , n4768 , n4774 );
and ( n4776 , n4760 , n4775 );
and ( n4777 , n4757 , n4759 );
or ( n4778 , n4776 , n4777 );
xor ( n4779 , n4742 , n4778 );
not ( n4780 , n3300 );
not ( n4781 , n547 );
not ( n4782 , n2698 );
or ( n4783 , n4781 , n4782 );
not ( n4784 , n2698 );
nand ( n4785 , n4784 , n2369 );
nand ( n4786 , n4783 , n4785 );
not ( n4787 , n4786 );
or ( n4788 , n4780 , n4787 );
not ( n4789 , n547 );
not ( n4790 , n3012 );
or ( n4791 , n4789 , n4790 );
buf ( n4792 , n3011 );
nand ( n4793 , n4792 , n2369 );
nand ( n4794 , n4791 , n4793 );
nand ( n4795 , n4794 , n3298 );
nand ( n4796 , n4788 , n4795 );
and ( n4797 , n4779 , n4796 );
and ( n4798 , n4742 , n4778 );
or ( n4799 , n4797 , n4798 );
and ( n4800 , n4740 , n4799 );
and ( n4801 , n4659 , n4739 );
or ( n4802 , n4800 , n4801 );
and ( n4803 , n4644 , n4802 );
and ( n4804 , n3294 , n4643 );
or ( n4805 , n4803 , n4804 );
not ( n4806 , n4020 );
not ( n4807 , n549 );
not ( n4808 , n455 );
not ( n4809 , n4486 );
not ( n4810 , n4354 );
or ( n4811 , n4809 , n4810 );
nand ( n4812 , n4811 , n4485 );
and ( n4813 , n517 , n489 );
not ( n4814 , n4443 );
not ( n4815 , n2028 );
or ( n4816 , n4814 , n4815 );
xor ( n4817 , n511 , n493 );
nand ( n4818 , n2031 , n4817 );
nand ( n4819 , n4816 , n4818 );
xor ( n4820 , n4813 , n4819 );
not ( n4821 , n4452 );
not ( n4822 , n2083 );
or ( n4823 , n4821 , n4822 );
xor ( n4824 , n507 , n497 );
nand ( n4825 , n2086 , n4824 );
nand ( n4826 , n4823 , n4825 );
not ( n4827 , n4826 );
and ( n4828 , n4820 , n4827 );
not ( n4829 , n4820 );
and ( n4830 , n4829 , n4826 );
or ( n4831 , n4828 , n4830 );
not ( n4832 , n4392 );
not ( n4833 , n3368 );
nand ( n4834 , n4833 , n3377 );
not ( n4835 , n4834 );
not ( n4836 , n4835 );
or ( n4837 , n4832 , n4836 );
xor ( n4838 , n490 , n491 );
xor ( n4839 , n515 , n489 );
nand ( n4840 , n4838 , n4839 );
nand ( n4841 , n4837 , n4840 );
not ( n4842 , n4433 );
not ( n4843 , n2455 );
or ( n4844 , n4842 , n4843 );
xor ( n4845 , n491 , n513 );
nand ( n4846 , n4845 , n2279 );
nand ( n4847 , n4844 , n4846 );
not ( n4848 , n4847 );
xor ( n4849 , n4841 , n4848 );
and ( n4850 , n4849 , n4399 );
not ( n4851 , n4849 );
and ( n4852 , n4851 , n4400 );
nor ( n4853 , n4850 , n4852 );
xor ( n4854 , n4831 , n4853 );
xor ( n4855 , n4394 , n4400 );
and ( n4856 , n4855 , n4284 );
and ( n4857 , n4394 , n4400 );
or ( n4858 , n4856 , n4857 );
not ( n4859 , n4858 );
and ( n4860 , n4854 , n4859 );
not ( n4861 , n4854 );
and ( n4862 , n4861 , n4858 );
nor ( n4863 , n4860 , n4862 );
not ( n4864 , n4424 );
not ( n4865 , n4431 );
not ( n4866 , n4865 );
not ( n4867 , n4866 );
or ( n4868 , n4864 , n4867 );
not ( n4869 , n4424 );
not ( n4870 , n4869 );
not ( n4871 , n4865 );
or ( n4872 , n4870 , n4871 );
nand ( n4873 , n4872 , n4455 );
nand ( n4874 , n4868 , n4873 );
not ( n4875 , n4874 );
not ( n4876 , n4438 );
not ( n4877 , n4876 );
not ( n4878 , n4446 );
or ( n4879 , n4877 , n4878 );
nand ( n4880 , n4879 , n4454 );
not ( n4881 , n4876 );
nand ( n4882 , n4881 , n4447 );
nand ( n4883 , n4880 , n4882 );
or ( n4884 , n4376 , n4380 );
nand ( n4885 , n4884 , n4368 );
nand ( n4886 , n4376 , n4380 );
nand ( n4887 , n4885 , n4886 );
and ( n4888 , n4883 , n4887 );
not ( n4889 , n4883 );
not ( n4890 , n4887 );
and ( n4891 , n4889 , n4890 );
nor ( n4892 , n4888 , n4891 );
not ( n4893 , n4370 );
not ( n4894 , n3339 );
or ( n4895 , n4893 , n4894 );
xor ( n4896 , n505 , n499 );
nand ( n4897 , n1634 , n4896 );
nand ( n4898 , n4895 , n4897 );
not ( n4899 , n4366 );
not ( n4900 , n1592 );
or ( n4901 , n4899 , n4900 );
xor ( n4902 , n509 , n495 );
nand ( n4903 , n1595 , n4902 );
nand ( n4904 , n4901 , n4903 );
xor ( n4905 , n4898 , n4904 );
not ( n4906 , n1889 );
not ( n4907 , n1573 );
or ( n4908 , n4906 , n4907 );
nand ( n4909 , n4908 , n501 );
xor ( n4910 , n4905 , n4909 );
and ( n4911 , n4892 , n4910 );
not ( n4912 , n4892 );
not ( n4913 , n4910 );
and ( n4914 , n4912 , n4913 );
nor ( n4915 , n4911 , n4914 );
and ( n4916 , n4875 , n4915 );
not ( n4917 , n4875 );
not ( n4918 , n4915 );
and ( n4919 , n4917 , n4918 );
nor ( n4920 , n4916 , n4919 );
not ( n4921 , n4383 );
nand ( n4922 , n4921 , n4403 );
not ( n4923 , n4922 );
not ( n4924 , n4387 );
or ( n4925 , n4923 , n4924 );
nand ( n4926 , n4402 , n4383 );
nand ( n4927 , n4925 , n4926 );
xor ( n4928 , n4920 , n4927 );
xor ( n4929 , n4863 , n4928 );
nand ( n4930 , n4416 , n4456 );
not ( n4931 , n4930 );
not ( n4932 , n4465 );
or ( n4933 , n4931 , n4932 );
not ( n4934 , n4456 );
nand ( n4935 , n4934 , n4415 );
nand ( n4936 , n4933 , n4935 );
xor ( n4937 , n4929 , n4936 );
not ( n4938 , n4937 );
not ( n4939 , n4466 );
not ( n4940 , n4404 );
or ( n4941 , n4939 , n4940 );
nand ( n4942 , n4941 , n4362 );
nand ( n4943 , n4467 , n4405 );
nand ( n4944 , n4942 , n4943 );
nand ( n4945 , n4938 , n4944 );
not ( n4946 , n4944 );
nand ( n4947 , n4937 , n4946 );
nand ( n4948 , n4945 , n4947 );
not ( n4949 , n4948 );
and ( n4950 , n4812 , n4949 );
not ( n4951 , n4812 );
and ( n4952 , n4951 , n4948 );
nor ( n4953 , n4950 , n4952 );
not ( n4954 , n4953 );
or ( n4955 , n4808 , n4954 );
not ( n4956 , n4625 );
or ( n4957 , n4956 , n4499 );
not ( n4958 , n4617 );
not ( n4959 , n4622 );
and ( n4960 , n4958 , n4959 );
nand ( n4961 , n4155 , n4161 );
and ( n4962 , n4626 , n4961 );
nor ( n4963 , n4960 , n4962 );
not ( n4964 , n4963 );
nand ( n4965 , n4957 , n4964 );
not ( n4966 , n3229 );
not ( n4967 , n489 );
nor ( n4968 , n4967 , n3565 );
not ( n4969 , n724 );
not ( n4970 , n493 );
not ( n4971 , n951 );
not ( n4972 , n4971 );
or ( n4973 , n4970 , n4972 );
not ( n4974 , n2576 );
nand ( n4975 , n4974 , n739 );
nand ( n4976 , n4973 , n4975 );
not ( n4977 , n4976 );
or ( n4978 , n4969 , n4977 );
nand ( n4979 , n4583 , n2966 );
nand ( n4980 , n4978 , n4979 );
xor ( n4981 , n4968 , n4980 );
not ( n4982 , n4593 );
not ( n4983 , n893 );
or ( n4984 , n4982 , n4983 );
not ( n4985 , n497 );
not ( n4986 , n4090 );
or ( n4987 , n4985 , n4986 );
or ( n4988 , n456 , n459 );
not ( n4989 , n475 );
nand ( n4990 , n4989 , n456 );
nand ( n4991 , n4988 , n4990 , n901 );
nand ( n4992 , n4987 , n4991 );
nand ( n4993 , n4992 , n912 );
nand ( n4994 , n4984 , n4993 );
xor ( n4995 , n4981 , n4994 );
not ( n4996 , n2624 );
not ( n4997 , n4606 );
or ( n4998 , n4996 , n4997 );
not ( n4999 , n873 );
and ( n5000 , n4999 , n491 );
not ( n5001 , n4999 );
and ( n5002 , n5001 , n2613 );
or ( n5003 , n5000 , n5002 );
nand ( n5004 , n5003 , n2606 );
nand ( n5005 , n4998 , n5004 );
not ( n5006 , n4545 );
not ( n5007 , n4056 );
or ( n5008 , n5006 , n5007 );
and ( n5009 , n489 , n2658 );
not ( n5010 , n489 );
and ( n5011 , n5010 , n989 );
or ( n5012 , n5009 , n5011 );
nand ( n5013 , n5012 , n4547 );
nand ( n5014 , n5008 , n5013 );
xor ( n5015 , n5005 , n5014 );
xor ( n5016 , n5015 , n4560 );
xor ( n5017 , n4995 , n5016 );
xor ( n5018 , n4555 , n4561 );
and ( n5019 , n5018 , n4563 );
and ( n5020 , n4555 , n4561 );
or ( n5021 , n5019 , n5020 );
xor ( n5022 , n5017 , n5021 );
xor ( n5023 , n4564 , n4610 );
and ( n5024 , n5023 , n4615 );
and ( n5025 , n4564 , n4610 );
or ( n5026 , n5024 , n5025 );
xor ( n5027 , n5022 , n5026 );
xor ( n5028 , n4587 , n4597 );
and ( n5029 , n5028 , n4608 );
and ( n5030 , n4587 , n4597 );
or ( n5031 , n5029 , n5030 );
xor ( n5032 , n4511 , n4512 );
and ( n5033 , n5032 , n4524 );
and ( n5034 , n4511 , n4512 );
or ( n5035 , n5033 , n5034 );
xor ( n5036 , n5031 , n5035 );
not ( n5037 , n1188 );
not ( n5038 , n857 );
or ( n5039 , n5037 , n5038 );
nand ( n5040 , n5039 , n501 );
not ( n5041 , n770 );
not ( n5042 , n4509 );
or ( n5043 , n5041 , n5042 );
not ( n5044 , n499 );
not ( n5045 , n4077 );
or ( n5046 , n5044 , n5045 );
nand ( n5047 , n4076 , n782 );
nand ( n5048 , n5046 , n5047 );
nand ( n5049 , n5048 , n1122 );
nand ( n5050 , n5043 , n5049 );
xor ( n5051 , n5040 , n5050 );
not ( n5052 , n1086 );
not ( n5053 , n4520 );
or ( n5054 , n5052 , n5053 );
not ( n5055 , n813 );
not ( n5056 , n1037 );
or ( n5057 , n5055 , n5056 );
nand ( n5058 , n1043 , n495 );
nand ( n5059 , n5057 , n5058 );
nand ( n5060 , n5059 , n1026 );
nand ( n5061 , n5054 , n5060 );
xor ( n5062 , n5051 , n5061 );
xor ( n5063 , n5036 , n5062 );
xor ( n5064 , n4568 , n4572 );
and ( n5065 , n5064 , n4609 );
and ( n5066 , n4568 , n4572 );
or ( n5067 , n5065 , n5066 );
xor ( n5068 , n5063 , n5067 );
xor ( n5069 , n4525 , n4529 );
and ( n5070 , n5069 , n4534 );
and ( n5071 , n4525 , n4529 );
or ( n5072 , n5070 , n5071 );
xor ( n5073 , n5068 , n5072 );
xor ( n5074 , n5027 , n5073 );
not ( n5075 , n5074 );
xor ( n5076 , n4535 , n4539 );
and ( n5077 , n5076 , n4616 );
and ( n5078 , n4535 , n4539 );
or ( n5079 , n5077 , n5078 );
not ( n5080 , n5079 );
nand ( n5081 , n5075 , n5080 );
buf ( n5082 , n5074 );
nand ( n5083 , n5082 , n5079 );
and ( n5084 , n5081 , n5083 );
nor ( n5085 , n4966 , n5084 );
and ( n5086 , n4965 , n5085 );
not ( n5087 , n4965 );
not ( n5088 , n455 );
and ( n5089 , n5084 , n5088 );
and ( n5090 , n5087 , n5089 );
nor ( n5091 , n5086 , n5090 );
nand ( n5092 , n4955 , n5091 );
buf ( n5093 , n5092 );
not ( n5094 , n5093 );
not ( n5095 , n5094 );
or ( n5096 , n4807 , n5095 );
nand ( n5097 , n5093 , n4013 );
nand ( n5098 , n5096 , n5097 );
not ( n5099 , n5098 );
or ( n5100 , n4806 , n5099 );
nand ( n5101 , n4022 , n4640 );
nand ( n5102 , n5100 , n5101 );
not ( n5103 , n552 );
not ( n5104 , n551 );
not ( n5105 , n1086 );
not ( n5106 , n5059 );
or ( n5107 , n5105 , n5106 );
not ( n5108 , n495 );
not ( n5109 , n2178 );
or ( n5110 , n5108 , n5109 );
nor ( n5111 , n456 , n460 );
not ( n5112 , n5111 );
not ( n5113 , n476 );
nand ( n5114 , n5113 , n456 );
nand ( n5115 , n5112 , n5114 , n813 );
nand ( n5116 , n5110 , n5115 );
nand ( n5117 , n5116 , n1026 );
nand ( n5118 , n5107 , n5117 );
not ( n5119 , n4547 );
xor ( n5120 , n489 , n778 );
not ( n5121 , n5120 );
or ( n5122 , n5119 , n5121 );
nand ( n5123 , n4056 , n5012 );
nand ( n5124 , n5122 , n5123 );
xor ( n5125 , n5118 , n5124 );
not ( n5126 , n489 );
nor ( n5127 , n5126 , n1263 );
xor ( n5128 , n5125 , n5127 );
not ( n5129 , n4992 );
not ( n5130 , n893 );
or ( n5131 , n5129 , n5130 );
not ( n5132 , n497 );
not ( n5133 , n3859 );
or ( n5134 , n5132 , n5133 );
nor ( n5135 , n456 , n458 );
not ( n5136 , n5135 );
not ( n5137 , n474 );
nand ( n5138 , n5137 , n456 );
nand ( n5139 , n5136 , n5138 , n901 );
nand ( n5140 , n5134 , n5139 );
nand ( n5141 , n5140 , n912 );
nand ( n5142 , n5131 , n5141 );
not ( n5143 , n2966 );
not ( n5144 , n4976 );
or ( n5145 , n5143 , n5144 );
not ( n5146 , n493 );
not ( n5147 , n2949 );
or ( n5148 , n5146 , n5147 );
nand ( n5149 , n739 , n4518 );
nand ( n5150 , n5148 , n5149 );
nand ( n5151 , n5150 , n2196 );
nand ( n5152 , n5145 , n5151 );
xor ( n5153 , n5142 , n5152 );
not ( n5154 , n3573 );
not ( n5155 , n5003 );
or ( n5156 , n5154 , n5155 );
not ( n5157 , n491 );
not ( n5158 , n3892 );
or ( n5159 , n5157 , n5158 );
not ( n5160 , n3892 );
nand ( n5161 , n5160 , n2613 );
nand ( n5162 , n5159 , n5161 );
nand ( n5163 , n5162 , n2606 );
nand ( n5164 , n5156 , n5163 );
xor ( n5165 , n5153 , n5164 );
xor ( n5166 , n5128 , n5165 );
xor ( n5167 , n5005 , n5014 );
and ( n5168 , n5167 , n4560 );
and ( n5169 , n5005 , n5014 );
or ( n5170 , n5168 , n5169 );
xor ( n5171 , n5166 , n5170 );
buf ( n5172 , n5048 );
and ( n5173 , n770 , n5172 );
not ( n5174 , n807 );
nor ( n5175 , n5174 , n782 );
nor ( n5176 , n5173 , n5175 );
xor ( n5177 , n5040 , n5050 );
and ( n5178 , n5177 , n5061 );
and ( n5179 , n5040 , n5050 );
or ( n5180 , n5178 , n5179 );
xor ( n5181 , n5176 , n5180 );
xor ( n5182 , n4968 , n4980 );
and ( n5183 , n5182 , n4994 );
and ( n5184 , n4968 , n4980 );
or ( n5185 , n5183 , n5184 );
xor ( n5186 , n5181 , n5185 );
xor ( n5187 , n5031 , n5035 );
and ( n5188 , n5187 , n5062 );
and ( n5189 , n5031 , n5035 );
or ( n5190 , n5188 , n5189 );
xor ( n5191 , n5186 , n5190 );
xor ( n5192 , n4995 , n5016 );
and ( n5193 , n5192 , n5021 );
and ( n5194 , n4995 , n5016 );
or ( n5195 , n5193 , n5194 );
xor ( n5196 , n5191 , n5195 );
xor ( n5197 , n5171 , n5196 );
xor ( n5198 , n5063 , n5067 );
and ( n5199 , n5198 , n5072 );
and ( n5200 , n5063 , n5067 );
or ( n5201 , n5199 , n5200 );
xor ( n5202 , n5197 , n5201 );
xor ( n5203 , n5022 , n5026 );
and ( n5204 , n5203 , n5073 );
and ( n5205 , n5022 , n5026 );
or ( n5206 , n5204 , n5205 );
nor ( n5207 , n5202 , n5206 );
not ( n5208 , n5207 );
not ( n5209 , n5208 );
or ( n5210 , n4155 , n4161 );
nand ( n5211 , n4624 , n5210 );
nor ( n5212 , n5074 , n5079 );
nor ( n5213 , n5211 , n5212 );
not ( n5214 , n5213 );
not ( n5215 , n4031 );
or ( n5216 , n5214 , n5215 );
not ( n5217 , n4963 );
not ( n5218 , n5081 );
or ( n5219 , n5217 , n5218 );
nand ( n5220 , n5219 , n5083 );
not ( n5221 , n5220 );
nand ( n5222 , n5216 , n5221 );
not ( n5223 , n5222 );
or ( n5224 , n5209 , n5223 );
nand ( n5225 , n5202 , n5206 );
buf ( n5226 , n5225 );
nand ( n5227 , n5224 , n5226 );
xor ( n5228 , n5118 , n5124 );
and ( n5229 , n5228 , n5127 );
and ( n5230 , n5118 , n5124 );
or ( n5231 , n5229 , n5230 );
not ( n5232 , n3573 );
not ( n5233 , n5162 );
or ( n5234 , n5232 , n5233 );
not ( n5235 , n491 );
not ( n5236 , n4971 );
or ( n5237 , n5235 , n5236 );
nand ( n5238 , n4974 , n2613 );
nand ( n5239 , n5237 , n5238 );
nand ( n5240 , n5239 , n2606 );
nand ( n5241 , n5234 , n5240 );
not ( n5242 , n1026 );
not ( n5243 , n813 );
not ( n5244 , n4093 );
or ( n5245 , n5243 , n5244 );
nand ( n5246 , n4090 , n495 );
nand ( n5247 , n5245 , n5246 );
not ( n5248 , n5247 );
or ( n5249 , n5242 , n5248 );
nand ( n5250 , n5116 , n1086 );
nand ( n5251 , n5249 , n5250 );
xor ( n5252 , n5241 , n5251 );
not ( n5253 , n4553 );
not ( n5254 , n5120 );
or ( n5255 , n5253 , n5254 );
not ( n5256 , n4999 );
xor ( n5257 , n489 , n5256 );
nand ( n5258 , n5257 , n4547 );
nand ( n5259 , n5255 , n5258 );
xor ( n5260 , n5252 , n5259 );
xor ( n5261 , n5231 , n5260 );
or ( n5262 , n807 , n770 );
nand ( n5263 , n5262 , n499 );
not ( n5264 , n5140 );
not ( n5265 , n893 );
or ( n5266 , n5264 , n5265 );
not ( n5267 , n497 );
not ( n5268 , n4077 );
or ( n5269 , n5267 , n5268 );
nand ( n5270 , n4076 , n901 );
nand ( n5271 , n5269 , n5270 );
nand ( n5272 , n5271 , n912 );
nand ( n5273 , n5266 , n5272 );
xor ( n5274 , n5263 , n5273 );
not ( n5275 , n2966 );
not ( n5276 , n5150 );
or ( n5277 , n5275 , n5276 );
not ( n5278 , n1043 );
not ( n5279 , n5278 );
not ( n5280 , n739 );
or ( n5281 , n5279 , n5280 );
nand ( n5282 , n1043 , n493 );
nand ( n5283 , n5281 , n5282 );
nand ( n5284 , n5283 , n2959 );
nand ( n5285 , n5277 , n5284 );
xor ( n5286 , n5274 , n5285 );
xor ( n5287 , n5261 , n5286 );
and ( n5288 , n982 , n489 );
not ( n5289 , n5176 );
xor ( n5290 , n5288 , n5289 );
xor ( n5291 , n5142 , n5152 );
and ( n5292 , n5291 , n5164 );
and ( n5293 , n5142 , n5152 );
or ( n5294 , n5292 , n5293 );
xor ( n5295 , n5290 , n5294 );
xor ( n5296 , n5176 , n5180 );
and ( n5297 , n5296 , n5185 );
and ( n5298 , n5176 , n5180 );
or ( n5299 , n5297 , n5298 );
xor ( n5300 , n5295 , n5299 );
xor ( n5301 , n5128 , n5165 );
and ( n5302 , n5301 , n5170 );
and ( n5303 , n5128 , n5165 );
or ( n5304 , n5302 , n5303 );
xor ( n5305 , n5300 , n5304 );
xor ( n5306 , n5287 , n5305 );
xor ( n5307 , n5186 , n5190 );
and ( n5308 , n5307 , n5195 );
and ( n5309 , n5186 , n5190 );
or ( n5310 , n5308 , n5309 );
xor ( n5311 , n5306 , n5310 );
xor ( n5312 , n5171 , n5196 );
and ( n5313 , n5312 , n5201 );
and ( n5314 , n5171 , n5196 );
or ( n5315 , n5313 , n5314 );
nand ( n5316 , n5311 , n5315 );
not ( n5317 , n5316 );
nor ( n5318 , n5315 , n5311 );
nor ( n5319 , n5317 , n5318 );
not ( n5320 , n455 );
and ( n5321 , n5319 , n5320 );
and ( n5322 , n5227 , n5321 );
not ( n5323 , n5227 );
not ( n5324 , n5315 );
not ( n5325 , n5311 );
nand ( n5326 , n5324 , n5325 );
nand ( n5327 , n5326 , n5316 );
and ( n5328 , n5327 , n5320 );
and ( n5329 , n5323 , n5328 );
nor ( n5330 , n5322 , n5329 );
not ( n5331 , n4910 );
nand ( n5332 , n4882 , n4880 );
or ( n5333 , n5332 , n4887 );
not ( n5334 , n5333 );
or ( n5335 , n5331 , n5334 );
nand ( n5336 , n4887 , n5332 );
nand ( n5337 , n5335 , n5336 );
not ( n5338 , n5337 );
not ( n5339 , n5338 );
not ( n5340 , n4896 );
not ( n5341 , n1630 );
or ( n5342 , n5340 , n5341 );
nand ( n5343 , n1634 , n499 );
nand ( n5344 , n5342 , n5343 );
xor ( n5345 , n4898 , n4904 );
and ( n5346 , n5345 , n4909 );
and ( n5347 , n4898 , n4904 );
or ( n5348 , n5346 , n5347 );
xor ( n5349 , n5344 , n5348 );
nor ( n5350 , n4819 , n4813 );
or ( n5351 , n5350 , n4827 );
nand ( n5352 , n4819 , n4813 );
nand ( n5353 , n5351 , n5352 );
xor ( n5354 , n5349 , n5353 );
not ( n5355 , n5354 );
not ( n5356 , n5355 );
or ( n5357 , n5339 , n5356 );
nand ( n5358 , n5354 , n5337 );
nand ( n5359 , n5357 , n5358 );
nand ( n5360 , n4918 , n4875 );
not ( n5361 , n5360 );
not ( n5362 , n4927 );
or ( n5363 , n5361 , n5362 );
not ( n5364 , n4918 );
nand ( n5365 , n5364 , n4874 );
nand ( n5366 , n5363 , n5365 );
not ( n5367 , n5366 );
xor ( n5368 , n5359 , n5367 );
not ( n5369 , n4859 );
not ( n5370 , n4853 );
or ( n5371 , n5369 , n5370 );
nand ( n5372 , n5371 , n4831 );
not ( n5373 , n4853 );
nand ( n5374 , n5373 , n4858 );
nand ( n5375 , n5372 , n5374 );
not ( n5376 , n5375 );
and ( n5377 , n516 , n489 );
not ( n5378 , n4839 );
not ( n5379 , n4835 );
or ( n5380 , n5378 , n5379 );
and ( n5381 , n514 , n489 );
not ( n5382 , n514 );
and ( n5383 , n5382 , n4046 );
nor ( n5384 , n5381 , n5383 );
nand ( n5385 , n2733 , n5384 );
nand ( n5386 , n5380 , n5385 );
xor ( n5387 , n5377 , n5386 );
not ( n5388 , n4902 );
buf ( n5389 , n1592 );
not ( n5390 , n5389 );
or ( n5391 , n5388 , n5390 );
buf ( n5392 , n1595 );
xor ( n5393 , n508 , n495 );
nand ( n5394 , n5392 , n5393 );
nand ( n5395 , n5391 , n5394 );
xor ( n5396 , n5387 , n5395 );
not ( n5397 , n4847 );
not ( n5398 , n4399 );
or ( n5399 , n5397 , n5398 );
not ( n5400 , n4848 );
not ( n5401 , n4400 );
or ( n5402 , n5400 , n5401 );
nand ( n5403 , n5402 , n4841 );
nand ( n5404 , n5399 , n5403 );
xor ( n5405 , n5396 , n5404 );
xor ( n5406 , n491 , n512 );
not ( n5407 , n5406 );
not ( n5408 , n2277 );
or ( n5409 , n5407 , n5408 );
nand ( n5410 , n2453 , n4845 , n3711 );
nand ( n5411 , n5409 , n5410 );
not ( n5412 , n4817 );
not ( n5413 , n2028 );
or ( n5414 , n5412 , n5413 );
xor ( n5415 , n510 , n493 );
nand ( n5416 , n5415 , n1561 );
nand ( n5417 , n5414 , n5416 );
xor ( n5418 , n5411 , n5417 );
not ( n5419 , n4824 );
not ( n5420 , n2083 );
or ( n5421 , n5419 , n5420 );
xor ( n5422 , n506 , n497 );
nand ( n5423 , n2086 , n5422 );
nand ( n5424 , n5421 , n5423 );
xor ( n5425 , n5418 , n5424 );
xor ( n5426 , n5405 , n5425 );
not ( n5427 , n5426 );
not ( n5428 , n5427 );
or ( n5429 , n5376 , n5428 );
not ( n5430 , n5375 );
nand ( n5431 , n5430 , n5426 );
nand ( n5432 , n5429 , n5431 );
xor ( n5433 , n5368 , n5432 );
not ( n5434 , n4928 );
or ( n5435 , n4936 , n4863 );
and ( n5436 , n5434 , n5435 );
and ( n5437 , n4936 , n4863 );
nor ( n5438 , n5436 , n5437 );
nand ( n5439 , n5433 , n5438 );
not ( n5440 , n5439 );
nand ( n5441 , n4937 , n4946 );
nand ( n5442 , n4352 , n5441 , n4486 );
nand ( n5443 , n3317 , n4347 , n4947 , n4486 );
not ( n5444 , n5441 );
not ( n5445 , n4484 );
or ( n5446 , n5444 , n5445 );
nand ( n5447 , n5446 , n4945 );
not ( n5448 , n5447 );
nand ( n5449 , n5442 , n5443 , n5448 );
not ( n5450 , n5449 );
or ( n5451 , n5440 , n5450 );
nor ( n5452 , n5433 , n5438 );
not ( n5453 , n5452 );
nand ( n5454 , n5451 , n5453 );
buf ( n5455 , n5354 );
not ( n5456 , n5455 );
not ( n5457 , n5456 );
not ( n5458 , n5426 );
or ( n5459 , n5457 , n5458 );
not ( n5460 , n5455 );
not ( n5461 , n5426 );
not ( n5462 , n5461 );
or ( n5463 , n5460 , n5462 );
nand ( n5464 , n5463 , n5337 );
nand ( n5465 , n5459 , n5464 );
not ( n5466 , n5465 );
not ( n5467 , n1718 );
not ( n5468 , n1630 );
not ( n5469 , n5468 );
or ( n5470 , n5467 , n5469 );
nand ( n5471 , n5470 , n499 );
not ( n5472 , n5415 );
not ( n5473 , n2028 );
or ( n5474 , n5472 , n5473 );
xor ( n5475 , n509 , n493 );
nand ( n5476 , n2031 , n5475 );
nand ( n5477 , n5474 , n5476 );
xor ( n5478 , n5471 , n5477 );
not ( n5479 , n5422 );
not ( n5480 , n2083 );
or ( n5481 , n5479 , n5480 );
xor ( n5482 , n505 , n497 );
nand ( n5483 , n2086 , n5482 );
nand ( n5484 , n5481 , n5483 );
xor ( n5485 , n5478 , n5484 );
not ( n5486 , n5406 );
buf ( n5487 , n2455 );
not ( n5488 , n5487 );
or ( n5489 , n5486 , n5488 );
xor ( n5490 , n491 , n511 );
nand ( n5491 , n2764 , n5490 );
nand ( n5492 , n5489 , n5491 );
not ( n5493 , n5384 );
not ( n5494 , n4835 );
or ( n5495 , n5493 , n5494 );
xor ( n5496 , n513 , n489 );
nand ( n5497 , n4838 , n5496 );
nand ( n5498 , n5495 , n5497 );
xor ( n5499 , n5492 , n5498 );
not ( n5500 , n5393 );
not ( n5501 , n5389 );
or ( n5502 , n5500 , n5501 );
xor ( n5503 , n507 , n495 );
nand ( n5504 , n5392 , n5503 );
nand ( n5505 , n5502 , n5504 );
xor ( n5506 , n5499 , n5505 );
xor ( n5507 , n5377 , n5386 );
and ( n5508 , n5507 , n5395 );
and ( n5509 , n5377 , n5386 );
or ( n5510 , n5508 , n5509 );
xor ( n5511 , n5506 , n5510 );
xnor ( n5512 , n5485 , n5511 );
not ( n5513 , n5512 );
not ( n5514 , n5513 );
xor ( n5515 , n5411 , n5417 );
and ( n5516 , n5515 , n5424 );
and ( n5517 , n5411 , n5417 );
or ( n5518 , n5516 , n5517 );
not ( n5519 , n5518 );
nand ( n5520 , n515 , n489 );
not ( n5521 , n5520 );
not ( n5522 , n5521 );
not ( n5523 , n5344 );
or ( n5524 , n5522 , n5523 );
or ( n5525 , n5521 , n5344 );
nand ( n5526 , n5524 , n5525 );
not ( n5527 , n5526 );
and ( n5528 , n5519 , n5527 );
and ( n5529 , n5518 , n5526 );
nor ( n5530 , n5528 , n5529 );
not ( n5531 , n5344 );
not ( n5532 , n5531 );
not ( n5533 , n5353 );
or ( n5534 , n5532 , n5533 );
or ( n5535 , n5353 , n5531 );
nand ( n5536 , n5535 , n5348 );
nand ( n5537 , n5534 , n5536 );
xor ( n5538 , n5530 , n5537 );
xor ( n5539 , n5396 , n5404 );
and ( n5540 , n5539 , n5425 );
and ( n5541 , n5396 , n5404 );
or ( n5542 , n5540 , n5541 );
xnor ( n5543 , n5538 , n5542 );
not ( n5544 , n5543 );
not ( n5545 , n5544 );
or ( n5546 , n5514 , n5545 );
nand ( n5547 , n5512 , n5543 );
nand ( n5548 , n5546 , n5547 );
not ( n5549 , n5548 );
or ( n5550 , n5466 , n5549 );
or ( n5551 , n5465 , n5548 );
nand ( n5552 , n5550 , n5551 );
not ( n5553 , n5552 );
not ( n5554 , n5430 );
not ( n5555 , n5427 );
not ( n5556 , n5359 );
not ( n5557 , n5556 );
or ( n5558 , n5555 , n5557 );
or ( n5559 , n5556 , n5461 );
nand ( n5560 , n5558 , n5559 );
not ( n5561 , n5560 );
or ( n5562 , n5554 , n5561 );
nand ( n5563 , n5562 , n5366 );
not ( n5564 , n5560 );
nand ( n5565 , n5564 , n5375 );
nand ( n5566 , n5563 , n5565 );
nand ( n5567 , n5553 , n5566 );
not ( n5568 , n5566 );
nand ( n5569 , n5568 , n5552 );
nand ( n5570 , n5567 , n5569 );
nor ( n5571 , n5570 , n5320 );
and ( n5572 , n5454 , n5571 );
not ( n5573 , n5454 );
and ( n5574 , n5570 , n455 );
and ( n5575 , n5573 , n5574 );
nor ( n5576 , n5572 , n5575 );
nand ( n5577 , n5330 , n5576 );
not ( n5578 , n5577 );
not ( n5579 , n5578 );
not ( n5580 , n5579 );
or ( n5581 , n5104 , n5580 );
not ( n5582 , n5577 );
nand ( n5583 , n5582 , n4018 );
nand ( n5584 , n5581 , n5583 );
not ( n5585 , n5584 );
or ( n5586 , n5103 , n5585 );
not ( n5587 , n551 );
not ( n5588 , n455 );
not ( n5589 , n5452 );
nand ( n5590 , n5589 , n5439 );
xnor ( n5591 , n5449 , n5590 );
not ( n5592 , n5591 );
or ( n5593 , n5588 , n5592 );
nand ( n5594 , n5208 , n5225 );
not ( n5595 , n5594 );
not ( n5596 , n5213 );
not ( n5597 , n4031 );
or ( n5598 , n5596 , n5597 );
nand ( n5599 , n5598 , n5221 );
not ( n5600 , n5599 );
or ( n5601 , n5595 , n5600 );
or ( n5602 , n5599 , n5594 );
nand ( n5603 , n5601 , n5602 );
not ( n5604 , n455 );
nand ( n5605 , n5603 , n5604 );
nand ( n5606 , n5593 , n5605 );
not ( n5607 , n5606 );
not ( n5608 , n5607 );
or ( n5609 , n5587 , n5608 );
not ( n5610 , n455 );
not ( n5611 , n5591 );
or ( n5612 , n5610 , n5611 );
nand ( n5613 , n5612 , n5605 );
buf ( n5614 , n5613 );
nand ( n5615 , n5614 , n4018 );
nand ( n5616 , n5609 , n5615 );
not ( n5617 , n552 );
nand ( n5618 , n5617 , n551 );
not ( n5619 , n5618 );
nand ( n5620 , n5616 , n5619 );
nand ( n5621 , n5586 , n5620 );
xor ( n5622 , n5102 , n5621 );
not ( n5623 , n2362 );
nand ( n5624 , n543 , n2698 );
nand ( n5625 , n2702 , n2123 );
nand ( n5626 , n5624 , n5625 );
not ( n5627 , n5626 );
or ( n5628 , n5623 , n5627 );
nand ( n5629 , n2360 , n714 );
nand ( n5630 , n5628 , n5629 );
not ( n5631 , n3017 );
not ( n5632 , n545 );
not ( n5633 , n3632 );
or ( n5634 , n5632 , n5633 );
nand ( n5635 , n3631 , n706 );
nand ( n5636 , n5634 , n5635 );
not ( n5637 , n5636 );
or ( n5638 , n5631 , n5637 );
nand ( n5639 , n3016 , n2376 );
nand ( n5640 , n5638 , n5639 );
xor ( n5641 , n5630 , n5640 );
xor ( n5642 , n3954 , n3989 );
and ( n5643 , n5642 , n4010 );
and ( n5644 , n3954 , n3989 );
or ( n5645 , n5643 , n5644 );
xor ( n5646 , n5641 , n5645 );
xor ( n5647 , n5622 , n5646 );
xor ( n5648 , n4805 , n5647 );
xor ( n5649 , n3950 , n4011 );
and ( n5650 , n5649 , n4642 );
and ( n5651 , n3950 , n4011 );
or ( n5652 , n5650 , n5651 );
not ( n5653 , n3298 );
not ( n5654 , n547 );
not ( n5655 , n4339 );
or ( n5656 , n5654 , n5655 );
nand ( n5657 , n4342 , n2369 );
nand ( n5658 , n5656 , n5657 );
not ( n5659 , n5658 );
or ( n5660 , n5653 , n5659 );
nand ( n5661 , n3948 , n3300 );
nand ( n5662 , n5660 , n5661 );
xor ( n5663 , n3991 , n3997 );
and ( n5664 , n5663 , n4009 );
and ( n5665 , n3991 , n3997 );
or ( n5666 , n5664 , n5665 );
not ( n5667 , n3955 );
not ( n5668 , n2122 );
not ( n5669 , n3023 );
or ( n5670 , n5668 , n5669 );
nand ( n5671 , n2125 , n541 );
nand ( n5672 , n5670 , n5671 );
not ( n5673 , n5672 );
or ( n5674 , n5667 , n5673 );
nand ( n5675 , n3985 , n3288 );
nand ( n5676 , n5674 , n5675 );
xor ( n5677 , n5666 , n5676 );
not ( n5678 , n3177 );
not ( n5679 , n3067 );
not ( n5680 , n5679 );
or ( n5681 , n5678 , n5680 );
nand ( n5682 , n537 , n3067 );
nand ( n5683 , n5681 , n5682 );
not ( n5684 , n5683 );
not ( n5685 , n3134 );
or ( n5686 , n5684 , n5685 );
nand ( n5687 , n3993 , n3182 );
nand ( n5688 , n5686 , n5687 );
and ( n5689 , n537 , n3149 );
xor ( n5690 , n5688 , n5689 );
not ( n5691 , n3026 );
not ( n5692 , n539 );
not ( n5693 , n3250 );
or ( n5694 , n5692 , n5693 );
not ( n5695 , n3249 );
not ( n5696 , n5695 );
nand ( n5697 , n5696 , n3069 );
nand ( n5698 , n5694 , n5697 );
not ( n5699 , n5698 );
or ( n5700 , n5691 , n5699 );
nand ( n5701 , n4005 , n3103 );
nand ( n5702 , n5700 , n5701 );
xor ( n5703 , n5690 , n5702 );
xor ( n5704 , n5677 , n5703 );
xor ( n5705 , n5662 , n5704 );
xor ( n5706 , n2364 , n3019 );
and ( n5707 , n5706 , n3293 );
and ( n5708 , n2364 , n3019 );
or ( n5709 , n5707 , n5708 );
xor ( n5710 , n5705 , n5709 );
xor ( n5711 , n5652 , n5710 );
xor ( n5712 , n4715 , n4726 );
and ( n5713 , n5712 , n4738 );
and ( n5714 , n4715 , n4726 );
or ( n5715 , n5713 , n5714 );
xor ( n5716 , n3105 , n3209 );
xor ( n5717 , n5716 , n3290 );
not ( n5718 , n3298 );
not ( n5719 , n3636 );
or ( n5720 , n5718 , n5719 );
nand ( n5721 , n4794 , n3300 );
nand ( n5722 , n5720 , n5721 );
xor ( n5723 , n5717 , n5722 );
not ( n5724 , n3214 );
not ( n5725 , n3284 );
or ( n5726 , n5724 , n5725 );
nand ( n5727 , n4748 , n3288 );
nand ( n5728 , n5726 , n5727 );
not ( n5729 , n714 );
not ( n5730 , n4766 );
or ( n5731 , n5729 , n5730 );
nand ( n5732 , n4724 , n2361 );
nand ( n5733 , n5731 , n5732 );
xor ( n5734 , n5728 , n5733 );
not ( n5735 , n2376 );
not ( n5736 , n545 );
not ( n5737 , n2122 );
not ( n5738 , n5737 );
or ( n5739 , n5736 , n5738 );
nand ( n5740 , n2122 , n706 );
nand ( n5741 , n5739 , n5740 );
not ( n5742 , n5741 );
or ( n5743 , n5735 , n5742 );
nand ( n5744 , n4736 , n3017 );
nand ( n5745 , n5743 , n5744 );
and ( n5746 , n5734 , n5745 );
and ( n5747 , n5728 , n5733 );
or ( n5748 , n5746 , n5747 );
and ( n5749 , n5723 , n5748 );
and ( n5750 , n5717 , n5722 );
or ( n5751 , n5749 , n5750 );
xor ( n5752 , n5715 , n5751 );
not ( n5753 , n5619 );
not ( n5754 , n5093 );
and ( n5755 , n5754 , n551 );
not ( n5756 , n5754 );
and ( n5757 , n5756 , n4018 );
or ( n5758 , n5755 , n5757 );
not ( n5759 , n5758 );
or ( n5760 , n5753 , n5759 );
nand ( n5761 , n5616 , n552 );
nand ( n5762 , n5760 , n5761 );
and ( n5763 , n5752 , n5762 );
and ( n5764 , n5715 , n5751 );
or ( n5765 , n5763 , n5764 );
xor ( n5766 , n5711 , n5765 );
xor ( n5767 , n5648 , n5766 );
xor ( n5768 , n5715 , n5751 );
xor ( n5769 , n5768 , n5762 );
not ( n5770 , n552 );
not ( n5771 , n5758 );
or ( n5772 , n5770 , n5771 );
and ( n5773 , n4635 , n551 );
not ( n5774 , n4635 );
and ( n5775 , n5774 , n4018 );
nor ( n5776 , n5773 , n5775 );
not ( n5777 , n5776 );
nand ( n5778 , n5777 , n5619 );
nand ( n5779 , n5772 , n5778 );
xor ( n5780 , n5717 , n5722 );
xor ( n5781 , n5780 , n5748 );
xor ( n5782 , n5779 , n5781 );
xor ( n5783 , n5728 , n5733 );
xor ( n5784 , n5783 , n5745 );
not ( n5785 , n4022 );
not ( n5786 , n549 );
not ( n5787 , n3632 );
or ( n5788 , n5786 , n5787 );
nand ( n5789 , n3631 , n4013 );
nand ( n5790 , n5788 , n5789 );
not ( n5791 , n5790 );
or ( n5792 , n5785 , n5791 );
nand ( n5793 , n4657 , n4020 );
nand ( n5794 , n5792 , n5793 );
xor ( n5795 , n5784 , n5794 );
not ( n5796 , n551 );
not ( n5797 , n4339 );
or ( n5798 , n5796 , n5797 );
buf ( n5799 , n4338 );
nand ( n5800 , n4018 , n5799 );
nand ( n5801 , n5798 , n5800 );
not ( n5802 , n5801 );
or ( n5803 , n5802 , n5618 );
or ( n5804 , n5776 , n5617 );
nand ( n5805 , n5803 , n5804 );
and ( n5806 , n5795 , n5805 );
and ( n5807 , n5784 , n5794 );
or ( n5808 , n5806 , n5807 );
and ( n5809 , n5782 , n5808 );
and ( n5810 , n5779 , n5781 );
or ( n5811 , n5809 , n5810 );
xor ( n5812 , n5769 , n5811 );
xor ( n5813 , n3294 , n4643 );
xor ( n5814 , n5813 , n4802 );
and ( n5815 , n5812 , n5814 );
and ( n5816 , n5769 , n5811 );
or ( n5817 , n5815 , n5816 );
nor ( n5818 , n5767 , n5817 );
not ( n5819 , n5818 );
nand ( n5820 , n5767 , n5817 );
nand ( n5821 , n5819 , n5820 );
not ( n5822 , n5821 );
xor ( n5823 , n5769 , n5811 );
xor ( n5824 , n5823 , n5814 );
xor ( n5825 , n4659 , n4739 );
xor ( n5826 , n5825 , n4799 );
not ( n5827 , n3017 );
not ( n5828 , n5741 );
or ( n5829 , n5827 , n5828 );
not ( n5830 , n545 );
not ( n5831 , n3979 );
buf ( n5832 , n5831 );
not ( n5833 , n5832 );
or ( n5834 , n5830 , n5833 );
nand ( n5835 , n3980 , n706 );
nand ( n5836 , n5834 , n5835 );
nand ( n5837 , n5836 , n2376 );
nand ( n5838 , n5829 , n5837 );
xor ( n5839 , n4696 , n4708 );
not ( n5840 , n3214 );
not ( n5841 , n4755 );
or ( n5842 , n5840 , n5841 );
and ( n5843 , n455 , n3137 );
not ( n5844 , n455 );
and ( n5845 , n5844 , n3147 );
nor ( n5846 , n5843 , n5845 );
and ( n5847 , n5846 , n541 );
not ( n5848 , n5846 );
and ( n5849 , n5848 , n3023 );
or ( n5850 , n5847 , n5849 );
nand ( n5851 , n5850 , n3288 );
nand ( n5852 , n5842 , n5851 );
xor ( n5853 , n5839 , n5852 );
and ( n5854 , n3128 , n3026 );
not ( n5855 , n3214 );
not ( n5856 , n5850 );
or ( n5857 , n5855 , n5856 );
not ( n5858 , n541 );
not ( n5859 , n3172 );
not ( n5860 , n5859 );
not ( n5861 , n5860 );
or ( n5862 , n5858 , n5861 );
nand ( n5863 , n5859 , n3023 );
nand ( n5864 , n5862 , n5863 );
nand ( n5865 , n5864 , n3288 );
nand ( n5866 , n5857 , n5865 );
xor ( n5867 , n5854 , n5866 );
not ( n5868 , n3214 );
not ( n5869 , n5864 );
or ( n5870 , n5868 , n5869 );
not ( n5871 , n541 );
not ( n5872 , n3190 );
or ( n5873 , n5871 , n5872 );
nand ( n5874 , n4704 , n3023 );
nand ( n5875 , n5873 , n5874 );
nand ( n5876 , n5875 , n3288 );
nand ( n5877 , n5870 , n5876 );
not ( n5878 , n542 );
nand ( n5879 , n5878 , n3203 );
and ( n5880 , n5879 , n543 );
not ( n5881 , n542 );
not ( n5882 , n3128 );
or ( n5883 , n5881 , n5882 );
nand ( n5884 , n5883 , n541 );
nor ( n5885 , n5880 , n5884 );
and ( n5886 , n5877 , n5885 );
and ( n5887 , n5867 , n5886 );
and ( n5888 , n5854 , n5866 );
or ( n5889 , n5887 , n5888 );
and ( n5890 , n5853 , n5889 );
and ( n5891 , n5839 , n5852 );
or ( n5892 , n5890 , n5891 );
xor ( n5893 , n5838 , n5892 );
xor ( n5894 , n4757 , n4759 );
xor ( n5895 , n5894 , n4775 );
and ( n5896 , n5893 , n5895 );
and ( n5897 , n5838 , n5892 );
or ( n5898 , n5896 , n5897 );
xor ( n5899 , n4742 , n4778 );
xor ( n5900 , n5899 , n4796 );
xor ( n5901 , n5898 , n5900 );
not ( n5902 , n3298 );
not ( n5903 , n4786 );
or ( n5904 , n5902 , n5903 );
not ( n5905 , n547 );
not ( n5906 , n2355 );
not ( n5907 , n5906 );
or ( n5908 , n5905 , n5907 );
not ( n5909 , n5906 );
nand ( n5910 , n5909 , n2369 );
nand ( n5911 , n5908 , n5910 );
nand ( n5912 , n5911 , n3300 );
nand ( n5913 , n5904 , n5912 );
not ( n5914 , n2361 );
not ( n5915 , n4773 );
or ( n5916 , n5914 , n5915 );
not ( n5917 , n543 );
not ( n5918 , n3067 );
or ( n5919 , n5917 , n5918 );
nand ( n5920 , n5679 , n2123 );
nand ( n5921 , n5919 , n5920 );
nand ( n5922 , n5921 , n714 );
nand ( n5923 , n5916 , n5922 );
not ( n5924 , n2376 );
not ( n5925 , n545 );
not ( n5926 , n3249 );
not ( n5927 , n5926 );
or ( n5928 , n5925 , n5927 );
nand ( n5929 , n3249 , n706 );
nand ( n5930 , n5928 , n5929 );
not ( n5931 , n5930 );
or ( n5932 , n5924 , n5931 );
nand ( n5933 , n5836 , n3017 );
nand ( n5934 , n5932 , n5933 );
xor ( n5935 , n5923 , n5934 );
xor ( n5936 , n5839 , n5852 );
xor ( n5937 , n5936 , n5889 );
and ( n5938 , n5935 , n5937 );
and ( n5939 , n5923 , n5934 );
or ( n5940 , n5938 , n5939 );
xor ( n5941 , n5913 , n5940 );
not ( n5942 , n4020 );
not ( n5943 , n5790 );
or ( n5944 , n5942 , n5943 );
not ( n5945 , n549 );
not ( n5946 , n3012 );
or ( n5947 , n5945 , n5946 );
nand ( n5948 , n4792 , n4013 );
nand ( n5949 , n5947 , n5948 );
nand ( n5950 , n5949 , n4022 );
nand ( n5951 , n5944 , n5950 );
and ( n5952 , n5941 , n5951 );
and ( n5953 , n5913 , n5940 );
or ( n5954 , n5952 , n5953 );
and ( n5955 , n5901 , n5954 );
and ( n5956 , n5898 , n5900 );
or ( n5957 , n5955 , n5956 );
xor ( n5958 , n5826 , n5957 );
xor ( n5959 , n5779 , n5781 );
xor ( n5960 , n5959 , n5808 );
and ( n5961 , n5958 , n5960 );
and ( n5962 , n5826 , n5957 );
or ( n5963 , n5961 , n5962 );
or ( n5964 , n5824 , n5963 );
not ( n5965 , n5964 );
xor ( n5966 , n5826 , n5957 );
xor ( n5967 , n5966 , n5960 );
buf ( n5968 , n5967 );
xor ( n5969 , n5784 , n5794 );
xor ( n5970 , n5969 , n5805 );
not ( n5971 , n552 );
not ( n5972 , n5801 );
or ( n5973 , n5971 , n5972 );
or ( n5974 , n551 , n3943 );
nand ( n5975 , n3943 , n551 );
nand ( n5976 , n5974 , n5975 );
nand ( n5977 , n5976 , n5619 );
nand ( n5978 , n5973 , n5977 );
xor ( n5979 , n5838 , n5892 );
xor ( n5980 , n5979 , n5895 );
xor ( n5981 , n5978 , n5980 );
not ( n5982 , n3300 );
not ( n5983 , n547 );
not ( n5984 , n2125 );
or ( n5985 , n5983 , n5984 );
nand ( n5986 , n2122 , n2369 );
nand ( n5987 , n5985 , n5986 );
not ( n5988 , n5987 );
or ( n5989 , n5982 , n5988 );
nand ( n5990 , n5911 , n3298 );
nand ( n5991 , n5989 , n5990 );
not ( n5992 , n2361 );
not ( n5993 , n5921 );
or ( n5994 , n5992 , n5993 );
not ( n5995 , n543 );
not ( n5996 , n3091 );
or ( n5997 , n5995 , n5996 );
nand ( n5998 , n3092 , n2123 );
nand ( n5999 , n5997 , n5998 );
nand ( n6000 , n5999 , n714 );
nand ( n6001 , n5994 , n6000 );
xor ( n6002 , n5854 , n5866 );
xor ( n6003 , n6002 , n5886 );
xor ( n6004 , n6001 , n6003 );
not ( n6005 , n3017 );
not ( n6006 , n5930 );
or ( n6007 , n6005 , n6006 );
not ( n6008 , n545 );
not ( n6009 , n4001 );
or ( n6010 , n6008 , n6009 );
nand ( n6011 , n3279 , n706 );
nand ( n6012 , n6010 , n6011 );
nand ( n6013 , n6012 , n2376 );
nand ( n6014 , n6007 , n6013 );
and ( n6015 , n6004 , n6014 );
and ( n6016 , n6001 , n6003 );
or ( n6017 , n6015 , n6016 );
xor ( n6018 , n5991 , n6017 );
not ( n6019 , n4020 );
not ( n6020 , n5949 );
or ( n6021 , n6019 , n6020 );
not ( n6022 , n549 );
not ( n6023 , n2697 );
not ( n6024 , n6023 );
or ( n6025 , n6022 , n6024 );
nand ( n6026 , n2697 , n4013 );
nand ( n6027 , n6025 , n6026 );
nand ( n6028 , n6027 , n4021 );
nand ( n6029 , n6021 , n6028 );
and ( n6030 , n6018 , n6029 );
and ( n6031 , n5991 , n6017 );
or ( n6032 , n6030 , n6031 );
and ( n6033 , n5981 , n6032 );
and ( n6034 , n5978 , n5980 );
or ( n6035 , n6033 , n6034 );
xor ( n6036 , n5970 , n6035 );
xor ( n6037 , n5898 , n5900 );
xor ( n6038 , n6037 , n5954 );
and ( n6039 , n6036 , n6038 );
and ( n6040 , n5970 , n6035 );
or ( n6041 , n6039 , n6040 );
nand ( n6042 , n5968 , n6041 );
xor ( n6043 , n5970 , n6035 );
xor ( n6044 , n6043 , n6038 );
xor ( n6045 , n5913 , n5940 );
xor ( n6046 , n6045 , n5951 );
not ( n6047 , n552 );
not ( n6048 , n5976 );
or ( n6049 , n6047 , n6048 );
buf ( n6050 , n5619 );
nand ( n6051 , n3632 , n6050 );
nand ( n6052 , n6049 , n6051 );
xor ( n6053 , n5923 , n5934 );
xor ( n6054 , n6053 , n5937 );
xor ( n6055 , n6052 , n6054 );
xor ( n6056 , n5885 , n5877 );
not ( n6057 , n2361 );
not ( n6058 , n5999 );
or ( n6059 , n6057 , n6058 );
not ( n6060 , n543 );
not ( n6061 , n5846 );
not ( n6062 , n6061 );
not ( n6063 , n6062 );
or ( n6064 , n6060 , n6063 );
nand ( n6065 , n3149 , n2123 );
nand ( n6066 , n6064 , n6065 );
nand ( n6067 , n6066 , n714 );
nand ( n6068 , n6059 , n6067 );
xor ( n6069 , n6056 , n6068 );
and ( n6070 , n3128 , n3214 );
not ( n6071 , n2361 );
not ( n6072 , n6066 );
or ( n6073 , n6071 , n6072 );
not ( n6074 , n543 );
not ( n6075 , n5860 );
or ( n6076 , n6074 , n6075 );
nand ( n6077 , n5859 , n2123 );
nand ( n6078 , n6076 , n6077 );
nand ( n6079 , n6078 , n714 );
nand ( n6080 , n6073 , n6079 );
xor ( n6081 , n6070 , n6080 );
not ( n6082 , n544 );
nand ( n6083 , n6082 , n3190 );
and ( n6084 , n6083 , n545 );
not ( n6085 , n544 );
not ( n6086 , n3199 );
or ( n6087 , n6085 , n6086 );
nand ( n6088 , n6087 , n543 );
nor ( n6089 , n6084 , n6088 );
not ( n6090 , n2361 );
not ( n6091 , n6078 );
or ( n6092 , n6090 , n6091 );
not ( n6093 , n543 );
not ( n6094 , n3190 );
or ( n6095 , n6093 , n6094 );
nand ( n6096 , n3199 , n2123 );
nand ( n6097 , n6095 , n6096 );
nand ( n6098 , n6097 , n714 );
nand ( n6099 , n6092 , n6098 );
and ( n6100 , n6089 , n6099 );
and ( n6101 , n6081 , n6100 );
and ( n6102 , n6070 , n6080 );
or ( n6103 , n6101 , n6102 );
and ( n6104 , n6069 , n6103 );
and ( n6105 , n6056 , n6068 );
or ( n6106 , n6104 , n6105 );
not ( n6107 , n3298 );
not ( n6108 , n5987 );
or ( n6109 , n6107 , n6108 );
not ( n6110 , n547 );
not ( n6111 , n4720 );
or ( n6112 , n6110 , n6111 );
not ( n6113 , n5832 );
nand ( n6114 , n6113 , n2369 );
nand ( n6115 , n6112 , n6114 );
nand ( n6116 , n6115 , n3299 );
nand ( n6117 , n6109 , n6116 );
xor ( n6118 , n6106 , n6117 );
xor ( n6119 , n6001 , n6003 );
xor ( n6120 , n6119 , n6014 );
and ( n6121 , n6118 , n6120 );
and ( n6122 , n6106 , n6117 );
or ( n6123 , n6121 , n6122 );
and ( n6124 , n6055 , n6123 );
and ( n6125 , n6052 , n6054 );
or ( n6126 , n6124 , n6125 );
xor ( n6127 , n6046 , n6126 );
xor ( n6128 , n5978 , n5980 );
xor ( n6129 , n6128 , n6032 );
and ( n6130 , n6127 , n6129 );
and ( n6131 , n6046 , n6126 );
or ( n6132 , n6130 , n6131 );
nand ( n6133 , n6044 , n6132 );
not ( n6134 , n6133 );
or ( n6135 , n5967 , n6041 );
nand ( n6136 , n6134 , n6135 );
xor ( n6137 , n6046 , n6126 );
xor ( n6138 , n6137 , n6129 );
not ( n6139 , n6138 );
not ( n6140 , n4020 );
not ( n6141 , n6027 );
or ( n6142 , n6140 , n6141 );
nand ( n6143 , n4732 , n549 );
not ( n6144 , n6143 );
nand ( n6145 , n2355 , n4013 );
not ( n6146 , n6145 );
or ( n6147 , n6144 , n6146 );
nand ( n6148 , n6147 , n4021 );
nand ( n6149 , n6142 , n6148 );
not ( n6150 , n551 );
not ( n6151 , n3012 );
or ( n6152 , n6150 , n6151 );
nand ( n6153 , n3011 , n4018 );
nand ( n6154 , n6152 , n6153 );
nand ( n6155 , n6154 , n5619 );
not ( n6156 , n3630 );
nor ( n6157 , n4018 , n5617 );
nand ( n6158 , n6156 , n6157 );
nor ( n6159 , n5617 , n551 );
nand ( n6160 , n3631 , n6159 );
nand ( n6161 , n6155 , n6158 , n6160 );
xor ( n6162 , n6149 , n6161 );
not ( n6163 , n3017 );
not ( n6164 , n6012 );
or ( n6165 , n6163 , n6164 );
not ( n6166 , n545 );
not ( n6167 , n3064 );
or ( n6168 , n6166 , n6167 );
nand ( n6169 , n5679 , n706 );
nand ( n6170 , n6168 , n6169 );
nand ( n6171 , n6170 , n2376 );
nand ( n6172 , n6165 , n6171 );
not ( n6173 , n3299 );
not ( n6174 , n547 );
not ( n6175 , n5695 );
or ( n6176 , n6174 , n6175 );
nand ( n6177 , n3249 , n2369 );
nand ( n6178 , n6176 , n6177 );
not ( n6179 , n6178 );
or ( n6180 , n6173 , n6179 );
nand ( n6181 , n6115 , n3298 );
nand ( n6182 , n6180 , n6181 );
xor ( n6183 , n6172 , n6182 );
xor ( n6184 , n6056 , n6068 );
xor ( n6185 , n6184 , n6103 );
and ( n6186 , n6183 , n6185 );
and ( n6187 , n6172 , n6182 );
or ( n6188 , n6186 , n6187 );
and ( n6189 , n6162 , n6188 );
and ( n6190 , n6149 , n6161 );
or ( n6191 , n6189 , n6190 );
xor ( n6192 , n5991 , n6017 );
xor ( n6193 , n6192 , n6029 );
xor ( n6194 , n6191 , n6193 );
xor ( n6195 , n6052 , n6054 );
xor ( n6196 , n6195 , n6123 );
and ( n6197 , n6194 , n6196 );
and ( n6198 , n6191 , n6193 );
or ( n6199 , n6197 , n6198 );
not ( n6200 , n6199 );
nand ( n6201 , n6139 , n6200 );
not ( n6202 , n6201 );
xor ( n6203 , n6191 , n6193 );
xor ( n6204 , n6203 , n6196 );
not ( n6205 , n6204 );
xor ( n6206 , n6106 , n6117 );
xor ( n6207 , n6206 , n6120 );
not ( n6208 , n4021 );
not ( n6209 , n2122 );
not ( n6210 , n4013 );
or ( n6211 , n6209 , n6210 );
not ( n6212 , n2122 );
nand ( n6213 , n6212 , n549 );
nand ( n6214 , n6211 , n6213 );
not ( n6215 , n6214 );
or ( n6216 , n6208 , n6215 );
not ( n6217 , n6143 );
not ( n6218 , n6145 );
or ( n6219 , n6217 , n6218 );
buf ( n6220 , n4020 );
nand ( n6221 , n6219 , n6220 );
nand ( n6222 , n6216 , n6221 );
not ( n6223 , n552 );
not ( n6224 , n6154 );
or ( n6225 , n6223 , n6224 );
not ( n6226 , n551 );
not ( n6227 , n6023 );
or ( n6228 , n6226 , n6227 );
nand ( n6229 , n2697 , n4018 );
nand ( n6230 , n6228 , n6229 );
nand ( n6231 , n6230 , n5619 );
nand ( n6232 , n6225 , n6231 );
xor ( n6233 , n6222 , n6232 );
not ( n6234 , n3017 );
not ( n6235 , n6170 );
or ( n6236 , n6234 , n6235 );
not ( n6237 , n545 );
not ( n6238 , n3093 );
or ( n6239 , n6237 , n6238 );
nand ( n6240 , n3092 , n706 );
nand ( n6241 , n6239 , n6240 );
nand ( n6242 , n6241 , n2376 );
nand ( n6243 , n6236 , n6242 );
xor ( n6244 , n6070 , n6080 );
xor ( n6245 , n6244 , n6100 );
xor ( n6246 , n6243 , n6245 );
not ( n6247 , n3298 );
not ( n6248 , n6178 );
or ( n6249 , n6247 , n6248 );
and ( n6250 , n3279 , n2369 );
not ( n6251 , n3279 );
and ( n6252 , n6251 , n547 );
or ( n6253 , n6250 , n6252 );
nand ( n6254 , n6253 , n3299 );
nand ( n6255 , n6249 , n6254 );
and ( n6256 , n6246 , n6255 );
and ( n6257 , n6243 , n6245 );
or ( n6258 , n6256 , n6257 );
and ( n6259 , n6233 , n6258 );
and ( n6260 , n6222 , n6232 );
or ( n6261 , n6259 , n6260 );
xor ( n6262 , n6207 , n6261 );
xor ( n6263 , n6149 , n6161 );
xor ( n6264 , n6263 , n6188 );
and ( n6265 , n6262 , n6264 );
and ( n6266 , n6207 , n6261 );
or ( n6267 , n6265 , n6266 );
not ( n6268 , n6267 );
nand ( n6269 , n6205 , n6268 );
xor ( n6270 , n6172 , n6182 );
xor ( n6271 , n6270 , n6185 );
xor ( n6272 , n6089 , n6099 );
not ( n6273 , n3017 );
not ( n6274 , n6241 );
or ( n6275 , n6273 , n6274 );
not ( n6276 , n545 );
not ( n6277 , n6062 );
or ( n6278 , n6276 , n6277 );
nand ( n6279 , n3149 , n706 );
nand ( n6280 , n6278 , n6279 );
nand ( n6281 , n6280 , n2376 );
nand ( n6282 , n6275 , n6281 );
xor ( n6283 , n6272 , n6282 );
not ( n6284 , n3298 );
not ( n6285 , n6253 );
or ( n6286 , n6284 , n6285 );
not ( n6287 , n547 );
not ( n6288 , n3064 );
or ( n6289 , n6287 , n6288 );
nand ( n6290 , n3063 , n2369 );
nand ( n6291 , n6289 , n6290 );
nand ( n6292 , n6291 , n3299 );
nand ( n6293 , n6286 , n6292 );
and ( n6294 , n6283 , n6293 );
and ( n6295 , n6272 , n6282 );
or ( n6296 , n6294 , n6295 );
not ( n6297 , n6214 );
not ( n6298 , n6220 );
or ( n6299 , n6297 , n6298 );
not ( n6300 , n549 );
not ( n6301 , n3979 );
not ( n6302 , n6301 );
or ( n6303 , n6300 , n6302 );
nand ( n6304 , n3980 , n4013 );
nand ( n6305 , n6303 , n6304 );
nand ( n6306 , n6305 , n4021 );
nand ( n6307 , n6299 , n6306 );
xor ( n6308 , n6296 , n6307 );
not ( n6309 , n552 );
not ( n6310 , n6230 );
or ( n6311 , n6309 , n6310 );
nand ( n6312 , n2356 , n6050 );
nand ( n6313 , n6311 , n6312 );
and ( n6314 , n6308 , n6313 );
and ( n6315 , n6296 , n6307 );
or ( n6316 , n6314 , n6315 );
xor ( n6317 , n6271 , n6316 );
xor ( n6318 , n6222 , n6232 );
xor ( n6319 , n6318 , n6258 );
xor ( n6320 , n6317 , n6319 );
not ( n6321 , n6320 );
xor ( n6322 , n6243 , n6245 );
xor ( n6323 , n6322 , n6255 );
and ( n6324 , n3128 , n2361 );
not ( n6325 , n3017 );
not ( n6326 , n6280 );
or ( n6327 , n6325 , n6326 );
not ( n6328 , n545 );
not ( n6329 , n5860 );
or ( n6330 , n6328 , n6329 );
nand ( n6331 , n5859 , n706 );
nand ( n6332 , n6330 , n6331 );
nand ( n6333 , n6332 , n2376 );
nand ( n6334 , n6327 , n6333 );
xor ( n6335 , n6324 , n6334 );
not ( n6336 , n545 );
not ( n6337 , n3190 );
or ( n6338 , n6336 , n6337 );
nand ( n6339 , n4704 , n706 );
nand ( n6340 , n6338 , n6339 );
nand ( n6341 , n6340 , n2376 );
nand ( n6342 , n6332 , n3017 );
nand ( n6343 , n6341 , n6342 );
nand ( n6344 , n2365 , n3203 );
and ( n6345 , n6344 , n547 );
not ( n6346 , n546 );
not ( n6347 , n4704 );
or ( n6348 , n6346 , n6347 );
nand ( n6349 , n6348 , n545 );
nor ( n6350 , n6345 , n6349 );
and ( n6351 , n6343 , n6350 );
and ( n6352 , n6335 , n6351 );
and ( n6353 , n6324 , n6334 );
or ( n6354 , n6352 , n6353 );
not ( n6355 , n4020 );
not ( n6356 , n6305 );
or ( n6357 , n6355 , n6356 );
and ( n6358 , n3249 , n4013 );
not ( n6359 , n3249 );
and ( n6360 , n6359 , n549 );
or ( n6361 , n6358 , n6360 );
nand ( n6362 , n6361 , n4021 );
nand ( n6363 , n6357 , n6362 );
xor ( n6364 , n6354 , n6363 );
not ( n6365 , n5619 );
not ( n6366 , n2125 );
or ( n6367 , n6365 , n6366 );
and ( n6368 , n2355 , n6159 );
not ( n6369 , n2355 );
and ( n6370 , n6369 , n6157 );
nor ( n6371 , n6368 , n6370 );
nand ( n6372 , n6367 , n6371 );
and ( n6373 , n6364 , n6372 );
and ( n6374 , n6354 , n6363 );
or ( n6375 , n6373 , n6374 );
xor ( n6376 , n6323 , n6375 );
xor ( n6377 , n6296 , n6307 );
xor ( n6378 , n6377 , n6313 );
and ( n6379 , n6376 , n6378 );
and ( n6380 , n6323 , n6375 );
or ( n6381 , n6379 , n6380 );
not ( n6382 , n6381 );
nand ( n6383 , n6321 , n6382 );
not ( n6384 , n6383 );
not ( n6385 , n4020 );
not ( n6386 , n549 );
not ( n6387 , n3280 );
or ( n6388 , n6386 , n6387 );
nand ( n6389 , n3279 , n4013 );
nand ( n6390 , n6388 , n6389 );
not ( n6391 , n6390 );
or ( n6392 , n6385 , n6391 );
and ( n6393 , n3063 , n4013 );
not ( n6394 , n3063 );
and ( n6395 , n6394 , n549 );
or ( n6396 , n6393 , n6395 );
nand ( n6397 , n6396 , n4021 );
nand ( n6398 , n6392 , n6397 );
not ( n6399 , n551 );
not ( n6400 , n5831 );
or ( n6401 , n6399 , n6400 );
nand ( n6402 , n4018 , n3979 );
nand ( n6403 , n6401 , n6402 );
not ( n6404 , n6403 );
not ( n6405 , n552 );
or ( n6406 , n6404 , n6405 );
nand ( n6407 , n5926 , n6050 );
nand ( n6408 , n6406 , n6407 );
xor ( n6409 , n6398 , n6408 );
xor ( n6410 , n6343 , n6350 );
not ( n6411 , n3298 );
not ( n6412 , n547 );
not ( n6413 , n3091 );
or ( n6414 , n6412 , n6413 );
nand ( n6415 , n2369 , n3092 );
nand ( n6416 , n6414 , n6415 );
not ( n6417 , n6416 );
or ( n6418 , n6411 , n6417 );
not ( n6419 , n2369 );
not ( n6420 , n6061 );
or ( n6421 , n6419 , n6420 );
nand ( n6422 , n5846 , n547 );
nand ( n6423 , n6421 , n6422 );
nand ( n6424 , n6423 , n3299 );
nand ( n6425 , n6418 , n6424 );
xor ( n6426 , n6410 , n6425 );
and ( n6427 , n3199 , n3017 );
not ( n6428 , n3298 );
not ( n6429 , n6423 );
or ( n6430 , n6428 , n6429 );
and ( n6431 , n5859 , n2369 );
not ( n6432 , n5859 );
and ( n6433 , n6432 , n547 );
or ( n6434 , n6431 , n6433 );
nand ( n6435 , n3299 , n6434 );
nand ( n6436 , n6430 , n6435 );
xor ( n6437 , n6427 , n6436 );
and ( n6438 , n6434 , n3298 );
nand ( n6439 , n2369 , n4704 );
nand ( n6440 , n4703 , n547 );
and ( n6441 , n6439 , n6440 );
not ( n6442 , n3299 );
nor ( n6443 , n6441 , n6442 );
nor ( n6444 , n6438 , n6443 );
and ( n6445 , n3128 , n548 );
nor ( n6446 , n6445 , n2369 );
not ( n6447 , n3295 );
not ( n6448 , n3190 );
or ( n6449 , n6447 , n6448 );
nand ( n6450 , n6449 , n549 );
nand ( n6451 , n6446 , n6450 );
nor ( n6452 , n6444 , n6451 );
and ( n6453 , n6437 , n6452 );
and ( n6454 , n6427 , n6436 );
or ( n6455 , n6453 , n6454 );
xor ( n6456 , n6426 , n6455 );
xor ( n6457 , n6409 , n6456 );
not ( n6458 , n4020 );
not ( n6459 , n6396 );
or ( n6460 , n6458 , n6459 );
and ( n6461 , n3092 , n4013 );
not ( n6462 , n3092 );
and ( n6463 , n6462 , n549 );
or ( n6464 , n6461 , n6463 );
nand ( n6465 , n6464 , n4021 );
nand ( n6466 , n6460 , n6465 );
xor ( n6467 , n6427 , n6436 );
xor ( n6468 , n6467 , n6452 );
xor ( n6469 , n6466 , n6468 );
nand ( n6470 , n4001 , n5619 );
nand ( n6471 , n5695 , n6157 );
nand ( n6472 , n3249 , n6159 );
nand ( n6473 , n6470 , n6471 , n6472 );
and ( n6474 , n6469 , n6473 );
and ( n6475 , n6466 , n6468 );
or ( n6476 , n6474 , n6475 );
or ( n6477 , n6457 , n6476 );
xor ( n6478 , n6466 , n6468 );
xor ( n6479 , n6478 , n6473 );
not ( n6480 , n6479 );
not ( n6481 , n6451 );
nor ( n6482 , n6444 , n6481 );
not ( n6483 , n6482 );
nand ( n6484 , n6481 , n6444 );
nand ( n6485 , n6483 , n6484 );
not ( n6486 , n4020 );
not ( n6487 , n6464 );
or ( n6488 , n6486 , n6487 );
and ( n6489 , n6062 , n549 );
not ( n6490 , n6062 );
and ( n6491 , n6490 , n4013 );
or ( n6492 , n6489 , n6491 );
nand ( n6493 , n6492 , n4021 );
nand ( n6494 , n6488 , n6493 );
xor ( n6495 , n6485 , n6494 );
not ( n6496 , n3279 );
nand ( n6497 , n6496 , n6157 );
and ( n6498 , n4018 , n3062 );
not ( n6499 , n4018 );
and ( n6500 , n6499 , n3063 );
nor ( n6501 , n6498 , n6500 );
nand ( n6502 , n6501 , n5619 );
nand ( n6503 , n3279 , n6159 );
nand ( n6504 , n6497 , n6502 , n6503 );
and ( n6505 , n6495 , n6504 );
and ( n6506 , n6485 , n6494 );
or ( n6507 , n6505 , n6506 );
not ( n6508 , n6507 );
nand ( n6509 , n6480 , n6508 );
not ( n6510 , n6509 );
xor ( n6511 , n6485 , n6494 );
xor ( n6512 , n6511 , n6504 );
and ( n6513 , n3128 , n3298 );
not ( n6514 , n4020 );
not ( n6515 , n6492 );
or ( n6516 , n6514 , n6515 );
not ( n6517 , n549 );
not ( n6518 , n3173 );
or ( n6519 , n6517 , n6518 );
not ( n6520 , n5860 );
nand ( n6521 , n6520 , n4013 );
nand ( n6522 , n6519 , n6521 );
nand ( n6523 , n6522 , n4021 );
nand ( n6524 , n6516 , n6523 );
xor ( n6525 , n6513 , n6524 );
not ( n6526 , n6220 );
not ( n6527 , n6522 );
or ( n6528 , n6526 , n6527 );
and ( n6529 , n4013 , n3199 );
not ( n6530 , n4013 );
and ( n6531 , n6530 , n4703 );
nor ( n6532 , n6529 , n6531 );
not ( n6533 , n4021 );
or ( n6534 , n6532 , n6533 );
nand ( n6535 , n6528 , n6534 );
not ( n6536 , n4014 );
not ( n6537 , n3203 );
or ( n6538 , n6536 , n6537 );
nand ( n6539 , n6538 , n551 );
and ( n6540 , n3199 , n550 );
nor ( n6541 , n6540 , n4013 );
and ( n6542 , n6539 , n6541 );
nand ( n6543 , n6535 , n6542 );
not ( n6544 , n6543 );
and ( n6545 , n6525 , n6544 );
and ( n6546 , n6513 , n6524 );
or ( n6547 , n6545 , n6546 );
or ( n6548 , n6512 , n6547 );
not ( n6549 , n6548 );
not ( n6550 , n552 );
not ( n6551 , n4018 );
nor ( n6552 , n6551 , n3093 );
not ( n6553 , n6552 );
or ( n6554 , n6550 , n6553 );
and ( n6555 , n3093 , n552 , n551 );
and ( n6556 , n4670 , n6050 );
nor ( n6557 , n6555 , n6556 );
nand ( n6558 , n6554 , n6557 );
not ( n6559 , n6558 );
or ( n6560 , n6542 , n6535 );
nand ( n6561 , n6560 , n6543 );
nand ( n6562 , n6559 , n6561 );
not ( n6563 , n6220 );
nor ( n6564 , n3190 , n6563 );
not ( n6565 , n551 );
not ( n6566 , n5860 );
or ( n6567 , n6565 , n6566 );
nand ( n6568 , n5859 , n4018 );
nand ( n6569 , n6567 , n6568 );
and ( n6570 , n6569 , n552 );
and ( n6571 , n3203 , n6050 );
nor ( n6572 , n6570 , n6571 );
nand ( n6573 , n3128 , n552 );
nand ( n6574 , n551 , n6573 );
nor ( n6575 , n6572 , n6574 );
xor ( n6576 , n6564 , n6575 );
nand ( n6577 , n4670 , n6157 );
nand ( n6578 , n3149 , n6159 );
nand ( n6579 , n6569 , n5619 );
nand ( n6580 , n6577 , n6578 , n6579 );
and ( n6581 , n6576 , n6580 );
or ( n6583 , n6581 , C0 );
and ( n6584 , n6562 , n6583 );
not ( n6585 , n6558 );
nor ( n6586 , n6585 , n6561 );
nor ( n6587 , n6584 , n6586 );
xor ( n6588 , n6513 , n6524 );
xor ( n6589 , n6588 , n6544 );
not ( n6590 , n552 );
not ( n6591 , n6501 );
or ( n6592 , n6590 , n6591 );
nand ( n6593 , n3093 , n6050 );
nand ( n6594 , n6592 , n6593 );
nor ( n6595 , n6589 , n6594 );
or ( n6596 , n6587 , n6595 );
nand ( n6597 , n6589 , n6594 );
nand ( n6598 , n6596 , n6597 );
not ( n6599 , n6598 );
or ( n6600 , n6549 , n6599 );
nand ( n6601 , n6512 , n6547 );
nand ( n6602 , n6600 , n6601 );
not ( n6603 , n6602 );
or ( n6604 , n6510 , n6603 );
nand ( n6605 , n6479 , n6507 );
nand ( n6606 , n6604 , n6605 );
and ( n6607 , n6477 , n6606 );
and ( n6608 , n6457 , n6476 );
nor ( n6609 , n6607 , n6608 );
not ( n6610 , n2122 );
nand ( n6611 , n6610 , n6157 );
not ( n6612 , n5737 );
nand ( n6613 , n6612 , n6159 );
nand ( n6614 , n6403 , n5619 );
nand ( n6615 , n6611 , n6613 , n6614 );
xor ( n6616 , n6410 , n6425 );
and ( n6617 , n6616 , n6455 );
and ( n6618 , n6410 , n6425 );
or ( n6619 , n6617 , n6618 );
xor ( n6620 , n6615 , n6619 );
not ( n6621 , n3298 );
not ( n6622 , n6291 );
or ( n6623 , n6621 , n6622 );
nand ( n6624 , n6416 , n3299 );
nand ( n6625 , n6623 , n6624 );
xor ( n6626 , n6324 , n6334 );
xor ( n6627 , n6626 , n6351 );
xor ( n6628 , n6625 , n6627 );
not ( n6629 , n4020 );
not ( n6630 , n6361 );
or ( n6631 , n6629 , n6630 );
nand ( n6632 , n6390 , n4021 );
nand ( n6633 , n6631 , n6632 );
xor ( n6634 , n6628 , n6633 );
xor ( n6635 , n6620 , n6634 );
xor ( n6636 , n6398 , n6408 );
and ( n6637 , n6636 , n6456 );
and ( n6638 , n6398 , n6408 );
or ( n6639 , n6637 , n6638 );
nor ( n6640 , n6635 , n6639 );
or ( n6641 , n6609 , n6640 );
nand ( n6642 , n6639 , n6635 );
nand ( n6643 , n6641 , n6642 );
xor ( n6644 , n6272 , n6282 );
xor ( n6645 , n6644 , n6293 );
xor ( n6646 , n6625 , n6627 );
and ( n6647 , n6646 , n6633 );
and ( n6648 , n6625 , n6627 );
or ( n6649 , n6647 , n6648 );
xor ( n6650 , n6645 , n6649 );
xor ( n6651 , n6354 , n6363 );
xor ( n6652 , n6651 , n6372 );
xor ( n6653 , n6650 , n6652 );
not ( n6654 , n6653 );
xor ( n6655 , n6615 , n6619 );
and ( n6656 , n6655 , n6634 );
and ( n6657 , n6615 , n6619 );
or ( n6658 , n6656 , n6657 );
not ( n6659 , n6658 );
nand ( n6660 , n6654 , n6659 );
and ( n6661 , n6643 , n6660 );
and ( n6662 , n6653 , n6658 );
nor ( n6663 , n6661 , n6662 );
xor ( n6664 , n6323 , n6375 );
xor ( n6665 , n6664 , n6378 );
xor ( n6666 , n6645 , n6649 );
and ( n6667 , n6666 , n6652 );
and ( n6668 , n6645 , n6649 );
or ( n6669 , n6667 , n6668 );
nor ( n6670 , n6665 , n6669 );
or ( n6671 , n6663 , n6670 );
nand ( n6672 , n6665 , n6669 );
nand ( n6673 , n6671 , n6672 );
not ( n6674 , n6673 );
or ( n6675 , n6384 , n6674 );
buf ( n6676 , n6320 );
nand ( n6677 , n6676 , n6381 );
nand ( n6678 , n6675 , n6677 );
xor ( n6679 , n6207 , n6261 );
xor ( n6680 , n6679 , n6264 );
not ( n6681 , n6680 );
xor ( n6682 , n6271 , n6316 );
and ( n6683 , n6682 , n6319 );
and ( n6684 , n6271 , n6316 );
or ( n6685 , n6683 , n6684 );
not ( n6686 , n6685 );
nand ( n6687 , n6681 , n6686 );
nand ( n6688 , n6269 , n6678 , n6687 );
not ( n6689 , n6204 );
nand ( n6690 , n6689 , n6268 );
not ( n6691 , n6680 );
nor ( n6692 , n6691 , n6686 );
nand ( n6693 , n6690 , n6692 );
buf ( n6694 , n6204 );
nand ( n6695 , n6694 , n6267 );
nand ( n6696 , n6688 , n6693 , n6695 );
not ( n6697 , n6696 );
or ( n6698 , n6202 , n6697 );
nand ( n6699 , n6199 , n6138 );
nand ( n6700 , n6698 , n6699 );
or ( n6701 , n6044 , n6132 );
nand ( n6702 , n6135 , n6700 , n6701 );
nand ( n6703 , n6042 , n6136 , n6702 );
not ( n6704 , n6703 );
or ( n6705 , n5965 , n6704 );
nand ( n6706 , n5824 , n5963 );
nand ( n6707 , n6705 , n6706 );
not ( n6708 , n6707 );
or ( n6709 , n5822 , n6708 );
or ( n6710 , n5821 , n6707 );
nand ( n6711 , n6709 , n6710 );
nand ( n6712 , n6711 , n454 );
not ( n6713 , n492 );
nand ( n6714 , n6713 , n493 );
and ( n6715 , n491 , n492 );
nor ( n6716 , n491 , n492 );
nor ( n6717 , n6715 , n6716 );
nand ( n6718 , n739 , n492 );
and ( n6719 , n6714 , n6717 , n6718 );
not ( n6720 , n6719 );
xor ( n6721 , n470 , n471 );
and ( n6722 , n6721 , n536 );
xor ( n6723 , n471 , n535 );
not ( n6724 , n6723 );
not ( n6725 , n472 );
nand ( n6726 , n6725 , n471 );
not ( n6727 , n6726 );
not ( n6728 , n6727 );
or ( n6729 , n6724 , n6728 );
xor ( n6730 , n534 , n471 );
nand ( n6731 , n6730 , n472 );
nand ( n6732 , n6729 , n6731 );
or ( n6733 , n6722 , n6732 );
not ( n6734 , n6733 );
not ( n6735 , n536 );
and ( n6736 , n471 , n6735 );
not ( n6737 , n471 );
and ( n6738 , n6737 , n536 );
or ( n6739 , n6736 , n6738 );
not ( n6740 , n6739 );
not ( n6741 , n6727 );
or ( n6742 , n6740 , n6741 );
nand ( n6743 , n6723 , n472 );
nand ( n6744 , n6742 , n6743 );
nand ( n6745 , n536 , n472 );
and ( n6746 , n6745 , n471 );
and ( n6747 , n6744 , n6746 );
not ( n6748 , n6747 );
or ( n6749 , n6734 , n6748 );
nand ( n6750 , n6732 , n6722 );
nand ( n6751 , n6749 , n6750 );
xor ( n6752 , n469 , n536 );
not ( n6753 , n6752 );
xor ( n6754 , n469 , n470 );
xor ( n6755 , n470 , n471 );
not ( n6756 , n6755 );
and ( n6757 , n6754 , n6756 );
not ( n6758 , n6757 );
or ( n6759 , n6753 , n6758 );
buf ( n6760 , n6755 );
xor ( n6761 , n469 , n535 );
nand ( n6762 , n6760 , n6761 );
nand ( n6763 , n6759 , n6762 );
not ( n6764 , n6763 );
nand ( n6765 , n536 , n470 );
or ( n6766 , n536 , n470 );
nand ( n6767 , n6766 , n471 );
and ( n6768 , n469 , n6765 , n6767 );
not ( n6769 , n6768 );
not ( n6770 , n471 );
nor ( n6771 , n6770 , n472 );
not ( n6772 , n6771 );
not ( n6773 , n6730 );
or ( n6774 , n6772 , n6773 );
xor ( n6775 , n533 , n471 );
nand ( n6776 , n6775 , n472 );
nand ( n6777 , n6774 , n6776 );
not ( n6778 , n6777 );
or ( n6779 , n6769 , n6778 );
or ( n6780 , n6777 , n6768 );
nand ( n6781 , n6779 , n6780 );
nand ( n6782 , n6764 , n6781 );
not ( n6783 , n6781 );
nand ( n6784 , n6783 , n6763 );
nand ( n6785 , n6782 , n6784 );
xor ( n6786 , n6751 , n6785 );
not ( n6787 , n6786 );
and ( n6788 , n491 , n6787 );
not ( n6789 , n491 );
not ( n6790 , n6787 );
and ( n6791 , n6789 , n6790 );
nor ( n6792 , n6788 , n6791 );
not ( n6793 , n6792 );
or ( n6794 , n6720 , n6793 );
not ( n6795 , n6754 );
nor ( n6796 , n6795 , n6755 );
and ( n6797 , n6761 , n6796 );
and ( n6798 , n469 , n534 );
not ( n6799 , n469 );
not ( n6800 , n534 );
and ( n6801 , n6799 , n6800 );
nor ( n6802 , n6798 , n6801 );
and ( n6803 , n6760 , n6802 );
nor ( n6804 , n6797 , n6803 );
xor ( n6805 , n468 , n469 );
not ( n6806 , n6805 );
not ( n6807 , n6806 );
nand ( n6808 , n6807 , n536 );
not ( n6809 , n6771 );
not ( n6810 , n6775 );
or ( n6811 , n6809 , n6810 );
xor ( n6812 , n532 , n471 );
nand ( n6813 , n6812 , n472 );
nand ( n6814 , n6811 , n6813 );
not ( n6815 , n6814 );
and ( n6816 , n6808 , n6815 );
not ( n6817 , n6808 );
and ( n6818 , n6817 , n6814 );
nor ( n6819 , n6816 , n6818 );
and ( n6820 , n6804 , n6819 );
not ( n6821 , n6804 );
not ( n6822 , n6819 );
and ( n6823 , n6821 , n6822 );
nor ( n6824 , n6820 , n6823 );
not ( n6825 , n6824 );
nand ( n6826 , n6777 , n6768 );
not ( n6827 , n6826 );
nand ( n6828 , n6825 , n6827 );
nand ( n6829 , n6824 , n6826 );
nand ( n6830 , n6828 , n6829 );
not ( n6831 , n6782 );
not ( n6832 , n6751 );
or ( n6833 , n6831 , n6832 );
nand ( n6834 , n6833 , n6784 );
buf ( n6835 , n6834 );
xnor ( n6836 , n6830 , n6835 );
not ( n6837 , n6836 );
and ( n6838 , n491 , n6837 );
not ( n6839 , n491 );
and ( n6840 , n6839 , n6836 );
nor ( n6841 , n6838 , n6840 );
nand ( n6842 , n6714 , n6718 );
not ( n6843 , n6842 );
or ( n6844 , n6841 , n6843 );
nand ( n6845 , n6794 , n6844 );
not ( n6846 , n6745 );
and ( n6847 , n489 , n6846 );
xor ( n6848 , n490 , n491 );
not ( n6849 , n6848 );
and ( n6850 , n6733 , n6750 );
not ( n6851 , n6850 );
and ( n6852 , n6747 , n6851 );
not ( n6853 , n6747 );
and ( n6854 , n6853 , n6850 );
or ( n6855 , n6852 , n6854 );
xor ( n6856 , n489 , n6855 );
not ( n6857 , n6856 );
or ( n6858 , n6849 , n6857 );
nor ( n6859 , n6744 , n6746 );
not ( n6860 , n6859 );
not ( n6861 , n6747 );
nand ( n6862 , n6860 , n6861 );
not ( n6863 , n6862 );
xor ( n6864 , n489 , n6863 );
and ( n6865 , n489 , n490 );
nor ( n6866 , n489 , n490 );
nor ( n6867 , n6865 , n6848 , n6866 );
nand ( n6868 , n6864 , n6867 );
nand ( n6869 , n6858 , n6868 );
xor ( n6870 , n6847 , n6869 );
or ( n6871 , n6846 , n490 );
nand ( n6872 , n6871 , n491 );
nand ( n6873 , n6846 , n490 );
and ( n6874 , n6872 , n6873 , n489 );
not ( n6875 , n6848 );
not ( n6876 , n6864 );
or ( n6877 , n6875 , n6876 );
xor ( n6878 , n489 , n6846 );
nand ( n6879 , n6878 , n6867 );
nand ( n6880 , n6877 , n6879 );
and ( n6881 , n6874 , n6880 );
xor ( n6882 , n6870 , n6881 );
xor ( n6883 , n6845 , n6882 );
xor ( n6884 , n6874 , n6880 );
not ( n6885 , n6842 );
not ( n6886 , n6792 );
or ( n6887 , n6885 , n6886 );
not ( n6888 , n491 );
not ( n6889 , n6855 );
not ( n6890 , n6889 );
or ( n6891 , n6888 , n6890 );
not ( n6892 , n491 );
nand ( n6893 , n6855 , n6892 );
nand ( n6894 , n6891 , n6893 );
nand ( n6895 , n6894 , n6719 );
nand ( n6896 , n6887 , n6895 );
xor ( n6897 , n6884 , n6896 );
not ( n6898 , n6848 );
nor ( n6899 , n6745 , n6898 );
not ( n6900 , n6842 );
not ( n6901 , n6894 );
or ( n6902 , n6900 , n6901 );
and ( n6903 , n491 , n6863 );
not ( n6904 , n491 );
and ( n6905 , n6904 , n6862 );
nor ( n6906 , n6903 , n6905 );
nand ( n6907 , n6906 , n6719 );
nand ( n6908 , n6902 , n6907 );
xor ( n6909 , n6899 , n6908 );
or ( n6910 , n6846 , n492 );
nand ( n6911 , n6910 , n493 );
and ( n6912 , n6846 , n492 );
nor ( n6913 , n6912 , n6892 );
and ( n6914 , n6911 , n6913 );
not ( n6915 , n6719 );
or ( n6916 , n6745 , n491 );
or ( n6917 , n6846 , n6892 );
nand ( n6918 , n6916 , n6917 );
not ( n6919 , n6918 );
or ( n6920 , n6915 , n6919 );
nand ( n6921 , n6906 , n6842 );
nand ( n6922 , n6920 , n6921 );
and ( n6923 , n6914 , n6922 );
and ( n6924 , n6909 , n6923 );
and ( n6925 , n6899 , n6908 );
or ( n6926 , n6924 , n6925 );
and ( n6927 , n6897 , n6926 );
and ( n6928 , n6884 , n6896 );
or ( n6929 , n6927 , n6928 );
and ( n6930 , n6883 , n6929 );
and ( n6931 , n6845 , n6882 );
or ( n6932 , n6930 , n6931 );
not ( n6933 , n496 );
not ( n6934 , n6933 );
not ( n6935 , n497 );
and ( n6936 , n6934 , n6935 );
nor ( n6937 , n1009 , n496 );
nor ( n6938 , n6936 , n6937 );
not ( n6939 , n6938 );
not ( n6940 , n6939 );
xor ( n6941 , n532 , n467 );
not ( n6942 , n6941 );
not ( n6943 , n467 );
not ( n6944 , n468 );
not ( n6945 , n6944 );
or ( n6946 , n6943 , n6945 );
nand ( n6947 , n980 , n468 );
nand ( n6948 , n6946 , n6947 );
not ( n6949 , n6805 );
nand ( n6950 , n6948 , n6949 );
not ( n6951 , n6950 );
buf ( n6952 , n6951 );
not ( n6953 , n6952 );
or ( n6954 , n6942 , n6953 );
xor ( n6955 , n468 , n469 );
xor ( n6956 , n531 , n467 );
nand ( n6957 , n6955 , n6956 );
nand ( n6958 , n6954 , n6957 );
xor ( n6959 , n464 , n465 );
and ( n6960 , n6959 , n536 );
xor ( n6961 , n471 , n529 );
not ( n6962 , n6961 );
not ( n6963 , n6771 );
or ( n6964 , n6962 , n6963 );
and ( n6965 , n528 , n471 );
not ( n6966 , n528 );
not ( n6967 , n471 );
and ( n6968 , n6966 , n6967 );
nor ( n6969 , n6965 , n6968 );
nand ( n6970 , n6969 , n472 );
nand ( n6971 , n6964 , n6970 );
xor ( n6972 , n6960 , n6971 );
xor ( n6973 , n465 , n535 );
not ( n6974 , n6973 );
not ( n6975 , n466 );
nand ( n6976 , n6975 , n465 );
not ( n6977 , n465 );
nand ( n6978 , n6977 , n466 );
nand ( n6979 , n6976 , n6978 );
xor ( n6980 , n466 , n467 );
not ( n6981 , n6980 );
nand ( n6982 , n6979 , n6981 );
not ( n6983 , n6982 );
not ( n6984 , n6983 );
or ( n6985 , n6974 , n6984 );
xor ( n6986 , n466 , n467 );
buf ( n6987 , n6986 );
xor ( n6988 , n534 , n465 );
nand ( n6989 , n6987 , n6988 );
nand ( n6990 , n6985 , n6989 );
and ( n6991 , n6972 , n6990 );
and ( n6992 , n6960 , n6971 );
or ( n6993 , n6991 , n6992 );
xor ( n6994 , n6958 , n6993 );
nand ( n6995 , n536 , n464 );
or ( n6996 , n536 , n464 );
nand ( n6997 , n6996 , n465 );
nand ( n6998 , n6995 , n463 , n6997 );
not ( n6999 , n6998 );
xor ( n7000 , n530 , n469 );
not ( n7001 , n7000 );
nand ( n7002 , n6756 , n6754 );
not ( n7003 , n7002 );
not ( n7004 , n7003 );
or ( n7005 , n7001 , n7004 );
xor ( n7006 , n529 , n469 );
nand ( n7007 , n6760 , n7006 );
nand ( n7008 , n7005 , n7007 );
not ( n7009 , n7008 );
or ( n7010 , n6999 , n7009 );
or ( n7011 , n7008 , n6998 );
nand ( n7012 , n7010 , n7011 );
xor ( n7013 , n6994 , n7012 );
not ( n7014 , n7013 );
xor ( n7015 , n536 , n463 );
not ( n7016 , n7015 );
not ( n7017 , n6959 );
and ( n7018 , n463 , n464 );
not ( n7019 , n463 );
not ( n7020 , n464 );
and ( n7021 , n7019 , n7020 );
nor ( n7022 , n7018 , n7021 );
and ( n7023 , n7017 , n7022 );
not ( n7024 , n7023 );
or ( n7025 , n7016 , n7024 );
xor ( n7026 , n464 , n465 );
xor ( n7027 , n535 , n463 );
nand ( n7028 , n7026 , n7027 );
nand ( n7029 , n7025 , n7028 );
not ( n7030 , n6988 );
not ( n7031 , n6978 );
not ( n7032 , n6976 );
or ( n7033 , n7031 , n7032 );
nand ( n7034 , n7033 , n6981 );
not ( n7035 , n7034 );
not ( n7036 , n7035 );
or ( n7037 , n7030 , n7036 );
xor ( n7038 , n533 , n465 );
nand ( n7039 , n6987 , n7038 );
nand ( n7040 , n7037 , n7039 );
not ( n7041 , n6969 );
not ( n7042 , n6727 );
or ( n7043 , n7041 , n7042 );
xor ( n7044 , n471 , n527 );
nand ( n7045 , n7044 , n472 );
nand ( n7046 , n7043 , n7045 );
nand ( n7047 , n7029 , n7040 , n7046 );
not ( n7048 , n7029 );
not ( n7049 , n7046 );
nand ( n7050 , n7048 , n7040 , n7049 );
not ( n7051 , n7040 );
nand ( n7052 , n7051 , n7048 , n7046 );
nand ( n7053 , n7051 , n7029 , n7049 );
nand ( n7054 , n7047 , n7050 , n7052 , n7053 );
nand ( n7055 , n536 , n466 );
nand ( n7056 , n7055 , n465 );
not ( n7057 , n7056 );
or ( n7058 , n536 , n466 );
nand ( n7059 , n7058 , n467 );
nand ( n7060 , n7057 , n7059 );
not ( n7061 , n7060 );
xor ( n7062 , n471 , n530 );
not ( n7063 , n7062 );
not ( n7064 , n6727 );
or ( n7065 , n7063 , n7064 );
nand ( n7066 , n6961 , n472 );
nand ( n7067 , n7065 , n7066 );
nand ( n7068 , n7061 , n7067 );
not ( n7069 , n7000 );
not ( n7070 , n6760 );
or ( n7071 , n7069 , n7070 );
and ( n7072 , n531 , n469 );
not ( n7073 , n531 );
not ( n7074 , n469 );
and ( n7075 , n7073 , n7074 );
nor ( n7076 , n7072 , n7075 );
nand ( n7077 , n6756 , n6754 , n7076 );
nand ( n7078 , n7071 , n7077 );
not ( n7079 , n7078 );
nand ( n7080 , n7068 , n7079 );
not ( n7081 , n7080 );
xor ( n7082 , n533 , n467 );
not ( n7083 , n7082 );
not ( n7084 , n6952 );
not ( n7085 , n7084 );
not ( n7086 , n7085 );
or ( n7087 , n7083 , n7086 );
buf ( n7088 , n6807 );
nand ( n7089 , n7088 , n6941 );
nand ( n7090 , n7087 , n7089 );
not ( n7091 , n7090 );
or ( n7092 , n7081 , n7091 );
or ( n7093 , n7068 , n7079 );
nand ( n7094 , n7092 , n7093 );
xor ( n7095 , n7054 , n7094 );
not ( n7096 , n7095 );
or ( n7097 , n7014 , n7096 );
or ( n7098 , n7095 , n7013 );
nand ( n7099 , n7097 , n7098 );
xor ( n7100 , n6960 , n6971 );
xor ( n7101 , n7100 , n6990 );
xor ( n7102 , n536 , n465 );
not ( n7103 , n7102 );
not ( n7104 , n6983 );
or ( n7105 , n7103 , n7104 );
nand ( n7106 , n6987 , n6973 );
nand ( n7107 , n7105 , n7106 );
xor ( n7108 , n469 , n532 );
not ( n7109 , n7108 );
not ( n7110 , n7003 );
or ( n7111 , n7109 , n7110 );
nand ( n7112 , n6760 , n7076 );
nand ( n7113 , n7111 , n7112 );
xor ( n7114 , n7107 , n7113 );
xor ( n7115 , n534 , n467 );
not ( n7116 , n7115 );
not ( n7117 , n7085 );
or ( n7118 , n7116 , n7117 );
nand ( n7119 , n7088 , n7082 );
nand ( n7120 , n7118 , n7119 );
and ( n7121 , n7114 , n7120 );
and ( n7122 , n7107 , n7113 );
or ( n7123 , n7121 , n7122 );
xor ( n7124 , n7101 , n7123 );
not ( n7125 , n7078 );
not ( n7126 , n7068 );
or ( n7127 , n7125 , n7126 );
or ( n7128 , n7068 , n7078 );
nand ( n7129 , n7127 , n7128 );
xor ( n7130 , n7090 , n7129 );
and ( n7131 , n7124 , n7130 );
and ( n7132 , n7101 , n7123 );
or ( n7133 , n7131 , n7132 );
not ( n7134 , n7133 );
nor ( n7135 , n7099 , n7134 );
not ( n7136 , n7135 );
nand ( n7137 , n7099 , n7134 );
nand ( n7138 , n7136 , n7137 );
not ( n7139 , n7060 );
not ( n7140 , n7139 );
not ( n7141 , n7067 );
or ( n7142 , n7140 , n7141 );
or ( n7143 , n7067 , n7139 );
nand ( n7144 , n7142 , n7143 );
xor ( n7145 , n533 , n469 );
not ( n7146 , n7145 );
not ( n7147 , n6757 );
or ( n7148 , n7146 , n7147 );
nand ( n7149 , n6721 , n7108 );
nand ( n7150 , n7148 , n7149 );
not ( n7151 , n7150 );
xor ( n7152 , n471 , n531 );
not ( n7153 , n7152 );
not ( n7154 , n6727 );
or ( n7155 , n7153 , n7154 );
nand ( n7156 , n7062 , n472 );
nand ( n7157 , n7155 , n7156 );
not ( n7158 , n7157 );
not ( n7159 , n6735 );
nand ( n7160 , n7159 , n6987 );
nand ( n7161 , n7158 , n7160 );
not ( n7162 , n7161 );
or ( n7163 , n7151 , n7162 );
not ( n7164 , n7160 );
nand ( n7165 , n7164 , n7157 );
nand ( n7166 , n7163 , n7165 );
xnor ( n7167 , n7144 , n7166 );
not ( n7168 , n7167 );
xor ( n7169 , n7107 , n7113 );
xor ( n7170 , n7169 , n7120 );
not ( n7171 , n7170 );
or ( n7172 , n7168 , n7171 );
or ( n7173 , n7170 , n7167 );
nand ( n7174 , n7172 , n7173 );
or ( n7175 , n536 , n468 );
nand ( n7176 , n7175 , n469 );
nand ( n7177 , n536 , n468 );
nand ( n7178 , n7176 , n7177 , n467 );
not ( n7179 , n7178 );
not ( n7180 , n6812 );
not ( n7181 , n6727 );
or ( n7182 , n7180 , n7181 );
nand ( n7183 , n7152 , n472 );
nand ( n7184 , n7182 , n7183 );
nand ( n7185 , n7179 , n7184 );
xor ( n7186 , n535 , n467 );
not ( n7187 , n7186 );
not ( n7188 , n6952 );
or ( n7189 , n7187 , n7188 );
nand ( n7190 , n7088 , n7115 );
nand ( n7191 , n7189 , n7190 );
not ( n7192 , n7191 );
nand ( n7193 , n7185 , n7192 );
not ( n7194 , n7193 );
not ( n7195 , n7157 );
not ( n7196 , n7160 );
and ( n7197 , n7195 , n7196 );
and ( n7198 , n7157 , n7160 );
nor ( n7199 , n7197 , n7198 );
xnor ( n7200 , n7199 , n7150 );
not ( n7201 , n7200 );
or ( n7202 , n7194 , n7201 );
not ( n7203 , n7185 );
nand ( n7204 , n7203 , n7191 );
nand ( n7205 , n7202 , n7204 );
not ( n7206 , n7205 );
nor ( n7207 , n7174 , n7206 );
not ( n7208 , n7207 );
not ( n7209 , n6829 );
not ( n7210 , n6834 );
or ( n7211 , n7209 , n7210 );
nand ( n7212 , n7211 , n6828 );
not ( n7213 , n6814 );
not ( n7214 , n6808 );
not ( n7215 , n7214 );
or ( n7216 , n7213 , n7215 );
nor ( n7217 , n6814 , n7214 );
or ( n7218 , n6804 , n7217 );
nand ( n7219 , n7216 , n7218 );
not ( n7220 , n7219 );
not ( n7221 , n6802 );
not ( n7222 , n6757 );
or ( n7223 , n7221 , n7222 );
nand ( n7224 , n6721 , n7145 );
nand ( n7225 , n7223 , n7224 );
not ( n7226 , n7225 );
and ( n7227 , n6955 , n7186 );
not ( n7228 , n6955 );
xor ( n7229 , n536 , n467 );
and ( n7230 , n7229 , n6948 );
and ( n7231 , n7228 , n7230 );
or ( n7232 , n7227 , n7231 );
xor ( n7233 , n7226 , n7232 );
not ( n7234 , n7184 );
not ( n7235 , n7178 );
and ( n7236 , n7234 , n7235 );
and ( n7237 , n7184 , n7178 );
nor ( n7238 , n7236 , n7237 );
xnor ( n7239 , n7233 , n7238 );
nand ( n7240 , n7220 , n7239 );
nand ( n7241 , n7212 , n7240 );
not ( n7242 , n7241 );
not ( n7243 , n7239 );
nand ( n7244 , n7243 , n7219 );
not ( n7245 , n7244 );
or ( n7246 , n7242 , n7245 );
not ( n7247 , n7226 );
not ( n7248 , n7238 );
or ( n7249 , n7247 , n7248 );
nand ( n7250 , n7249 , n7232 );
not ( n7251 , n7238 );
nand ( n7252 , n7251 , n7225 );
nand ( n7253 , n7250 , n7252 );
not ( n7254 , n7253 );
not ( n7255 , n7203 );
not ( n7256 , n7192 );
and ( n7257 , n7255 , n7256 );
and ( n7258 , n7203 , n7192 );
nor ( n7259 , n7257 , n7258 );
not ( n7260 , n7259 );
not ( n7261 , n7200 );
and ( n7262 , n7260 , n7261 );
and ( n7263 , n7200 , n7259 );
nor ( n7264 , n7262 , n7263 );
nand ( n7265 , n7254 , n7264 );
nand ( n7266 , n7246 , n7265 );
not ( n7267 , n7253 );
nor ( n7268 , n7267 , n7264 );
not ( n7269 , n7268 );
nand ( n7270 , n7208 , n7266 , n7269 );
not ( n7271 , n7270 );
xor ( n7272 , n7101 , n7123 );
xor ( n7273 , n7272 , n7130 );
not ( n7274 , n7273 );
not ( n7275 , n7166 );
nand ( n7276 , n7275 , n7144 );
not ( n7277 , n7276 );
not ( n7278 , n7170 );
or ( n7279 , n7277 , n7278 );
not ( n7280 , n7144 );
nand ( n7281 , n7280 , n7166 );
nand ( n7282 , n7279 , n7281 );
not ( n7283 , n7282 );
and ( n7284 , n7274 , n7283 );
not ( n7285 , n7170 );
not ( n7286 , n7167 );
and ( n7287 , n7285 , n7286 );
not ( n7288 , n7285 );
and ( n7289 , n7288 , n7167 );
nor ( n7290 , n7287 , n7289 );
nor ( n7291 , n7290 , n7205 );
nor ( n7292 , n7284 , n7291 );
not ( n7293 , n7292 );
or ( n7294 , n7271 , n7293 );
nand ( n7295 , n7273 , n7282 );
nand ( n7296 , n7294 , n7295 );
xnor ( n7297 , n7138 , n7296 );
not ( n7298 , n7297 );
and ( n7299 , n495 , n7298 );
not ( n7300 , n495 );
buf ( n7301 , n7297 );
and ( n7302 , n7300 , n7301 );
or ( n7303 , n7299 , n7302 );
not ( n7304 , n7303 );
or ( n7305 , n6940 , n7304 );
or ( n7306 , n7273 , n7282 );
nand ( n7307 , n7306 , n7295 );
not ( n7308 , n7206 );
not ( n7309 , n7290 );
not ( n7310 , n7309 );
or ( n7311 , n7308 , n7310 );
nand ( n7312 , n7311 , n7270 );
not ( n7313 , n7312 );
not ( n7314 , n7313 );
and ( n7315 , n7307 , n7314 );
not ( n7316 , n7307 );
buf ( n7317 , n7313 );
and ( n7318 , n7316 , n7317 );
nor ( n7319 , n7315 , n7318 );
not ( n7320 , n7319 );
not ( n7321 , n7320 );
xor ( n7322 , n495 , n7321 );
and ( n7323 , n495 , n496 );
nor ( n7324 , n495 , n496 );
nor ( n7325 , n7323 , n7324 );
and ( n7326 , n7325 , n6938 );
nand ( n7327 , n7322 , n7326 );
nand ( n7328 , n7305 , n7327 );
xor ( n7329 , n6932 , n7328 );
not ( n7330 , n6842 );
not ( n7331 , n491 );
nand ( n7332 , n7244 , n7240 );
not ( n7333 , n7332 );
not ( n7334 , n7333 );
not ( n7335 , n7212 );
not ( n7336 , n7335 );
or ( n7337 , n7334 , n7336 );
nand ( n7338 , n7332 , n7212 );
nand ( n7339 , n7337 , n7338 );
not ( n7340 , n7339 );
not ( n7341 , n7340 );
or ( n7342 , n7331 , n7341 );
nand ( n7343 , n7339 , n6892 );
nand ( n7344 , n7342 , n7343 );
not ( n7345 , n7344 );
or ( n7346 , n7330 , n7345 );
not ( n7347 , n6841 );
nand ( n7348 , n7347 , n6719 );
nand ( n7349 , n7346 , n7348 );
and ( n7350 , n489 , n6863 );
not ( n7351 , n6848 );
xor ( n7352 , n489 , n6787 );
not ( n7353 , n7352 );
or ( n7354 , n7351 , n7353 );
not ( n7355 , n6867 );
not ( n7356 , n7355 );
nand ( n7357 , n7356 , n6856 );
nand ( n7358 , n7354 , n7357 );
xor ( n7359 , n7350 , n7358 );
xor ( n7360 , n6847 , n6869 );
and ( n7361 , n7360 , n6881 );
and ( n7362 , n6847 , n6869 );
or ( n7363 , n7361 , n7362 );
xor ( n7364 , n7359 , n7363 );
xor ( n7365 , n7349 , n7364 );
and ( n7366 , n494 , n1554 );
not ( n7367 , n494 );
and ( n7368 , n7367 , n495 );
or ( n7369 , n7366 , n7368 );
not ( n7370 , n7369 );
not ( n7371 , n7370 );
not ( n7372 , n7371 );
not ( n7373 , n7207 );
not ( n7374 , n7373 );
nand ( n7375 , n7309 , n7206 );
not ( n7376 , n7375 );
or ( n7377 , n7374 , n7376 );
nand ( n7378 , n7266 , n7269 );
nand ( n7379 , n7377 , n7378 );
not ( n7380 , n7378 );
nand ( n7381 , n7380 , n7375 , n7373 );
nand ( n7382 , n7379 , n7381 );
buf ( n7383 , n7382 );
not ( n7384 , n7383 );
and ( n7385 , n493 , n7384 );
not ( n7386 , n493 );
and ( n7387 , n7386 , n7383 );
or ( n7388 , n7385 , n7387 );
not ( n7389 , n7388 );
or ( n7390 , n7372 , n7389 );
not ( n7391 , n7265 );
nor ( n7392 , n7391 , n7268 );
nand ( n7393 , n7241 , n7244 );
xor ( n7394 , n7392 , n7393 );
buf ( n7395 , n7394 );
not ( n7396 , n7395 );
and ( n7397 , n493 , n7396 );
not ( n7398 , n493 );
and ( n7399 , n7398 , n7395 );
or ( n7400 , n7397 , n7399 );
or ( n7401 , n493 , n494 );
nand ( n7402 , n493 , n494 );
nand ( n7403 , n7401 , n7402 );
nor ( n7404 , n7369 , n7403 );
buf ( n7405 , n7404 );
nand ( n7406 , n7400 , n7405 );
nand ( n7407 , n7390 , n7406 );
xor ( n7408 , n7365 , n7407 );
xor ( n7409 , n7329 , n7408 );
xor ( n7410 , n498 , n499 );
not ( n7411 , n7410 );
not ( n7412 , n7411 );
xnor ( n7413 , n497 , n498 );
nor ( n7414 , n7412 , n7413 );
buf ( n7415 , n7414 );
not ( n7416 , n7415 );
not ( n7417 , n1009 );
not ( n7418 , n7301 );
or ( n7419 , n7417 , n7418 );
or ( n7420 , n7301 , n1009 );
nand ( n7421 , n7419 , n7420 );
not ( n7422 , n7421 );
or ( n7423 , n7416 , n7422 );
and ( n7424 , n7273 , n7282 , n7137 );
nor ( n7425 , n7134 , n7099 );
nor ( n7426 , n7424 , n7425 );
nand ( n7427 , n7313 , n7137 , n7306 );
nand ( n7428 , n7426 , n7427 );
nand ( n7429 , n7027 , n7022 );
buf ( n7430 , n6959 );
or ( n7431 , n7429 , n7430 );
xor ( n7432 , n534 , n463 );
nand ( n7433 , n7430 , n7432 );
nand ( n7434 , n7431 , n7433 );
not ( n7435 , n7434 );
not ( n7436 , n7044 );
not ( n7437 , n6727 );
or ( n7438 , n7436 , n7437 );
xor ( n7439 , n471 , n526 );
nand ( n7440 , n7439 , n472 );
nand ( n7441 , n7438 , n7440 );
and ( n7442 , n7435 , n7441 );
not ( n7443 , n7435 );
not ( n7444 , n7441 );
and ( n7445 , n7443 , n7444 );
nor ( n7446 , n7442 , n7445 );
not ( n7447 , n6956 );
not ( n7448 , n6950 );
buf ( n7449 , n7448 );
not ( n7450 , n7449 );
or ( n7451 , n7447 , n7450 );
xor ( n7452 , n530 , n467 );
nand ( n7453 , n6955 , n7452 );
nand ( n7454 , n7451 , n7453 );
xor ( n7455 , n7446 , n7454 );
not ( n7456 , n7455 );
xor ( n7457 , n6958 , n6993 );
and ( n7458 , n7457 , n7012 );
and ( n7459 , n6958 , n6993 );
or ( n7460 , n7458 , n7459 );
not ( n7461 , n7460 );
or ( n7462 , n7456 , n7461 );
or ( n7463 , n7460 , n7455 );
nand ( n7464 , n7462 , n7463 );
not ( n7465 , n6998 );
nand ( n7466 , n7465 , n7008 );
not ( n7467 , n7049 );
not ( n7468 , n7051 );
or ( n7469 , n7467 , n7468 );
nand ( n7470 , n7469 , n7029 );
nand ( n7471 , n7040 , n7046 );
nand ( n7472 , n7470 , n7471 );
xor ( n7473 , n7466 , n7472 );
xor ( n7474 , n462 , n463 );
buf ( n7475 , n7474 );
and ( n7476 , n7475 , n536 );
not ( n7477 , n7038 );
not ( n7478 , n6983 );
or ( n7479 , n7477 , n7478 );
xor ( n7480 , n532 , n465 );
nand ( n7481 , n6987 , n7480 );
nand ( n7482 , n7479 , n7481 );
not ( n7483 , n7482 );
xor ( n7484 , n7476 , n7483 );
not ( n7485 , n7006 );
not ( n7486 , n6757 );
or ( n7487 , n7485 , n7486 );
xor ( n7488 , n528 , n469 );
nand ( n7489 , n6721 , n7488 );
nand ( n7490 , n7487 , n7489 );
not ( n7491 , n7490 );
xnor ( n7492 , n7484 , n7491 );
xnor ( n7493 , n7473 , n7492 );
and ( n7494 , n7464 , n7493 );
not ( n7495 , n7464 );
not ( n7496 , n7493 );
and ( n7497 , n7495 , n7496 );
nor ( n7498 , n7494 , n7497 );
not ( n7499 , n7498 );
not ( n7500 , n7013 );
or ( n7501 , n7054 , n7094 );
not ( n7502 , n7501 );
or ( n7503 , n7500 , n7502 );
nand ( n7504 , n7054 , n7094 );
nand ( n7505 , n7503 , n7504 );
nand ( n7506 , n7499 , n7505 );
not ( n7507 , n7505 );
nand ( n7508 , n7498 , n7507 );
nand ( n7509 , n7506 , n7508 );
xnor ( n7510 , n7428 , n7509 );
buf ( n7511 , n7510 );
not ( n7512 , n7511 );
and ( n7513 , n497 , n7512 );
not ( n7514 , n497 );
and ( n7515 , n7514 , n7511 );
or ( n7516 , n7513 , n7515 );
not ( n7517 , n7411 );
nand ( n7518 , n7516 , n7517 );
nand ( n7519 , n7423 , n7518 );
not ( n7520 , n7369 );
and ( n7521 , n493 , n7339 );
not ( n7522 , n493 );
and ( n7523 , n7522 , n7340 );
nor ( n7524 , n7521 , n7523 );
not ( n7525 , n7524 );
or ( n7526 , n7520 , n7525 );
and ( n7527 , n493 , n6836 );
not ( n7528 , n493 );
and ( n7529 , n7528 , n6837 );
nor ( n7530 , n7527 , n7529 );
nand ( n7531 , n7530 , n7405 );
nand ( n7532 , n7526 , n7531 );
xor ( n7533 , n6884 , n6896 );
xor ( n7534 , n7533 , n6926 );
xor ( n7535 , n7532 , n7534 );
not ( n7536 , n6939 );
and ( n7537 , n495 , n7384 );
not ( n7538 , n495 );
and ( n7539 , n7538 , n7383 );
or ( n7540 , n7537 , n7539 );
not ( n7541 , n7540 );
or ( n7542 , n7536 , n7541 );
and ( n7543 , n495 , n7396 );
not ( n7544 , n495 );
and ( n7545 , n7544 , n7395 );
or ( n7546 , n7543 , n7545 );
nand ( n7547 , n7546 , n7326 );
nand ( n7548 , n7542 , n7547 );
and ( n7549 , n7535 , n7548 );
and ( n7550 , n7532 , n7534 );
or ( n7551 , n7549 , n7550 );
xor ( n7552 , n7519 , n7551 );
not ( n7553 , n1122 );
and ( n7554 , n499 , n500 );
nor ( n7555 , n499 , n500 );
nor ( n7556 , n7554 , n7555 );
nand ( n7557 , n7553 , n7556 );
not ( n7558 , n7557 );
not ( n7559 , n7558 );
buf ( n7560 , n7507 );
not ( n7561 , n7499 );
and ( n7562 , n7560 , n7561 );
not ( n7563 , n7137 );
nor ( n7564 , n7562 , n7563 );
nand ( n7565 , n7564 , n7296 );
not ( n7566 , n7508 );
not ( n7567 , n7135 );
or ( n7568 , n7566 , n7567 );
nand ( n7569 , n7568 , n7506 );
not ( n7570 , n7569 );
nand ( n7571 , n7565 , n7570 );
not ( n7572 , n7455 );
buf ( n7573 , n7460 );
not ( n7574 , n7573 );
not ( n7575 , n7574 );
or ( n7576 , n7572 , n7575 );
nand ( n7577 , n7576 , n7496 );
not ( n7578 , n7455 );
nand ( n7579 , n7578 , n7573 );
nand ( n7580 , n7577 , n7579 );
xor ( n7581 , n536 , n461 );
not ( n7582 , n7581 );
xnor ( n7583 , n461 , n462 );
nor ( n7584 , n7583 , n7474 );
buf ( n7585 , n7584 );
not ( n7586 , n7585 );
or ( n7587 , n7582 , n7586 );
xor ( n7588 , n535 , n461 );
nand ( n7589 , n7588 , n7475 );
nand ( n7590 , n7587 , n7589 );
not ( n7591 , n7590 );
not ( n7592 , n7452 );
not ( n7593 , n7449 );
or ( n7594 , n7592 , n7593 );
xor ( n7595 , n529 , n467 );
nand ( n7596 , n6955 , n7595 );
nand ( n7597 , n7594 , n7596 );
xor ( n7598 , n7591 , n7597 );
not ( n7599 , n7488 );
not ( n7600 , n7003 );
or ( n7601 , n7599 , n7600 );
xor ( n7602 , n527 , n469 );
nand ( n7603 , n6721 , n7602 );
nand ( n7604 , n7601 , n7603 );
or ( n7605 , n536 , n462 );
nand ( n7606 , n7605 , n463 );
nand ( n7607 , n536 , n462 );
nand ( n7608 , n7606 , n7607 , n461 );
not ( n7609 , n7608 );
and ( n7610 , n7604 , n7609 );
not ( n7611 , n7604 );
and ( n7612 , n7611 , n7608 );
nor ( n7613 , n7610 , n7612 );
xnor ( n7614 , n7598 , n7613 );
or ( n7615 , n7466 , n7492 );
not ( n7616 , n7466 );
not ( n7617 , n7492 );
or ( n7618 , n7616 , n7617 );
nand ( n7619 , n7471 , n7470 );
nand ( n7620 , n7618 , n7619 );
nand ( n7621 , n7615 , n7620 );
xor ( n7622 , n7614 , n7621 );
not ( n7623 , n7435 );
not ( n7624 , n7444 );
or ( n7625 , n7623 , n7624 );
nand ( n7626 , n7625 , n7454 );
nand ( n7627 , n7441 , n7434 );
nand ( n7628 , n7626 , n7627 );
not ( n7629 , n7628 );
not ( n7630 , n7629 );
not ( n7631 , n7476 );
not ( n7632 , n7490 );
or ( n7633 , n7631 , n7632 );
or ( n7634 , n7490 , n7476 );
nand ( n7635 , n7634 , n7482 );
nand ( n7636 , n7633 , n7635 );
not ( n7637 , n7636 );
and ( n7638 , n7630 , n7637 );
and ( n7639 , n7629 , n7636 );
nor ( n7640 , n7638 , n7639 );
nand ( n7641 , n7432 , n7022 );
not ( n7642 , n7017 );
or ( n7643 , n7641 , n7642 );
xor ( n7644 , n533 , n463 );
nand ( n7645 , n7644 , n7026 );
nand ( n7646 , n7643 , n7645 );
not ( n7647 , n7480 );
not ( n7648 , n7035 );
or ( n7649 , n7647 , n7648 );
xor ( n7650 , n531 , n465 );
nand ( n7651 , n6987 , n7650 );
nand ( n7652 , n7649 , n7651 );
xor ( n7653 , n7646 , n7652 );
not ( n7654 , n7439 );
not ( n7655 , n6727 );
or ( n7656 , n7654 , n7655 );
xor ( n7657 , n525 , n471 );
nand ( n7658 , n7657 , n472 );
nand ( n7659 , n7656 , n7658 );
xnor ( n7660 , n7653 , n7659 );
not ( n7661 , n7660 );
not ( n7662 , n7661 );
and ( n7663 , n7640 , n7662 );
not ( n7664 , n7640 );
and ( n7665 , n7664 , n7661 );
nor ( n7666 , n7663 , n7665 );
xor ( n7667 , n7622 , n7666 );
nand ( n7668 , n7580 , n7667 );
not ( n7669 , n7668 );
not ( n7670 , n7669 );
not ( n7671 , n7580 );
not ( n7672 , n7667 );
nand ( n7673 , n7671 , n7672 );
nand ( n7674 , n7670 , n7673 );
not ( n7675 , n7674 );
xor ( n7676 , n7571 , n7675 );
buf ( n7677 , n7676 );
not ( n7678 , n7677 );
and ( n7679 , n499 , n7678 );
not ( n7680 , n499 );
and ( n7681 , n7680 , n7677 );
or ( n7682 , n7679 , n7681 );
not ( n7683 , n7682 );
or ( n7684 , n7559 , n7683 );
not ( n7685 , n7565 );
not ( n7686 , n7570 );
or ( n7687 , n7685 , n7686 );
nand ( n7688 , n7687 , n7673 );
not ( n7689 , n7669 );
nand ( n7690 , n7688 , n7689 );
xor ( n7691 , n7614 , n7621 );
and ( n7692 , n7691 , n7666 );
and ( n7693 , n7614 , n7621 );
or ( n7694 , n7692 , n7693 );
not ( n7695 , n7694 );
and ( n7696 , n7604 , n7609 );
not ( n7697 , n7696 );
not ( n7698 , n7697 );
not ( n7699 , n7595 );
not ( n7700 , n7449 );
or ( n7701 , n7699 , n7700 );
xor ( n7702 , n528 , n467 );
nand ( n7703 , n7088 , n7702 );
nand ( n7704 , n7701 , n7703 );
not ( n7705 , n7704 );
or ( n7706 , n7698 , n7705 );
not ( n7707 , n7704 );
nand ( n7708 , n7707 , n7696 );
nand ( n7709 , n7706 , n7708 );
buf ( n7710 , n7646 );
not ( n7711 , n7710 );
not ( n7712 , n7659 );
or ( n7713 , n7711 , n7712 );
or ( n7714 , n7710 , n7659 );
nand ( n7715 , n7714 , n7652 );
nand ( n7716 , n7713 , n7715 );
not ( n7717 , n7716 );
and ( n7718 , n7709 , n7717 );
not ( n7719 , n7709 );
and ( n7720 , n7719 , n7716 );
or ( n7721 , n7718 , n7720 );
not ( n7722 , n7628 );
not ( n7723 , n7661 );
or ( n7724 , n7722 , n7723 );
not ( n7725 , n7629 );
not ( n7726 , n7660 );
or ( n7727 , n7725 , n7726 );
nand ( n7728 , n7727 , n7636 );
nand ( n7729 , n7724 , n7728 );
and ( n7730 , n7721 , n7729 );
not ( n7731 , n7721 );
not ( n7732 , n7729 );
and ( n7733 , n7731 , n7732 );
nor ( n7734 , n7730 , n7733 );
not ( n7735 , n461 );
and ( n7736 , n460 , n7735 );
not ( n7737 , n460 );
and ( n7738 , n7737 , n461 );
or ( n7739 , n7736 , n7738 );
and ( n7740 , n7739 , n536 );
not ( n7741 , n7602 );
not ( n7742 , n470 );
and ( n7743 , n471 , n7742 );
not ( n7744 , n471 );
and ( n7745 , n7744 , n470 );
nor ( n7746 , n7743 , n7745 );
and ( n7747 , n7746 , n6754 );
not ( n7748 , n7747 );
or ( n7749 , n7741 , n7748 );
xor ( n7750 , n526 , n469 );
nand ( n7751 , n6755 , n7750 );
nand ( n7752 , n7749 , n7751 );
xor ( n7753 , n7740 , n7752 );
not ( n7754 , n7650 );
not ( n7755 , n7035 );
or ( n7756 , n7754 , n7755 );
and ( n7757 , n530 , n465 );
not ( n7758 , n530 );
not ( n7759 , n465 );
and ( n7760 , n7758 , n7759 );
nor ( n7761 , n7757 , n7760 );
nand ( n7762 , n6987 , n7761 );
nand ( n7763 , n7756 , n7762 );
not ( n7764 , n7763 );
xnor ( n7765 , n7753 , n7764 );
not ( n7766 , n7657 );
not ( n7767 , n6727 );
or ( n7768 , n7766 , n7767 );
xor ( n7769 , n524 , n471 );
nand ( n7770 , n7769 , n472 );
nand ( n7771 , n7768 , n7770 );
not ( n7772 , n7644 );
not ( n7773 , n7023 );
or ( n7774 , n7772 , n7773 );
xor ( n7775 , n532 , n463 );
nand ( n7776 , n7430 , n7775 );
nand ( n7777 , n7774 , n7776 );
xor ( n7778 , n7771 , n7777 );
not ( n7779 , n7588 );
not ( n7780 , n7585 );
or ( n7781 , n7779 , n7780 );
xor ( n7782 , n461 , n534 );
nand ( n7783 , n7475 , n7782 );
nand ( n7784 , n7781 , n7783 );
xor ( n7785 , n7778 , n7784 );
xor ( n7786 , n7765 , n7785 );
not ( n7787 , n7613 );
not ( n7788 , n7597 );
nand ( n7789 , n7788 , n7591 );
not ( n7790 , n7789 );
or ( n7791 , n7787 , n7790 );
nand ( n7792 , n7597 , n7590 );
nand ( n7793 , n7791 , n7792 );
xor ( n7794 , n7786 , n7793 );
and ( n7795 , n7734 , n7794 );
not ( n7796 , n7734 );
not ( n7797 , n7794 );
and ( n7798 , n7796 , n7797 );
nor ( n7799 , n7795 , n7798 );
not ( n7800 , n7799 );
or ( n7801 , n7695 , n7800 );
not ( n7802 , n7799 );
not ( n7803 , n7694 );
nand ( n7804 , n7802 , n7803 );
nand ( n7805 , n7801 , n7804 );
and ( n7806 , n7690 , n7805 );
not ( n7807 , n7690 );
not ( n7808 , n7805 );
and ( n7809 , n7807 , n7808 );
nor ( n7810 , n7806 , n7809 );
not ( n7811 , n7810 );
buf ( n7812 , n7811 );
buf ( n7813 , n1122 );
not ( n7814 , n7813 );
nor ( n7815 , n7814 , n499 );
and ( n7816 , n7812 , n7815 );
not ( n7817 , n7812 );
nand ( n7818 , n7813 , n499 );
not ( n7819 , n7818 );
and ( n7820 , n7817 , n7819 );
nor ( n7821 , n7816 , n7820 );
nand ( n7822 , n7684 , n7821 );
and ( n7823 , n7552 , n7822 );
and ( n7824 , n7519 , n7551 );
or ( n7825 , n7823 , n7824 );
xor ( n7826 , n7409 , n7825 );
xor ( n7827 , n503 , n502 );
buf ( n7828 , n7827 );
not ( n7829 , n7828 );
not ( n7830 , n501 );
nand ( n7831 , n7761 , n6979 );
or ( n7832 , n7831 , n6986 );
and ( n7833 , n529 , n465 );
not ( n7834 , n529 );
and ( n7835 , n7834 , n7759 );
nor ( n7836 , n7833 , n7835 );
nand ( n7837 , n6986 , n7836 );
nand ( n7838 , n7832 , n7837 );
not ( n7839 , n7750 );
not ( n7840 , n7747 );
or ( n7841 , n7839 , n7840 );
xor ( n7842 , n525 , n469 );
nand ( n7843 , n6721 , n7842 );
nand ( n7844 , n7841 , n7843 );
or ( n7845 , n7838 , n7844 );
not ( n7846 , n7775 );
not ( n7847 , n7023 );
or ( n7848 , n7846 , n7847 );
xor ( n7849 , n531 , n463 );
nand ( n7850 , n7430 , n7849 );
nand ( n7851 , n7848 , n7850 );
nand ( n7852 , n7845 , n7851 );
nand ( n7853 , n7838 , n7844 );
nand ( n7854 , n7852 , n7853 );
not ( n7855 , n7854 );
not ( n7856 , n7855 );
not ( n7857 , n7782 );
not ( n7858 , n7584 );
or ( n7859 , n7857 , n7858 );
xor ( n7860 , n461 , n533 );
nand ( n7861 , n7475 , n7860 );
nand ( n7862 , n7859 , n7861 );
not ( n7863 , n7862 );
not ( n7864 , n7863 );
not ( n7865 , n7702 );
not ( n7866 , n6951 );
or ( n7867 , n7865 , n7866 );
xor ( n7868 , n527 , n467 );
nand ( n7869 , n6807 , n7868 );
nand ( n7870 , n7867 , n7869 );
not ( n7871 , n7870 );
not ( n7872 , n7871 );
or ( n7873 , n7864 , n7872 );
xor ( n7874 , n536 , n459 );
not ( n7875 , n7874 );
not ( n7876 , n460 );
nand ( n7877 , n7735 , n7876 , n459 );
not ( n7878 , n459 );
nand ( n7879 , n7878 , n460 , n461 );
nand ( n7880 , n7877 , n7879 );
buf ( n7881 , n7880 );
not ( n7882 , n7881 );
or ( n7883 , n7875 , n7882 );
nand ( n7884 , n7735 , n460 );
not ( n7885 , n460 );
nand ( n7886 , n7885 , n461 );
nand ( n7887 , n7884 , n7886 );
buf ( n7888 , n7887 );
xor ( n7889 , n535 , n459 );
nand ( n7890 , n7888 , n7889 );
nand ( n7891 , n7883 , n7890 );
nand ( n7892 , n7873 , n7891 );
nand ( n7893 , n7870 , n7862 );
nand ( n7894 , n7892 , n7893 );
not ( n7895 , n7894 );
and ( n7896 , n7856 , n7895 );
and ( n7897 , n7855 , n7894 );
nor ( n7898 , n7896 , n7897 );
not ( n7899 , n472 );
xor ( n7900 , n471 , n522 );
not ( n7901 , n7900 );
or ( n7902 , n7899 , n7901 );
not ( n7903 , n471 );
nor ( n7904 , n7903 , n472 );
xor ( n7905 , n471 , n523 );
nand ( n7906 , n7904 , n7905 );
nand ( n7907 , n7902 , n7906 );
xor ( n7908 , n458 , n459 );
and ( n7909 , n7908 , n536 );
xor ( n7910 , n7907 , n7909 );
not ( n7911 , n7842 );
not ( n7912 , n7003 );
or ( n7913 , n7911 , n7912 );
xor ( n7914 , n524 , n469 );
nand ( n7915 , n6721 , n7914 );
nand ( n7916 , n7913 , n7915 );
xor ( n7917 , n7910 , n7916 );
buf ( n7918 , n7917 );
not ( n7919 , n7918 );
and ( n7920 , n7898 , n7919 );
not ( n7921 , n7898 );
and ( n7922 , n7921 , n7918 );
nor ( n7923 , n7920 , n7922 );
not ( n7924 , n7923 );
not ( n7925 , n7924 );
xor ( n7926 , n532 , n461 );
not ( n7927 , n7926 );
not ( n7928 , n7475 );
or ( n7929 , n7927 , n7928 );
nand ( n7930 , n7860 , n7584 );
nand ( n7931 , n7929 , n7930 );
not ( n7932 , n7889 );
not ( n7933 , n7880 );
or ( n7934 , n7932 , n7933 );
and ( n7935 , n459 , n534 );
not ( n7936 , n459 );
and ( n7937 , n7936 , n6800 );
nor ( n7938 , n7935 , n7937 );
nand ( n7939 , n7887 , n7938 );
nand ( n7940 , n7934 , n7939 );
not ( n7941 , n7940 );
xor ( n7942 , n7931 , n7941 );
not ( n7943 , n6727 );
not ( n7944 , n7769 );
or ( n7945 , n7943 , n7944 );
nand ( n7946 , n7905 , n472 );
nand ( n7947 , n7945 , n7946 );
or ( n7948 , n536 , n460 );
nand ( n7949 , n7948 , n461 );
nand ( n7950 , n536 , n460 );
nand ( n7951 , n7949 , n7950 , n459 );
not ( n7952 , n7951 );
nand ( n7953 , n7947 , n7952 );
not ( n7954 , n7953 );
xnor ( n7955 , n7942 , n7954 );
not ( n7956 , n7836 );
not ( n7957 , n7035 );
or ( n7958 , n7956 , n7957 );
xor ( n7959 , n528 , n465 );
nand ( n7960 , n6987 , n7959 );
nand ( n7961 , n7958 , n7960 );
not ( n7962 , n7849 );
not ( n7963 , n7023 );
or ( n7964 , n7962 , n7963 );
xor ( n7965 , n530 , n463 );
nand ( n7966 , n7430 , n7965 );
nand ( n7967 , n7964 , n7966 );
xor ( n7968 , n7961 , n7967 );
not ( n7969 , n7868 );
not ( n7970 , n7449 );
or ( n7971 , n7969 , n7970 );
xor ( n7972 , n526 , n467 );
nand ( n7973 , n6955 , n7972 );
nand ( n7974 , n7971 , n7973 );
xor ( n7975 , n7968 , n7974 );
not ( n7976 , n7975 );
xor ( n7977 , n7955 , n7976 );
and ( n7978 , n7947 , n7951 );
not ( n7979 , n7947 );
and ( n7980 , n7979 , n7952 );
or ( n7981 , n7978 , n7980 );
not ( n7982 , n7763 );
or ( n7983 , n7752 , n7740 );
not ( n7984 , n7983 );
or ( n7985 , n7982 , n7984 );
nand ( n7986 , n7752 , n7740 );
nand ( n7987 , n7985 , n7986 );
or ( n7988 , n7981 , n7987 );
xor ( n7989 , n7771 , n7777 );
and ( n7990 , n7989 , n7784 );
and ( n7991 , n7771 , n7777 );
or ( n7992 , n7990 , n7991 );
nand ( n7993 , n7988 , n7992 );
nand ( n7994 , n7987 , n7981 );
nand ( n7995 , n7993 , n7994 );
xnor ( n7996 , n7977 , n7995 );
not ( n7997 , n7996 );
not ( n7998 , n7997 );
or ( n7999 , n7925 , n7998 );
xor ( n8000 , n7838 , n7851 );
xnor ( n8001 , n8000 , n7844 );
not ( n8002 , n8001 );
not ( n8003 , n7863 );
not ( n8004 , n7870 );
or ( n8005 , n8003 , n8004 );
or ( n8006 , n7870 , n7863 );
nand ( n8007 , n8005 , n8006 );
not ( n8008 , n7891 );
and ( n8009 , n8007 , n8008 );
not ( n8010 , n8007 );
and ( n8011 , n8010 , n7891 );
nor ( n8012 , n8009 , n8011 );
not ( n8013 , n8012 );
or ( n8014 , n8002 , n8013 );
not ( n8015 , n7704 );
not ( n8016 , n7696 );
or ( n8017 , n8015 , n8016 );
not ( n8018 , n7707 );
not ( n8019 , n7697 );
or ( n8020 , n8018 , n8019 );
nand ( n8021 , n8020 , n7716 );
nand ( n8022 , n8017 , n8021 );
nand ( n8023 , n8014 , n8022 );
not ( n8024 , n8001 );
not ( n8025 , n8012 );
nand ( n8026 , n8024 , n8025 );
nand ( n8027 , n8023 , n8026 );
nand ( n8028 , n7999 , n8027 );
nand ( n8029 , n7996 , n7923 );
nand ( n8030 , n8028 , n8029 );
not ( n8031 , n8030 );
not ( n8032 , n7975 );
not ( n8033 , n7955 );
nand ( n8034 , n8032 , n8033 );
not ( n8035 , n8034 );
not ( n8036 , n7995 );
or ( n8037 , n8035 , n8036 );
not ( n8038 , n8033 );
nand ( n8039 , n8038 , n7975 );
nand ( n8040 , n8037 , n8039 );
not ( n8041 , n8040 );
not ( n8042 , n7961 );
not ( n8043 , n7967 );
or ( n8044 , n8042 , n8043 );
or ( n8045 , n7967 , n7961 );
nand ( n8046 , n8045 , n7974 );
nand ( n8047 , n8044 , n8046 );
not ( n8048 , n8047 );
not ( n8049 , n7972 );
not ( n8050 , n6951 );
or ( n8051 , n8049 , n8050 );
xor ( n8052 , n525 , n467 );
nand ( n8053 , n6807 , n8052 );
nand ( n8054 , n8051 , n8053 );
not ( n8055 , n7965 );
not ( n8056 , n7023 );
or ( n8057 , n8055 , n8056 );
xor ( n8058 , n529 , n463 );
nand ( n8059 , n7026 , n8058 );
nand ( n8060 , n8057 , n8059 );
xor ( n8061 , n8054 , n8060 );
not ( n8062 , n7926 );
not ( n8063 , n7585 );
or ( n8064 , n8062 , n8063 );
xor ( n8065 , n461 , n531 );
nand ( n8066 , n7475 , n8065 );
nand ( n8067 , n8064 , n8066 );
not ( n8068 , n8067 );
and ( n8069 , n8061 , n8068 );
not ( n8070 , n8061 );
and ( n8071 , n8070 , n8067 );
nor ( n8072 , n8069 , n8071 );
not ( n8073 , n8072 );
or ( n8074 , n8048 , n8073 );
or ( n8075 , n8047 , n8072 );
nand ( n8076 , n8074 , n8075 );
not ( n8077 , n7959 );
not ( n8078 , n7035 );
or ( n8079 , n8077 , n8078 );
xor ( n8080 , n527 , n465 );
nand ( n8081 , n6987 , n8080 );
nand ( n8082 , n8079 , n8081 );
not ( n8083 , n8082 );
not ( n8084 , n7914 );
not ( n8085 , n7003 );
or ( n8086 , n8084 , n8085 );
xor ( n8087 , n523 , n469 );
nand ( n8088 , n6721 , n8087 );
nand ( n8089 , n8086 , n8088 );
not ( n8090 , n8089 );
not ( n8091 , n8090 );
or ( n8092 , n8083 , n8091 );
or ( n8093 , n8090 , n8082 );
nand ( n8094 , n8092 , n8093 );
xnor ( n8095 , n458 , n459 );
xor ( n8096 , n536 , n457 );
xor ( n8097 , n457 , n458 );
and ( n8098 , n8096 , n8097 );
and ( n8099 , n8095 , n8098 );
not ( n8100 , n8095 );
xor ( n8101 , n535 , n457 );
and ( n8102 , n8100 , n8101 );
or ( n8103 , n8099 , n8102 );
not ( n8104 , n8103 );
xor ( n8105 , n8094 , n8104 );
and ( n8106 , n8076 , n8105 );
not ( n8107 , n8076 );
not ( n8108 , n8105 );
and ( n8109 , n8107 , n8108 );
nor ( n8110 , n8106 , n8109 );
not ( n8111 , n8110 );
and ( n8112 , n8041 , n8111 );
and ( n8113 , n8040 , n8110 );
nor ( n8114 , n8112 , n8113 );
xor ( n8115 , n533 , n459 );
not ( n8116 , n8115 );
not ( n8117 , n7887 );
or ( n8118 , n8116 , n8117 );
not ( n8119 , n7879 );
not ( n8120 , n7877 );
or ( n8121 , n8119 , n8120 );
nand ( n8122 , n8121 , n7938 );
nand ( n8123 , n8118 , n8122 );
not ( n8124 , n8123 );
not ( n8125 , n7900 );
not ( n8126 , n6771 );
or ( n8127 , n8125 , n8126 );
xor ( n8128 , n471 , n521 );
nand ( n8129 , n8128 , n472 );
nand ( n8130 , n8127 , n8129 );
not ( n8131 , n8130 );
nand ( n8132 , n536 , n458 );
or ( n8133 , n536 , n458 );
nand ( n8134 , n8133 , n459 );
nand ( n8135 , n8132 , n457 , n8134 );
not ( n8136 , n8135 );
and ( n8137 , n8131 , n8136 );
and ( n8138 , n8130 , n8135 );
nor ( n8139 , n8137 , n8138 );
not ( n8140 , n8139 );
not ( n8141 , n8140 );
or ( n8142 , n8124 , n8141 );
not ( n8143 , n8123 );
nand ( n8144 , n8143 , n8139 );
nand ( n8145 , n8142 , n8144 );
xor ( n8146 , n7907 , n7909 );
and ( n8147 , n8146 , n7916 );
and ( n8148 , n7907 , n7909 );
or ( n8149 , n8147 , n8148 );
and ( n8150 , n8145 , n8149 );
not ( n8151 , n8145 );
not ( n8152 , n8149 );
and ( n8153 , n8151 , n8152 );
nor ( n8154 , n8150 , n8153 );
not ( n8155 , n8154 );
not ( n8156 , n7953 );
not ( n8157 , n7941 );
or ( n8158 , n8156 , n8157 );
nand ( n8159 , n8158 , n7931 );
nand ( n8160 , n7954 , n7940 );
nand ( n8161 , n8159 , n8160 );
buf ( n8162 , n8161 );
not ( n8163 , n8162 );
and ( n8164 , n8155 , n8163 );
not ( n8165 , n8155 );
and ( n8166 , n8165 , n8162 );
nor ( n8167 , n8164 , n8166 );
not ( n8168 , n7917 );
not ( n8169 , n8168 );
not ( n8170 , n7855 );
or ( n8171 , n8169 , n8170 );
nand ( n8172 , n8171 , n7894 );
nand ( n8173 , n7854 , n7917 );
nand ( n8174 , n8172 , n8173 );
xor ( n8175 , n8167 , n8174 );
and ( n8176 , n8114 , n8175 );
not ( n8177 , n8114 );
not ( n8178 , n8175 );
and ( n8179 , n8177 , n8178 );
nor ( n8180 , n8176 , n8179 );
not ( n8181 , n8180 );
nand ( n8182 , n8031 , n8181 );
nand ( n8183 , n8030 , n8180 );
buf ( n8184 , n8183 );
nand ( n8185 , n8182 , n8184 );
xor ( n8186 , n7981 , n7992 );
xnor ( n8187 , n8186 , n7987 );
xor ( n8188 , n7765 , n7785 );
and ( n8189 , n8188 , n7793 );
and ( n8190 , n7765 , n7785 );
or ( n8191 , n8189 , n8190 );
not ( n8192 , n8191 );
xor ( n8193 , n8187 , n8192 );
not ( n8194 , n8001 );
not ( n8195 , n8025 );
or ( n8196 , n8194 , n8195 );
nand ( n8197 , n8012 , n8024 );
nand ( n8198 , n8196 , n8197 );
not ( n8199 , n8022 );
and ( n8200 , n8198 , n8199 );
not ( n8201 , n8198 );
and ( n8202 , n8201 , n8022 );
nor ( n8203 , n8200 , n8202 );
and ( n8204 , n8193 , n8203 );
and ( n8205 , n8187 , n8192 );
or ( n8206 , n8204 , n8205 );
not ( n8207 , n8206 );
and ( n8208 , n7923 , n8027 );
not ( n8209 , n7923 );
not ( n8210 , n8027 );
and ( n8211 , n8209 , n8210 );
nor ( n8212 , n8208 , n8211 );
xnor ( n8213 , n7996 , n8212 );
not ( n8214 , n8213 );
or ( n8215 , n8207 , n8214 );
not ( n8216 , n7797 );
not ( n8217 , n7721 );
not ( n8218 , n8217 );
and ( n8219 , n8216 , n8218 );
nand ( n8220 , n7797 , n8217 );
buf ( n8221 , n7729 );
and ( n8222 , n8220 , n8221 );
nor ( n8223 , n8219 , n8222 );
xor ( n8224 , n8187 , n8192 );
xor ( n8225 , n8224 , n8203 );
nand ( n8226 , n8223 , n8225 );
nand ( n8227 , n8215 , n8226 );
not ( n8228 , n8227 );
not ( n8229 , n7672 );
not ( n8230 , n7671 );
or ( n8231 , n8229 , n8230 );
nand ( n8232 , n8231 , n7804 );
not ( n8233 , n8232 );
nand ( n8234 , n8228 , n7571 , n8233 );
not ( n8235 , n8206 );
not ( n8236 , n8213 );
nor ( n8237 , n8235 , n8236 );
not ( n8238 , n8223 );
not ( n8239 , n8225 );
nand ( n8240 , n8238 , n8239 );
or ( n8241 , n8237 , n8240 );
nand ( n8242 , n8235 , n8236 );
nand ( n8243 , n8241 , n8242 );
not ( n8244 , n8243 );
not ( n8245 , n7694 );
not ( n8246 , n7799 );
or ( n8247 , n8245 , n8246 );
nand ( n8248 , n8247 , n7668 );
nand ( n8249 , n7804 , n8248 );
not ( n8250 , n8249 );
nand ( n8251 , n8250 , n8228 );
nand ( n8252 , n8234 , n8244 , n8251 );
xnor ( n8253 , n8185 , n8252 );
buf ( n8254 , n8253 );
not ( n8255 , n8254 );
not ( n8256 , n8255 );
or ( n8257 , n7830 , n8256 );
not ( n8258 , n8253 );
not ( n8259 , n8258 );
not ( n8260 , n501 );
nand ( n8261 , n8259 , n8260 );
nand ( n8262 , n8257 , n8261 );
not ( n8263 , n8262 );
or ( n8264 , n7829 , n8263 );
not ( n8265 , n501 );
not ( n8266 , n8233 );
not ( n8267 , n7571 );
or ( n8268 , n8266 , n8267 );
nand ( n8269 , n8268 , n8249 );
buf ( n8270 , n8226 );
nand ( n8271 , n8269 , n8270 );
not ( n8272 , n8271 );
buf ( n8273 , n8240 );
not ( n8274 , n8273 );
or ( n8275 , n8272 , n8274 );
not ( n8276 , n8237 );
nand ( n8277 , n8276 , n8242 );
nand ( n8278 , n8275 , n8277 );
not ( n8279 , n8277 );
nand ( n8280 , n8279 , n8271 , n8273 );
nand ( n8281 , n8278 , n8280 );
not ( n8282 , n8281 );
not ( n8283 , n8282 );
or ( n8284 , n8265 , n8283 );
not ( n8285 , n8281 );
not ( n8286 , n8285 );
nand ( n8287 , n8286 , n8260 );
nand ( n8288 , n8284 , n8287 );
not ( n8289 , n2914 );
not ( n8290 , n502 );
not ( n8291 , n8290 );
or ( n8292 , n8289 , n8291 );
or ( n8293 , n8290 , n2914 );
nand ( n8294 , n8292 , n8293 );
nor ( n8295 , n8294 , n7827 );
not ( n8296 , n8295 );
not ( n8297 , n8296 );
nand ( n8298 , n8288 , n8297 );
nand ( n8299 , n8264 , n8298 );
xor ( n8300 , n7826 , n8299 );
xor ( n8301 , n7519 , n7551 );
xor ( n8302 , n8301 , n7822 );
not ( n8303 , n504 );
nand ( n8304 , n8303 , n503 );
not ( n8305 , n8304 );
buf ( n8306 , n8305 );
not ( n8307 , n8306 );
and ( n8308 , n503 , n8258 );
not ( n8309 , n503 );
and ( n8310 , n8309 , n8254 );
or ( n8311 , n8308 , n8310 );
not ( n8312 , n8311 );
or ( n8313 , n8307 , n8312 );
not ( n8314 , n8182 );
nand ( n8315 , n8234 , n8244 , n8251 );
not ( n8316 , n8315 );
or ( n8317 , n8314 , n8316 );
nand ( n8318 , n8317 , n8184 );
not ( n8319 , n8080 );
not ( n8320 , n7035 );
or ( n8321 , n8319 , n8320 );
xor ( n8322 , n526 , n465 );
nand ( n8323 , n6987 , n8322 );
nand ( n8324 , n8321 , n8323 );
not ( n8325 , n8058 );
nand ( n8326 , n7017 , n7022 );
not ( n8327 , n8326 );
not ( n8328 , n8327 );
or ( n8329 , n8325 , n8328 );
xor ( n8330 , n528 , n463 );
nand ( n8331 , n7026 , n8330 );
nand ( n8332 , n8329 , n8331 );
xnor ( n8333 , n8324 , n8332 );
not ( n8334 , n8101 );
xnor ( n8335 , n458 , n459 );
nand ( n8336 , n8335 , n8097 );
not ( n8337 , n8336 );
not ( n8338 , n8337 );
or ( n8339 , n8334 , n8338 );
xor ( n8340 , n534 , n457 );
nand ( n8341 , n7908 , n8340 );
nand ( n8342 , n8339 , n8341 );
not ( n8343 , n8342 );
and ( n8344 , n8333 , n8343 );
not ( n8345 , n8333 );
and ( n8346 , n8345 , n8342 );
nor ( n8347 , n8344 , n8346 );
not ( n8348 , n8347 );
not ( n8349 , n8348 );
not ( n8350 , n8065 );
nor ( n8351 , n7583 , n7474 );
not ( n8352 , n8351 );
or ( n8353 , n8350 , n8352 );
xor ( n8354 , n461 , n530 );
nand ( n8355 , n7474 , n8354 );
nand ( n8356 , n8353 , n8355 );
not ( n8357 , n8356 );
not ( n8358 , n8052 );
not ( n8359 , n7448 );
or ( n8360 , n8358 , n8359 );
xor ( n8361 , n524 , n467 );
nand ( n8362 , n6955 , n8361 );
nand ( n8363 , n8360 , n8362 );
and ( n8364 , n8357 , n8363 );
not ( n8365 , n8357 );
not ( n8366 , n8363 );
and ( n8367 , n8365 , n8366 );
nor ( n8368 , n8364 , n8367 );
not ( n8369 , n7880 );
not ( n8370 , n8115 );
or ( n8371 , n8369 , n8370 );
not ( n8372 , n7886 );
not ( n8373 , n7884 );
or ( n8374 , n8372 , n8373 );
xor ( n8375 , n532 , n459 );
nand ( n8376 , n8374 , n8375 );
nand ( n8377 , n8371 , n8376 );
not ( n8378 , n8377 );
xnor ( n8379 , n8368 , n8378 );
not ( n8380 , n8379 );
and ( n8381 , n536 , n457 );
not ( n8382 , n6727 );
not ( n8383 , n8128 );
or ( n8384 , n8382 , n8383 );
nand ( n8385 , n471 , n472 );
nand ( n8386 , n8384 , n8385 );
xor ( n8387 , n8381 , n8386 );
not ( n8388 , n8087 );
not ( n8389 , n7747 );
or ( n8390 , n8388 , n8389 );
xor ( n8391 , n522 , n469 );
nand ( n8392 , n6721 , n8391 );
nand ( n8393 , n8390 , n8392 );
xor ( n8394 , n8387 , n8393 );
not ( n8395 , n8394 );
and ( n8396 , n8380 , n8395 );
and ( n8397 , n8379 , n8394 );
nor ( n8398 , n8396 , n8397 );
not ( n8399 , n8398 );
not ( n8400 , n8399 );
or ( n8401 , n8349 , n8400 );
nand ( n8402 , n8347 , n8398 );
nand ( n8403 , n8401 , n8402 );
not ( n8404 , n8174 );
not ( n8405 , n8161 );
nand ( n8406 , n8405 , n8154 );
not ( n8407 , n8406 );
or ( n8408 , n8404 , n8407 );
not ( n8409 , n8154 );
nand ( n8410 , n8409 , n8161 );
nand ( n8411 , n8408 , n8410 );
and ( n8412 , n8403 , n8411 );
not ( n8413 , n8403 );
not ( n8414 , n8411 );
and ( n8415 , n8413 , n8414 );
nor ( n8416 , n8412 , n8415 );
not ( n8417 , n8144 );
not ( n8418 , n8149 );
or ( n8419 , n8417 , n8418 );
not ( n8420 , n8139 );
nand ( n8421 , n8420 , n8123 );
nand ( n8422 , n8419 , n8421 );
not ( n8423 , n8130 );
nor ( n8424 , n8423 , n8135 );
not ( n8425 , n8060 );
not ( n8426 , n8054 );
or ( n8427 , n8425 , n8426 );
or ( n8428 , n8054 , n8060 );
nand ( n8429 , n8428 , n8067 );
nand ( n8430 , n8427 , n8429 );
xor ( n8431 , n8424 , n8430 );
not ( n8432 , n8104 );
not ( n8433 , n8090 );
or ( n8434 , n8432 , n8433 );
nand ( n8435 , n8434 , n8082 );
nand ( n8436 , n8089 , n8103 );
nand ( n8437 , n8435 , n8436 );
xor ( n8438 , n8431 , n8437 );
xor ( n8439 , n8422 , n8438 );
not ( n8440 , n8047 );
not ( n8441 , n8108 );
or ( n8442 , n8440 , n8441 );
not ( n8443 , n8105 );
not ( n8444 , n8047 );
not ( n8445 , n8444 );
or ( n8446 , n8443 , n8445 );
not ( n8447 , n8072 );
nand ( n8448 , n8446 , n8447 );
nand ( n8449 , n8442 , n8448 );
xor ( n8450 , n8439 , n8449 );
and ( n8451 , n8416 , n8450 );
not ( n8452 , n8416 );
not ( n8453 , n8450 );
and ( n8454 , n8452 , n8453 );
nor ( n8455 , n8451 , n8454 );
not ( n8456 , n8455 );
not ( n8457 , n8110 );
not ( n8458 , n8457 );
not ( n8459 , n8178 );
or ( n8460 , n8458 , n8459 );
not ( n8461 , n8110 );
not ( n8462 , n8175 );
or ( n8463 , n8461 , n8462 );
nand ( n8464 , n8463 , n8040 );
nand ( n8465 , n8460 , n8464 );
not ( n8466 , n8465 );
nand ( n8467 , n8456 , n8466 );
nand ( n8468 , n8455 , n8465 );
nand ( n8469 , n8467 , n8468 );
and ( n8470 , n8318 , n8469 );
not ( n8471 , n8318 );
not ( n8472 , n8469 );
and ( n8473 , n8471 , n8472 );
nor ( n8474 , n8470 , n8473 );
not ( n8475 , n8474 );
and ( n8476 , n503 , n8475 );
not ( n8477 , n503 );
not ( n8478 , n8474 );
not ( n8479 , n8478 );
and ( n8480 , n8477 , n8479 );
nor ( n8481 , n8476 , n8480 );
nand ( n8482 , n8481 , n504 );
nand ( n8483 , n8313 , n8482 );
xor ( n8484 , n8302 , n8483 );
not ( n8485 , n6939 );
not ( n8486 , n7546 );
or ( n8487 , n8485 , n8486 );
and ( n8488 , n495 , n7339 );
not ( n8489 , n495 );
and ( n8490 , n8489 , n7340 );
nor ( n8491 , n8488 , n8490 );
nand ( n8492 , n8491 , n7326 );
nand ( n8493 , n8487 , n8492 );
not ( n8494 , n7410 );
not ( n8495 , n7321 );
and ( n8496 , n497 , n8495 );
not ( n8497 , n497 );
not ( n8498 , n7320 );
and ( n8499 , n8497 , n8498 );
or ( n8500 , n8496 , n8499 );
not ( n8501 , n8500 );
or ( n8502 , n8494 , n8501 );
and ( n8503 , n497 , n7384 );
not ( n8504 , n497 );
and ( n8505 , n8504 , n7383 );
or ( n8506 , n8503 , n8505 );
nand ( n8507 , n8506 , n7415 );
nand ( n8508 , n8502 , n8507 );
xor ( n8509 , n8493 , n8508 );
not ( n8510 , n7369 );
not ( n8511 , n7530 );
or ( n8512 , n8510 , n8511 );
and ( n8513 , n493 , n6787 );
not ( n8514 , n493 );
and ( n8515 , n8514 , n6790 );
nor ( n8516 , n8513 , n8515 );
nand ( n8517 , n8516 , n7405 );
nand ( n8518 , n8512 , n8517 );
xor ( n8519 , n6899 , n6908 );
xor ( n8520 , n8519 , n6923 );
xor ( n8521 , n8518 , n8520 );
xor ( n8522 , n6914 , n6922 );
not ( n8523 , n7369 );
not ( n8524 , n8516 );
or ( n8525 , n8523 , n8524 );
and ( n8526 , n493 , n6889 );
not ( n8527 , n493 );
and ( n8528 , n8527 , n6855 );
or ( n8529 , n8526 , n8528 );
nand ( n8530 , n8529 , n7405 );
nand ( n8531 , n8525 , n8530 );
xor ( n8532 , n8522 , n8531 );
nor ( n8533 , n6745 , n6843 );
and ( n8534 , n493 , n6862 );
not ( n8535 , n493 );
and ( n8536 , n8535 , n6863 );
or ( n8537 , n8534 , n8536 );
and ( n8538 , n8537 , n7369 );
not ( n8539 , n7405 );
and ( n8540 , n493 , n6745 );
not ( n8541 , n493 );
and ( n8542 , n8541 , n6846 );
nor ( n8543 , n8540 , n8542 );
nor ( n8544 , n8539 , n8543 );
nor ( n8545 , n8538 , n8544 );
or ( n8546 , n6846 , n494 );
nand ( n8547 , n8546 , n495 );
and ( n8548 , n6846 , n494 );
nor ( n8549 , n8548 , n739 );
nand ( n8550 , n8547 , n8549 );
nor ( n8551 , n8545 , n8550 );
xor ( n8552 , n8533 , n8551 );
not ( n8553 , n7405 );
not ( n8554 , n8537 );
or ( n8555 , n8553 , n8554 );
nand ( n8556 , n8529 , n7369 );
nand ( n8557 , n8555 , n8556 );
and ( n8558 , n8552 , n8557 );
or ( n8560 , n8558 , C0 );
and ( n8561 , n8532 , n8560 );
and ( n8562 , n8522 , n8531 );
or ( n8563 , n8561 , n8562 );
xor ( n8564 , n8521 , n8563 );
and ( n8565 , n8509 , n8564 );
and ( n8566 , n8493 , n8508 );
or ( n8567 , n8565 , n8566 );
not ( n8568 , n7813 );
not ( n8569 , n7682 );
or ( n8570 , n8568 , n8569 );
and ( n8571 , n499 , n7512 );
not ( n8572 , n499 );
and ( n8573 , n8572 , n7511 );
or ( n8574 , n8571 , n8573 );
nand ( n8575 , n8574 , n7558 );
nand ( n8576 , n8570 , n8575 );
xor ( n8577 , n8567 , n8576 );
not ( n8578 , n7828 );
nand ( n8579 , n8270 , n8273 );
xnor ( n8580 , n8269 , n8579 );
buf ( n8581 , n8580 );
and ( n8582 , n8581 , n8260 );
not ( n8583 , n8581 );
and ( n8584 , n8583 , n501 );
or ( n8585 , n8582 , n8584 );
not ( n8586 , n8585 );
or ( n8587 , n8578 , n8586 );
not ( n8588 , n501 );
not ( n8589 , n7811 );
not ( n8590 , n8589 );
or ( n8591 , n8588 , n8590 );
nand ( n8592 , n7812 , n8260 );
nand ( n8593 , n8591 , n8592 );
not ( n8594 , n8296 );
nand ( n8595 , n8593 , n8594 );
nand ( n8596 , n8587 , n8595 );
and ( n8597 , n8577 , n8596 );
and ( n8598 , n8567 , n8576 );
or ( n8599 , n8597 , n8598 );
and ( n8600 , n8484 , n8599 );
and ( n8601 , n8302 , n8483 );
or ( n8602 , n8600 , n8601 );
xor ( n8603 , n8300 , n8602 );
not ( n8604 , n7369 );
not ( n8605 , n7400 );
or ( n8606 , n8604 , n8605 );
not ( n8607 , n7524 );
not ( n8608 , n7405 );
or ( n8609 , n8607 , n8608 );
nand ( n8610 , n8606 , n8609 );
not ( n8611 , n6939 );
not ( n8612 , n7322 );
or ( n8613 , n8611 , n8612 );
nand ( n8614 , n7540 , n7326 );
nand ( n8615 , n8613 , n8614 );
xor ( n8616 , n8610 , n8615 );
xor ( n8617 , n6845 , n6882 );
xor ( n8618 , n8617 , n6929 );
and ( n8619 , n8616 , n8618 );
and ( n8620 , n8610 , n8615 );
or ( n8621 , n8619 , n8620 );
not ( n8622 , n7517 );
and ( n8623 , n497 , n7677 );
not ( n8624 , n497 );
not ( n8625 , n7677 );
and ( n8626 , n8624 , n8625 );
nor ( n8627 , n8623 , n8626 );
not ( n8628 , n8627 );
or ( n8629 , n8622 , n8628 );
nand ( n8630 , n7516 , n7415 );
nand ( n8631 , n8629 , n8630 );
xor ( n8632 , n8621 , n8631 );
not ( n8633 , n7813 );
xor ( n8634 , n499 , n8581 );
not ( n8635 , n8634 );
or ( n8636 , n8633 , n8635 );
xnor ( n8637 , n499 , n8589 );
nand ( n8638 , n8637 , n7558 );
nand ( n8639 , n8636 , n8638 );
xor ( n8640 , n8632 , n8639 );
not ( n8641 , n504 );
nand ( n8642 , n8234 , n8244 , n8251 );
not ( n8643 , n8642 );
not ( n8644 , n8643 );
nand ( n8645 , n8467 , n8182 );
not ( n8646 , n8645 );
and ( n8647 , n8644 , n8646 );
not ( n8648 , n8183 );
not ( n8649 , n8468 );
or ( n8650 , n8648 , n8649 );
nand ( n8651 , n8650 , n8467 );
not ( n8652 , n8651 );
nor ( n8653 , n8647 , n8652 );
not ( n8654 , n8403 );
nand ( n8655 , n8414 , n8654 );
not ( n8656 , n8655 );
not ( n8657 , n8450 );
or ( n8658 , n8656 , n8657 );
nand ( n8659 , n8411 , n8403 );
nand ( n8660 , n8658 , n8659 );
not ( n8661 , n8660 );
xor ( n8662 , n8422 , n8438 );
and ( n8663 , n8662 , n8449 );
and ( n8664 , n8422 , n8438 );
or ( n8665 , n8663 , n8664 );
not ( n8666 , n8665 );
xor ( n8667 , n8424 , n8430 );
and ( n8668 , n8667 , n8437 );
and ( n8669 , n8424 , n8430 );
or ( n8670 , n8668 , n8669 );
nand ( n8671 , n535 , n457 );
xor ( n8672 , n6967 , n8671 );
not ( n8673 , n8340 );
and ( n8674 , n8097 , n8335 );
not ( n8675 , n8674 );
or ( n8676 , n8673 , n8675 );
xor ( n8677 , n533 , n457 );
nand ( n8678 , n7908 , n8677 );
nand ( n8679 , n8676 , n8678 );
xor ( n8680 , n8672 , n8679 );
not ( n8681 , n8680 );
not ( n8682 , n8361 );
not ( n8683 , n6951 );
or ( n8684 , n8682 , n8683 );
xor ( n8685 , n523 , n467 );
nand ( n8686 , n6955 , n8685 );
nand ( n8687 , n8684 , n8686 );
not ( n8688 , n8391 );
not ( n8689 , n7747 );
or ( n8690 , n8688 , n8689 );
xor ( n8691 , n521 , n469 );
nand ( n8692 , n6721 , n8691 );
nand ( n8693 , n8690 , n8692 );
xor ( n8694 , n8687 , n8693 );
not ( n8695 , n8330 );
not ( n8696 , n8327 );
or ( n8697 , n8695 , n8696 );
xor ( n8698 , n527 , n463 );
nand ( n8699 , n7642 , n8698 );
nand ( n8700 , n8697 , n8699 );
xor ( n8701 , n8694 , n8700 );
not ( n8702 , n8701 );
or ( n8703 , n8681 , n8702 );
or ( n8704 , n8701 , n8680 );
nand ( n8705 , n8703 , n8704 );
xnor ( n8706 , n8670 , n8705 );
not ( n8707 , n8706 );
and ( n8708 , n8666 , n8707 );
and ( n8709 , n8665 , n8706 );
nor ( n8710 , n8708 , n8709 );
not ( n8711 , n8375 );
not ( n8712 , n7881 );
or ( n8713 , n8711 , n8712 );
xor ( n8714 , n531 , n459 );
nand ( n8715 , n7888 , n8714 );
nand ( n8716 , n8713 , n8715 );
not ( n8717 , n8716 );
not ( n8718 , n8354 );
buf ( n8719 , n7585 );
not ( n8720 , n8719 );
or ( n8721 , n8718 , n8720 );
xor ( n8722 , n461 , n529 );
nand ( n8723 , n7475 , n8722 );
nand ( n8724 , n8721 , n8723 );
not ( n8725 , n8724 );
xor ( n8726 , n8717 , n8725 );
not ( n8727 , n8322 );
buf ( n8728 , n6983 );
not ( n8729 , n8728 );
or ( n8730 , n8727 , n8729 );
xnor ( n8731 , n465 , n525 );
not ( n8732 , n8731 );
nand ( n8733 , n8732 , n6987 );
nand ( n8734 , n8730 , n8733 );
not ( n8735 , n8734 );
xor ( n8736 , n8726 , n8735 );
not ( n8737 , n8394 );
not ( n8738 , n8379 );
not ( n8739 , n8738 );
or ( n8740 , n8737 , n8739 );
not ( n8741 , n8394 );
not ( n8742 , n8741 );
not ( n8743 , n8379 );
or ( n8744 , n8742 , n8743 );
nand ( n8745 , n8744 , n8347 );
nand ( n8746 , n8740 , n8745 );
xor ( n8747 , n8736 , n8746 );
not ( n8748 , n8324 );
not ( n8749 , n8342 );
or ( n8750 , n8748 , n8749 );
or ( n8751 , n8324 , n8342 );
nand ( n8752 , n8751 , n8332 );
nand ( n8753 , n8750 , n8752 );
not ( n8754 , n8377 );
not ( n8755 , n8356 );
or ( n8756 , n8754 , n8755 );
not ( n8757 , n8378 );
not ( n8758 , n8357 );
or ( n8759 , n8757 , n8758 );
nand ( n8760 , n8759 , n8363 );
nand ( n8761 , n8756 , n8760 );
xor ( n8762 , n8381 , n8386 );
and ( n8763 , n8762 , n8393 );
and ( n8764 , n8381 , n8386 );
or ( n8765 , n8763 , n8764 );
xor ( n8766 , n8761 , n8765 );
not ( n8767 , n8766 );
and ( n8768 , n8753 , n8767 );
not ( n8769 , n8753 );
and ( n8770 , n8769 , n8766 );
nor ( n8771 , n8768 , n8770 );
xor ( n8772 , n8747 , n8771 );
nand ( n8773 , n8661 , n8710 , n8772 );
not ( n8774 , n8710 );
not ( n8775 , n8772 );
nand ( n8776 , n8774 , n8661 , n8775 );
nand ( n8777 , n8773 , n8776 );
not ( n8778 , n8777 );
nand ( n8779 , n8710 , n8775 );
not ( n8780 , n8779 );
not ( n8781 , n8775 );
nand ( n8782 , n8781 , n8774 );
not ( n8783 , n8782 );
or ( n8784 , n8780 , n8783 );
nand ( n8785 , n8784 , n8660 );
nand ( n8786 , n8778 , n8785 );
and ( n8787 , n8653 , n8786 );
not ( n8788 , n8653 );
not ( n8789 , n8786 );
and ( n8790 , n8788 , n8789 );
nor ( n8791 , n8787 , n8790 );
buf ( n8792 , n8791 );
and ( n8793 , n503 , n8792 );
not ( n8794 , n503 );
not ( n8795 , n8791 );
and ( n8796 , n8794 , n8795 );
nor ( n8797 , n8793 , n8796 );
not ( n8798 , n8797 );
or ( n8799 , n8641 , n8798 );
nand ( n8800 , n8481 , n8306 );
nand ( n8801 , n8799 , n8800 );
xor ( n8802 , n8640 , n8801 );
xor ( n8803 , n8610 , n8615 );
xor ( n8804 , n8803 , n8618 );
xor ( n8805 , n8518 , n8520 );
and ( n8806 , n8805 , n8563 );
and ( n8807 , n8518 , n8520 );
or ( n8808 , n8806 , n8807 );
not ( n8809 , n7517 );
not ( n8810 , n7421 );
or ( n8811 , n8809 , n8810 );
nand ( n8812 , n8500 , n7415 );
nand ( n8813 , n8811 , n8812 );
xor ( n8814 , n8808 , n8813 );
xor ( n8815 , n7532 , n7534 );
xor ( n8816 , n8815 , n7548 );
and ( n8817 , n8814 , n8816 );
and ( n8818 , n8808 , n8813 );
or ( n8819 , n8817 , n8818 );
xor ( n8820 , n8804 , n8819 );
not ( n8821 , n7828 );
not ( n8822 , n8288 );
or ( n8823 , n8821 , n8822 );
nand ( n8824 , n8585 , n8594 );
nand ( n8825 , n8823 , n8824 );
and ( n8826 , n8820 , n8825 );
and ( n8827 , n8804 , n8819 );
or ( n8828 , n8826 , n8827 );
xor ( n8829 , n8802 , n8828 );
and ( n8830 , n8603 , n8829 );
and ( n8831 , n8300 , n8602 );
or ( n8832 , n8830 , n8831 );
xor ( n8833 , n8640 , n8801 );
and ( n8834 , n8833 , n8828 );
and ( n8835 , n8640 , n8801 );
or ( n8836 , n8834 , n8835 );
xor ( n8837 , n7349 , n7364 );
and ( n8838 , n8837 , n7407 );
and ( n8839 , n7349 , n7364 );
or ( n8840 , n8838 , n8839 );
buf ( n8841 , n6939 );
not ( n8842 , n8841 );
not ( n8843 , n7511 );
and ( n8844 , n495 , n8843 );
not ( n8845 , n495 );
and ( n8846 , n8845 , n7511 );
or ( n8847 , n8844 , n8846 );
not ( n8848 , n8847 );
or ( n8849 , n8842 , n8848 );
nand ( n8850 , n7303 , n7326 );
nand ( n8851 , n8849 , n8850 );
xor ( n8852 , n8840 , n8851 );
not ( n8853 , n7415 );
not ( n8854 , n8627 );
or ( n8855 , n8853 , n8854 );
not ( n8856 , n497 );
not ( n8857 , n8589 );
or ( n8858 , n8856 , n8857 );
or ( n8859 , n8589 , n497 );
nand ( n8860 , n8858 , n8859 );
nand ( n8861 , n8860 , n7517 );
nand ( n8862 , n8855 , n8861 );
xor ( n8863 , n8852 , n8862 );
not ( n8864 , n7828 );
not ( n8865 , n501 );
not ( n8866 , n8475 );
not ( n8867 , n8866 );
or ( n8868 , n8865 , n8867 );
buf ( n8869 , n8475 );
nand ( n8870 , n8869 , n8260 );
nand ( n8871 , n8868 , n8870 );
not ( n8872 , n8871 );
or ( n8873 , n8864 , n8872 );
nand ( n8874 , n8262 , n8297 );
nand ( n8875 , n8873 , n8874 );
xor ( n8876 , n8863 , n8875 );
not ( n8877 , n8306 );
not ( n8878 , n8797 );
or ( n8879 , n8877 , n8878 );
not ( n8880 , n503 );
nand ( n8881 , n534 , n457 );
not ( n8882 , n6806 );
and ( n8883 , n8685 , n6948 );
not ( n8884 , n8883 );
or ( n8885 , n8882 , n8884 );
xor ( n8886 , n522 , n467 );
nand ( n8887 , n6955 , n8886 );
nand ( n8888 , n8885 , n8887 );
xor ( n8889 , n8881 , n8888 );
and ( n8890 , n8698 , n8327 );
xor ( n8891 , n526 , n463 );
and ( n8892 , n7642 , n8891 );
nor ( n8893 , n8890 , n8892 );
xnor ( n8894 , n8889 , n8893 );
not ( n8895 , n8894 );
not ( n8896 , n8691 );
not ( n8897 , n7747 );
or ( n8898 , n8896 , n8897 );
nand ( n8899 , n6721 , n469 );
nand ( n8900 , n8898 , n8899 );
not ( n8901 , n8900 );
not ( n8902 , n8901 );
not ( n8903 , n8677 );
not ( n8904 , n8674 );
or ( n8905 , n8903 , n8904 );
xor ( n8906 , n532 , n457 );
nand ( n8907 , n7908 , n8906 );
nand ( n8908 , n8905 , n8907 );
not ( n8909 , n8908 );
not ( n8910 , n8909 );
or ( n8911 , n8902 , n8910 );
nand ( n8912 , n8908 , n8900 );
nand ( n8913 , n8911 , n8912 );
and ( n8914 , n8913 , n8735 );
not ( n8915 , n8913 );
and ( n8916 , n8915 , n8734 );
nor ( n8917 , n8914 , n8916 );
not ( n8918 , n8917 );
and ( n8919 , n8895 , n8918 );
not ( n8920 , n8895 );
and ( n8921 , n8920 , n8917 );
nor ( n8922 , n8919 , n8921 );
or ( n8923 , n8761 , n8765 );
nand ( n8924 , n8923 , n8753 );
nand ( n8925 , n8761 , n8765 );
nand ( n8926 , n8924 , n8925 );
buf ( n8927 , n8926 );
xor ( n8928 , n8922 , n8927 );
not ( n8929 , n8928 );
not ( n8930 , n8746 );
not ( n8931 , n8736 );
not ( n8932 , n8931 );
not ( n8933 , n8932 );
or ( n8934 , n8930 , n8933 );
not ( n8935 , n8931 );
not ( n8936 , n8746 );
not ( n8937 , n8936 );
or ( n8938 , n8935 , n8937 );
not ( n8939 , n8771 );
nand ( n8940 , n8938 , n8939 );
nand ( n8941 , n8934 , n8940 );
not ( n8942 , n8941 );
or ( n8943 , n8929 , n8942 );
or ( n8944 , n8928 , n8941 );
nand ( n8945 , n8943 , n8944 );
not ( n8946 , n8717 );
not ( n8947 , n8946 );
not ( n8948 , n8725 );
not ( n8949 , n8948 );
or ( n8950 , n8947 , n8949 );
or ( n8951 , n8948 , n8946 );
nand ( n8952 , n8951 , n8735 );
nand ( n8953 , n8950 , n8952 );
nand ( n8954 , n8671 , n471 );
not ( n8955 , n8954 );
not ( n8956 , n8679 );
or ( n8957 , n8955 , n8956 );
or ( n8958 , n8671 , n471 );
nand ( n8959 , n8957 , n8958 );
not ( n8960 , n8693 );
not ( n8961 , n8687 );
or ( n8962 , n8960 , n8961 );
nor ( n8963 , n8693 , n8687 );
not ( n8964 , n8700 );
or ( n8965 , n8963 , n8964 );
nand ( n8966 , n8962 , n8965 );
not ( n8967 , n8966 );
xor ( n8968 , n8959 , n8967 );
xor ( n8969 , n530 , n459 );
and ( n8970 , n7887 , n8969 );
not ( n8971 , n7887 );
not ( n8972 , n8714 );
xnor ( n8973 , n459 , n460 );
nor ( n8974 , n8972 , n8973 );
and ( n8975 , n8971 , n8974 );
or ( n8976 , n8970 , n8975 );
not ( n8977 , n8722 );
not ( n8978 , n7585 );
or ( n8979 , n8977 , n8978 );
xor ( n8980 , n528 , n461 );
nand ( n8981 , n7475 , n8980 );
nand ( n8982 , n8979 , n8981 );
xor ( n8983 , n8976 , n8982 );
not ( n8984 , n6986 );
not ( n8985 , n8984 );
not ( n8986 , n6979 );
nor ( n8987 , n8986 , n8731 );
not ( n8988 , n8987 );
or ( n8989 , n8985 , n8988 );
xor ( n8990 , n524 , n465 );
nand ( n8991 , n6987 , n8990 );
nand ( n8992 , n8989 , n8991 );
xor ( n8993 , n8983 , n8992 );
xnor ( n8994 , n8968 , n8993 );
xor ( n8995 , n8953 , n8994 );
not ( n8996 , n8701 );
nand ( n8997 , n8996 , n8680 );
not ( n8998 , n8997 );
not ( n8999 , n8670 );
or ( n9000 , n8998 , n8999 );
not ( n9001 , n8680 );
nand ( n9002 , n9001 , n8701 );
nand ( n9003 , n9000 , n9002 );
xor ( n9004 , n8995 , n9003 );
not ( n9005 , n9004 );
nand ( n9006 , n8945 , n9005 );
not ( n9007 , n9006 );
not ( n9008 , n8945 );
not ( n9009 , n9005 );
nand ( n9010 , n9008 , n9009 );
not ( n9011 , n9010 );
or ( n9012 , n9007 , n9011 );
not ( n9013 , n8772 );
not ( n9014 , n8706 );
nand ( n9015 , n9013 , n9014 );
or ( n9016 , n8775 , n9014 );
nand ( n9017 , n9016 , n8665 );
nand ( n9018 , n9015 , n9017 );
not ( n9019 , n9018 );
nand ( n9020 , n9012 , n9019 );
not ( n9021 , n9020 );
not ( n9022 , n9021 );
nand ( n9023 , n9009 , n9008 );
nand ( n9024 , n9023 , n9018 , n9006 );
not ( n9025 , n9024 );
not ( n9026 , n9025 );
nand ( n9027 , n9022 , n9026 );
not ( n9028 , n9027 );
not ( n9029 , n9028 );
nand ( n9030 , n8467 , n8182 );
nor ( n9031 , n8777 , n9030 );
not ( n9032 , n9031 );
not ( n9033 , n8642 );
or ( n9034 , n9032 , n9033 );
or ( n9035 , n8651 , n8777 );
nand ( n9036 , n9035 , n8785 );
not ( n9037 , n9036 );
nand ( n9038 , n9034 , n9037 );
not ( n9039 , n9038 );
not ( n9040 , n9039 );
or ( n9041 , n9029 , n9040 );
not ( n9042 , n9039 );
nand ( n9043 , n9042 , n9027 );
nand ( n9044 , n9041 , n9043 );
not ( n9045 , n9044 );
not ( n9046 , n9045 );
and ( n9047 , n8880 , n9046 );
not ( n9048 , n8880 );
buf ( n9049 , n9044 );
not ( n9050 , n9049 );
and ( n9051 , n9048 , n9050 );
nor ( n9052 , n9047 , n9051 );
or ( n9053 , n9052 , n8303 );
nand ( n9054 , n8879 , n9053 );
xor ( n9055 , n8876 , n9054 );
xor ( n9056 , n8836 , n9055 );
xor ( n9057 , n8621 , n8631 );
and ( n9058 , n9057 , n8639 );
and ( n9059 , n8621 , n8631 );
or ( n9060 , n9058 , n9059 );
xor ( n9061 , n7350 , n7358 );
and ( n9062 , n9061 , n7363 );
and ( n9063 , n7350 , n7358 );
or ( n9064 , n9062 , n9063 );
not ( n9065 , n7369 );
xor ( n9066 , n493 , n7321 );
not ( n9067 , n9066 );
or ( n9068 , n9065 , n9067 );
nand ( n9069 , n7388 , n7405 );
nand ( n9070 , n9068 , n9069 );
xor ( n9071 , n9064 , n9070 );
and ( n9072 , n489 , n6855 );
not ( n9073 , n6848 );
xor ( n9074 , n489 , n6836 );
not ( n9075 , n9074 );
or ( n9076 , n9073 , n9075 );
nand ( n9077 , n7352 , n6867 );
nand ( n9078 , n9076 , n9077 );
xor ( n9079 , n9072 , n9078 );
not ( n9080 , n6842 );
not ( n9081 , n491 );
not ( n9082 , n7396 );
or ( n9083 , n9081 , n9082 );
nand ( n9084 , n7395 , n6892 );
nand ( n9085 , n9083 , n9084 );
not ( n9086 , n9085 );
or ( n9087 , n9080 , n9086 );
nand ( n9088 , n7344 , n6719 );
nand ( n9089 , n9087 , n9088 );
xor ( n9090 , n9079 , n9089 );
xor ( n9091 , n9071 , n9090 );
not ( n9092 , n7558 );
not ( n9093 , n8634 );
or ( n9094 , n9092 , n9093 );
not ( n9095 , n499 );
not ( n9096 , n8282 );
or ( n9097 , n9095 , n9096 );
not ( n9098 , n499 );
nand ( n9099 , n9098 , n8281 );
nand ( n9100 , n9097 , n9099 );
nand ( n9101 , n9100 , n7813 );
nand ( n9102 , n9094 , n9101 );
xor ( n9103 , n9091 , n9102 );
xor ( n9104 , n6932 , n7328 );
and ( n9105 , n9104 , n7408 );
and ( n9106 , n6932 , n7328 );
or ( n9107 , n9105 , n9106 );
xor ( n9108 , n9103 , n9107 );
xor ( n9109 , n9060 , n9108 );
xor ( n9110 , n7409 , n7825 );
and ( n9111 , n9110 , n8299 );
and ( n9112 , n7409 , n7825 );
or ( n9113 , n9111 , n9112 );
xor ( n9114 , n9109 , n9113 );
xor ( n9115 , n9056 , n9114 );
xor ( n9116 , n8832 , n9115 );
xor ( n9117 , n8300 , n8602 );
xor ( n9118 , n9117 , n8829 );
xor ( n9119 , n8804 , n8819 );
xor ( n9120 , n9119 , n8825 );
xor ( n9121 , n8808 , n8813 );
xor ( n9122 , n9121 , n8816 );
not ( n9123 , n6939 );
not ( n9124 , n8491 );
or ( n9125 , n9123 , n9124 );
and ( n9126 , n495 , n6836 );
not ( n9127 , n495 );
and ( n9128 , n9127 , n6837 );
nor ( n9129 , n9126 , n9128 );
nand ( n9130 , n7326 , n9129 );
nand ( n9131 , n9125 , n9130 );
xor ( n9132 , n8522 , n8531 );
xor ( n9133 , n9132 , n8560 );
xor ( n9134 , n9131 , n9133 );
not ( n9135 , n7410 );
not ( n9136 , n8506 );
or ( n9137 , n9135 , n9136 );
and ( n9138 , n497 , n7395 );
not ( n9139 , n497 );
and ( n9140 , n9139 , n7396 );
nor ( n9141 , n9138 , n9140 );
nand ( n9142 , n9141 , n7415 );
nand ( n9143 , n9137 , n9142 );
and ( n9144 , n9134 , n9143 );
and ( n9145 , n9131 , n9133 );
or ( n9146 , n9144 , n9145 );
not ( n9147 , n7813 );
not ( n9148 , n8574 );
or ( n9149 , n9147 , n9148 );
and ( n9150 , n499 , n7298 );
not ( n9151 , n499 );
and ( n9152 , n9151 , n7301 );
or ( n9153 , n9150 , n9152 );
nand ( n9154 , n9153 , n7558 );
nand ( n9155 , n9149 , n9154 );
xor ( n9156 , n9146 , n9155 );
xor ( n9157 , n8493 , n8508 );
xor ( n9158 , n9157 , n8564 );
and ( n9159 , n9156 , n9158 );
and ( n9160 , n9146 , n9155 );
or ( n9161 , n9159 , n9160 );
xor ( n9162 , n9122 , n9161 );
not ( n9163 , n8306 );
not ( n9164 , n503 );
not ( n9165 , n8285 );
or ( n9166 , n9164 , n9165 );
buf ( n9167 , n8281 );
nand ( n9168 , n9167 , n8880 );
nand ( n9169 , n9166 , n9168 );
not ( n9170 , n9169 );
or ( n9171 , n9163 , n9170 );
nand ( n9172 , n8311 , n504 );
nand ( n9173 , n9171 , n9172 );
and ( n9174 , n9162 , n9173 );
and ( n9175 , n9122 , n9161 );
or ( n9176 , n9174 , n9175 );
xor ( n9177 , n9120 , n9176 );
xor ( n9178 , n8302 , n8483 );
xor ( n9179 , n9178 , n8599 );
and ( n9180 , n9177 , n9179 );
and ( n9181 , n9120 , n9176 );
or ( n9182 , n9180 , n9181 );
or ( n9183 , n9118 , n9182 );
not ( n9184 , n9183 );
xor ( n9185 , n9120 , n9176 );
xor ( n9186 , n9185 , n9179 );
not ( n9187 , n8594 );
and ( n9188 , n501 , n7677 );
not ( n9189 , n501 );
and ( n9190 , n9189 , n8625 );
nor ( n9191 , n9188 , n9190 );
not ( n9192 , n9191 );
or ( n9193 , n9187 , n9192 );
nand ( n9194 , n8593 , n7828 );
nand ( n9195 , n9193 , n9194 );
not ( n9196 , n6939 );
not ( n9197 , n9129 );
or ( n9198 , n9196 , n9197 );
and ( n9199 , n495 , n6790 );
not ( n9200 , n495 );
and ( n9201 , n9200 , n6787 );
or ( n9202 , n9199 , n9201 );
nand ( n9203 , n9202 , n7326 );
nand ( n9204 , n9198 , n9203 );
xor ( n9205 , n8533 , n8551 );
xor ( n9206 , n9205 , n8557 );
xor ( n9207 , n9204 , n9206 );
not ( n9208 , n8550 );
not ( n9209 , n8545 );
not ( n9210 , n9209 );
or ( n9211 , n9208 , n9210 );
or ( n9212 , n9209 , n8550 );
nand ( n9213 , n9211 , n9212 );
not ( n9214 , n6939 );
not ( n9215 , n9202 );
or ( n9216 , n9214 , n9215 );
and ( n9217 , n495 , n6889 );
not ( n9218 , n495 );
and ( n9219 , n9218 , n6855 );
or ( n9220 , n9217 , n9219 );
nand ( n9221 , n9220 , n7326 );
nand ( n9222 , n9216 , n9221 );
xor ( n9223 , n9213 , n9222 );
nor ( n9224 , n6745 , n7370 );
not ( n9225 , n7326 );
and ( n9226 , n495 , n6863 );
not ( n9227 , n495 );
and ( n9228 , n9227 , n6862 );
nor ( n9229 , n9226 , n9228 );
not ( n9230 , n9229 );
or ( n9231 , n9225 , n9230 );
nand ( n9232 , n9220 , n6939 );
nand ( n9233 , n9231 , n9232 );
xor ( n9234 , n9224 , n9233 );
and ( n9235 , n6846 , n496 );
and ( n9236 , n6745 , n6933 );
not ( n9237 , n497 );
nor ( n9238 , n9236 , n9237 );
nor ( n9239 , n9235 , n9238 , n1554 );
not ( n9240 , n7326 );
and ( n9241 , n495 , n6846 );
not ( n9242 , n495 );
and ( n116794 , n9242 , n6745 );
nor ( n9243 , n9241 , n116794 );
not ( n9244 , n9243 );
or ( n9245 , n9240 , n9244 );
nand ( n9246 , n9229 , n6939 );
nand ( n9247 , n9245 , n9246 );
and ( n9248 , n9239 , n9247 );
and ( n9249 , n9234 , n9248 );
and ( n9250 , n9224 , n9233 );
or ( n9251 , n9249 , n9250 );
and ( n9252 , n9223 , n9251 );
and ( n9253 , n9213 , n9222 );
or ( n9254 , n9252 , n9253 );
and ( n9255 , n9207 , n9254 );
and ( n9256 , n9204 , n9206 );
or ( n9257 , n9255 , n9256 );
xor ( n9258 , n9131 , n9133 );
xor ( n9259 , n9258 , n9143 );
xor ( n9260 , n9257 , n9259 );
and ( n9261 , n499 , n8495 );
not ( n9262 , n499 );
not ( n9263 , n7320 );
and ( n9264 , n9262 , n9263 );
or ( n9265 , n9261 , n9264 );
not ( n9266 , n9265 );
not ( n9267 , n7558 );
or ( n9268 , n9266 , n9267 );
not ( n9269 , n9153 );
or ( n9270 , n9269 , n7814 );
nand ( n9271 , n9268 , n9270 );
and ( n9272 , n9260 , n9271 );
and ( n9273 , n9257 , n9259 );
or ( n9274 , n9272 , n9273 );
xor ( n9275 , n9195 , n9274 );
not ( n9276 , n8306 );
not ( n9277 , n503 );
not ( n9278 , n8581 );
not ( n9279 , n9278 );
or ( n9280 , n9277 , n9279 );
nand ( n9281 , n8581 , n8880 );
nand ( n9282 , n9280 , n9281 );
not ( n9283 , n9282 );
or ( n9284 , n9276 , n9283 );
nand ( n9285 , n9169 , n504 );
nand ( n9286 , n9284 , n9285 );
and ( n9287 , n9275 , n9286 );
and ( n9288 , n9195 , n9274 );
or ( n9289 , n9287 , n9288 );
xor ( n9290 , n8567 , n8576 );
xor ( n9291 , n9290 , n8596 );
xor ( n9292 , n9289 , n9291 );
xor ( n9293 , n9122 , n9161 );
xor ( n9294 , n9293 , n9173 );
and ( n9295 , n9292 , n9294 );
and ( n9296 , n9289 , n9291 );
or ( n9297 , n9295 , n9296 );
nor ( n9298 , n9186 , n9297 );
xor ( n9299 , n9289 , n9291 );
xor ( n9300 , n9299 , n9294 );
xor ( n9301 , n9146 , n9155 );
xor ( n9302 , n9301 , n9158 );
not ( n9303 , n7410 );
not ( n9304 , n9141 );
or ( n9305 , n9303 , n9304 );
and ( n9306 , n497 , n7339 );
not ( n9307 , n497 );
and ( n9308 , n9307 , n7340 );
nor ( n9309 , n9306 , n9308 );
nand ( n9310 , n9309 , n7415 );
nand ( n9311 , n9305 , n9310 );
not ( n9312 , n7813 );
not ( n9313 , n9265 );
or ( n9314 , n9312 , n9313 );
and ( n9315 , n499 , n7384 );
not ( n9316 , n499 );
and ( n9317 , n9316 , n7383 );
or ( n9318 , n9315 , n9317 );
nand ( n9319 , n9318 , n7558 );
nand ( n9320 , n9314 , n9319 );
xor ( n9321 , n9311 , n9320 );
xor ( n9322 , n9204 , n9206 );
xor ( n9323 , n9322 , n9254 );
and ( n9324 , n9321 , n9323 );
and ( n9325 , n9311 , n9320 );
or ( n9326 , n9324 , n9325 );
not ( n9327 , n7828 );
not ( n9328 , n9191 );
or ( n9329 , n9327 , n9328 );
not ( n9330 , n501 );
not ( n9331 , n7512 );
or ( n9332 , n9330 , n9331 );
nand ( n9333 , n7511 , n8260 );
nand ( n9334 , n9332 , n9333 );
nand ( n9335 , n9334 , n8594 );
nand ( n9336 , n9329 , n9335 );
xor ( n9337 , n9326 , n9336 );
not ( n9338 , n504 );
not ( n9339 , n9282 );
or ( n9340 , n9338 , n9339 );
xnor ( n9341 , n503 , n8589 );
nand ( n9342 , n9341 , n8306 );
nand ( n9343 , n9340 , n9342 );
and ( n9344 , n9337 , n9343 );
and ( n9345 , n9326 , n9336 );
or ( n9346 , n9344 , n9345 );
xor ( n9347 , n9302 , n9346 );
xor ( n9348 , n9195 , n9274 );
xor ( n9349 , n9348 , n9286 );
and ( n9350 , n9347 , n9349 );
and ( n9351 , n9302 , n9346 );
or ( n9352 , n9350 , n9351 );
nor ( n9353 , n9300 , n9352 );
nor ( n9354 , n9298 , n9353 );
not ( n9355 , n9354 );
not ( n9356 , n7813 );
and ( n9357 , n499 , n7395 );
not ( n9358 , n499 );
and ( n9359 , n9358 , n7396 );
nor ( n9360 , n9357 , n9359 );
not ( n9361 , n9360 );
or ( n9362 , n9356 , n9361 );
and ( n9363 , n499 , n7339 );
not ( n9364 , n499 );
and ( n9365 , n9364 , n7340 );
nor ( n9366 , n9363 , n9365 );
not ( n9367 , n9366 );
or ( n9368 , n9367 , n7557 );
nand ( n9369 , n9362 , n9368 );
not ( n9370 , n7415 );
and ( n9371 , n497 , n6787 );
not ( n9372 , n497 );
and ( n9373 , n9372 , n6790 );
nor ( n9374 , n9371 , n9373 );
not ( n9375 , n9374 );
or ( n9376 , n9370 , n9375 );
and ( n9377 , n497 , n6836 );
not ( n9378 , n497 );
and ( n9379 , n9378 , n6837 );
nor ( n9380 , n9377 , n9379 );
nand ( n9381 , n7410 , n9380 );
nand ( n9382 , n9376 , n9381 );
xor ( n9383 , n9224 , n9233 );
xor ( n9384 , n9383 , n9248 );
xor ( n9385 , n9382 , n9384 );
xor ( n9386 , n9239 , n9247 );
not ( n9387 , n7410 );
not ( n9388 , n9374 );
or ( n9389 , n9387 , n9388 );
and ( n9390 , n497 , n6889 );
not ( n9391 , n497 );
not ( n9392 , n6889 );
and ( n9393 , n9391 , n9392 );
or ( n9394 , n9390 , n9393 );
nand ( n9395 , n9394 , n7415 );
nand ( n9396 , n9389 , n9395 );
xor ( n9397 , n9386 , n9396 );
nor ( n9398 , n6938 , n6745 );
not ( n9399 , n7415 );
and ( n9400 , n497 , n6863 );
not ( n9401 , n497 );
and ( n9402 , n9401 , n6862 );
nor ( n9403 , n9400 , n9402 );
not ( n9404 , n9403 );
or ( n9405 , n9399 , n9404 );
nand ( n9406 , n9394 , n7410 );
nand ( n9407 , n9405 , n9406 );
xor ( n9408 , n9398 , n9407 );
or ( n9409 , n6846 , n498 );
nand ( n9410 , n9409 , n499 );
and ( n9411 , n6846 , n498 );
nor ( n9412 , n9411 , n1009 );
and ( n9413 , n9410 , n9412 );
not ( n9414 , n7415 );
and ( n9415 , n497 , n6846 );
not ( n9416 , n497 );
and ( n9417 , n9416 , n6745 );
nor ( n9418 , n9415 , n9417 );
not ( n9419 , n9418 );
or ( n9420 , n9414 , n9419 );
nand ( n9421 , n9403 , n7410 );
nand ( n9422 , n9420 , n9421 );
and ( n9423 , n9413 , n9422 );
and ( n9424 , n9408 , n9423 );
and ( n9425 , n9398 , n9407 );
or ( n9426 , n9424 , n9425 );
and ( n9427 , n9397 , n9426 );
and ( n9428 , n9386 , n9396 );
or ( n9429 , n9427 , n9428 );
xor ( n9430 , n9385 , n9429 );
xor ( n9431 , n9369 , n9430 );
not ( n9432 , n7828 );
xor ( n9433 , n501 , n9263 );
not ( n9434 , n9433 );
or ( n9435 , n9432 , n9434 );
and ( n9436 , n8295 , n8260 );
and ( n9437 , n7383 , n9436 );
and ( n9438 , n8290 , n8880 , n501 );
and ( n9439 , n7384 , n9438 );
nor ( n9440 , n9437 , n9439 );
nand ( n9441 , n9435 , n9440 );
and ( n9442 , n9431 , n9441 );
and ( n9443 , n9369 , n9430 );
or ( n9444 , n9442 , n9443 );
not ( n9445 , n504 );
and ( n9446 , n503 , n7677 );
not ( n9447 , n503 );
and ( n9448 , n9447 , n8625 );
nor ( n9449 , n9446 , n9448 );
not ( n9450 , n9449 );
or ( n9451 , n9445 , n9450 );
and ( n9452 , n503 , n7511 );
not ( n9453 , n503 );
and ( n9454 , n9453 , n7512 );
nor ( n9455 , n9452 , n9454 );
nand ( n9456 , n9455 , n8306 );
nand ( n9457 , n9451 , n9456 );
xor ( n9458 , n9444 , n9457 );
xor ( n9459 , n9382 , n9384 );
and ( n9460 , n9459 , n9429 );
and ( n9461 , n9382 , n9384 );
or ( n9462 , n9460 , n9461 );
not ( n9463 , n7410 );
not ( n9464 , n9309 );
or ( n9465 , n9463 , n9464 );
not ( n9466 , n9380 );
not ( n9467 , n7414 );
or ( n9468 , n9466 , n9467 );
nand ( n9469 , n9465 , n9468 );
xor ( n9470 , n9213 , n9222 );
xor ( n9471 , n9470 , n9251 );
xor ( n9472 , n9469 , n9471 );
not ( n9473 , n7813 );
not ( n9474 , n9318 );
or ( n9475 , n9473 , n9474 );
nand ( n9476 , n9360 , n7558 );
nand ( n9477 , n9475 , n9476 );
xor ( n9478 , n9472 , n9477 );
xor ( n9479 , n9462 , n9478 );
not ( n9480 , n8594 );
not ( n9481 , n9433 );
or ( n9482 , n9480 , n9481 );
and ( n9483 , n501 , n7301 );
not ( n9484 , n501 );
and ( n9485 , n9484 , n7298 );
nor ( n9486 , n9483 , n9485 );
nand ( n9487 , n9486 , n7828 );
nand ( n9488 , n9482 , n9487 );
xor ( n9489 , n9479 , n9488 );
xor ( n9490 , n9458 , n9489 );
not ( n9491 , n8306 );
not ( n9492 , n503 );
not ( n9493 , n7298 );
or ( n9494 , n9492 , n9493 );
nand ( n9495 , n7301 , n8880 );
nand ( n9496 , n9494 , n9495 );
not ( n9497 , n9496 );
or ( n9498 , n9491 , n9497 );
nand ( n9499 , n9455 , n504 );
nand ( n9500 , n9498 , n9499 );
not ( n9501 , n7813 );
not ( n9502 , n9366 );
or ( n9503 , n9501 , n9502 );
and ( n9504 , n499 , n6836 );
not ( n9505 , n499 );
and ( n9506 , n9505 , n6837 );
nor ( n9507 , n9504 , n9506 );
nand ( n9508 , n7558 , n9507 );
nand ( n9509 , n9503 , n9508 );
xor ( n9510 , n9386 , n9396 );
xor ( n9511 , n9510 , n9426 );
xor ( n9512 , n9509 , n9511 );
and ( n9513 , n501 , n7383 );
not ( n9514 , n501 );
and ( n9515 , n9514 , n7384 );
nor ( n9516 , n9513 , n9515 );
not ( n9517 , n9516 );
not ( n9518 , n7828 );
or ( n9519 , n9517 , n9518 );
and ( n9520 , n7395 , n9436 );
not ( n9521 , n7395 );
and ( n9522 , n9521 , n9438 );
nor ( n9523 , n9520 , n9522 );
nand ( n9524 , n9519 , n9523 );
and ( n9525 , n9512 , n9524 );
and ( n9526 , n9509 , n9511 );
or ( n9527 , n9525 , n9526 );
xor ( n9528 , n9500 , n9527 );
xor ( n9529 , n9369 , n9430 );
xor ( n9530 , n9529 , n9441 );
and ( n9531 , n9528 , n9530 );
and ( n9532 , n9500 , n9527 );
or ( n9533 , n9531 , n9532 );
or ( n9534 , n9490 , n9533 );
not ( n9535 , n7813 );
not ( n9536 , n9507 );
or ( n9537 , n9535 , n9536 );
and ( n9538 , n499 , n6787 );
not ( n9539 , n499 );
and ( n9540 , n9539 , n6790 );
nor ( n9541 , n9538 , n9540 );
nand ( n9542 , n9541 , n7558 );
nand ( n9543 , n9537 , n9542 );
xor ( n9544 , n9398 , n9407 );
xor ( n9545 , n9544 , n9423 );
xor ( n9546 , n9543 , n9545 );
not ( n9547 , n7827 );
and ( n9548 , n501 , n7395 );
not ( n9549 , n501 );
not ( n9550 , n7394 );
and ( n9551 , n9549 , n9550 );
nor ( n9552 , n9548 , n9551 );
not ( n9553 , n9552 );
or ( n9554 , n9547 , n9553 );
and ( n9555 , n501 , n7339 );
not ( n9556 , n501 );
and ( n9557 , n9556 , n7340 );
nor ( n9558 , n9555 , n9557 );
nand ( n9559 , n9558 , n8594 );
nand ( n9560 , n9554 , n9559 );
and ( n9561 , n9546 , n9560 );
and ( n9562 , n9543 , n9545 );
or ( n9563 , n9561 , n9562 );
xor ( n9564 , n9509 , n9511 );
xor ( n9565 , n9564 , n9524 );
xor ( n9566 , n9563 , n9565 );
not ( n9567 , n504 );
not ( n9568 , n9496 );
or ( n9569 , n9567 , n9568 );
not ( n9570 , n7321 );
nand ( n9571 , n9570 , n8305 );
nand ( n9572 , n9569 , n9571 );
and ( n9573 , n9566 , n9572 );
and ( n9574 , n9563 , n9565 );
or ( n9575 , n9573 , n9574 );
xor ( n9576 , n9500 , n9527 );
xor ( n9577 , n9576 , n9530 );
xor ( n9578 , n9575 , n9577 );
xor ( n9579 , n9413 , n9422 );
not ( n9580 , n7813 );
not ( n9581 , n9541 );
or ( n9582 , n9580 , n9581 );
and ( n9583 , n499 , n6889 );
not ( n9584 , n499 );
and ( n9585 , n9584 , n9392 );
or ( n9586 , n9583 , n9585 );
nand ( n9587 , n9586 , n7558 );
nand ( n9588 , n9582 , n9587 );
xor ( n9589 , n9579 , n9588 );
nor ( n9590 , n6745 , n7411 );
not ( n9591 , n7813 );
not ( n9592 , n9586 );
or ( n9593 , n9591 , n9592 );
and ( n9594 , n499 , n6863 );
not ( n9595 , n499 );
and ( n9596 , n9595 , n6862 );
nor ( n9597 , n9594 , n9596 );
nand ( n9598 , n9597 , n7558 );
nand ( n9599 , n9593 , n9598 );
xor ( n9600 , n9590 , n9599 );
or ( n9601 , n6846 , n500 );
nand ( n9602 , n9601 , n501 );
and ( n9603 , n6846 , n500 );
nor ( n9604 , n9603 , n1808 );
and ( n9605 , n9602 , n9604 );
not ( n9606 , n7813 );
not ( n9607 , n9597 );
or ( n9608 , n9606 , n9607 );
and ( n9609 , n499 , n6846 );
not ( n9610 , n499 );
and ( n9611 , n9610 , n6745 );
nor ( n9612 , n9609 , n9611 );
nand ( n9613 , n9612 , n7558 );
nand ( n9614 , n9608 , n9613 );
and ( n9615 , n9605 , n9614 );
and ( n9616 , n9600 , n9615 );
and ( n9617 , n9590 , n9599 );
or ( n9618 , n9616 , n9617 );
and ( n9619 , n9589 , n9618 );
and ( n9620 , n9579 , n9588 );
or ( n9621 , n9619 , n9620 );
xor ( n9622 , n9543 , n9545 );
xor ( n9623 , n9622 , n9560 );
xor ( n9624 , n9621 , n9623 );
nand ( n9625 , n503 , n504 );
or ( n9626 , n9625 , n9263 );
nor ( n9627 , n8303 , n503 );
nand ( n9628 , n9263 , n9627 );
and ( n9629 , n7384 , n880 );
not ( n9630 , n7384 );
and ( n9631 , n9630 , n503 );
nor ( n9632 , n9629 , n9631 );
nand ( n9633 , n9632 , n8306 );
nand ( n9634 , n9626 , n9628 , n9633 );
xor ( n9635 , n9624 , n9634 );
not ( n9636 , n9635 );
not ( n9637 , n8594 );
and ( n9638 , n6836 , n501 );
not ( n9639 , n6836 );
and ( n9640 , n9639 , n8260 );
nor ( n9641 , n9638 , n9640 );
not ( n9642 , n9641 );
or ( n9643 , n9637 , n9642 );
nand ( n9644 , n9558 , n7827 );
nand ( n9645 , n9643 , n9644 );
xor ( n9646 , n9579 , n9588 );
xor ( n9647 , n9646 , n9618 );
xor ( n9648 , n9645 , n9647 );
not ( n9649 , n8306 );
and ( n9650 , n503 , n7394 );
not ( n9651 , n503 );
and ( n9652 , n9651 , n9550 );
nor ( n9653 , n9650 , n9652 );
not ( n9654 , n9653 );
or ( n9655 , n9649 , n9654 );
nand ( n9656 , n9632 , n504 );
nand ( n9657 , n9655 , n9656 );
and ( n9658 , n9648 , n9657 );
and ( n9659 , n9645 , n9647 );
or ( n9660 , n9658 , n9659 );
not ( n9661 , n9660 );
nand ( n9662 , n9636 , n9661 );
not ( n9663 , n8295 );
and ( n9664 , n6787 , n501 );
not ( n9665 , n6787 );
and ( n9666 , n9665 , n8260 );
nor ( n9667 , n9664 , n9666 );
not ( n9668 , n9667 );
or ( n9669 , n9663 , n9668 );
nand ( n9670 , n9641 , n7827 );
nand ( n9671 , n9669 , n9670 );
xor ( n9672 , n9590 , n9599 );
xor ( n9673 , n9672 , n9615 );
xor ( n9674 , n9671 , n9673 );
not ( n9675 , n8306 );
not ( n9676 , n503 );
not ( n9677 , n7340 );
or ( n9678 , n9676 , n9677 );
nand ( n9679 , n7339 , n8880 );
nand ( n9680 , n9678 , n9679 );
not ( n9681 , n9680 );
or ( n9682 , n9675 , n9681 );
nand ( n9683 , n9653 , n504 );
nand ( n9684 , n9682 , n9683 );
and ( n9685 , n9674 , n9684 );
and ( n9686 , n9671 , n9673 );
or ( n9687 , n9685 , n9686 );
xor ( n9688 , n9645 , n9647 );
xor ( n9689 , n9688 , n9657 );
xor ( n9690 , n9687 , n9689 );
xor ( n9691 , n9605 , n9614 );
not ( n9692 , n7827 );
not ( n9693 , n9667 );
or ( n9694 , n9692 , n9693 );
not ( n9695 , n501 );
not ( n9696 , n6889 );
or ( n9697 , n9695 , n9696 );
nand ( n9698 , n9392 , n8260 );
nand ( n9699 , n9697 , n9698 );
nand ( n9700 , n9699 , n8295 );
nand ( n9701 , n9694 , n9700 );
xor ( n9702 , n9691 , n9701 );
and ( n9703 , n6846 , n7813 );
not ( n9704 , n7827 );
or ( n9705 , n6862 , n501 );
or ( n9706 , n6747 , n6859 );
nand ( n9707 , n9706 , n501 );
nand ( n9708 , n9705 , n9707 );
not ( n9709 , n9708 );
or ( n9710 , n9704 , n9709 );
and ( n9711 , n9436 , n6846 );
and ( n9712 , n9438 , n6745 );
nor ( n9713 , n9711 , n9712 );
nand ( n9714 , n9710 , n9713 );
not ( n9715 , n9714 );
or ( n9716 , n6846 , n502 );
nand ( n9717 , n9716 , n503 );
and ( n9718 , n6846 , n502 );
nor ( n9719 , n9718 , n8260 );
nand ( n9720 , n9717 , n9719 );
nor ( n9721 , n9715 , n9720 );
xor ( n9722 , n9703 , n9721 );
not ( n9723 , n7827 );
not ( n9724 , n9699 );
or ( n9725 , n9723 , n9724 );
nand ( n9726 , n8295 , n9708 );
nand ( n9727 , n9725 , n9726 );
and ( n9728 , n9722 , n9727 );
or ( n9730 , n9728 , C0 );
and ( n9731 , n9702 , n9730 );
and ( n9732 , n9691 , n9701 );
or ( n9733 , n9731 , n9732 );
xor ( n9734 , n9691 , n9701 );
xor ( n9735 , n9734 , n9730 );
not ( n9736 , n9680 );
or ( n9737 , n9736 , n8303 );
and ( n9738 , n503 , n6837 );
not ( n9739 , n503 );
and ( n9740 , n9739 , n6836 );
nor ( n9741 , n9738 , n9740 );
or ( n9742 , n9741 , n8304 );
nand ( n9743 , n9737 , n9742 );
or ( n9744 , n9735 , n9743 );
not ( n9745 , n6790 );
not ( n9746 , n503 );
or ( n9747 , n9745 , n9746 );
nand ( n9748 , n6787 , n8880 );
nand ( n9749 , n9747 , n9748 );
not ( n9750 , n9749 );
not ( n9751 , n8306 );
or ( n9752 , n9750 , n9751 );
or ( n9753 , n9741 , n8303 );
nand ( n9754 , n9752 , n9753 );
xor ( n9755 , n9703 , n9721 );
xor ( n9756 , n9755 , n9727 );
nor ( n9757 , n9754 , n9756 );
and ( n9758 , n8880 , n9392 );
not ( n9759 , n8880 );
and ( n9760 , n9759 , n6889 );
nor ( n9761 , n9758 , n9760 );
not ( n9762 , n9761 );
not ( n9763 , n8304 );
and ( n9764 , n9762 , n9763 );
and ( n9765 , n9749 , n504 );
nor ( n9766 , n9764 , n9765 );
xor ( n9767 , n9714 , n9720 );
nand ( n9768 , n9766 , n9767 );
not ( n9769 , n7827 );
nor ( n9770 , n9769 , n6745 );
not ( n9771 , n8304 );
not ( n9772 , n6846 );
and ( n9773 , n9771 , n9772 );
not ( n9774 , n503 );
not ( n9775 , n6862 );
or ( n9776 , n9774 , n9775 );
nand ( n9777 , n6863 , n8880 );
nand ( n9778 , n9776 , n9777 );
and ( n9779 , n9778 , n504 );
nor ( n9780 , n9773 , n9779 );
and ( n9781 , n6846 , n504 );
or ( n9782 , n9781 , n8880 );
nor ( n9783 , n9780 , n9782 );
xor ( n9784 , n9770 , n9783 );
not ( n9785 , n8305 );
not ( n9786 , n9778 );
or ( n9787 , n9785 , n9786 );
or ( n9788 , n9761 , n8303 );
nand ( n9789 , n9787 , n9788 );
and ( n9790 , n9784 , n9789 );
or ( n9792 , n9790 , C0 );
and ( n9793 , n9768 , n9792 );
nor ( n9794 , n9766 , n9767 );
nor ( n9795 , n9793 , n9794 );
or ( n9796 , n9757 , n9795 );
nand ( n9797 , n9754 , n9756 );
nand ( n9798 , n9796 , n9797 );
nand ( n9799 , n9744 , n9798 );
nand ( n9800 , n9735 , n9743 );
nand ( n9801 , n9799 , n9800 );
xor ( n9802 , n9733 , n9801 );
xor ( n9803 , n9671 , n9673 );
xor ( n9804 , n9803 , n9684 );
and ( n9805 , n9802 , n9804 );
and ( n9806 , n9733 , n9801 );
or ( n9807 , n9805 , n9806 );
and ( n9808 , n9690 , n9807 );
and ( n9809 , n9687 , n9689 );
or ( n9810 , n9808 , n9809 );
and ( n9811 , n9662 , n9810 );
nor ( n9812 , n9636 , n9661 );
nor ( n9813 , n9811 , n9812 );
xor ( n9814 , n9563 , n9565 );
xor ( n9815 , n9814 , n9572 );
xor ( n9816 , n9621 , n9623 );
and ( n9817 , n9816 , n9634 );
and ( n9818 , n9621 , n9623 );
or ( n9819 , n9817 , n9818 );
nor ( n9820 , n9815 , n9819 );
or ( n9821 , n9813 , n9820 );
nand ( n9822 , n9815 , n9819 );
nand ( n9823 , n9821 , n9822 );
and ( n9824 , n9578 , n9823 );
and ( n9825 , n9575 , n9577 );
or ( n9826 , n9824 , n9825 );
and ( n9827 , n9534 , n9826 );
and ( n9828 , n9490 , n9533 );
nor ( n9829 , n9827 , n9828 );
xor ( n9830 , n9311 , n9320 );
xor ( n9831 , n9830 , n9323 );
xor ( n9832 , n9462 , n9478 );
and ( n9833 , n9832 , n9488 );
and ( n9834 , n9462 , n9478 );
or ( n9835 , n9833 , n9834 );
xor ( n9836 , n9831 , n9835 );
not ( n9837 , n7828 );
not ( n9838 , n9334 );
or ( n9839 , n9837 , n9838 );
nand ( n9840 , n9486 , n8594 );
nand ( n9841 , n9839 , n9840 );
xor ( n9842 , n9469 , n9471 );
and ( n9843 , n9842 , n9477 );
and ( n9844 , n9469 , n9471 );
or ( n9845 , n9843 , n9844 );
xor ( n9846 , n9841 , n9845 );
not ( n9847 , n8306 );
not ( n9848 , n9449 );
or ( n9849 , n9847 , n9848 );
nand ( n9850 , n9341 , n504 );
nand ( n9851 , n9849 , n9850 );
xor ( n9852 , n9846 , n9851 );
xor ( n9853 , n9836 , n9852 );
xor ( n9854 , n9444 , n9457 );
and ( n9855 , n9854 , n9489 );
and ( n9856 , n9444 , n9457 );
or ( n9857 , n9855 , n9856 );
nor ( n9858 , n9853 , n9857 );
or ( n9859 , n9829 , n9858 );
nand ( n9860 , n9853 , n9857 );
nand ( n9861 , n9859 , n9860 );
not ( n9862 , n9861 );
xor ( n9863 , n9302 , n9346 );
xor ( n9864 , n9863 , n9349 );
xor ( n9865 , n9257 , n9259 );
xor ( n9866 , n9865 , n9271 );
xor ( n9867 , n9841 , n9845 );
and ( n9868 , n9867 , n9851 );
and ( n9869 , n9841 , n9845 );
or ( n9870 , n9868 , n9869 );
xor ( n9871 , n9866 , n9870 );
xor ( n9872 , n9326 , n9336 );
xor ( n9873 , n9872 , n9343 );
and ( n9874 , n9871 , n9873 );
and ( n9875 , n9866 , n9870 );
or ( n9876 , n9874 , n9875 );
nor ( n9877 , n9864 , n9876 );
xor ( n9878 , n9866 , n9870 );
xor ( n9879 , n9878 , n9873 );
xor ( n9880 , n9831 , n9835 );
and ( n9881 , n9880 , n9852 );
and ( n9882 , n9831 , n9835 );
or ( n9883 , n9881 , n9882 );
nor ( n9884 , n9879 , n9883 );
nor ( n9885 , n9877 , n9884 );
not ( n9886 , n9885 );
or ( n9887 , n9862 , n9886 );
not ( n9888 , n9877 );
and ( n9889 , n9879 , n9883 );
and ( n9890 , n9888 , n9889 );
and ( n9891 , n9864 , n9876 );
nor ( n9892 , n9890 , n9891 );
nand ( n9893 , n9887 , n9892 );
not ( n9894 , n9893 );
or ( n9895 , n9355 , n9894 );
not ( n9896 , n9298 );
and ( n9897 , n9300 , n9352 );
and ( n9898 , n9896 , n9897 );
and ( n9899 , n9186 , n9297 );
nor ( n9900 , n9898 , n9899 );
nand ( n9901 , n9895 , n9900 );
not ( n9902 , n9901 );
or ( n9903 , n9184 , n9902 );
nand ( n9904 , n9118 , n9182 );
nand ( n9905 , n9903 , n9904 );
xor ( n9906 , n9116 , n9905 );
not ( n9907 , n454 );
nand ( n9908 , n9906 , n9907 );
nand ( n9909 , n6712 , n9908 );
nand ( n9910 , n5964 , n6706 );
not ( n9911 , n9910 );
and ( n9912 , n6703 , n9911 );
not ( n9913 , n6703 );
and ( n9914 , n9913 , n9910 );
nor ( n9915 , n9912 , n9914 );
nand ( n9916 , n9915 , n454 );
nand ( n9917 , n9183 , n9904 );
xnor ( n9918 , n9901 , n9917 );
nand ( n9919 , n9918 , n9907 );
nand ( n9920 , n9916 , n9919 );
not ( n9921 , n454 );
nand ( n9922 , n6701 , n6133 );
buf ( n9923 , n6700 );
not ( n9924 , n9923 );
and ( n9925 , n9922 , n9924 );
not ( n9926 , n9922 );
and ( n9927 , n9926 , n9923 );
nor ( n9928 , n9925 , n9927 );
not ( n9929 , n9928 );
or ( n9930 , n9921 , n9929 );
not ( n9931 , n9353 );
not ( n9932 , n9897 );
nand ( n9933 , n9931 , n9932 );
buf ( n9934 , n9893 );
xnor ( n9935 , n9933 , n9934 );
nand ( n9936 , n9935 , n9907 );
nand ( n9937 , n9930 , n9936 );
not ( n9938 , n9907 );
not ( n9939 , n9858 );
nand ( n9940 , n9939 , n9860 );
xor ( n9941 , n9940 , n9829 );
not ( n9942 , n9941 );
or ( n9943 , n9938 , n9942 );
buf ( n9944 , n6678 );
not ( n9945 , n6692 );
nand ( n9946 , n9945 , n6687 );
not ( n9947 , n9946 );
and ( n9948 , n9944 , n9947 );
not ( n9949 , n9944 );
and ( n9950 , n9949 , n9946 );
nor ( n9951 , n9948 , n9950 );
nand ( n9952 , n9951 , n454 );
nand ( n9953 , n9943 , n9952 );
nand ( n9954 , n6677 , n6383 );
buf ( n9955 , n6673 );
not ( n9956 , n9955 );
and ( n9957 , n9954 , n9956 );
not ( n9958 , n9954 );
and ( n9959 , n9958 , n9955 );
nor ( n9960 , n9957 , n9959 );
nand ( n9961 , n9960 , n454 );
buf ( n9962 , n9826 );
not ( n9963 , n9962 );
not ( n9964 , n9828 );
nand ( n9965 , n9964 , n9534 );
not ( n9966 , n9965 );
or ( n9967 , n9963 , n9966 );
or ( n9968 , n9965 , n9962 );
nand ( n9969 , n9967 , n9968 );
nand ( n9970 , n9969 , n9907 );
nand ( n9971 , n9961 , n9970 );
buf ( n9972 , n6663 );
not ( n9973 , n9972 );
not ( n9974 , n9973 );
not ( n9975 , n6670 );
nand ( n9976 , n9975 , n6672 );
not ( n9977 , n9976 );
not ( n9978 , n9977 );
or ( n9979 , n9974 , n9978 );
and ( n9980 , n9976 , n9972 );
not ( n9981 , n454 );
nor ( n9982 , n9980 , n9981 );
nand ( n9983 , n9979 , n9982 );
xor ( n9984 , n9575 , n9577 );
xor ( n9985 , n9984 , n9823 );
nand ( n9986 , n9985 , n9907 );
nand ( n9987 , n9983 , n9986 );
not ( n9988 , n6662 );
nand ( n9989 , n9988 , n6660 );
buf ( n9990 , n6643 );
not ( n9991 , n9990 );
and ( n9992 , n9989 , n9991 );
not ( n9993 , n9989 );
and ( n9994 , n9993 , n9990 );
nor ( n9995 , n9992 , n9994 );
nand ( n9996 , n9995 , n454 );
and ( n9997 , n9662 , n9810 );
nor ( n9998 , n9997 , n9812 );
not ( n9999 , n9998 );
not ( n10000 , n9999 );
not ( n10001 , n9820 );
nand ( n10002 , n10001 , n9822 );
not ( n10003 , n10002 );
or ( n10004 , n10000 , n10003 );
or ( n10005 , n10002 , n9999 );
nand ( n10006 , n10004 , n10005 );
nand ( n10007 , n10006 , n9907 );
nand ( n10008 , n9996 , n10007 );
buf ( n10009 , n6609 );
not ( n10010 , n10009 );
not ( n10011 , n10010 );
not ( n10012 , n6640 );
nand ( n10013 , n10012 , n6642 );
not ( n10014 , n10013 );
not ( n10015 , n10014 );
or ( n10016 , n10011 , n10015 );
and ( n10017 , n10013 , n10009 );
nor ( n10018 , n10017 , n9981 );
nand ( n10019 , n10016 , n10018 );
not ( n10020 , n9810 );
not ( n10021 , n9812 );
nand ( n10022 , n10021 , n9662 );
not ( n10023 , n10022 );
or ( n10024 , n10020 , n10023 );
or ( n10025 , n10022 , n9810 );
nand ( n10026 , n10024 , n10025 );
nand ( n10027 , n10026 , n9907 );
nand ( n10028 , n10019 , n10027 );
not ( n10029 , n552 );
not ( n10030 , n551 );
not ( n10031 , n716 );
xor ( n10032 , n5241 , n5251 );
and ( n10033 , n10032 , n5259 );
and ( n10034 , n5241 , n5251 );
or ( n10035 , n10033 , n10034 );
xor ( n10036 , n5263 , n5273 );
and ( n10037 , n10036 , n5285 );
and ( n10038 , n5263 , n5273 );
or ( n10039 , n10037 , n10038 );
xor ( n10040 , n10035 , n10039 );
not ( n10041 , n3573 );
not ( n10042 , n5239 );
or ( n10043 , n10041 , n10042 );
not ( n10044 , n491 );
not ( n10045 , n2949 );
or ( n10046 , n10044 , n10045 );
nand ( n10047 , n2613 , n2948 );
nand ( n10048 , n10046 , n10047 );
nand ( n10049 , n10048 , n2606 );
nand ( n10050 , n10043 , n10049 );
not ( n10051 , n4553 );
not ( n10052 , n5257 );
or ( n10053 , n10051 , n10052 );
and ( n10054 , n456 , n480 );
not ( n10055 , n456 );
and ( n10056 , n10055 , n464 );
nor ( n10057 , n10054 , n10056 );
and ( n10058 , n489 , n10057 );
not ( n10059 , n489 );
and ( n10060 , n10059 , n5160 );
or ( n10061 , n10058 , n10060 );
nand ( n10062 , n10061 , n4547 );
nand ( n10063 , n10053 , n10062 );
xor ( n10064 , n10050 , n10063 );
not ( n10065 , n5271 );
not ( n10066 , n893 );
or ( n10067 , n10065 , n10066 );
nand ( n10068 , n912 , n497 );
nand ( n10069 , n10067 , n10068 );
xor ( n10070 , n10064 , n10069 );
and ( n10071 , n10040 , n10070 );
and ( n10072 , n10035 , n10039 );
or ( n10073 , n10071 , n10072 );
or ( n10074 , n912 , n893 );
nand ( n10075 , n10074 , n497 );
not ( n10076 , n1026 );
not ( n10077 , n495 );
not ( n10078 , n4077 );
or ( n10079 , n10077 , n10078 );
nand ( n10080 , n4076 , n813 );
nand ( n10081 , n10079 , n10080 );
not ( n10082 , n10081 );
or ( n10083 , n10076 , n10082 );
not ( n10084 , n495 );
not ( n10085 , n3859 );
or ( n10086 , n10084 , n10085 );
nand ( n10087 , n3858 , n813 );
nand ( n10088 , n10086 , n10087 );
nand ( n10089 , n10088 , n1086 );
nand ( n10090 , n10083 , n10089 );
xor ( n10091 , n10075 , n10090 );
not ( n10092 , n2606 );
not ( n10093 , n491 );
not ( n10094 , n1043 );
or ( n10095 , n10093 , n10094 );
nand ( n10096 , n5278 , n2613 );
nand ( n10097 , n10095 , n10096 );
not ( n10098 , n10097 );
or ( n10099 , n10092 , n10098 );
nand ( n10100 , n10048 , n3573 );
nand ( n10101 , n10099 , n10100 );
xor ( n10102 , n10091 , n10101 );
and ( n10103 , n489 , n778 );
not ( n10104 , n2959 );
not ( n10105 , n493 );
not ( n10106 , n2178 );
or ( n10107 , n10105 , n10106 );
not ( n10108 , n2178 );
nand ( n10109 , n10108 , n739 );
nand ( n10110 , n10107 , n10109 );
not ( n10111 , n10110 );
or ( n10112 , n10104 , n10111 );
nand ( n10113 , n5283 , n2967 );
nand ( n10114 , n10112 , n10113 );
xor ( n10115 , n10103 , n10114 );
not ( n10116 , n1086 );
not ( n10117 , n5247 );
or ( n10118 , n10116 , n10117 );
nand ( n10119 , n10088 , n1026 );
nand ( n10120 , n10118 , n10119 );
not ( n10121 , n10120 );
and ( n10122 , n10115 , n10121 );
and ( n10123 , n10103 , n10114 );
or ( n10124 , n10122 , n10123 );
xor ( n10125 , n10102 , n10124 );
xor ( n10126 , n10050 , n10063 );
and ( n10127 , n10126 , n10069 );
and ( n10128 , n10050 , n10063 );
or ( n10129 , n10127 , n10128 );
xor ( n10130 , n10120 , n10129 );
not ( n10131 , n4547 );
not ( n10132 , n489 );
not ( n10133 , n4971 );
or ( n10134 , n10132 , n10133 );
not ( n10135 , n489 );
nand ( n10136 , n10135 , n951 );
nand ( n10137 , n10134 , n10136 );
not ( n10138 , n10137 );
or ( n10139 , n10131 , n10138 );
nand ( n10140 , n10061 , n4553 );
nand ( n10141 , n10139 , n10140 );
not ( n10142 , n2967 );
not ( n10143 , n10110 );
or ( n10144 , n10142 , n10143 );
not ( n10145 , n493 );
not ( n10146 , n2547 );
not ( n10147 , n10146 );
or ( n10148 , n10145 , n10147 );
nand ( n10149 , n4093 , n739 );
nand ( n10150 , n10148 , n10149 );
nand ( n10151 , n10150 , n724 );
nand ( n10152 , n10144 , n10151 );
xor ( n10153 , n10141 , n10152 );
not ( n10154 , n4999 );
and ( n10155 , n489 , n10154 );
xor ( n10156 , n10153 , n10155 );
xor ( n10157 , n10130 , n10156 );
xor ( n10158 , n10125 , n10157 );
xor ( n10159 , n10073 , n10158 );
xor ( n10160 , n10103 , n10114 );
xor ( n10161 , n10160 , n10121 );
xor ( n10162 , n5288 , n5289 );
and ( n10163 , n10162 , n5294 );
and ( n10164 , n5288 , n5289 );
or ( n10165 , n10163 , n10164 );
xor ( n10166 , n10161 , n10165 );
xor ( n10167 , n5231 , n5260 );
and ( n10168 , n10167 , n5286 );
and ( n10169 , n5231 , n5260 );
or ( n10170 , n10168 , n10169 );
and ( n10171 , n10166 , n10170 );
and ( n10172 , n10161 , n10165 );
or ( n10173 , n10171 , n10172 );
xor ( n10174 , n10159 , n10173 );
not ( n10175 , n10174 );
xor ( n10176 , n10035 , n10039 );
xor ( n10177 , n10176 , n10070 );
xor ( n10178 , n10161 , n10165 );
xor ( n10179 , n10178 , n10170 );
xor ( n10180 , n10177 , n10179 );
xor ( n10181 , n5295 , n5299 );
and ( n10182 , n10181 , n5304 );
and ( n10183 , n5295 , n5299 );
or ( n10184 , n10182 , n10183 );
and ( n10185 , n10180 , n10184 );
and ( n10186 , n10177 , n10179 );
or ( n10187 , n10185 , n10186 );
not ( n10188 , n10187 );
nand ( n10189 , n10175 , n10188 );
not ( n10190 , n10175 );
not ( n10191 , n10188 );
nand ( n10192 , n10190 , n10191 );
and ( n10193 , n10189 , n10192 );
xor ( n10194 , n10177 , n10179 );
xor ( n10195 , n10194 , n10184 );
buf ( n10196 , n10195 );
xor ( n10197 , n5287 , n5305 );
and ( n10198 , n10197 , n5310 );
and ( n10199 , n5287 , n5305 );
or ( n10200 , n10198 , n10199 );
buf ( n10201 , n10200 );
nand ( n10202 , n10196 , n10201 );
nand ( n10203 , n10193 , n10202 );
not ( n10204 , n5315 );
not ( n10205 , n5311 );
and ( n10206 , n10204 , n10205 );
nor ( n10207 , n5202 , n5206 );
nor ( n10208 , n10206 , n10207 );
not ( n10209 , n10208 );
not ( n10210 , n5222 );
or ( n10211 , n10209 , n10210 );
not ( n10212 , n5326 );
not ( n10213 , n5202 );
not ( n10214 , n5206 );
nor ( n10215 , n10213 , n10214 );
not ( n10216 , n10215 );
or ( n10217 , n10212 , n10216 );
nand ( n10218 , n10217 , n5316 );
not ( n10219 , n10218 );
nand ( n10220 , n10211 , n10219 );
or ( n10221 , n10203 , n10220 );
or ( n10222 , n10196 , n10201 );
not ( n10223 , n10222 );
nor ( n10224 , n10223 , n10193 );
nand ( n10225 , n10220 , n10224 );
not ( n10226 , n10202 );
nor ( n10227 , n10226 , n10222 );
and ( n10228 , n10193 , n10227 );
nor ( n10229 , n10202 , n10193 );
nor ( n10230 , n10228 , n10229 );
nand ( n10231 , n10221 , n10225 , n10230 );
not ( n10232 , n10231 );
or ( n10233 , n10031 , n10232 );
xor ( n10234 , n5471 , n5477 );
and ( n10235 , n10234 , n5484 );
and ( n10236 , n5471 , n5477 );
or ( n10237 , n10235 , n10236 );
xor ( n10238 , n5492 , n5498 );
and ( n10239 , n10238 , n5505 );
and ( n10240 , n5492 , n5498 );
or ( n10241 , n10239 , n10240 );
xor ( n10242 , n10237 , n10241 );
not ( n10243 , n5496 );
not ( n10244 , n4835 );
or ( n10245 , n10243 , n10244 );
xor ( n10246 , n512 , n489 );
nand ( n10247 , n4838 , n10246 );
nand ( n10248 , n10245 , n10247 );
not ( n10249 , n5482 );
not ( n10250 , n2083 );
or ( n10251 , n10249 , n10250 );
nand ( n10252 , n2086 , n497 );
nand ( n10253 , n10251 , n10252 );
xor ( n10254 , n10248 , n10253 );
not ( n10255 , n5490 );
not ( n10256 , n5487 );
or ( n10257 , n10255 , n10256 );
xor ( n10258 , n491 , n510 );
nand ( n10259 , n2764 , n10258 );
nand ( n10260 , n10257 , n10259 );
xor ( n10261 , n10254 , n10260 );
xnor ( n10262 , n10242 , n10261 );
or ( n10263 , n5485 , n5510 );
nand ( n10264 , n10263 , n5506 );
nand ( n10265 , n5485 , n5510 );
nand ( n10266 , n10264 , n10265 );
not ( n10267 , n10266 );
not ( n10268 , n10267 );
nand ( n10269 , n514 , n489 );
not ( n10270 , n5475 );
not ( n10271 , n2028 );
or ( n10272 , n10270 , n10271 );
xor ( n10273 , n508 , n493 );
nand ( n10274 , n2031 , n10273 );
nand ( n10275 , n10272 , n10274 );
xor ( n10276 , n10269 , n10275 );
not ( n10277 , n5503 );
not ( n10278 , n5389 );
or ( n10279 , n10277 , n10278 );
xor ( n10280 , n506 , n495 );
nand ( n10281 , n5392 , n10280 );
nand ( n10282 , n10279 , n10281 );
not ( n10283 , n10282 );
xnor ( n10284 , n10276 , n10283 );
not ( n10285 , n10284 );
nand ( n10286 , n5531 , n5520 );
not ( n10287 , n10286 );
not ( n10288 , n5518 );
or ( n10289 , n10287 , n10288 );
nand ( n10290 , n5521 , n5344 );
nand ( n10291 , n10289 , n10290 );
and ( n10292 , n10285 , n10291 );
not ( n10293 , n10285 );
not ( n10294 , n10291 );
and ( n10295 , n10293 , n10294 );
nor ( n10296 , n10292 , n10295 );
not ( n10297 , n10296 );
not ( n10298 , n10297 );
or ( n10299 , n10268 , n10298 );
nand ( n10300 , n10296 , n10266 );
nand ( n10301 , n10299 , n10300 );
xor ( n10302 , n10262 , n10301 );
not ( n10303 , n5542 );
buf ( n10304 , n5530 );
or ( n10305 , n10303 , n10304 );
not ( n10306 , n10304 );
not ( n10307 , n10303 );
or ( n10308 , n10306 , n10307 );
nand ( n10309 , n10308 , n5537 );
nand ( n10310 , n10305 , n10309 );
xnor ( n10311 , n10302 , n10310 );
not ( n10312 , n5513 );
not ( n10313 , n5543 );
or ( n10314 , n10312 , n10313 );
not ( n10315 , n5512 );
not ( n10316 , n5544 );
or ( n10317 , n10315 , n10316 );
nand ( n10318 , n10317 , n5465 );
nand ( n10319 , n10314 , n10318 );
nor ( n10320 , n10311 , n10319 );
not ( n10321 , n10320 );
not ( n10322 , n10321 );
not ( n10323 , n4354 );
and ( n10324 , n5569 , n5439 , n4947 , n4486 );
not ( n10325 , n10324 );
or ( n10326 , n10323 , n10325 );
and ( n10327 , n5569 , n5439 );
not ( n10328 , n5448 );
and ( n10329 , n10327 , n10328 );
not ( n10330 , n5452 );
not ( n10331 , n5569 );
or ( n10332 , n10330 , n10331 );
nand ( n10333 , n10332 , n5567 );
nor ( n10334 , n10329 , n10333 );
nand ( n10335 , n10326 , n10334 );
not ( n10336 , n10335 );
or ( n10337 , n10322 , n10336 );
nand ( n10338 , n10319 , n10311 );
buf ( n10339 , n10338 );
nand ( n10340 , n10337 , n10339 );
not ( n10341 , n10261 );
or ( n10342 , n10241 , n10237 );
not ( n10343 , n10342 );
or ( n10344 , n10341 , n10343 );
nand ( n10345 , n10241 , n10237 );
nand ( n10346 , n10344 , n10345 );
not ( n10347 , n10269 );
not ( n10348 , n10347 );
not ( n10349 , n10283 );
or ( n10350 , n10348 , n10349 );
not ( n10351 , n10269 );
not ( n10352 , n10282 );
or ( n10353 , n10351 , n10352 );
nand ( n10354 , n10353 , n10275 );
nand ( n10355 , n10350 , n10354 );
not ( n10356 , n10355 );
not ( n10357 , n10356 );
not ( n10358 , n2086 );
not ( n10359 , n10358 );
not ( n10360 , n2082 );
or ( n10361 , n10359 , n10360 );
nand ( n10362 , n10361 , n497 );
not ( n10363 , n10280 );
not ( n10364 , n5389 );
or ( n10365 , n10363 , n10364 );
xor ( n10366 , n505 , n495 );
nand ( n10367 , n5392 , n10366 );
nand ( n10368 , n10365 , n10367 );
xor ( n10369 , n10362 , n10368 );
not ( n10370 , n10258 );
not ( n10371 , n5487 );
or ( n10372 , n10370 , n10371 );
xor ( n10373 , n491 , n509 );
nand ( n10374 , n2764 , n10373 );
nand ( n10375 , n10372 , n10374 );
xnor ( n10376 , n10369 , n10375 );
not ( n10377 , n10376 );
not ( n10378 , n10377 );
or ( n10379 , n10357 , n10378 );
nand ( n10380 , n10376 , n10355 );
nand ( n10381 , n10379 , n10380 );
not ( n10382 , n10248 );
not ( n10383 , n10260 );
or ( n10384 , n10382 , n10383 );
or ( n10385 , n10260 , n10248 );
nand ( n10386 , n10385 , n10253 );
nand ( n10387 , n10384 , n10386 );
xor ( n10388 , n10283 , n10387 );
and ( n10389 , n513 , n489 );
not ( n10390 , n10273 );
not ( n10391 , n2028 );
or ( n10392 , n10390 , n10391 );
xor ( n10393 , n507 , n493 );
nand ( n10394 , n2031 , n10393 );
nand ( n10395 , n10392 , n10394 );
not ( n10396 , n10395 );
and ( n10397 , n10389 , n10396 );
not ( n10398 , n10389 );
and ( n10399 , n10398 , n10395 );
or ( n10400 , n10397 , n10399 );
not ( n10401 , n10246 );
not ( n10402 , n4835 );
or ( n10403 , n10401 , n10402 );
xor ( n10404 , n511 , n489 );
nand ( n10405 , n4838 , n10404 );
nand ( n10406 , n10403 , n10405 );
xor ( n10407 , n10400 , n10406 );
xnor ( n10408 , n10388 , n10407 );
xor ( n10409 , n10381 , n10408 );
xor ( n10410 , n10346 , n10409 );
nand ( n10411 , n10285 , n10294 );
not ( n10412 , n10411 );
not ( n10413 , n10266 );
or ( n10414 , n10412 , n10413 );
nand ( n10415 , n10284 , n10291 );
nand ( n10416 , n10414 , n10415 );
xor ( n10417 , n10410 , n10416 );
not ( n10418 , n10301 );
buf ( n10419 , n10262 );
nand ( n10420 , n10418 , n10419 );
not ( n10421 , n10420 );
not ( n10422 , n10310 );
or ( n10423 , n10421 , n10422 );
not ( n10424 , n10419 );
nand ( n10425 , n10424 , n10301 );
nand ( n10426 , n10423 , n10425 );
nor ( n10427 , n10417 , n10426 );
not ( n10428 , n10427 );
nand ( n10429 , n10426 , n10417 );
nand ( n10430 , n10428 , n10429 );
not ( n10431 , n10430 );
and ( n10432 , n10340 , n10431 );
not ( n10433 , n10340 );
and ( n10434 , n10433 , n10430 );
nor ( n10435 , n10432 , n10434 );
nand ( n10436 , n10435 , n455 );
nand ( n10437 , n10233 , n10436 );
buf ( n10438 , n10437 );
not ( n10439 , n10438 );
not ( n10440 , n10439 );
or ( n10441 , n10030 , n10440 );
nand ( n10442 , n4018 , n10438 );
nand ( n10443 , n10441 , n10442 );
not ( n10444 , n10443 );
or ( n10445 , n10029 , n10444 );
not ( n10446 , n551 );
not ( n10447 , n716 );
not ( n10448 , n10208 );
and ( n10449 , n4031 , n5213 );
not ( n10450 , n10449 );
or ( n10451 , n10448 , n10450 );
not ( n10452 , n5081 );
not ( n10453 , n4963 );
or ( n10454 , n10452 , n10453 );
nand ( n10455 , n10454 , n5083 );
nor ( n10456 , n5318 , n5207 );
and ( n10457 , n10455 , n10456 );
nor ( n10458 , n10457 , n10218 );
nand ( n10459 , n10451 , n10458 );
nand ( n10460 , n10222 , n10202 );
xnor ( n10461 , n10459 , n10460 );
not ( n10462 , n10461 );
or ( n10463 , n10447 , n10462 );
nand ( n10464 , n10321 , n10338 );
not ( n10465 , n10464 );
not ( n10466 , n10335 );
or ( n10467 , n10465 , n10466 );
or ( n10468 , n10335 , n10464 );
nand ( n10469 , n10467 , n10468 );
nand ( n10470 , n10469 , n455 );
nand ( n10471 , n10463 , n10470 );
buf ( n10472 , n10471 );
not ( n10473 , n10472 );
not ( n10474 , n10473 );
or ( n10475 , n10446 , n10474 );
nand ( n10476 , n10472 , n4018 );
nand ( n10477 , n10475 , n10476 );
nand ( n10478 , n10477 , n5619 );
nand ( n10479 , n10445 , n10478 );
not ( n10480 , n3134 );
not ( n10481 , n537 );
not ( n10482 , n3280 );
or ( n10483 , n10481 , n10482 );
nand ( n10484 , n3279 , n3177 );
nand ( n10485 , n10483 , n10484 );
not ( n10486 , n10485 );
or ( n10487 , n10480 , n10486 );
nand ( n10488 , n5683 , n3182 );
nand ( n10489 , n10487 , n10488 );
and ( n10490 , n537 , n3096 );
xor ( n10491 , n10489 , n10490 );
not ( n10492 , n3026 );
and ( n10493 , n3980 , n3069 );
not ( n10494 , n3980 );
and ( n10495 , n10494 , n539 );
or ( n10496 , n10493 , n10495 );
not ( n10497 , n10496 );
or ( n10498 , n10492 , n10497 );
not ( n10499 , n5698 );
or ( n10500 , n10499 , n3102 );
nand ( n10501 , n10498 , n10500 );
xor ( n10502 , n10491 , n10501 );
not ( n10503 , n5636 );
not ( n10504 , n2376 );
or ( n10505 , n10503 , n10504 );
not ( n10506 , n545 );
not ( n10507 , n4653 );
or ( n10508 , n10506 , n10507 );
nand ( n10509 , n4652 , n706 );
nand ( n10510 , n10508 , n10509 );
not ( n10511 , n10510 );
not ( n10512 , n3017 );
or ( n10513 , n10511 , n10512 );
nand ( n10514 , n10505 , n10513 );
xor ( n10515 , n10502 , n10514 );
not ( n10516 , n3298 );
not ( n10517 , n547 );
not ( n10518 , n4635 );
or ( n10519 , n10517 , n10518 );
nand ( n10520 , n4638 , n2369 );
nand ( n10521 , n10519 , n10520 );
not ( n10522 , n10521 );
or ( n10523 , n10516 , n10522 );
nand ( n10524 , n5658 , n3300 );
nand ( n10525 , n10523 , n10524 );
and ( n10526 , n10515 , n10525 );
and ( n10527 , n10502 , n10514 );
or ( n10528 , n10526 , n10527 );
xor ( n10529 , n10479 , n10528 );
xor ( n10530 , n5666 , n5676 );
and ( n10531 , n10530 , n5703 );
and ( n10532 , n5666 , n5676 );
or ( n10533 , n10531 , n10532 );
not ( n10534 , n3288 );
not ( n10535 , n5672 );
or ( n10536 , n10534 , n10535 );
not ( n10537 , n541 );
not ( n10538 , n5906 );
or ( n10539 , n10537 , n10538 );
not ( n10540 , n6369 );
nand ( n10541 , n10540 , n3023 );
nand ( n10542 , n10539 , n10541 );
nand ( n10543 , n10542 , n3955 );
nand ( n10544 , n10536 , n10543 );
xor ( n10545 , n5688 , n5689 );
and ( n10546 , n10545 , n5702 );
and ( n10547 , n5688 , n5689 );
or ( n10548 , n10546 , n10547 );
xor ( n10549 , n10544 , n10548 );
not ( n10550 , n714 );
not ( n10551 , n5626 );
or ( n10552 , n10550 , n10551 );
not ( n10553 , n543 );
not ( n10554 , n4792 );
not ( n10555 , n10554 );
or ( n10556 , n10553 , n10555 );
nand ( n10557 , n4792 , n2123 );
nand ( n10558 , n10556 , n10557 );
nand ( n10559 , n2362 , n10558 );
nand ( n10560 , n10552 , n10559 );
xor ( n10561 , n10549 , n10560 );
xor ( n10562 , n10533 , n10561 );
not ( n10563 , n4022 );
not ( n10564 , n5098 );
or ( n10565 , n10563 , n10564 );
not ( n10566 , n549 );
not ( n10567 , n5607 );
or ( n10568 , n10566 , n10567 );
nand ( n10569 , n5614 , n4013 );
nand ( n10570 , n10568 , n10569 );
nand ( n10571 , n10570 , n6220 );
nand ( n10572 , n10565 , n10571 );
and ( n10573 , n10562 , n10572 );
and ( n10574 , n10533 , n10561 );
or ( n10575 , n10573 , n10574 );
xor ( n10576 , n10529 , n10575 );
xor ( n10577 , n10502 , n10514 );
xor ( n10578 , n10577 , n10525 );
xor ( n10579 , n10533 , n10561 );
xor ( n10580 , n10579 , n10572 );
xor ( n10581 , n10578 , n10580 );
xor ( n10582 , n5102 , n5621 );
and ( n10583 , n10582 , n5646 );
and ( n10584 , n5102 , n5621 );
or ( n10585 , n10583 , n10584 );
and ( n10586 , n10581 , n10585 );
and ( n10587 , n10578 , n10580 );
or ( n10588 , n10586 , n10587 );
xor ( n10589 , n10576 , n10588 );
not ( n10590 , n10485 );
not ( n10591 , n3182 );
or ( n10592 , n10590 , n10591 );
and ( n10593 , n3249 , n3177 );
not ( n10594 , n3249 );
and ( n10595 , n10594 , n537 );
or ( n10596 , n10593 , n10595 );
not ( n10597 , n10596 );
not ( n10598 , n3134 );
or ( n10599 , n10597 , n10598 );
nand ( n10600 , n10592 , n10599 );
not ( n10601 , n10496 );
not ( n10602 , n3103 );
or ( n10603 , n10601 , n10602 );
not ( n10604 , n5737 );
not ( n10605 , n539 );
and ( n10606 , n10604 , n10605 );
and ( n10607 , n6212 , n539 );
nor ( n10608 , n10606 , n10607 );
not ( n10609 , n3026 );
or ( n10610 , n10608 , n10609 );
nand ( n10611 , n10603 , n10610 );
xor ( n10612 , n10600 , n10611 );
nor ( n10613 , n3064 , n3177 );
xor ( n10614 , n10612 , n10613 );
not ( n10615 , n5799 );
and ( n10616 , n545 , n10615 );
not ( n10617 , n545 );
and ( n10618 , n10617 , n4342 );
nor ( n10619 , n10616 , n10618 );
or ( n10620 , n10512 , n10619 );
nand ( n10621 , n10510 , n2376 );
nand ( n10622 , n10620 , n10621 );
xor ( n10623 , n10614 , n10622 );
xor ( n10624 , n10544 , n10548 );
and ( n10625 , n10624 , n10560 );
and ( n10626 , n10544 , n10548 );
or ( n10627 , n10625 , n10626 );
xor ( n10628 , n10623 , n10627 );
not ( n10629 , n3298 );
not ( n10630 , n547 );
not ( n10631 , n5093 );
not ( n10632 , n10631 );
or ( n10633 , n10630 , n10632 );
nand ( n10634 , n5093 , n2369 );
nand ( n10635 , n10633 , n10634 );
not ( n10636 , n10635 );
or ( n10637 , n10629 , n10636 );
nand ( n10638 , n10521 , n3300 );
nand ( n10639 , n10637 , n10638 );
xor ( n10640 , n10489 , n10490 );
and ( n10641 , n10640 , n10501 );
and ( n10642 , n10489 , n10490 );
or ( n10643 , n10641 , n10642 );
not ( n10644 , n10542 );
not ( n10645 , n3288 );
or ( n10646 , n10644 , n10645 );
and ( n10647 , n541 , n2701 );
not ( n10648 , n541 );
not ( n10649 , n2697 );
not ( n10650 , n10649 );
and ( n10651 , n10648 , n10650 );
nor ( n10652 , n10647 , n10651 );
not ( n10653 , n10652 );
nand ( n10654 , n10653 , n3955 );
nand ( n10655 , n10646 , n10654 );
xor ( n10656 , n10643 , n10655 );
not ( n10657 , n2362 );
not ( n10658 , n543 );
not ( n10659 , n3632 );
or ( n10660 , n10658 , n10659 );
not ( n10661 , n6156 );
nand ( n10662 , n10661 , n2123 );
nand ( n10663 , n10660 , n10662 );
not ( n10664 , n10663 );
or ( n10665 , n10657 , n10664 );
nand ( n10666 , n10558 , n714 );
nand ( n10667 , n10665 , n10666 );
xor ( n10668 , n10656 , n10667 );
xor ( n10669 , n10639 , n10668 );
not ( n10670 , n6220 );
not ( n10671 , n549 );
not ( n10672 , n5582 );
not ( n10673 , n10672 );
or ( n10674 , n10671 , n10673 );
nand ( n10675 , n5582 , n4013 );
nand ( n10676 , n10674 , n10675 );
not ( n10677 , n10676 );
or ( n10678 , n10670 , n10677 );
nand ( n10679 , n10570 , n4022 );
nand ( n10680 , n10678 , n10679 );
xor ( n10681 , n10669 , n10680 );
xor ( n10682 , n10628 , n10681 );
xor ( n10683 , n5630 , n5640 );
and ( n10684 , n10683 , n5645 );
and ( n10685 , n5630 , n5640 );
or ( n10686 , n10684 , n10685 );
not ( n10687 , n5619 );
not ( n10688 , n5584 );
or ( n10689 , n10687 , n10688 );
nand ( n10690 , n552 , n10477 );
nand ( n10691 , n10689 , n10690 );
xor ( n10692 , n10686 , n10691 );
xor ( n10693 , n5662 , n5704 );
and ( n10694 , n10693 , n5709 );
and ( n10695 , n5662 , n5704 );
or ( n10696 , n10694 , n10695 );
and ( n10697 , n10692 , n10696 );
and ( n10698 , n10686 , n10691 );
or ( n10699 , n10697 , n10698 );
xor ( n10700 , n10682 , n10699 );
xor ( n10701 , n10589 , n10700 );
not ( n10702 , n10701 );
xor ( n10703 , n10686 , n10691 );
xor ( n10704 , n10703 , n10696 );
xor ( n10705 , n5652 , n5710 );
and ( n10706 , n10705 , n5765 );
and ( n10707 , n5652 , n5710 );
or ( n10708 , n10706 , n10707 );
xor ( n10709 , n10704 , n10708 );
xor ( n10710 , n10578 , n10580 );
xor ( n10711 , n10710 , n10585 );
and ( n10712 , n10709 , n10711 );
and ( n10713 , n10704 , n10708 );
or ( n10714 , n10712 , n10713 );
not ( n10715 , n10714 );
and ( n10716 , n10702 , n10715 );
xor ( n10717 , n10704 , n10708 );
xor ( n10718 , n10717 , n10711 );
not ( n10719 , n10718 );
xor ( n10720 , n4805 , n5647 );
and ( n10721 , n10720 , n5766 );
and ( n10722 , n4805 , n5647 );
or ( n10723 , n10721 , n10722 );
not ( n10724 , n10723 );
and ( n10725 , n10719 , n10724 );
nor ( n10726 , n10716 , n10725 );
not ( n10727 , n10726 );
nand ( n10728 , n6702 , n6042 , n6136 );
nand ( n10729 , n10728 , n5819 , n5964 );
not ( n10730 , n6706 );
nand ( n10731 , n5819 , n10730 );
nand ( n10732 , n10729 , n10731 , n5820 );
not ( n10733 , n10732 );
or ( n10734 , n10727 , n10733 );
nor ( n10735 , n10701 , n10714 );
not ( n10736 , n10735 );
and ( n10737 , n10718 , n10723 );
and ( n10738 , n10736 , n10737 );
and ( n10739 , n10701 , n10714 );
nor ( n10740 , n10738 , n10739 );
nand ( n10741 , n10734 , n10740 );
not ( n10742 , n5619 );
not ( n10743 , n10443 );
or ( n10744 , n10742 , n10743 );
not ( n10745 , n10174 );
not ( n10746 , n10187 );
and ( n10747 , n10745 , n10746 );
not ( n10748 , n10195 );
not ( n10749 , n10200 );
and ( n10750 , n10748 , n10749 );
nor ( n10751 , n10747 , n10750 );
buf ( n10752 , n10751 );
not ( n10753 , n10752 );
nand ( n10754 , n10195 , n10200 );
not ( n10755 , n10754 );
not ( n10756 , n10755 );
not ( n10757 , n10189 );
or ( n10758 , n10756 , n10757 );
nand ( n10759 , n10758 , n10192 );
not ( n10760 , n10759 );
buf ( n10761 , n10760 );
nand ( n10762 , n10753 , n10761 );
not ( n10763 , n10762 );
xor ( n10764 , n10073 , n10158 );
and ( n10765 , n10764 , n10173 );
and ( n10766 , n10073 , n10158 );
or ( n10767 , n10765 , n10766 );
not ( n10768 , n10767 );
xor ( n10769 , n10120 , n10129 );
and ( n10770 , n10769 , n10156 );
and ( n10771 , n10120 , n10129 );
or ( n10772 , n10770 , n10771 );
xor ( n10773 , n10075 , n10090 );
and ( n10774 , n10773 , n10101 );
and ( n10775 , n10075 , n10090 );
or ( n10776 , n10774 , n10775 );
not ( n10777 , n4553 );
not ( n10778 , n10137 );
or ( n10779 , n10777 , n10778 );
not ( n10780 , n489 );
not ( n10781 , n2949 );
or ( n10782 , n10780 , n10781 );
not ( n10783 , n489 );
nand ( n10784 , n10783 , n2948 );
nand ( n10785 , n10782 , n10784 );
nand ( n10786 , n10785 , n4547 );
nand ( n10787 , n10779 , n10786 );
not ( n10788 , n489 );
nor ( n10789 , n10788 , n10057 );
xor ( n10790 , n10787 , n10789 );
not ( n10791 , n1086 );
not ( n10792 , n10081 );
or ( n10793 , n10791 , n10792 );
nand ( n10794 , n1026 , n495 );
nand ( n10795 , n10793 , n10794 );
xor ( n10796 , n10790 , n10795 );
xor ( n10797 , n10776 , n10796 );
not ( n10798 , n3573 );
not ( n10799 , n10097 );
or ( n10800 , n10798 , n10799 );
not ( n10801 , n491 );
not ( n10802 , n2178 );
or ( n10803 , n10801 , n10802 );
nand ( n10804 , n2613 , n10108 );
nand ( n10805 , n10803 , n10804 );
nand ( n10806 , n10805 , n2606 );
nand ( n10807 , n10800 , n10806 );
not ( n10808 , n2966 );
not ( n10809 , n10150 );
or ( n10810 , n10808 , n10809 );
not ( n10811 , n493 );
not ( n10812 , n3859 );
or ( n10813 , n10811 , n10812 );
nand ( n10814 , n3858 , n739 );
nand ( n10815 , n10813 , n10814 );
nand ( n10816 , n10815 , n2959 );
nand ( n10817 , n10810 , n10816 );
not ( n10818 , n10817 );
xor ( n10819 , n10807 , n10818 );
xor ( n10820 , n10141 , n10152 );
and ( n10821 , n10820 , n10155 );
and ( n10822 , n10141 , n10152 );
or ( n10823 , n10821 , n10822 );
xor ( n10824 , n10819 , n10823 );
xor ( n10825 , n10797 , n10824 );
xor ( n10826 , n10772 , n10825 );
xor ( n10827 , n10102 , n10124 );
and ( n10828 , n10827 , n10157 );
and ( n10829 , n10102 , n10124 );
or ( n10830 , n10828 , n10829 );
xor ( n10831 , n10826 , n10830 );
not ( n10832 , n10831 );
nand ( n10833 , n10768 , n10832 );
nand ( n10834 , n10767 , n10831 );
buf ( n10835 , n10834 );
nand ( n10836 , n10833 , n10835 );
and ( n10837 , n10836 , n5320 );
not ( n10838 , n10837 );
and ( n10839 , n10763 , n10838 );
not ( n10840 , n10220 );
not ( n10841 , n10761 );
nor ( n10842 , n10841 , n10837 );
and ( n10843 , n10840 , n10842 );
nor ( n10844 , n10839 , n10843 );
not ( n10845 , n10844 );
not ( n10846 , n10761 );
not ( n10847 , n10840 );
or ( n10848 , n10846 , n10847 );
not ( n10849 , n10762 );
not ( n10850 , n10836 );
and ( n10851 , n10850 , n5320 );
nor ( n10852 , n10849 , n10851 );
nand ( n10853 , n10848 , n10852 );
not ( n10854 , n10853 );
or ( n10855 , n10845 , n10854 );
not ( n10856 , n10417 );
not ( n10857 , n10426 );
and ( n10858 , n10856 , n10857 );
nor ( n10859 , n10858 , n10320 );
not ( n10860 , n10859 );
not ( n10861 , n10335 );
or ( n10862 , n10860 , n10861 );
or ( n10863 , n10338 , n10427 );
nand ( n10864 , n10863 , n10429 );
not ( n10865 , n10864 );
nand ( n10866 , n10862 , n10865 );
xor ( n10867 , n10346 , n10409 );
and ( n10868 , n10867 , n10416 );
and ( n10869 , n10346 , n10409 );
or ( n10870 , n10868 , n10869 );
not ( n10871 , n10870 );
not ( n10872 , n10283 );
not ( n10873 , n10407 );
not ( n10874 , n10873 );
or ( n10875 , n10872 , n10874 );
nand ( n10876 , n10875 , n10387 );
nand ( n10877 , n10407 , n10282 );
nand ( n10878 , n10876 , n10877 );
not ( n10879 , n10878 );
and ( n10880 , n512 , n489 );
not ( n10881 , n10366 );
not ( n10882 , n5389 );
or ( n10883 , n10881 , n10882 );
nand ( n10884 , n5392 , n495 );
nand ( n10885 , n10883 , n10884 );
xor ( n10886 , n10880 , n10885 );
not ( n10887 , n10404 );
not ( n10888 , n4835 );
or ( n10889 , n10887 , n10888 );
xor ( n10890 , n489 , n510 );
nand ( n10891 , n4838 , n10890 );
nand ( n10892 , n10889 , n10891 );
xor ( n10893 , n10886 , n10892 );
not ( n10894 , n10368 );
not ( n10895 , n10375 );
or ( n10896 , n10894 , n10895 );
or ( n10897 , n10375 , n10368 );
nand ( n10898 , n10897 , n10362 );
nand ( n10899 , n10896 , n10898 );
xor ( n10900 , n10893 , n10899 );
not ( n10901 , n10389 );
nand ( n10902 , n10901 , n10396 );
not ( n10903 , n10902 );
not ( n10904 , n10406 );
or ( n10905 , n10903 , n10904 );
not ( n10906 , n10396 );
nand ( n10907 , n10906 , n10389 );
nand ( n10908 , n10905 , n10907 );
not ( n10909 , n10908 );
not ( n10910 , n10393 );
not ( n10911 , n2028 );
or ( n10912 , n10910 , n10911 );
xor ( n10913 , n493 , n506 );
nand ( n10914 , n2031 , n10913 );
nand ( n10915 , n10912 , n10914 );
not ( n10916 , n10373 );
not ( n10917 , n5487 );
or ( n10918 , n10916 , n10917 );
xor ( n10919 , n491 , n508 );
nand ( n10920 , n2764 , n10919 );
nand ( n10921 , n10918 , n10920 );
xor ( n10922 , n10915 , n10921 );
not ( n10923 , n10922 );
or ( n10924 , n10909 , n10923 );
or ( n10925 , n10908 , n10922 );
nand ( n10926 , n10924 , n10925 );
xor ( n10927 , n10900 , n10926 );
xor ( n10928 , n10879 , n10927 );
nand ( n10929 , n10376 , n10356 );
not ( n10930 , n10929 );
not ( n10931 , n10408 );
or ( n10932 , n10930 , n10931 );
nand ( n10933 , n10377 , n10355 );
nand ( n10934 , n10932 , n10933 );
xor ( n10935 , n10928 , n10934 );
nor ( n10936 , n10871 , n10935 );
not ( n10937 , n10936 );
not ( n10938 , n10870 );
nand ( n10939 , n10938 , n10935 );
nand ( n10940 , n10937 , n10939 );
nor ( n10941 , n10940 , n5320 );
and ( n10942 , n10866 , n10941 );
not ( n10943 , n10866 );
not ( n10944 , n10940 );
nor ( n10945 , n10944 , n5320 );
and ( n10946 , n10943 , n10945 );
nor ( n10947 , n10942 , n10946 );
nand ( n10948 , n10855 , n10947 );
not ( n10949 , n10948 );
and ( n10950 , n10949 , n4018 );
not ( n10951 , n10949 );
and ( n10952 , n10951 , n551 );
or ( n10953 , n10950 , n10952 );
nand ( n10954 , n10953 , n552 );
nand ( n10955 , n10744 , n10954 );
xor ( n10956 , n10614 , n10622 );
and ( n10957 , n10956 , n10627 );
and ( n10958 , n10614 , n10622 );
or ( n10959 , n10957 , n10958 );
xor ( n10960 , n10955 , n10959 );
not ( n10961 , n3182 );
not ( n10962 , n10596 );
or ( n10963 , n10961 , n10962 );
and ( n10964 , n6301 , n537 );
not ( n10965 , n6301 );
and ( n10966 , n10965 , n3177 );
or ( n10967 , n10964 , n10966 );
nand ( n10968 , n10967 , n3134 );
nand ( n10969 , n10963 , n10968 );
nand ( n10970 , n3279 , n537 );
xor ( n10971 , n10969 , n10970 );
not ( n10972 , n10971 );
not ( n10973 , n3103 );
not ( n10974 , n10608 );
not ( n10975 , n10974 );
or ( n10976 , n10973 , n10975 );
nand ( n10977 , n5906 , n539 );
not ( n10978 , n10977 );
nand ( n10979 , n10540 , n3069 );
not ( n10980 , n10979 );
or ( n10981 , n10978 , n10980 );
nand ( n10982 , n10981 , n3026 );
nand ( n10983 , n10976 , n10982 );
not ( n10984 , n10983 );
or ( n10985 , n10972 , n10984 );
or ( n10986 , n10983 , n10971 );
nand ( n10987 , n10985 , n10986 );
not ( n10988 , n2376 );
not ( n10989 , n10619 );
not ( n10990 , n10989 );
or ( n10991 , n10988 , n10990 );
not ( n10992 , n706 );
not ( n10993 , n4638 );
or ( n10994 , n10992 , n10993 );
not ( n10995 , n4638 );
nand ( n10996 , n10995 , n545 );
nand ( n10997 , n10994 , n10996 );
nand ( n10998 , n10997 , n3017 );
nand ( n10999 , n10991 , n10998 );
xor ( n11000 , n10987 , n10999 );
not ( n11001 , n3300 );
not ( n11002 , n10635 );
or ( n11003 , n11001 , n11002 );
and ( n11004 , n2369 , n5607 );
not ( n11005 , n2369 );
and ( n11006 , n11005 , n5614 );
nor ( n11007 , n11004 , n11006 );
nand ( n11008 , n11007 , n3298 );
nand ( n11009 , n11003 , n11008 );
xor ( n11010 , n11000 , n11009 );
xor ( n11011 , n10960 , n11010 );
xor ( n11012 , n10628 , n10681 );
and ( n11013 , n11012 , n10699 );
and ( n11014 , n10628 , n10681 );
or ( n11015 , n11013 , n11014 );
xor ( n11016 , n11011 , n11015 );
xor ( n11017 , n10639 , n10668 );
and ( n11018 , n11017 , n10680 );
and ( n11019 , n10639 , n10668 );
or ( n11020 , n11018 , n11019 );
xor ( n11021 , n10643 , n10655 );
and ( n11022 , n11021 , n10667 );
and ( n11023 , n10643 , n10655 );
or ( n11024 , n11022 , n11023 );
not ( n11025 , n3288 );
or ( n11026 , n10652 , n11025 );
not ( n11027 , n3012 );
not ( n11028 , n541 );
and ( n11029 , n11027 , n11028 );
and ( n11030 , n10554 , n541 );
nor ( n11031 , n11029 , n11030 );
not ( n11032 , n3955 );
or ( n11033 , n11031 , n11032 );
nand ( n11034 , n11026 , n11033 );
xor ( n11035 , n10600 , n10611 );
and ( n11036 , n11035 , n10613 );
and ( n11037 , n10600 , n10611 );
or ( n11038 , n11036 , n11037 );
xor ( n11039 , n11034 , n11038 );
not ( n11040 , n714 );
not ( n11041 , n10663 );
or ( n11042 , n11040 , n11041 );
not ( n11043 , n543 );
not ( n11044 , n4653 );
or ( n11045 , n11043 , n11044 );
nand ( n11046 , n4652 , n2123 );
nand ( n11047 , n11045 , n11046 );
nand ( n11048 , n11047 , n2362 );
nand ( n11049 , n11042 , n11048 );
xor ( n11050 , n11039 , n11049 );
xor ( n11051 , n11024 , n11050 );
not ( n11052 , n4022 );
not ( n11053 , n10676 );
or ( n11054 , n11052 , n11053 );
not ( n11055 , n10471 );
and ( n11056 , n11055 , n549 );
not ( n11057 , n11055 );
and ( n11058 , n11057 , n4013 );
or ( n11059 , n11056 , n11058 );
nand ( n11060 , n11059 , n6220 );
nand ( n11061 , n11054 , n11060 );
xor ( n11062 , n11051 , n11061 );
xor ( n11063 , n11020 , n11062 );
xor ( n11064 , n10479 , n10528 );
and ( n11065 , n11064 , n10575 );
and ( n11066 , n10479 , n10528 );
or ( n11067 , n11065 , n11066 );
xor ( n11068 , n11063 , n11067 );
and ( n11069 , n11016 , n11068 );
and ( n11070 , n11011 , n11015 );
or ( n11071 , n11069 , n11070 );
not ( n11072 , n552 );
not ( n11073 , n716 );
xor ( n11074 , n10772 , n10825 );
and ( n11075 , n11074 , n10830 );
and ( n11076 , n10772 , n10825 );
or ( n11077 , n11075 , n11076 );
xor ( n11078 , n10807 , n10818 );
and ( n11079 , n11078 , n10823 );
and ( n11080 , n10807 , n10818 );
or ( n11081 , n11079 , n11080 );
xor ( n11082 , n10787 , n10789 );
and ( n11083 , n11082 , n10795 );
and ( n11084 , n10787 , n10789 );
or ( n11085 , n11083 , n11084 );
or ( n11086 , n1026 , n1086 );
nand ( n11087 , n11086 , n495 );
not ( n11088 , n2959 );
not ( n11089 , n493 );
not ( n11090 , n4077 );
or ( n11091 , n11089 , n11090 );
nand ( n11092 , n4076 , n739 );
nand ( n11093 , n11091 , n11092 );
not ( n11094 , n11093 );
or ( n11095 , n11088 , n11094 );
nand ( n11096 , n10815 , n2967 );
nand ( n11097 , n11095 , n11096 );
xor ( n11098 , n11087 , n11097 );
not ( n11099 , n4547 );
xor ( n11100 , n489 , n5278 );
not ( n11101 , n11100 );
or ( n11102 , n11099 , n11101 );
nand ( n11103 , n4553 , n10785 );
nand ( n11104 , n11102 , n11103 );
xor ( n11105 , n11098 , n11104 );
xor ( n11106 , n11085 , n11105 );
buf ( n11107 , n844 );
not ( n11108 , n11107 );
and ( n11109 , n11108 , n489 );
not ( n11110 , n3573 );
not ( n11111 , n10805 );
or ( n11112 , n11110 , n11111 );
not ( n11113 , n491 );
not ( n11114 , n4090 );
or ( n11115 , n11113 , n11114 );
nand ( n11116 , n4093 , n2613 );
nand ( n11117 , n11115 , n11116 );
nand ( n11118 , n11117 , n2606 );
nand ( n11119 , n11112 , n11118 );
xor ( n11120 , n11109 , n11119 );
xor ( n11121 , n11120 , n10817 );
xor ( n11122 , n11106 , n11121 );
xor ( n11123 , n11081 , n11122 );
xor ( n11124 , n10776 , n10796 );
and ( n11125 , n11124 , n10824 );
and ( n11126 , n10776 , n10796 );
or ( n11127 , n11125 , n11126 );
xor ( n11128 , n11123 , n11127 );
nand ( n11129 , n11077 , n11128 );
not ( n11130 , n11077 );
not ( n11131 , n11128 );
nand ( n11132 , n11130 , n11131 );
nand ( n11133 , n11129 , n11132 );
not ( n11134 , n10835 );
or ( n11135 , n11133 , n11134 );
and ( n11136 , n10752 , n10208 );
not ( n11137 , n11136 );
not ( n11138 , n5222 );
or ( n11139 , n11137 , n11138 );
not ( n11140 , n10752 );
not ( n11141 , n5326 );
not ( n11142 , n10215 );
or ( n11143 , n11141 , n11142 );
nand ( n11144 , n11143 , n5316 );
not ( n11145 , n11144 );
or ( n11146 , n11140 , n11145 );
nand ( n11147 , n11146 , n10760 );
not ( n11148 , n11147 );
nand ( n11149 , n11139 , n11148 );
or ( n11150 , n11135 , n11149 );
and ( n11151 , n11133 , n10833 );
nand ( n11152 , n11149 , n11151 );
and ( n11153 , n11133 , n11134 );
nor ( n11154 , n11133 , n10833 , n11134 );
nor ( n11155 , n11153 , n11154 );
nand ( n11156 , n11150 , n11152 , n11155 );
not ( n11157 , n11156 );
or ( n11158 , n11073 , n11157 );
buf ( n11159 , n10859 );
buf ( n11160 , n10939 );
and ( n11161 , n11159 , n11160 );
not ( n11162 , n11161 );
not ( n11163 , n10335 );
or ( n11164 , n11162 , n11163 );
and ( n11165 , n10939 , n10864 );
nor ( n11166 , n11165 , n10936 );
nand ( n11167 , n11164 , n11166 );
not ( n11168 , n10879 );
not ( n11169 , n10927 );
not ( n11170 , n11169 );
or ( n11171 , n11168 , n11170 );
nand ( n11172 , n11171 , n10934 );
not ( n11173 , n11169 );
nand ( n11174 , n11173 , n10878 );
nand ( n11175 , n11172 , n11174 );
not ( n11176 , n10921 );
nand ( n11177 , n11176 , n10915 );
not ( n11178 , n11177 );
not ( n11179 , n10908 );
or ( n11180 , n11178 , n11179 );
not ( n11181 , n10915 );
nand ( n11182 , n11181 , n10921 );
nand ( n11183 , n11180 , n11182 );
xor ( n11184 , n10893 , n10899 );
and ( n11185 , n11184 , n10926 );
and ( n11186 , n10893 , n10899 );
or ( n11187 , n11185 , n11186 );
xor ( n11188 , n11183 , n11187 );
and ( n11189 , n511 , n489 );
xor ( n11190 , n11189 , n10915 );
not ( n11191 , n10919 );
not ( n11192 , n5487 );
or ( n11193 , n11191 , n11192 );
xor ( n11194 , n507 , n491 );
nand ( n11195 , n2764 , n11194 );
nand ( n11196 , n11193 , n11195 );
xor ( n11197 , n11190 , n11196 );
buf ( n11198 , n11197 );
not ( n11199 , n11198 );
not ( n11200 , n10913 );
not ( n11201 , n2028 );
or ( n11202 , n11200 , n11201 );
xor ( n11203 , n505 , n493 );
nand ( n11204 , n2031 , n11203 );
nand ( n11205 , n11202 , n11204 );
not ( n11206 , n10890 );
not ( n11207 , n4835 );
or ( n11208 , n11206 , n11207 );
xor ( n11209 , n489 , n509 );
nand ( n11210 , n4838 , n11209 );
nand ( n11211 , n11208 , n11210 );
xor ( n11212 , n11205 , n11211 );
or ( n11213 , n5392 , n5389 );
nand ( n11214 , n11213 , n495 );
xor ( n11215 , n11212 , n11214 );
buf ( n11216 , n11215 );
not ( n11217 , n11216 );
xor ( n11218 , n10880 , n10885 );
and ( n11219 , n11218 , n10892 );
and ( n11220 , n10880 , n10885 );
or ( n11221 , n11219 , n11220 );
nand ( n11222 , n11199 , n11217 , n11221 );
not ( n11223 , n11221 );
nand ( n11224 , n11198 , n11217 , n11223 );
nand ( n11225 , n11199 , n11216 , n11223 );
nand ( n11226 , n11198 , n11216 , n11221 );
nand ( n11227 , n11222 , n11224 , n11225 , n11226 );
xor ( n11228 , n11188 , n11227 );
and ( n11229 , n11175 , n11228 );
not ( n11230 , n11229 );
nor ( n11231 , n11175 , n11228 );
not ( n11232 , n11231 );
nand ( n11233 , n11230 , n11232 );
not ( n11234 , n11233 );
and ( n11235 , n11167 , n11234 );
not ( n11236 , n11167 );
and ( n11237 , n11236 , n11233 );
nor ( n11238 , n11235 , n11237 );
nand ( n11239 , n11238 , n455 );
nand ( n11240 , n11158 , n11239 );
buf ( n11241 , n11240 );
and ( n11242 , n11241 , n4018 );
not ( n11243 , n11241 );
and ( n11244 , n11243 , n551 );
or ( n11245 , n11242 , n11244 );
not ( n11246 , n11245 );
or ( n11247 , n11072 , n11246 );
nand ( n11248 , n5619 , n10953 );
nand ( n11249 , n11247 , n11248 );
xor ( n11250 , n10987 , n10999 );
and ( n11251 , n11250 , n11009 );
and ( n11252 , n10987 , n10999 );
or ( n11253 , n11251 , n11252 );
xor ( n11254 , n11249 , n11253 );
xor ( n11255 , n11024 , n11050 );
and ( n11256 , n11255 , n11061 );
and ( n11257 , n11024 , n11050 );
or ( n11258 , n11256 , n11257 );
xor ( n11259 , n11254 , n11258 );
xor ( n11260 , n11020 , n11062 );
and ( n11261 , n11260 , n11067 );
and ( n11262 , n11020 , n11062 );
or ( n11263 , n11261 , n11262 );
xor ( n11264 , n11259 , n11263 );
nand ( n11265 , n3017 , n545 );
not ( n11266 , n11265 );
nand ( n11267 , n11266 , n5094 );
nand ( n11268 , n10997 , n2376 );
not ( n11269 , n10631 );
not ( n11270 , n3017 );
nor ( n11271 , n11270 , n545 );
nand ( n11272 , n11269 , n11271 );
nand ( n11273 , n11267 , n11268 , n11272 );
xor ( n11274 , n11034 , n11038 );
and ( n11275 , n11274 , n11049 );
and ( n11276 , n11034 , n11038 );
or ( n11277 , n11275 , n11276 );
xor ( n11278 , n11273 , n11277 );
not ( n11279 , n10969 );
nor ( n11280 , n11279 , n10970 );
not ( n11281 , n3103 );
nand ( n11282 , n10979 , n10977 );
not ( n11283 , n11282 );
or ( n11284 , n11281 , n11283 );
not ( n11285 , n539 );
not ( n11286 , n10649 );
or ( n11287 , n11285 , n11286 );
nand ( n11288 , n2697 , n3069 );
nand ( n11289 , n11287 , n11288 );
nand ( n11290 , n11289 , n3026 );
nand ( n11291 , n11284 , n11290 );
xor ( n11292 , n11280 , n11291 );
not ( n11293 , n537 );
nor ( n11294 , n11293 , n3250 );
not ( n11295 , n3186 );
or ( n11296 , n2122 , n3177 );
nand ( n11297 , n2122 , n3177 );
nand ( n11298 , n11296 , n11297 );
not ( n11299 , n11298 );
or ( n11300 , n11295 , n11299 );
nand ( n11301 , n10967 , n3182 );
nand ( n11302 , n11300 , n11301 );
xor ( n11303 , n11294 , n11302 );
xor ( n11304 , n11292 , n11303 );
xor ( n11305 , n11278 , n11304 );
not ( n11306 , n3298 );
and ( n11307 , n547 , n5579 );
not ( n11308 , n547 );
and ( n11309 , n11308 , n5578 );
or ( n11310 , n11307 , n11309 );
not ( n11311 , n11310 );
or ( n11312 , n11306 , n11311 );
nand ( n11313 , n11007 , n3300 );
nand ( n11314 , n11312 , n11313 );
not ( n11315 , n549 );
not ( n11316 , n10439 );
or ( n11317 , n11315 , n11316 );
nand ( n11318 , n10438 , n4013 );
nand ( n11319 , n11317 , n11318 );
not ( n11320 , n11319 );
not ( n11321 , n4020 );
or ( n11322 , n11320 , n11321 );
nand ( n11323 , n4022 , n11059 );
nand ( n11324 , n11322 , n11323 );
xor ( n11325 , n11314 , n11324 );
not ( n11326 , n3955 );
not ( n11327 , n541 );
not ( n11328 , n3632 );
or ( n11329 , n11327 , n11328 );
nand ( n11330 , n10661 , n3023 );
nand ( n11331 , n11329 , n11330 );
not ( n11332 , n11331 );
or ( n11333 , n11326 , n11332 );
not ( n11334 , n11031 );
nand ( n11335 , n11334 , n3288 );
nand ( n11336 , n11333 , n11335 );
not ( n11337 , n10983 );
nor ( n11338 , n11337 , n10971 );
xor ( n11339 , n11336 , n11338 );
not ( n11340 , n2362 );
not ( n11341 , n543 );
not ( n11342 , n10615 );
or ( n11343 , n11341 , n11342 );
nand ( n11344 , n4342 , n2123 );
nand ( n11345 , n11343 , n11344 );
not ( n11346 , n11345 );
or ( n11347 , n11340 , n11346 );
nand ( n11348 , n11047 , n714 );
nand ( n11349 , n11347 , n11348 );
xor ( n11350 , n11339 , n11349 );
xor ( n11351 , n11325 , n11350 );
xor ( n11352 , n11305 , n11351 );
xor ( n11353 , n10955 , n10959 );
and ( n11354 , n11353 , n11010 );
and ( n11355 , n10955 , n10959 );
or ( n11356 , n11354 , n11355 );
xor ( n11357 , n11352 , n11356 );
xor ( n11358 , n11264 , n11357 );
nor ( n11359 , n11071 , n11358 );
xor ( n11360 , n11011 , n11015 );
xor ( n11361 , n11360 , n11068 );
xor ( n11362 , n10576 , n10588 );
and ( n11363 , n11362 , n10700 );
and ( n11364 , n10576 , n10588 );
or ( n11365 , n11363 , n11364 );
nor ( n11366 , n11361 , n11365 );
nor ( n11367 , n11359 , n11366 );
not ( n11368 , n3955 );
not ( n11369 , n541 );
not ( n11370 , n3943 );
or ( n11371 , n11369 , n11370 );
nand ( n11372 , n4652 , n3023 );
nand ( n11373 , n11371 , n11372 );
not ( n11374 , n11373 );
or ( n11375 , n11368 , n11374 );
nand ( n11376 , n11331 , n3288 );
nand ( n11377 , n11375 , n11376 );
xor ( n11378 , n11280 , n11291 );
and ( n11379 , n11378 , n11303 );
and ( n11380 , n11280 , n11291 );
or ( n11381 , n11379 , n11380 );
xor ( n11382 , n11377 , n11381 );
not ( n11383 , n2362 );
not ( n11384 , n543 );
not ( n11385 , n4635 );
or ( n11386 , n11384 , n11385 );
not ( n11387 , n4635 );
nand ( n11388 , n11387 , n2123 );
nand ( n11389 , n11386 , n11388 );
not ( n11390 , n11389 );
or ( n11391 , n11383 , n11390 );
nand ( n11392 , n11345 , n714 );
nand ( n11393 , n11391 , n11392 );
xor ( n11394 , n11382 , n11393 );
xor ( n11395 , n11273 , n11277 );
and ( n11396 , n11395 , n11304 );
and ( n11397 , n11273 , n11277 );
or ( n11398 , n11396 , n11397 );
xor ( n11399 , n11394 , n11398 );
not ( n11400 , n2376 );
not ( n11401 , n545 );
not ( n11402 , n5754 );
or ( n11403 , n11401 , n11402 );
nand ( n11404 , n5093 , n706 );
nand ( n11405 , n11403 , n11404 );
not ( n11406 , n11405 );
or ( n11407 , n11400 , n11406 );
not ( n11408 , n545 );
not ( n11409 , n5607 );
or ( n11410 , n11408 , n11409 );
nand ( n11411 , n5614 , n706 );
nand ( n11412 , n11410 , n11411 );
nand ( n11413 , n11412 , n3017 );
nand ( n11414 , n11407 , n11413 );
not ( n11415 , n3011 );
nor ( n11416 , n10609 , n3069 );
nand ( n11417 , n11415 , n11416 );
nand ( n11418 , n2697 , n4699 );
nor ( n11419 , n10609 , n539 );
nand ( n11420 , n3011 , n11419 );
not ( n11421 , n2697 );
nand ( n11422 , n11421 , n4701 );
nand ( n11423 , n11417 , n11418 , n11420 , n11422 );
and ( n11424 , n11302 , n11294 );
xor ( n11425 , n11423 , n11424 );
nand ( n11426 , n3981 , n537 );
not ( n11427 , n11426 );
not ( n11428 , n537 );
not ( n11429 , n4732 );
or ( n11430 , n11428 , n11429 );
nand ( n11431 , n2355 , n3177 );
nand ( n11432 , n11430 , n11431 );
nand ( n11433 , n11432 , n3134 );
not ( n11434 , n11298 );
nor ( n11435 , n11434 , n3194 );
not ( n11436 , n11435 );
nand ( n11437 , n11433 , n11436 );
not ( n11438 , n11437 );
or ( n11439 , n11427 , n11438 );
nor ( n11440 , n11435 , n11426 );
nand ( n11441 , n11433 , n11440 );
nand ( n11442 , n11439 , n11441 );
xor ( n11443 , n11425 , n11442 );
xor ( n11444 , n11414 , n11443 );
not ( n11445 , n3298 );
not ( n11446 , n547 );
not ( n11447 , n10472 );
not ( n11448 , n11447 );
or ( n11449 , n11446 , n11448 );
nand ( n11450 , n10472 , n2369 );
nand ( n11451 , n11449 , n11450 );
not ( n11452 , n11451 );
or ( n11453 , n11445 , n11452 );
nand ( n11454 , n11310 , n3300 );
nand ( n11455 , n11453 , n11454 );
xor ( n11456 , n11444 , n11455 );
xor ( n11457 , n11399 , n11456 );
xor ( n11458 , n11305 , n11351 );
and ( n11459 , n11458 , n11356 );
and ( n11460 , n11305 , n11351 );
or ( n11461 , n11459 , n11460 );
xor ( n11462 , n11457 , n11461 );
xor ( n11463 , n11314 , n11324 );
and ( n11464 , n11463 , n11350 );
and ( n11465 , n11314 , n11324 );
or ( n11466 , n11464 , n11465 );
xor ( n11467 , n11336 , n11338 );
and ( n11468 , n11467 , n11349 );
and ( n11469 , n11336 , n11338 );
or ( n11470 , n11468 , n11469 );
not ( n11471 , n4022 );
not ( n11472 , n11319 );
or ( n11473 , n11471 , n11472 );
not ( n11474 , n549 );
not ( n11475 , n10949 );
not ( n11476 , n11475 );
or ( n11477 , n11474 , n11476 );
buf ( n11478 , n10949 );
nand ( n11479 , n11478 , n4013 );
nand ( n11480 , n11477 , n11479 );
nand ( n11481 , n11480 , n4020 );
nand ( n11482 , n11473 , n11481 );
xor ( n11483 , n11470 , n11482 );
not ( n11484 , n5619 );
not ( n11485 , n11245 );
or ( n11486 , n11484 , n11485 );
not ( n11487 , n551 );
not ( n11488 , n3229 );
xor ( n11489 , n11081 , n11122 );
and ( n11490 , n11489 , n11127 );
and ( n11491 , n11081 , n11122 );
or ( n11492 , n11490 , n11491 );
xor ( n11493 , n11109 , n11119 );
and ( n11494 , n11493 , n10817 );
and ( n11495 , n11109 , n11119 );
or ( n11496 , n11494 , n11495 );
and ( n11497 , n11093 , n2966 );
and ( n11498 , n758 , n493 );
nor ( n11499 , n11497 , n11498 );
xor ( n11500 , n11087 , n11097 );
and ( n11501 , n11500 , n11104 );
and ( n11502 , n11087 , n11097 );
or ( n11503 , n11501 , n11502 );
xor ( n11504 , n11499 , n11503 );
and ( n11505 , n2948 , n489 );
not ( n11506 , n3573 );
not ( n11507 , n11117 );
or ( n11508 , n11506 , n11507 );
not ( n11509 , n491 );
not ( n11510 , n3859 );
or ( n11511 , n11509 , n11510 );
nand ( n11512 , n3858 , n2613 );
nand ( n11513 , n11511 , n11512 );
nand ( n11514 , n11513 , n2606 );
nand ( n11515 , n11508 , n11514 );
xor ( n11516 , n11505 , n11515 );
not ( n11517 , n4547 );
xor ( n11518 , n489 , n10108 );
not ( n11519 , n11518 );
or ( n11520 , n11517 , n11519 );
nand ( n11521 , n11100 , n4056 );
nand ( n11522 , n11520 , n11521 );
xor ( n11523 , n11516 , n11522 );
xor ( n11524 , n11504 , n11523 );
xor ( n11525 , n11496 , n11524 );
xor ( n11526 , n11085 , n11105 );
and ( n11527 , n11526 , n11121 );
and ( n11528 , n11085 , n11105 );
or ( n11529 , n11527 , n11528 );
xor ( n11530 , n11525 , n11529 );
or ( n11531 , n11492 , n11530 );
nand ( n11532 , n11492 , n11530 );
nand ( n11533 , n11531 , n11532 );
not ( n11534 , n10752 );
nand ( n11535 , n11130 , n11131 );
nand ( n11536 , n10833 , n11535 );
nor ( n11537 , n11534 , n11536 );
not ( n11538 , n11537 );
not ( n11539 , n10459 );
or ( n11540 , n11538 , n11539 );
not ( n11541 , n10832 );
not ( n11542 , n10767 );
not ( n11543 , n11542 );
or ( n11544 , n11541 , n11543 );
nand ( n11545 , n11544 , n11535 );
not ( n11546 , n11545 );
and ( n11547 , n10759 , n11546 );
nand ( n11548 , n11130 , n11131 );
not ( n11549 , n11548 );
not ( n11550 , n10834 );
not ( n11551 , n11550 );
or ( n11552 , n11549 , n11551 );
nand ( n11553 , n11552 , n11129 );
nor ( n11554 , n11547 , n11553 );
buf ( n11555 , n11554 );
nand ( n11556 , n11540 , n11555 );
or ( n11557 , n11533 , n11556 );
nand ( n11558 , n11556 , n11533 );
nand ( n11559 , n11557 , n11558 );
not ( n11560 , n11559 );
or ( n11561 , n11488 , n11560 );
xor ( n11562 , n11183 , n11187 );
and ( n11563 , n11562 , n11227 );
and ( n11564 , n11183 , n11187 );
or ( n11565 , n11563 , n11564 );
not ( n11566 , n11198 );
not ( n11567 , n11221 );
or ( n11568 , n11566 , n11567 );
not ( n11569 , n11223 );
not ( n11570 , n11199 );
or ( n11571 , n11569 , n11570 );
nand ( n11572 , n11571 , n11216 );
nand ( n11573 , n11568 , n11572 );
xor ( n11574 , n11189 , n10915 );
and ( n11575 , n11574 , n11196 );
and ( n11576 , n11189 , n10915 );
or ( n11577 , n11575 , n11576 );
xor ( n11578 , n11573 , n11577 );
not ( n11579 , n11203 );
not ( n11580 , n2028 );
or ( n11581 , n11579 , n11580 );
not ( n11582 , n2473 );
nand ( n11583 , n11582 , n493 );
nand ( n11584 , n11581 , n11583 );
not ( n11585 , n11584 );
not ( n11586 , n11209 );
not ( n11587 , n4835 );
or ( n11588 , n11586 , n11587 );
xor ( n11589 , n489 , n508 );
nand ( n11590 , n4838 , n11589 );
nand ( n11591 , n11588 , n11590 );
nand ( n11592 , n489 , n510 );
xor ( n11593 , n11591 , n11592 );
not ( n11594 , n11194 );
not ( n11595 , n5487 );
or ( n11596 , n11594 , n11595 );
xor ( n11597 , n491 , n506 );
nand ( n11598 , n2764 , n11597 );
nand ( n11599 , n11596 , n11598 );
xnor ( n11600 , n11593 , n11599 );
xor ( n11601 , n11585 , n11600 );
xor ( n11602 , n11205 , n11211 );
and ( n11603 , n11602 , n11214 );
and ( n11604 , n11205 , n11211 );
or ( n11605 , n11603 , n11604 );
xor ( n11606 , n11601 , n11605 );
xor ( n11607 , n11578 , n11606 );
nor ( n11608 , n11565 , n11607 );
not ( n11609 , n11608 );
nand ( n11610 , n11565 , n11607 );
and ( n11611 , n11609 , n11610 );
not ( n11612 , n5449 );
nand ( n11613 , n10327 , n11159 , n11160 , n11232 );
not ( n11614 , n11613 );
not ( n11615 , n11614 );
or ( n11616 , n11612 , n11615 );
not ( n11617 , n10333 );
not ( n11618 , n10859 );
nand ( n11619 , n11232 , n10939 );
nor ( n11620 , n11618 , n11619 );
not ( n11621 , n11620 );
or ( n11622 , n11617 , n11621 );
not ( n11623 , n11619 );
not ( n11624 , n11623 );
not ( n11625 , n10864 );
or ( n11626 , n11624 , n11625 );
not ( n11627 , n11232 );
not ( n11628 , n10936 );
or ( n11629 , n11627 , n11628 );
not ( n11630 , n11229 );
nand ( n11631 , n11629 , n11630 );
not ( n11632 , n11631 );
nand ( n11633 , n11626 , n11632 );
not ( n11634 , n11633 );
nand ( n11635 , n11622 , n11634 );
not ( n11636 , n11635 );
nand ( n11637 , n11616 , n11636 );
xor ( n11638 , n11611 , n11637 );
nand ( n11639 , n11638 , n455 );
nand ( n11640 , n11561 , n11639 );
not ( n11641 , n11640 );
not ( n11642 , n11641 );
or ( n11643 , n11487 , n11642 );
not ( n11644 , n11641 );
nand ( n11645 , n11644 , n4018 );
nand ( n11646 , n11643 , n11645 );
nand ( n11647 , n11646 , n552 );
nand ( n11648 , n11486 , n11647 );
xor ( n11649 , n11483 , n11648 );
xor ( n11650 , n11466 , n11649 );
xor ( n11651 , n11249 , n11253 );
and ( n11652 , n11651 , n11258 );
and ( n11653 , n11249 , n11253 );
or ( n11654 , n11652 , n11653 );
xor ( n11655 , n11650 , n11654 );
xor ( n11656 , n11462 , n11655 );
not ( n11657 , n11656 );
xor ( n11658 , n11259 , n11263 );
and ( n11659 , n11658 , n11357 );
and ( n11660 , n11259 , n11263 );
or ( n11661 , n11659 , n11660 );
not ( n11662 , n11661 );
nand ( n11663 , n11657 , n11662 );
and ( n11664 , n11367 , n11663 );
xor ( n11665 , n11423 , n11424 );
and ( n11666 , n11665 , n11442 );
and ( n11667 , n11423 , n11424 );
or ( n11668 , n11666 , n11667 );
not ( n11669 , n3955 );
not ( n11670 , n541 );
not ( n11671 , n10615 );
or ( n11672 , n11670 , n11671 );
nand ( n11673 , n4342 , n3023 );
nand ( n11674 , n11672 , n11673 );
not ( n11675 , n11674 );
or ( n11676 , n11669 , n11675 );
nand ( n11677 , n11373 , n3288 );
nand ( n11678 , n11676 , n11677 );
xor ( n11679 , n11668 , n11678 );
not ( n11680 , n2362 );
and ( n11681 , n5093 , n2123 );
not ( n11682 , n5093 );
and ( n11683 , n11682 , n543 );
or ( n11684 , n11681 , n11683 );
not ( n11685 , n11684 );
or ( n11686 , n11680 , n11685 );
nand ( n11687 , n11389 , n714 );
nand ( n11688 , n11686 , n11687 );
xor ( n11689 , n11679 , n11688 );
xor ( n11690 , n11414 , n11443 );
and ( n11691 , n11690 , n11455 );
and ( n11692 , n11414 , n11443 );
or ( n11693 , n11691 , n11692 );
xor ( n11694 , n11689 , n11693 );
not ( n11695 , n3017 );
not ( n11696 , n545 );
not ( n11697 , n5579 );
or ( n11698 , n11696 , n11697 );
nand ( n11699 , n5578 , n706 );
nand ( n11700 , n11698 , n11699 );
not ( n11701 , n11700 );
or ( n11702 , n11695 , n11701 );
nand ( n11703 , n11412 , n2376 );
nand ( n11704 , n11702 , n11703 );
and ( n11705 , n11433 , n11436 );
nor ( n11706 , n11705 , n11426 );
not ( n11707 , n3026 );
and ( n11708 , n3630 , n539 );
not ( n11709 , n3630 );
and ( n11710 , n11709 , n3069 );
nor ( n11711 , n11708 , n11710 );
not ( n11712 , n11711 );
or ( n11713 , n11707 , n11712 );
and ( n11714 , n3012 , n4701 );
not ( n11715 , n3012 );
and ( n11716 , n11715 , n4699 );
nor ( n11717 , n11714 , n11716 );
nand ( n11718 , n11713 , n11717 );
xor ( n11719 , n11706 , n11718 );
not ( n11720 , n2125 );
nand ( n11721 , n11720 , n537 );
not ( n11722 , n11721 );
not ( n11723 , n3134 );
or ( n11724 , n2697 , n3177 );
nand ( n11725 , n2697 , n3177 );
nand ( n11726 , n11724 , n11725 );
not ( n11727 , n11726 );
or ( n11728 , n11723 , n11727 );
buf ( n11729 , n3182 );
nand ( n11730 , n11432 , n11729 );
nand ( n11731 , n11728 , n11730 );
not ( n11732 , n11731 );
or ( n11733 , n11722 , n11732 );
or ( n11734 , n11731 , n11721 );
nand ( n11735 , n11733 , n11734 );
xor ( n11736 , n11719 , n11735 );
xor ( n11737 , n11704 , n11736 );
not ( n11738 , n3300 );
not ( n11739 , n11451 );
or ( n11740 , n11738 , n11739 );
not ( n11741 , n10438 );
and ( n11742 , n547 , n11741 );
not ( n11743 , n547 );
not ( n11744 , n10439 );
and ( n11745 , n11743 , n11744 );
nor ( n11746 , n11742 , n11745 );
not ( n11747 , n3298 );
or ( n11748 , n11746 , n11747 );
nand ( n11749 , n11740 , n11748 );
xor ( n11750 , n11737 , n11749 );
xor ( n11751 , n11694 , n11750 );
xor ( n11752 , n11466 , n11649 );
and ( n11753 , n11752 , n11654 );
and ( n11754 , n11466 , n11649 );
or ( n11755 , n11753 , n11754 );
xor ( n11756 , n11751 , n11755 );
xor ( n11757 , n11470 , n11482 );
and ( n11758 , n11757 , n11648 );
and ( n11759 , n11470 , n11482 );
or ( n11760 , n11758 , n11759 );
xor ( n11761 , n11394 , n11398 );
and ( n11762 , n11761 , n11456 );
and ( n11763 , n11394 , n11398 );
or ( n11764 , n11762 , n11763 );
xor ( n11765 , n11760 , n11764 );
xor ( n11766 , n11377 , n11381 );
and ( n11767 , n11766 , n11393 );
and ( n11768 , n11377 , n11381 );
or ( n11769 , n11767 , n11768 );
not ( n11770 , n4020 );
and ( n11771 , n11241 , n549 );
not ( n11772 , n11241 );
and ( n11773 , n11772 , n4013 );
nor ( n11774 , n11771 , n11773 );
not ( n11775 , n11774 );
or ( n11776 , n11770 , n11775 );
nand ( n11777 , n11480 , n4022 );
nand ( n11778 , n11776 , n11777 );
xor ( n11779 , n11769 , n11778 );
not ( n11780 , n552 );
not ( n11781 , n551 );
not ( n11782 , n11609 );
not ( n11783 , n11637 );
or ( n11784 , n11782 , n11783 );
nand ( n11785 , n11784 , n11610 );
not ( n11786 , n11591 );
nand ( n11787 , n11786 , n11592 );
not ( n11788 , n11787 );
not ( n11789 , n11599 );
or ( n11790 , n11788 , n11789 );
not ( n11791 , n11592 );
nand ( n11792 , n11791 , n11591 );
nand ( n11793 , n11790 , n11792 );
nand ( n11794 , n2473 , n2027 );
nand ( n11795 , n11794 , n493 );
and ( n11796 , n489 , n509 );
xor ( n11797 , n11795 , n11796 );
not ( n11798 , n11597 );
not ( n11799 , n5487 );
or ( n11800 , n11798 , n11799 );
and ( n11801 , n491 , n505 );
not ( n11802 , n491 );
not ( n11803 , n505 );
and ( n11804 , n11802 , n11803 );
nor ( n11805 , n11801 , n11804 );
nand ( n11806 , n2764 , n11805 );
nand ( n11807 , n11800 , n11806 );
xor ( n11808 , n11797 , n11807 );
xor ( n11809 , n11793 , n11808 );
not ( n11810 , n11589 );
not ( n11811 , n4835 );
or ( n11812 , n11810 , n11811 );
xnor ( n11813 , n489 , n507 );
not ( n11814 , n11813 );
nand ( n11815 , n11814 , n4838 );
nand ( n11816 , n11812 , n11815 );
and ( n11817 , n11816 , n11584 );
not ( n11818 , n11816 );
and ( n11819 , n11818 , n11585 );
nor ( n11820 , n11817 , n11819 );
xor ( n11821 , n11809 , n11820 );
not ( n11822 , n11821 );
xor ( n11823 , n11585 , n11600 );
and ( n11824 , n11823 , n11605 );
and ( n11825 , n11585 , n11600 );
or ( n11826 , n11824 , n11825 );
not ( n11827 , n11826 );
not ( n11828 , n11827 );
or ( n11829 , n11822 , n11828 );
or ( n11830 , n11827 , n11821 );
nand ( n11831 , n11829 , n11830 );
or ( n11832 , n11573 , n11577 );
not ( n11833 , n11832 );
not ( n11834 , n11606 );
or ( n11835 , n11833 , n11834 );
nand ( n11836 , n11573 , n11577 );
nand ( n11837 , n11835 , n11836 );
nor ( n11838 , n11831 , n11837 );
not ( n11839 , n11838 );
nand ( n11840 , n11831 , n11837 );
nand ( n11841 , n11839 , n11840 );
not ( n11842 , n11841 );
and ( n11843 , n11785 , n11842 );
not ( n11844 , n11785 );
and ( n11845 , n11844 , n11841 );
nor ( n11846 , n11843 , n11845 );
nand ( n11847 , n11846 , n455 );
not ( n11848 , n11556 );
xor ( n11849 , n11496 , n11524 );
and ( n11850 , n11849 , n11529 );
and ( n11851 , n11496 , n11524 );
or ( n11852 , n11850 , n11851 );
or ( n11853 , n2966 , n2196 );
nand ( n11854 , n11853 , n493 );
not ( n11855 , n2606 );
not ( n11856 , n491 );
not ( n11857 , n4077 );
or ( n11858 , n11856 , n11857 );
nand ( n11859 , n4076 , n2613 );
nand ( n11860 , n11858 , n11859 );
not ( n11861 , n11860 );
or ( n11862 , n11855 , n11861 );
nand ( n11863 , n11513 , n3573 );
nand ( n11864 , n11862 , n11863 );
xor ( n11865 , n11854 , n11864 );
and ( n11866 , n489 , n5278 );
xor ( n11867 , n11865 , n11866 );
not ( n11868 , n4056 );
not ( n11869 , n11518 );
or ( n11870 , n11868 , n11869 );
xor ( n11871 , n489 , n4093 );
nand ( n11872 , n11871 , n4547 );
nand ( n11873 , n11870 , n11872 );
not ( n11874 , n11499 );
xor ( n11875 , n11873 , n11874 );
xor ( n11876 , n11505 , n11515 );
and ( n11877 , n11876 , n11522 );
and ( n11878 , n11505 , n11515 );
or ( n11879 , n11877 , n11878 );
xor ( n11880 , n11875 , n11879 );
xor ( n11881 , n11867 , n11880 );
xor ( n11882 , n11499 , n11503 );
and ( n11883 , n11882 , n11523 );
and ( n11884 , n11499 , n11503 );
or ( n11885 , n11883 , n11884 );
xor ( n11886 , n11881 , n11885 );
nand ( n11887 , n11852 , n11886 );
not ( n11888 , n11887 );
nor ( n11889 , n11886 , n11852 );
nor ( n11890 , n11888 , n11889 );
nand ( n11891 , n11890 , n716 );
nand ( n11892 , n11848 , n11891 , n11532 );
not ( n11893 , n716 );
nor ( n11894 , n11893 , n11890 );
not ( n11895 , n11531 );
nor ( n11896 , n11894 , n11895 );
nand ( n11897 , n11556 , n11896 );
and ( n11898 , n11891 , n11895 , n11532 );
nor ( n11899 , n11894 , n11532 );
nor ( n11900 , n11898 , n11899 );
nand ( n11901 , n11892 , n11897 , n11900 );
nand ( n11902 , n11847 , n11901 );
not ( n11903 , n11902 );
not ( n11904 , n11903 );
or ( n11905 , n11781 , n11904 );
nand ( n11906 , n11847 , n11901 );
not ( n11907 , n11906 );
not ( n11908 , n11907 );
nand ( n11909 , n11908 , n4018 );
nand ( n11910 , n11905 , n11909 );
not ( n11911 , n11910 );
or ( n11912 , n11780 , n11911 );
nand ( n11913 , n11646 , n5619 );
nand ( n11914 , n11912 , n11913 );
xor ( n11915 , n11779 , n11914 );
xor ( n11916 , n11765 , n11915 );
xor ( n11917 , n11756 , n11916 );
xor ( n11918 , n11457 , n11461 );
and ( n11919 , n11918 , n11655 );
and ( n11920 , n11457 , n11461 );
or ( n11921 , n11919 , n11920 );
nor ( n11922 , n11917 , n11921 );
not ( n11923 , n11922 );
nand ( n11924 , n10741 , n11664 , n11923 );
not ( n11925 , n11662 );
not ( n11926 , n11656 );
not ( n11927 , n11926 );
or ( n11928 , n11925 , n11927 );
nor ( n11929 , n11358 , n11071 );
nand ( n11930 , n11361 , n11365 );
or ( n11931 , n11929 , n11930 );
nand ( n11932 , n11358 , n11071 );
nand ( n11933 , n11931 , n11932 );
nand ( n11934 , n11928 , n11933 );
not ( n11935 , n11934 );
not ( n11936 , n11921 );
not ( n11937 , n11917 );
or ( n11938 , n11936 , n11937 );
nand ( n11939 , n11656 , n11661 );
nand ( n11940 , n11938 , n11939 );
or ( n11941 , n11935 , n11940 );
nand ( n11942 , n11941 , n11923 );
nand ( n11943 , n11924 , n11942 );
buf ( n11944 , n11943 );
xor ( n11945 , n11751 , n11755 );
and ( n11946 , n11945 , n11916 );
and ( n11947 , n11751 , n11755 );
or ( n11948 , n11946 , n11947 );
not ( n11949 , n3288 );
not ( n11950 , n11674 );
or ( n11951 , n11949 , n11950 );
nand ( n11952 , n541 , n10995 );
not ( n11953 , n11952 );
nand ( n11954 , n4638 , n3023 );
not ( n11955 , n11954 );
or ( n11956 , n11953 , n11955 );
nand ( n11957 , n11956 , n3214 );
nand ( n11958 , n11951 , n11957 );
not ( n11959 , n714 );
not ( n11960 , n11684 );
or ( n11961 , n11959 , n11960 );
and ( n11962 , n2123 , n5607 );
not ( n11963 , n2123 );
and ( n11964 , n11963 , n5614 );
nor ( n11965 , n11962 , n11964 );
nand ( n11966 , n11965 , n2362 );
nand ( n11967 , n11961 , n11966 );
xor ( n11968 , n11958 , n11967 );
not ( n11969 , n3017 );
not ( n11970 , n545 );
not ( n11971 , n11055 );
or ( n11972 , n11970 , n11971 );
nand ( n11973 , n706 , n10471 );
nand ( n11974 , n11972 , n11973 );
not ( n11975 , n11974 );
or ( n11976 , n11969 , n11975 );
nand ( n11977 , n11700 , n2376 );
nand ( n11978 , n11976 , n11977 );
xor ( n11979 , n11968 , n11978 );
xor ( n11980 , n11704 , n11736 );
and ( n11981 , n11980 , n11749 );
and ( n11982 , n11704 , n11736 );
or ( n11983 , n11981 , n11982 );
xor ( n11984 , n11979 , n11983 );
xor ( n11985 , n11706 , n11718 );
and ( n11986 , n11985 , n11735 );
and ( n11987 , n11706 , n11718 );
or ( n11988 , n11986 , n11987 );
not ( n11989 , n3298 );
and ( n11990 , n10949 , n2369 );
not ( n11991 , n10949 );
and ( n11992 , n11991 , n547 );
or ( n11993 , n11990 , n11992 );
not ( n11994 , n11993 );
or ( n11995 , n11989 , n11994 );
not ( n11996 , n3300 );
nor ( n11997 , n11996 , n2369 );
and ( n11998 , n11741 , n11997 );
nor ( n11999 , n11996 , n547 );
and ( n12000 , n10438 , n11999 );
nor ( n12001 , n11998 , n12000 );
nand ( n12002 , n11995 , n12001 );
xor ( n12003 , n11988 , n12002 );
not ( n12004 , n539 );
not ( n12005 , n3943 );
or ( n12006 , n12004 , n12005 );
nand ( n12007 , n4652 , n3069 );
nand ( n12008 , n12006 , n12007 );
not ( n12009 , n12008 );
not ( n12010 , n3026 );
or ( n12011 , n12009 , n12010 );
nand ( n12012 , n3103 , n11711 );
nand ( n12013 , n12011 , n12012 );
not ( n12014 , n11731 );
nor ( n12015 , n12014 , n11721 );
xor ( n12016 , n12013 , n12015 );
not ( n12017 , n11729 );
not ( n12018 , n11726 );
or ( n12019 , n12017 , n12018 );
not ( n12020 , n537 );
or ( n12021 , n716 , n2850 );
nand ( n12022 , n12021 , n3009 );
not ( n12023 , n12022 );
or ( n12024 , n12020 , n12023 );
nand ( n12025 , n3011 , n3177 );
nand ( n12026 , n12024 , n12025 );
nand ( n12027 , n12026 , n3134 );
nand ( n12028 , n12019 , n12027 );
not ( n12029 , n2356 );
nand ( n12030 , n12029 , n537 );
xnor ( n12031 , n12028 , n12030 );
xor ( n12032 , n12016 , n12031 );
xor ( n12033 , n12003 , n12032 );
xor ( n12034 , n11984 , n12033 );
xor ( n12035 , n11760 , n11764 );
and ( n12036 , n12035 , n11915 );
and ( n12037 , n11760 , n11764 );
or ( n12038 , n12036 , n12037 );
xor ( n12039 , n12034 , n12038 );
xor ( n12040 , n11769 , n11778 );
and ( n12041 , n12040 , n11914 );
and ( n12042 , n11769 , n11778 );
or ( n12043 , n12041 , n12042 );
not ( n12044 , n4022 );
not ( n12045 , n11774 );
or ( n12046 , n12044 , n12045 );
not ( n12047 , n3229 );
not ( n12048 , n11559 );
or ( n12049 , n12047 , n12048 );
nand ( n12050 , n12049 , n11639 );
and ( n12051 , n12050 , n4013 );
not ( n12052 , n12050 );
and ( n12053 , n12052 , n549 );
or ( n12054 , n12051 , n12053 );
nand ( n12055 , n12054 , n6220 );
nand ( n12056 , n12046 , n12055 );
xor ( n12057 , n11668 , n11678 );
and ( n12058 , n12057 , n11688 );
and ( n12059 , n11668 , n11678 );
or ( n12060 , n12058 , n12059 );
xor ( n12061 , n12056 , n12060 );
not ( n12062 , n5619 );
not ( n12063 , n11910 );
or ( n12064 , n12062 , n12063 );
not ( n12065 , n551 );
not ( n12066 , n716 );
or ( n12067 , n11852 , n11886 );
nand ( n12068 , n11531 , n12067 );
nor ( n12069 , n11545 , n12068 );
not ( n12070 , n12069 );
xor ( n12071 , n11867 , n11880 );
and ( n12072 , n12071 , n11885 );
and ( n12073 , n11867 , n11880 );
or ( n12074 , n12072 , n12073 );
not ( n12075 , n12074 );
xor ( n12076 , n11854 , n11864 );
and ( n12077 , n12076 , n11866 );
and ( n12078 , n11854 , n11864 );
or ( n12079 , n12077 , n12078 );
not ( n12080 , n4547 );
and ( n12081 , n489 , n3859 );
not ( n12082 , n489 );
and ( n12083 , n12082 , n3858 );
or ( n12084 , n12081 , n12083 );
not ( n12085 , n12084 );
or ( n12086 , n12080 , n12085 );
nand ( n12087 , n11871 , n4056 );
nand ( n12088 , n12086 , n12087 );
and ( n12089 , n489 , n10108 );
xor ( n12090 , n12088 , n12089 );
and ( n12091 , n3573 , n11860 );
nor ( n12092 , n2200 , n2613 );
nor ( n12093 , n12091 , n12092 );
xor ( n12094 , n12090 , n12093 );
xor ( n12095 , n12079 , n12094 );
xor ( n12096 , n11873 , n11874 );
and ( n12097 , n12096 , n11879 );
and ( n12098 , n11873 , n11874 );
or ( n12099 , n12097 , n12098 );
xor ( n12100 , n12095 , n12099 );
not ( n12101 , n12100 );
nand ( n12102 , n12075 , n12101 );
not ( n12103 , n12102 );
not ( n12104 , n12100 );
nor ( n12105 , n12104 , n12075 );
nor ( n12106 , n12103 , n12105 );
nor ( n12107 , n12070 , n12106 );
not ( n12108 , n12107 );
not ( n12109 , n11149 );
or ( n12110 , n12108 , n12109 );
not ( n12111 , n12068 );
and ( n12112 , n12111 , n11553 );
or ( n12113 , n11532 , n11889 );
nand ( n12114 , n12113 , n11887 );
nor ( n12115 , n12112 , n12114 );
or ( n12116 , n12115 , n12106 );
nand ( n12117 , n12110 , n12116 );
not ( n12118 , n12117 );
not ( n12119 , n11149 );
and ( n12120 , n12115 , n12106 );
and ( n12121 , n12119 , n12120 );
not ( n12122 , n12106 );
nor ( n12123 , n12122 , n12069 );
and ( n12124 , n12123 , n12115 );
nor ( n12125 , n12121 , n12124 );
nand ( n12126 , n12118 , n12125 );
not ( n12127 , n12126 );
or ( n12128 , n12066 , n12127 );
nor ( n12129 , n11608 , n11838 );
not ( n12130 , n12129 );
not ( n12131 , n11637 );
or ( n12132 , n12130 , n12131 );
or ( n12133 , n11838 , n11610 );
nand ( n12134 , n12133 , n11840 );
not ( n12135 , n12134 );
nand ( n12136 , n12132 , n12135 );
not ( n12137 , n11826 );
not ( n12138 , n11808 );
xnor ( n12139 , n11820 , n11793 );
nand ( n12140 , n12138 , n12139 );
not ( n12141 , n12140 );
or ( n12142 , n12137 , n12141 );
not ( n12143 , n12139 );
nand ( n12144 , n12143 , n11808 );
nand ( n12145 , n12142 , n12144 );
xor ( n12146 , n11795 , n11796 );
and ( n12147 , n12146 , n11807 );
and ( n12148 , n11795 , n11796 );
or ( n12149 , n12147 , n12148 );
and ( n12150 , n489 , n508 );
not ( n12151 , n11805 );
not ( n12152 , n5487 );
or ( n12153 , n12151 , n12152 );
nand ( n12154 , n2764 , n491 );
nand ( n12155 , n12153 , n12154 );
not ( n12156 , n12155 );
xor ( n12157 , n12150 , n12156 );
not ( n12158 , n4835 );
or ( n12159 , n12158 , n11813 );
not ( n12160 , n4838 );
and ( n12161 , n506 , n4046 );
not ( n12162 , n506 );
and ( n12163 , n12162 , n489 );
nor ( n12164 , n12161 , n12163 );
or ( n12165 , n12160 , n12164 );
nand ( n12166 , n12159 , n12165 );
xor ( n12167 , n12157 , n12166 );
xor ( n12168 , n12149 , n12167 );
not ( n12169 , n11793 );
not ( n12170 , n11816 );
nand ( n12171 , n12170 , n11585 );
not ( n12172 , n12171 );
or ( n12173 , n12169 , n12172 );
nand ( n12174 , n11584 , n11816 );
nand ( n12175 , n12173 , n12174 );
xor ( n12176 , n12168 , n12175 );
or ( n12177 , n12145 , n12176 );
nand ( n12178 , n12145 , n12176 );
nand ( n12179 , n12177 , n12178 );
not ( n12180 , n12179 );
and ( n12181 , n12136 , n12180 );
not ( n12182 , n12136 );
and ( n12183 , n12182 , n12179 );
nor ( n12184 , n12181 , n12183 );
nand ( n12185 , n12184 , n455 );
nand ( n12186 , n12128 , n12185 );
not ( n12187 , n12186 );
not ( n12188 , n12187 );
or ( n12189 , n12065 , n12188 );
not ( n12190 , n12187 );
nand ( n12191 , n12190 , n4018 );
nand ( n12192 , n12189 , n12191 );
nand ( n12193 , n12192 , n552 );
nand ( n12194 , n12064 , n12193 );
xor ( n12195 , n12061 , n12194 );
xor ( n12196 , n12043 , n12195 );
xor ( n12197 , n11689 , n11693 );
and ( n12198 , n12197 , n11750 );
and ( n12199 , n11689 , n11693 );
or ( n12200 , n12198 , n12199 );
xor ( n12201 , n12196 , n12200 );
xor ( n12202 , n12039 , n12201 );
or ( n12203 , n11948 , n12202 );
nand ( n12204 , n12202 , n11948 );
buf ( n12205 , n12204 );
nand ( n12206 , n12203 , n12205 );
not ( n12207 , n12206 );
and ( n12208 , n11944 , n12207 );
not ( n12209 , n11944 );
and ( n12210 , n12209 , n12206 );
nor ( n12211 , n12208 , n12210 );
nand ( n12212 , n12211 , n454 );
not ( n12213 , n8980 );
not ( n12214 , n7585 );
or ( n12215 , n12213 , n12214 );
xor ( n12216 , n527 , n461 );
nand ( n12217 , n7475 , n12216 );
nand ( n12218 , n12215 , n12217 );
not ( n12219 , n12218 );
nand ( n12220 , n533 , n457 );
not ( n12221 , n12220 );
and ( n12222 , n12219 , n12221 );
and ( n12223 , n12218 , n12220 );
nor ( n12224 , n12222 , n12223 );
not ( n12225 , n8990 );
not ( n12226 , n8728 );
or ( n12227 , n12225 , n12226 );
xor ( n12228 , n523 , n465 );
nand ( n12229 , n6987 , n12228 );
nand ( n12230 , n12227 , n12229 );
not ( n12231 , n12230 );
and ( n12232 , n12224 , n12231 );
not ( n12233 , n12224 );
and ( n12234 , n12233 , n12230 );
nor ( n12235 , n12232 , n12234 );
not ( n12236 , n8969 );
not ( n12237 , n7881 );
or ( n12238 , n12236 , n12237 );
xor ( n12239 , n529 , n459 );
nand ( n12240 , n7888 , n12239 );
nand ( n12241 , n12238 , n12240 );
xor ( n12242 , n8900 , n12241 );
not ( n12243 , n8906 );
not ( n12244 , n8337 );
or ( n12245 , n12243 , n12244 );
xor ( n12246 , n531 , n457 );
nand ( n12247 , n7908 , n12246 );
nand ( n12248 , n12245 , n12247 );
not ( n12249 , n12248 );
xnor ( n12250 , n12242 , n12249 );
xor ( n12251 , n12235 , n12250 );
nand ( n12252 , n8734 , n8901 );
or ( n12253 , n8734 , n8901 );
nand ( n12254 , n12253 , n8908 );
nand ( n12255 , n12252 , n12254 );
and ( n12256 , n12251 , n12255 );
and ( n12257 , n12235 , n12250 );
or ( n12258 , n12256 , n12257 );
not ( n12259 , n12258 );
not ( n12260 , n12248 );
not ( n12261 , n8900 );
or ( n12262 , n12260 , n12261 );
not ( n12263 , n8901 );
not ( n12264 , n12249 );
or ( n12265 , n12263 , n12264 );
nand ( n12266 , n12265 , n12241 );
nand ( n12267 , n12262 , n12266 );
not ( n12268 , n12267 );
not ( n12269 , n12228 );
not ( n12270 , n7035 );
or ( n12271 , n12269 , n12270 );
xor ( n12272 , n522 , n465 );
nand ( n12273 , n6987 , n12272 );
nand ( n12274 , n12271 , n12273 );
not ( n12275 , n12274 );
not ( n12276 , n12275 );
not ( n12277 , n12216 );
not ( n12278 , n8351 );
or ( n12279 , n12277 , n12278 );
xor ( n12280 , n526 , n461 );
nand ( n12281 , n7475 , n12280 );
nand ( n12282 , n12279 , n12281 );
not ( n12283 , n12282 );
or ( n12284 , n12276 , n12283 );
not ( n12285 , n12282 );
nand ( n12286 , n12285 , n12274 );
nand ( n12287 , n12284 , n12286 );
not ( n12288 , n12239 );
not ( n12289 , n7881 );
or ( n12290 , n12288 , n12289 );
xor ( n12291 , n528 , n459 );
nand ( n12292 , n7888 , n12291 );
nand ( n12293 , n12290 , n12292 );
not ( n12294 , n12293 );
and ( n12295 , n12287 , n12294 );
not ( n12296 , n12287 );
and ( n12297 , n12296 , n12293 );
nor ( n12298 , n12295 , n12297 );
and ( n12299 , n12268 , n12298 );
not ( n12300 , n12268 );
not ( n12301 , n12298 );
and ( n12302 , n12300 , n12301 );
nor ( n12303 , n12299 , n12302 );
nand ( n12304 , n532 , n457 );
not ( n12305 , n12246 );
not ( n12306 , n8674 );
or ( n12307 , n12305 , n12306 );
xor ( n12308 , n530 , n457 );
nand ( n12309 , n7908 , n12308 );
nand ( n12310 , n12307 , n12309 );
xor ( n12311 , n12304 , n12310 );
xor ( n12312 , n525 , n463 );
not ( n12313 , n12312 );
not ( n12314 , n8327 );
nor ( n12315 , n12313 , n12314 );
xor ( n12316 , n524 , n463 );
and ( n12317 , n7642 , n12316 );
nor ( n12318 , n12315 , n12317 );
xor ( n12319 , n12311 , n12318 );
not ( n12320 , n12319 );
and ( n12321 , n12303 , n12320 );
not ( n12322 , n12303 );
not ( n12323 , n12320 );
and ( n12324 , n12322 , n12323 );
nor ( n12325 , n12321 , n12324 );
not ( n12326 , n12325 );
not ( n12327 , n12326 );
not ( n12328 , n8888 );
not ( n12329 , n8881 );
not ( n12330 , n12329 );
or ( n12331 , n12328 , n12330 );
nor ( n12332 , n8888 , n12329 );
or ( n12333 , n8893 , n12332 );
nand ( n12334 , n12331 , n12333 );
not ( n12335 , n8976 );
not ( n12336 , n8992 );
or ( n12337 , n12335 , n12336 );
or ( n12338 , n8976 , n8992 );
nand ( n12339 , n12338 , n8982 );
nand ( n12340 , n12337 , n12339 );
xor ( n12341 , n12334 , n12340 );
not ( n12342 , n8891 );
not ( n12343 , n8327 );
or ( n12344 , n12342 , n12343 );
nand ( n12345 , n7026 , n12312 );
nand ( n12346 , n12344 , n12345 );
not ( n12347 , n7746 );
not ( n12348 , n6754 );
not ( n12349 , n12348 );
or ( n12350 , n12347 , n12349 );
nand ( n12351 , n12350 , n469 );
not ( n12352 , n12351 );
not ( n12353 , n12352 );
and ( n12354 , n8886 , n6948 );
nand ( n12355 , n6806 , n12354 );
not ( n12356 , n6806 );
xor ( n12357 , n521 , n467 );
nand ( n12358 , n12356 , n12357 );
nand ( n12359 , n12355 , n12358 );
not ( n12360 , n12359 );
or ( n12361 , n12353 , n12360 );
or ( n12362 , n12359 , n12352 );
nand ( n12363 , n12361 , n12362 );
xor ( n12364 , n12346 , n12363 );
and ( n12365 , n12341 , n12364 );
and ( n12366 , n12334 , n12340 );
or ( n12367 , n12365 , n12366 );
not ( n12368 , n12367 );
not ( n12369 , n12351 );
not ( n12370 , n12359 );
or ( n12371 , n12369 , n12370 );
nand ( n12372 , n12358 , n12352 , n12355 );
nand ( n12373 , n12346 , n12372 );
nand ( n12374 , n12371 , n12373 );
not ( n12375 , n12374 );
not ( n12376 , n12357 );
not ( n12377 , n7449 );
or ( n12378 , n12376 , n12377 );
nand ( n12379 , n7088 , n467 );
nand ( n12380 , n12378 , n12379 );
not ( n12381 , n12380 );
and ( n12382 , n12375 , n12381 );
not ( n12383 , n12359 );
not ( n12384 , n12351 );
or ( n12385 , n12383 , n12384 );
not ( n12386 , n12346 );
and ( n12387 , n12352 , n12358 , n12355 );
or ( n12388 , n12386 , n12387 );
nand ( n12389 , n12385 , n12388 );
not ( n12390 , n12380 );
not ( n12391 , n12390 );
and ( n12392 , n12389 , n12391 );
nor ( n12393 , n12382 , n12392 );
not ( n12394 , n12220 );
not ( n12395 , n12394 );
not ( n12396 , n12218 );
or ( n12397 , n12395 , n12396 );
or ( n12398 , n12218 , n12394 );
nand ( n12399 , n12398 , n12230 );
nand ( n12400 , n12397 , n12399 );
and ( n12401 , n12393 , n12400 );
not ( n12402 , n12393 );
not ( n12403 , n12400 );
and ( n12404 , n12402 , n12403 );
nor ( n12405 , n12401 , n12404 );
not ( n12406 , n12405 );
or ( n12407 , n12368 , n12406 );
or ( n12408 , n12367 , n12405 );
nand ( n12409 , n12407 , n12408 );
not ( n12410 , n12409 );
not ( n12411 , n12410 );
or ( n12412 , n12327 , n12411 );
nand ( n12413 , n12409 , n12325 );
nand ( n12414 , n12412 , n12413 );
not ( n12415 , n12414 );
or ( n12416 , n12259 , n12415 );
not ( n12417 , n12258 );
not ( n12418 , n12417 );
not ( n12419 , n12414 );
not ( n12420 , n12419 );
or ( n12421 , n12418 , n12420 );
not ( n12422 , n8959 );
nand ( n12423 , n12422 , n8967 );
not ( n12424 , n12423 );
not ( n12425 , n8993 );
or ( n12426 , n12424 , n12425 );
nand ( n12427 , n8966 , n8959 );
nand ( n12428 , n12426 , n12427 );
xor ( n12429 , n12334 , n12340 );
xor ( n12430 , n12429 , n12364 );
xor ( n12431 , n12428 , n12430 );
not ( n12432 , n8894 );
not ( n12433 , n8917 );
or ( n12434 , n12432 , n12433 );
nand ( n12435 , n12434 , n8926 );
nand ( n12436 , n8918 , n8895 );
nand ( n12437 , n12435 , n12436 );
and ( n12438 , n12431 , n12437 );
and ( n12439 , n12428 , n12430 );
or ( n12440 , n12438 , n12439 );
nand ( n12441 , n12421 , n12440 );
nand ( n12442 , n12416 , n12441 );
not ( n12443 , n12442 );
not ( n12444 , n6955 );
not ( n12445 , n12444 );
not ( n12446 , n7084 );
or ( n12447 , n12445 , n12446 );
nand ( n12448 , n12447 , n467 );
not ( n12449 , n12272 );
not ( n12450 , n8728 );
or ( n12451 , n12449 , n12450 );
xor ( n12452 , n521 , n465 );
nand ( n12453 , n6987 , n12452 );
nand ( n12454 , n12451 , n12453 );
xor ( n12455 , n12448 , n12454 );
not ( n12456 , n12280 );
not ( n12457 , n8719 );
or ( n12458 , n12456 , n12457 );
xor ( n12459 , n525 , n461 );
nand ( n12460 , n7475 , n12459 );
nand ( n12461 , n12458 , n12460 );
xor ( n12462 , n12455 , n12461 );
buf ( n12463 , n12462 );
not ( n12464 , n12463 );
or ( n12465 , n12318 , n12304 );
not ( n12466 , n12310 );
nand ( n12467 , n12465 , n12466 );
nand ( n12468 , n12318 , n12304 );
nand ( n12469 , n12467 , n12468 );
not ( n12470 , n12469 );
not ( n12471 , n12291 );
not ( n12472 , n7881 );
or ( n12473 , n12471 , n12472 );
xor ( n12474 , n527 , n459 );
nand ( n12475 , n7887 , n12474 );
nand ( n12476 , n12473 , n12475 );
not ( n12477 , n12476 );
not ( n12478 , n12316 );
not ( n12479 , n8327 );
or ( n12480 , n12478 , n12479 );
xor ( n12481 , n523 , n463 );
nand ( n12482 , n7642 , n12481 );
nand ( n12483 , n12480 , n12482 );
not ( n12484 , n12483 );
not ( n12485 , n12484 );
or ( n12486 , n12477 , n12485 );
not ( n12487 , n12483 );
or ( n12488 , n12487 , n12476 );
nand ( n12489 , n12486 , n12488 );
not ( n12490 , n12308 );
not ( n12491 , n8337 );
or ( n12492 , n12490 , n12491 );
xor ( n12493 , n529 , n457 );
nand ( n12494 , n7908 , n12493 );
nand ( n12495 , n12492 , n12494 );
not ( n12496 , n12495 );
and ( n12497 , n12489 , n12496 );
not ( n12498 , n12489 );
and ( n12499 , n12498 , n12495 );
nor ( n12500 , n12497 , n12499 );
not ( n12501 , n12500 );
not ( n12502 , n12501 );
or ( n12503 , n12470 , n12502 );
not ( n12504 , n12469 );
nand ( n12505 , n12500 , n12504 );
nand ( n12506 , n12503 , n12505 );
not ( n12507 , n12506 );
or ( n12508 , n12464 , n12507 );
or ( n12509 , n12506 , n12463 );
nand ( n12510 , n12508 , n12509 );
not ( n12511 , n12510 );
not ( n12512 , n12275 );
not ( n12513 , n12285 );
or ( n12514 , n12512 , n12513 );
nand ( n12515 , n12514 , n12293 );
nand ( n12516 , n12282 , n12274 );
nand ( n12517 , n12515 , n12516 );
not ( n12518 , n12390 );
nand ( n12519 , n531 , n457 );
not ( n12520 , n12519 );
not ( n12521 , n12520 );
and ( n12522 , n12518 , n12521 );
and ( n12523 , n12390 , n12520 );
nor ( n12524 , n12522 , n12523 );
or ( n12525 , n12517 , n12524 );
nand ( n12526 , n12524 , n12517 );
nand ( n12527 , n12525 , n12526 );
not ( n12528 , n12400 );
not ( n12529 , n12391 );
not ( n12530 , n12529 );
or ( n12531 , n12528 , n12530 );
or ( n12532 , n12529 , n12400 );
nand ( n12533 , n12532 , n12374 );
nand ( n12534 , n12531 , n12533 );
xor ( n12535 , n12527 , n12534 );
not ( n12536 , n12267 );
not ( n12537 , n12319 );
or ( n12538 , n12536 , n12537 );
not ( n12539 , n12320 );
not ( n12540 , n12268 );
or ( n12541 , n12539 , n12540 );
nand ( n12542 , n12541 , n12301 );
nand ( n12543 , n12538 , n12542 );
xor ( n12544 , n12535 , n12543 );
not ( n12545 , n12544 );
or ( n12546 , n12511 , n12545 );
or ( n12547 , n12544 , n12510 );
nand ( n12548 , n12546 , n12547 );
not ( n12549 , n12548 );
buf ( n12550 , n12367 );
not ( n12551 , n12550 );
nand ( n12552 , n12551 , n12405 );
not ( n12553 , n12552 );
not ( n12554 , n12326 );
or ( n12555 , n12553 , n12554 );
not ( n12556 , n12405 );
nand ( n12557 , n12556 , n12550 );
nand ( n12558 , n12555 , n12557 );
not ( n12559 , n12558 );
nand ( n12560 , n12549 , n12559 );
nand ( n12561 , n12558 , n12548 );
nand ( n12562 , n12560 , n12561 );
nand ( n12563 , n12443 , n12562 );
xor ( n12564 , n8953 , n8994 );
and ( n12565 , n12564 , n9003 );
and ( n12566 , n8953 , n8994 );
or ( n12567 , n12565 , n12566 );
xor ( n12568 , n12235 , n12250 );
xor ( n12569 , n12568 , n12255 );
or ( n12570 , n12567 , n12569 );
xor ( n12571 , n12428 , n12430 );
xor ( n12572 , n12571 , n12437 );
buf ( n12573 , n12572 );
nand ( n12574 , n12570 , n12573 );
nand ( n12575 , n12567 , n12569 );
nand ( n12576 , n12574 , n12575 );
not ( n12577 , n12576 );
not ( n12578 , n12326 );
not ( n12579 , n12410 );
or ( n12580 , n12578 , n12579 );
nand ( n12581 , n12580 , n12413 );
xor ( n12582 , n12258 , n12581 );
xnor ( n12583 , n12582 , n12440 );
nand ( n12584 , n12577 , n12583 );
nand ( n12585 , n12563 , n12584 );
not ( n12586 , n12585 );
buf ( n12587 , n12586 );
not ( n12588 , n12587 );
xor ( n12589 , n12569 , n12572 );
xnor ( n12590 , n12589 , n12567 );
not ( n12591 , n8928 );
not ( n12592 , n9004 );
or ( n12593 , n12591 , n12592 );
or ( n12594 , n8928 , n9004 );
buf ( n12595 , n8941 );
nand ( n12596 , n12594 , n12595 );
nand ( n12597 , n12593 , n12596 );
not ( n12598 , n12597 );
nand ( n12599 , n12590 , n12598 );
and ( n12600 , n12599 , n9020 );
and ( n12601 , n8642 , n12600 , n9031 );
not ( n12602 , n12601 );
nand ( n12603 , n12590 , n12598 );
nand ( n12604 , n12603 , n9020 );
not ( n12605 , n12604 );
nand ( n12606 , n12605 , n9036 );
not ( n12607 , n9025 );
not ( n12608 , n12603 );
or ( n12609 , n12607 , n12608 );
not ( n12610 , n12590 );
nand ( n12611 , n12610 , n12597 );
nand ( n12612 , n12609 , n12611 );
not ( n12613 , n12612 );
nand ( n12614 , n12606 , n12613 );
not ( n12615 , n12614 );
nand ( n12616 , n12602 , n12615 );
not ( n12617 , n12616 );
or ( n12618 , n12588 , n12617 );
buf ( n12619 , n12560 );
and ( n12620 , n12619 , n12561 );
nor ( n12621 , n12620 , n12442 );
not ( n12622 , n12583 );
nand ( n12623 , n12622 , n12576 );
or ( n12624 , n12621 , n12623 );
not ( n12625 , n12562 );
nand ( n12626 , n12625 , n12442 );
nand ( n12627 , n12624 , n12626 );
not ( n12628 , n12627 );
nand ( n12629 , n12618 , n12628 );
not ( n12630 , n12510 );
not ( n12631 , n12630 );
not ( n12632 , n12544 );
or ( n12633 , n12631 , n12632 );
not ( n12634 , n12510 );
not ( n12635 , n12544 );
not ( n12636 , n12635 );
or ( n12637 , n12634 , n12636 );
nand ( n12638 , n12637 , n12558 );
nand ( n12639 , n12633 , n12638 );
not ( n12640 , n12476 );
not ( n12641 , n12640 );
not ( n12642 , n12487 );
or ( n12643 , n12641 , n12642 );
nand ( n12644 , n12643 , n12495 );
or ( n12645 , n12487 , n12640 );
nand ( n12646 , n12644 , n12645 );
xor ( n12647 , n12448 , n12454 );
and ( n12648 , n12647 , n12461 );
and ( n12649 , n12448 , n12454 );
or ( n12650 , n12648 , n12649 );
xor ( n12651 , n12646 , n12650 );
not ( n12652 , n12493 );
not ( n12653 , n8674 );
or ( n12654 , n12652 , n12653 );
xor ( n12655 , n528 , n457 );
nand ( n12656 , n12655 , n7908 );
nand ( n12657 , n12654 , n12656 );
not ( n12658 , n12657 );
not ( n12659 , n12452 );
not ( n12660 , n7035 );
or ( n12661 , n12659 , n12660 );
not ( n12662 , n8984 );
nand ( n12663 , n12662 , n465 );
nand ( n12664 , n12661 , n12663 );
not ( n12665 , n12664 );
not ( n12666 , n12474 );
not ( n12667 , n7880 );
or ( n12668 , n12666 , n12667 );
xor ( n12669 , n526 , n459 );
nand ( n12670 , n7887 , n12669 );
nand ( n12671 , n12668 , n12670 );
not ( n12672 , n12671 );
not ( n12673 , n12672 );
and ( n12674 , n12665 , n12673 );
and ( n12675 , n12664 , n12672 );
nor ( n12676 , n12674 , n12675 );
not ( n12677 , n12676 );
or ( n12678 , n12658 , n12677 );
or ( n12679 , n12676 , n12657 );
nand ( n12680 , n12678 , n12679 );
xor ( n12681 , n12651 , n12680 );
xor ( n12682 , n12527 , n12534 );
and ( n12683 , n12682 , n12543 );
and ( n12684 , n12527 , n12534 );
or ( n12685 , n12683 , n12684 );
xor ( n12686 , n12681 , n12685 );
not ( n12687 , n12469 );
not ( n12688 , n12500 );
or ( n12689 , n12687 , n12688 );
nand ( n12690 , n12689 , n12462 );
nand ( n12691 , n12501 , n12504 );
nand ( n12692 , n12690 , n12691 );
not ( n12693 , n12692 );
nand ( n12694 , n12390 , n12519 );
not ( n12695 , n12694 );
not ( n12696 , n12517 );
or ( n12697 , n12695 , n12696 );
nand ( n12698 , n12391 , n12520 );
nand ( n12699 , n12697 , n12698 );
nand ( n12700 , n530 , n457 );
not ( n12701 , n12700 );
not ( n12702 , n12701 );
not ( n12703 , n12481 );
not ( n12704 , n8327 );
or ( n12705 , n12703 , n12704 );
xor ( n12706 , n522 , n463 );
nand ( n12707 , n7026 , n12706 );
nand ( n12708 , n12705 , n12707 );
not ( n12709 , n12708 );
or ( n12710 , n12702 , n12709 );
not ( n12711 , n12708 );
nand ( n12712 , n12711 , n12700 );
nand ( n12713 , n12710 , n12712 );
not ( n12714 , n12459 );
not ( n12715 , n8719 );
or ( n12716 , n12714 , n12715 );
xor ( n12717 , n524 , n461 );
nand ( n12718 , n7475 , n12717 );
nand ( n12719 , n12716 , n12718 );
not ( n12720 , n12719 );
xor ( n12721 , n12713 , n12720 );
xor ( n12722 , n12699 , n12721 );
not ( n12723 , n12722 );
or ( n12724 , n12693 , n12723 );
or ( n12725 , n12692 , n12722 );
nand ( n12726 , n12724 , n12725 );
xor ( n12727 , n12686 , n12726 );
nor ( n12728 , n12639 , n12727 );
not ( n12729 , n12728 );
nand ( n12730 , n12727 , n12639 );
nand ( n12731 , n12729 , n12730 );
not ( n12732 , n12731 );
and ( n12733 , n12629 , n12732 );
not ( n12734 , n12629 );
and ( n12735 , n12734 , n12731 );
nor ( n12736 , n12733 , n12735 );
buf ( n12737 , n12736 );
not ( n12738 , n12737 );
nand ( n12739 , n12738 , n8305 );
not ( n12740 , n9625 );
not ( n12741 , n12601 );
nand ( n12742 , n12586 , n12729 );
not ( n12743 , n12742 );
not ( n12744 , n12743 );
or ( n12745 , n12741 , n12744 );
not ( n12746 , n12606 );
nand ( n12747 , n12746 , n12743 );
nand ( n12748 , n12745 , n12747 );
not ( n12749 , n12748 );
not ( n12750 , n12612 );
not ( n12751 , n12750 );
not ( n12752 , n12742 );
and ( n12753 , n12751 , n12752 );
xor ( n12754 , n12646 , n12650 );
and ( n12755 , n12754 , n12680 );
and ( n12756 , n12646 , n12650 );
or ( n12757 , n12755 , n12756 );
not ( n12758 , n12757 );
not ( n12759 , n12758 );
not ( n12760 , n12672 );
not ( n12761 , n12657 );
not ( n12762 , n12761 );
or ( n12763 , n12760 , n12762 );
nand ( n12764 , n12763 , n12664 );
nand ( n12765 , n12671 , n12657 );
nand ( n12766 , n12764 , n12765 );
not ( n12767 , n12766 );
not ( n12768 , n12708 );
or ( n12769 , n12767 , n12768 );
not ( n12770 , n12708 );
nand ( n12771 , n12770 , n12764 , n12765 );
nand ( n12772 , n12769 , n12771 );
nand ( n12773 , n529 , n457 );
not ( n12774 , n12773 );
not ( n12775 , n12655 );
not ( n12776 , n8674 );
or ( n12777 , n12775 , n12776 );
xor ( n12778 , n527 , n457 );
nand ( n12779 , n7908 , n12778 );
nand ( n12780 , n12777 , n12779 );
xor ( n12781 , n12774 , n12780 );
not ( n12782 , n12717 );
not ( n12783 , n7585 );
or ( n12784 , n12782 , n12783 );
xor ( n12785 , n523 , n461 );
nand ( n12786 , n7475 , n12785 );
nand ( n12787 , n12784 , n12786 );
xnor ( n12788 , n12781 , n12787 );
and ( n12789 , n12772 , n12788 );
not ( n12790 , n12772 );
not ( n12791 , n12788 );
and ( n12792 , n12790 , n12791 );
nor ( n12793 , n12789 , n12792 );
nand ( n12794 , n12711 , n12701 );
not ( n12795 , n12794 );
not ( n12796 , n12720 );
or ( n12797 , n12795 , n12796 );
nand ( n12798 , n12700 , n12708 );
nand ( n12799 , n12797 , n12798 );
not ( n12800 , n12706 );
not ( n12801 , n8327 );
or ( n12802 , n12800 , n12801 );
xor ( n12803 , n521 , n463 );
nand ( n12804 , n7642 , n12803 );
nand ( n12805 , n12802 , n12804 );
not ( n12806 , n12669 );
not ( n12807 , n7881 );
or ( n12808 , n12806 , n12807 );
xor ( n12809 , n525 , n459 );
nand ( n12810 , n7888 , n12809 );
nand ( n12811 , n12808 , n12810 );
xor ( n12812 , n12805 , n12811 );
or ( n12813 , n6987 , n8728 );
nand ( n12814 , n12813 , n465 );
xor ( n12815 , n12812 , n12814 );
and ( n12816 , n12799 , n12815 );
not ( n12817 , n12799 );
not ( n12818 , n12815 );
and ( n12819 , n12817 , n12818 );
nor ( n12820 , n12816 , n12819 );
and ( n12821 , n12793 , n12820 );
not ( n12822 , n12793 );
not ( n12823 , n12820 );
and ( n12824 , n12822 , n12823 );
nor ( n12825 , n12821 , n12824 );
not ( n12826 , n12825 );
not ( n12827 , n12826 );
or ( n12828 , n12759 , n12827 );
nand ( n12829 , n12825 , n12757 );
nand ( n12830 , n12828 , n12829 );
not ( n12831 , n12699 );
nand ( n12832 , n12831 , n12721 );
not ( n12833 , n12832 );
not ( n12834 , n12692 );
or ( n12835 , n12833 , n12834 );
not ( n12836 , n12721 );
nand ( n12837 , n12836 , n12699 );
nand ( n12838 , n12835 , n12837 );
not ( n12839 , n12838 );
and ( n12840 , n12830 , n12839 );
not ( n12841 , n12830 );
and ( n12842 , n12841 , n12838 );
nor ( n12843 , n12840 , n12842 );
not ( n12844 , n12843 );
xor ( n12845 , n12681 , n12685 );
and ( n12846 , n12845 , n12726 );
and ( n12847 , n12681 , n12685 );
or ( n12848 , n12846 , n12847 );
nand ( n12849 , n12844 , n12848 );
not ( n12850 , n12848 );
nand ( n12851 , n12843 , n12850 );
nand ( n12852 , n12849 , n12851 );
nor ( n12853 , n12753 , n12852 );
not ( n12854 , n12729 );
not ( n12855 , n12627 );
or ( n12856 , n12854 , n12855 );
nand ( n12857 , n12856 , n12730 );
not ( n12858 , n12857 );
nand ( n12859 , n12749 , n12853 , n12858 );
not ( n12860 , n12750 );
nand ( n12861 , n12860 , n12743 );
nand ( n12862 , n12861 , n12858 );
or ( n12863 , n12862 , n12748 );
nand ( n12864 , n12863 , n12852 );
nand ( n12865 , n12859 , n12864 );
not ( n12866 , n12865 );
nand ( n12867 , n12740 , n12866 );
not ( n12868 , n12866 );
nand ( n12869 , n12868 , n9627 );
nand ( n12870 , n12739 , n12867 , n12869 );
not ( n12871 , n6848 );
not ( n12872 , n489 );
not ( n12873 , n9570 );
or ( n12874 , n12872 , n12873 );
nand ( n12875 , n8498 , n4046 );
nand ( n12876 , n12874 , n12875 );
not ( n12877 , n12876 );
or ( n12878 , n12871 , n12877 );
xor ( n12879 , n489 , n7383 );
nand ( n12880 , n12879 , n6867 );
nand ( n12881 , n12878 , n12880 );
and ( n12882 , n489 , n7395 );
xor ( n12883 , n12881 , n12882 );
not ( n12884 , n6842 );
not ( n12885 , n491 );
not ( n12886 , n8843 );
or ( n12887 , n12885 , n12886 );
nand ( n12888 , n7511 , n6892 );
nand ( n12889 , n12887 , n12888 );
not ( n12890 , n12889 );
or ( n12891 , n12884 , n12890 );
not ( n12892 , n491 );
not ( n12893 , n7298 );
or ( n12894 , n12892 , n12893 );
nand ( n12895 , n7301 , n6892 );
nand ( n12896 , n12894 , n12895 );
nand ( n12897 , n12896 , n6719 );
nand ( n12898 , n12891 , n12897 );
xor ( n12899 , n12883 , n12898 );
not ( n12900 , n8258 );
and ( n12901 , n497 , n12900 );
not ( n12902 , n497 );
and ( n12903 , n12902 , n8258 );
nor ( n12904 , n12901 , n12903 );
not ( n12905 , n12904 );
or ( n12906 , n12905 , n9467 );
not ( n12907 , n497 );
not ( n12908 , n8475 );
or ( n12909 , n12907 , n12908 );
or ( n12910 , n8475 , n497 );
nand ( n12911 , n12909 , n12910 );
or ( n12912 , n12911 , n7411 );
nand ( n12913 , n12906 , n12912 );
xor ( n12914 , n12899 , n12913 );
and ( n12915 , n499 , n8795 );
not ( n12916 , n499 );
and ( n12917 , n12916 , n8792 );
nor ( n12918 , n12915 , n12917 );
or ( n12919 , n12918 , n7557 );
and ( n12920 , n499 , n9049 );
not ( n12921 , n499 );
and ( n12922 , n12921 , n9045 );
nor ( n12923 , n12920 , n12922 );
not ( n12924 , n12923 );
or ( n12925 , n12924 , n7814 );
nand ( n12926 , n12919 , n12925 );
and ( n12927 , n12914 , n12926 );
and ( n12928 , n12899 , n12913 );
or ( n12929 , n12927 , n12928 );
xor ( n12930 , n12870 , n12929 );
and ( n12931 , n495 , n8282 );
not ( n12932 , n495 );
and ( n12933 , n12932 , n8286 );
or ( n12934 , n12931 , n12933 );
not ( n12935 , n12934 );
not ( n12936 , n7326 );
or ( n12937 , n12935 , n12936 );
and ( n12938 , n495 , n8255 );
not ( n12939 , n495 );
and ( n12940 , n12939 , n12900 );
or ( n12941 , n12938 , n12940 );
nand ( n12942 , n6939 , n12941 );
nand ( n12943 , n12937 , n12942 );
not ( n12944 , n7517 );
and ( n12945 , n497 , n8795 );
not ( n12946 , n497 );
and ( n12947 , n12946 , n8792 );
or ( n12948 , n12945 , n12947 );
not ( n12949 , n12948 );
or ( n12950 , n12944 , n12949 );
not ( n12951 , n12911 );
nand ( n12952 , n12951 , n7415 );
nand ( n12953 , n12950 , n12952 );
xor ( n12954 , n12943 , n12953 );
not ( n12955 , n7405 );
and ( n12956 , n493 , n7677 );
not ( n12957 , n493 );
and ( n12958 , n12957 , n8625 );
nor ( n12959 , n12956 , n12958 );
not ( n12960 , n12959 );
or ( n12961 , n12955 , n12960 );
and ( n12962 , n493 , n8589 );
not ( n12963 , n493 );
and ( n12964 , n12963 , n7812 );
or ( n12965 , n12962 , n12964 );
nand ( n12966 , n12965 , n7371 );
nand ( n12967 , n12961 , n12966 );
not ( n12968 , n6848 );
not ( n12969 , n12879 );
or ( n12970 , n12968 , n12969 );
xor ( n12971 , n489 , n7395 );
nand ( n12972 , n12971 , n6867 );
nand ( n12973 , n12970 , n12972 );
and ( n12974 , n489 , n7339 );
xor ( n12975 , n12973 , n12974 );
nand ( n12976 , n6842 , n491 );
not ( n12977 , n12976 );
nand ( n12978 , n12977 , n7298 );
nor ( n12979 , n6843 , n491 );
nand ( n12980 , n7301 , n12979 );
and ( n12981 , n8498 , n6892 );
not ( n12982 , n8498 );
and ( n12983 , n12982 , n491 );
or ( n12984 , n12981 , n12983 );
nand ( n12985 , n12984 , n6719 );
nand ( n12986 , n12978 , n12980 , n12985 );
and ( n12987 , n12975 , n12986 );
and ( n12988 , n12973 , n12974 );
or ( n12989 , n12987 , n12988 );
xor ( n12990 , n12967 , n12989 );
not ( n12991 , n6939 );
not ( n12992 , n12934 );
or ( n12993 , n12991 , n12992 );
xor ( n12994 , n495 , n8581 );
nand ( n12995 , n12994 , n7326 );
nand ( n12996 , n12993 , n12995 );
and ( n12997 , n12990 , n12996 );
and ( n12998 , n12967 , n12989 );
or ( n12999 , n12997 , n12998 );
xor ( n13000 , n12954 , n12999 );
xor ( n13001 , n12930 , n13000 );
xor ( n13002 , n12899 , n12913 );
xor ( n13003 , n13002 , n12926 );
not ( n13004 , n6848 );
not ( n13005 , n12971 );
or ( n13006 , n13004 , n13005 );
xor ( n13007 , n489 , n7339 );
nand ( n13008 , n13007 , n6867 );
nand ( n13009 , n13006 , n13008 );
and ( n13010 , n489 , n6836 );
xor ( n13011 , n13009 , n13010 );
not ( n13012 , n6842 );
not ( n13013 , n12984 );
or ( n13014 , n13012 , n13013 );
not ( n13015 , n491 );
not ( n13016 , n7384 );
or ( n13017 , n13015 , n13016 );
nand ( n13018 , n7383 , n6892 );
nand ( n13019 , n13017 , n13018 );
nand ( n13020 , n13019 , n6719 );
nand ( n13021 , n13014 , n13020 );
and ( n13022 , n13011 , n13021 );
and ( n13023 , n13009 , n13010 );
or ( n13024 , n13022 , n13023 );
not ( n13025 , n493 );
not ( n13026 , n8843 );
or ( n13027 , n13025 , n13026 );
not ( n13028 , n493 );
nand ( n13029 , n13028 , n7511 );
nand ( n13030 , n13027 , n13029 );
nand ( n13031 , n13030 , n7405 );
nand ( n13032 , n7369 , n493 );
or ( n13033 , n7677 , n13032 );
nor ( n13034 , n7370 , n493 );
nand ( n13035 , n7677 , n13034 );
nand ( n13036 , n13031 , n13033 , n13035 );
xor ( n13037 , n13024 , n13036 );
xor ( n13038 , n12973 , n12974 );
xor ( n13039 , n13038 , n12986 );
and ( n13040 , n13037 , n13039 );
and ( n13041 , n13024 , n13036 );
or ( n13042 , n13040 , n13041 );
xor ( n13043 , n12967 , n12989 );
xor ( n13044 , n13043 , n12996 );
xor ( n13045 , n13042 , n13044 );
not ( n13046 , n8297 );
not ( n13047 , n9021 );
not ( n13048 , n13047 );
not ( n13049 , n9038 );
or ( n13050 , n13048 , n13049 );
nand ( n13051 , n13050 , n9026 );
not ( n13052 , n13051 );
nand ( n13053 , n12611 , n12599 );
not ( n13054 , n13053 );
and ( n13055 , n13052 , n13054 );
and ( n13056 , n13051 , n13053 );
nor ( n13057 , n13055 , n13056 );
not ( n13058 , n13057 );
not ( n13059 , n13058 );
not ( n13060 , n13059 );
and ( n13061 , n501 , n13060 );
not ( n13062 , n501 );
not ( n13063 , n13058 );
and ( n13064 , n13062 , n13063 );
nor ( n13065 , n13061 , n13064 );
not ( n13066 , n13065 );
or ( n13067 , n13046 , n13066 );
not ( n13068 , n501 );
buf ( n13069 , n12623 );
nand ( n13070 , n12584 , n13069 );
not ( n13071 , n13070 );
not ( n13072 , n12601 );
nand ( n13073 , n13072 , n12615 );
not ( n13074 , n13073 );
or ( n13075 , n13071 , n13074 );
not ( n13076 , n12616 );
not ( n13077 , n13070 );
nand ( n13078 , n13076 , n13077 );
nand ( n13079 , n13075 , n13078 );
not ( n13080 , n13079 );
not ( n13081 , n13080 );
or ( n13082 , n13068 , n13081 );
not ( n13083 , n13079 );
not ( n13084 , n13083 );
nand ( n13085 , n13084 , n8260 );
nand ( n13086 , n13082 , n13085 );
nand ( n13087 , n13086 , n7828 );
nand ( n13088 , n13067 , n13087 );
xor ( n13089 , n13045 , n13088 );
xor ( n13090 , n13003 , n13089 );
not ( n13091 , n8841 );
not ( n13092 , n12994 );
or ( n13093 , n13091 , n13092 );
and ( n13094 , n7811 , n495 );
not ( n13095 , n7811 );
and ( n13096 , n13095 , n719 );
nor ( n13097 , n13094 , n13096 );
nand ( n13098 , n13097 , n7326 );
nand ( n13099 , n13093 , n13098 );
and ( n13100 , n489 , n6787 );
not ( n13101 , n6848 );
not ( n13102 , n13007 );
or ( n13103 , n13101 , n13102 );
nand ( n13104 , n9074 , n6867 );
nand ( n13105 , n13103 , n13104 );
xor ( n13106 , n13100 , n13105 );
not ( n13107 , n9085 );
not ( n13108 , n6719 );
or ( n13109 , n13107 , n13108 );
not ( n13110 , n13019 );
or ( n13111 , n13110 , n6843 );
nand ( n13112 , n13109 , n13111 );
and ( n13113 , n13106 , n13112 );
and ( n13114 , n13100 , n13105 );
or ( n13115 , n13113 , n13114 );
not ( n13116 , n7371 );
not ( n13117 , n13030 );
or ( n13118 , n13116 , n13117 );
xor ( n13119 , n493 , n7301 );
nand ( n13120 , n13119 , n7405 );
nand ( n13121 , n13118 , n13120 );
xor ( n13122 , n13115 , n13121 );
xor ( n13123 , n13009 , n13010 );
xor ( n13124 , n13123 , n13021 );
and ( n13125 , n13122 , n13124 );
and ( n13126 , n13115 , n13121 );
or ( n13127 , n13125 , n13126 );
xor ( n13128 , n13099 , n13127 );
not ( n13129 , n7415 );
and ( n13130 , n497 , n9167 );
not ( n13131 , n497 );
and ( n13132 , n13131 , n8282 );
nor ( n13133 , n13130 , n13132 );
not ( n13134 , n13133 );
or ( n13135 , n13129 , n13134 );
nand ( n13136 , n7517 , n12904 );
nand ( n13137 , n13135 , n13136 );
xor ( n13138 , n13128 , n13137 );
not ( n13139 , n7828 );
not ( n13140 , n13065 );
or ( n13141 , n13139 , n13140 );
not ( n13142 , n501 );
not ( n13143 , n9045 );
or ( n13144 , n13142 , n13143 );
nand ( n13145 , n9046 , n8260 );
nand ( n13146 , n13144 , n13145 );
nand ( n13147 , n13146 , n8297 );
nand ( n13148 , n13141 , n13147 );
xor ( n13149 , n13138 , n13148 );
not ( n13150 , n504 );
not ( n13151 , n13073 );
not ( n13152 , n13069 );
and ( n13153 , n12626 , n12563 );
not ( n13154 , n13153 );
nor ( n13155 , n13152 , n13154 );
nand ( n13156 , n13151 , n13155 );
not ( n13157 , n12584 );
nor ( n13158 , n13153 , n13157 );
nand ( n13159 , n13073 , n13158 );
not ( n13160 , n13153 );
not ( n13161 , n13069 );
and ( n13162 , n13160 , n13161 );
nand ( n13163 , n13069 , n13157 );
nor ( n13164 , n13163 , n13154 );
nor ( n13165 , n13162 , n13164 );
nand ( n13166 , n13156 , n13159 , n13165 );
buf ( n13167 , n13166 );
not ( n13168 , n13167 );
and ( n13169 , n8880 , n13168 );
not ( n13170 , n8880 );
and ( n13171 , n13170 , n13167 );
or ( n13172 , n13169 , n13171 );
not ( n13173 , n13172 );
not ( n13174 , n13173 );
or ( n13175 , n13150 , n13174 );
not ( n13176 , n503 );
not ( n13177 , n13080 );
or ( n13178 , n13176 , n13177 );
not ( n13179 , n13079 );
not ( n13180 , n13179 );
nand ( n13181 , n13180 , n8880 );
nand ( n13182 , n13178 , n13181 );
nand ( n13183 , n13182 , n8306 );
nand ( n13184 , n13175 , n13183 );
and ( n13185 , n13149 , n13184 );
and ( n13186 , n13138 , n13148 );
or ( n13187 , n13185 , n13186 );
and ( n13188 , n13090 , n13187 );
and ( n13189 , n13003 , n13089 );
or ( n13190 , n13188 , n13189 );
xor ( n13191 , n13001 , n13190 );
xor ( n13192 , n13042 , n13044 );
and ( n13193 , n13192 , n13088 );
and ( n13194 , n13042 , n13044 );
or ( n13195 , n13193 , n13194 );
xor ( n13196 , n13099 , n13127 );
and ( n13197 , n13196 , n13137 );
and ( n13198 , n13099 , n13127 );
or ( n13199 , n13197 , n13198 );
nor ( n13200 , n8792 , n7818 );
not ( n13201 , n13200 );
not ( n13202 , n8478 );
nand ( n13203 , n7558 , n499 );
not ( n13204 , n13203 );
and ( n13205 , n13202 , n13204 );
nor ( n13206 , n7557 , n499 );
and ( n13207 , n8478 , n13206 );
nor ( n13208 , n13205 , n13207 );
nand ( n13209 , n8792 , n7815 );
nand ( n13210 , n13201 , n13208 , n13209 );
xor ( n13211 , n13024 , n13036 );
xor ( n13212 , n13211 , n13039 );
xor ( n13213 , n13210 , n13212 );
not ( n13214 , n6939 );
not ( n13215 , n13097 );
or ( n13216 , n13214 , n13215 );
and ( n13217 , n495 , n7678 );
not ( n13218 , n495 );
and ( n13219 , n13218 , n7677 );
nor ( n13220 , n13217 , n13219 );
not ( n13221 , n7326 );
or ( n13222 , n13220 , n13221 );
nand ( n13223 , n13216 , n13222 );
nor ( n13224 , n9467 , n497 );
not ( n13225 , n13224 );
not ( n13226 , n8581 );
or ( n13227 , n13225 , n13226 );
nor ( n13228 , n7411 , n497 );
nand ( n13229 , n8281 , n13228 );
nand ( n13230 , n13227 , n13229 );
not ( n13231 , n13230 );
not ( n13232 , n8581 );
nand ( n13233 , n7415 , n497 );
not ( n13234 , n13233 );
and ( n13235 , n13232 , n13234 );
nand ( n13236 , n7410 , n497 );
nor ( n13237 , n9167 , n13236 );
nor ( n13238 , n13235 , n13237 );
nand ( n13239 , n13231 , n13238 );
xor ( n13240 , n13223 , n13239 );
xor ( n13241 , n9072 , n9078 );
and ( n13242 , n13241 , n9089 );
and ( n13243 , n9072 , n9078 );
or ( n13244 , n13242 , n13243 );
not ( n13245 , n9066 );
not ( n13246 , n7405 );
or ( n13247 , n13245 , n13246 );
not ( n13248 , n13119 );
or ( n13249 , n13248 , n7370 );
nand ( n13250 , n13247 , n13249 );
xor ( n13251 , n13244 , n13250 );
xor ( n13252 , n13100 , n13105 );
xor ( n13253 , n13252 , n13112 );
and ( n13254 , n13251 , n13253 );
and ( n13255 , n13244 , n13250 );
or ( n13256 , n13254 , n13255 );
and ( n13257 , n13240 , n13256 );
and ( n13258 , n13223 , n13239 );
or ( n13259 , n13257 , n13258 );
and ( n13260 , n13213 , n13259 );
and ( n13261 , n13210 , n13212 );
or ( n13262 , n13260 , n13261 );
xor ( n13263 , n13199 , n13262 );
or ( n13264 , n13172 , n8304 );
and ( n13265 , n12737 , n503 );
not ( n13266 , n12737 );
and ( n13267 , n13266 , n8880 );
or ( n13268 , n13265 , n13267 );
or ( n13269 , n13268 , n8303 );
nand ( n13270 , n13264 , n13269 );
and ( n13271 , n13263 , n13270 );
and ( n13272 , n13199 , n13262 );
or ( n13273 , n13271 , n13272 );
xor ( n13274 , n13195 , n13273 );
not ( n13275 , n13058 );
nand ( n13276 , n13275 , n7819 );
not ( n13277 , n13275 );
nand ( n13278 , n13277 , n7815 );
nand ( n13279 , n12923 , n7558 );
nand ( n13280 , n13276 , n13278 , n13279 );
xor ( n13281 , n12881 , n12882 );
and ( n13282 , n13281 , n12898 );
and ( n13283 , n12881 , n12882 );
or ( n13284 , n13282 , n13283 );
not ( n13285 , n7371 );
and ( n13286 , n493 , n9278 );
not ( n13287 , n493 );
and ( n13288 , n13287 , n8581 );
or ( n13289 , n13286 , n13288 );
not ( n13290 , n13289 );
or ( n13291 , n13285 , n13290 );
nand ( n13292 , n12965 , n7405 );
nand ( n13293 , n13291 , n13292 );
xor ( n13294 , n13284 , n13293 );
not ( n13295 , n6848 );
xor ( n13296 , n489 , n7301 );
not ( n13297 , n13296 );
or ( n13298 , n13295 , n13297 );
nand ( n13299 , n12876 , n6867 );
nand ( n13300 , n13298 , n13299 );
and ( n13301 , n489 , n7383 );
xor ( n13302 , n13300 , n13301 );
not ( n13303 , n6842 );
not ( n13304 , n491 );
not ( n13305 , n7678 );
or ( n13306 , n13304 , n13305 );
nand ( n13307 , n7677 , n6892 );
nand ( n13308 , n13306 , n13307 );
not ( n13309 , n13308 );
or ( n13310 , n13303 , n13309 );
nand ( n13311 , n12889 , n6719 );
nand ( n13312 , n13310 , n13311 );
xor ( n13313 , n13302 , n13312 );
xor ( n13314 , n13294 , n13313 );
xor ( n13315 , n13280 , n13314 );
not ( n13316 , n7828 );
not ( n13317 , n501 );
not ( n13318 , n13168 );
or ( n13319 , n13317 , n13318 );
nand ( n13320 , n13167 , n8260 );
nand ( n13321 , n13319 , n13320 );
not ( n13322 , n13321 );
or ( n13323 , n13316 , n13322 );
nand ( n13324 , n13086 , n8297 );
nand ( n13325 , n13323 , n13324 );
xor ( n13326 , n13315 , n13325 );
xor ( n13327 , n13274 , n13326 );
xor ( n13328 , n13191 , n13327 );
xor ( n13329 , n13199 , n13262 );
xor ( n13330 , n13329 , n13270 );
xor ( n13331 , n13115 , n13121 );
xor ( n13332 , n13331 , n13124 );
not ( n13333 , n7558 );
and ( n13334 , n499 , n8255 );
not ( n13335 , n499 );
and ( n13336 , n13335 , n8259 );
or ( n13337 , n13334 , n13336 );
not ( n13338 , n13337 );
or ( n13339 , n13333 , n13338 );
and ( n13340 , n499 , n8869 );
not ( n13341 , n499 );
and ( n13342 , n13341 , n8866 );
nor ( n13343 , n13340 , n13342 );
nand ( n13344 , n13343 , n7813 );
nand ( n13345 , n13339 , n13344 );
xor ( n13346 , n13332 , n13345 );
not ( n13347 , n501 );
not ( n13348 , n8795 );
or ( n13349 , n13347 , n13348 );
nand ( n13350 , n8792 , n8260 );
nand ( n13351 , n13349 , n13350 );
not ( n13352 , n13351 );
not ( n13353 , n8594 );
or ( n13354 , n13352 , n13353 );
nand ( n13355 , n13146 , n7828 );
nand ( n13356 , n13354 , n13355 );
and ( n13357 , n13346 , n13356 );
and ( n13358 , n13332 , n13345 );
or ( n13359 , n13357 , n13358 );
xor ( n13360 , n13210 , n13212 );
xor ( n13361 , n13360 , n13259 );
xor ( n13362 , n13359 , n13361 );
xor ( n13363 , n9064 , n9070 );
and ( n13364 , n13363 , n9090 );
and ( n13365 , n9064 , n9070 );
or ( n13366 , n13364 , n13365 );
not ( n13367 , n6939 );
not ( n13368 , n13220 );
not ( n13369 , n13368 );
or ( n13370 , n13367 , n13369 );
nand ( n13371 , n8847 , n7326 );
nand ( n13372 , n13370 , n13371 );
xor ( n13373 , n13366 , n13372 );
not ( n13374 , n7517 );
and ( n13375 , n497 , n9278 );
not ( n13376 , n497 );
and ( n13377 , n13376 , n8581 );
or ( n13378 , n13375 , n13377 );
not ( n13379 , n13378 );
or ( n13380 , n13374 , n13379 );
nand ( n13381 , n7415 , n8860 );
nand ( n13382 , n13380 , n13381 );
and ( n13383 , n13373 , n13382 );
and ( n13384 , n13366 , n13372 );
or ( n13385 , n13383 , n13384 );
xor ( n13386 , n13223 , n13239 );
xor ( n13387 , n13386 , n13256 );
xor ( n13388 , n13385 , n13387 );
xor ( n13389 , n13244 , n13250 );
xor ( n13390 , n13389 , n13253 );
not ( n13391 , n7813 );
not ( n13392 , n13337 );
or ( n13393 , n13391 , n13392 );
nand ( n13394 , n9100 , n7558 );
nand ( n13395 , n13393 , n13394 );
xor ( n13396 , n13390 , n13395 );
xor ( n13397 , n8840 , n8851 );
and ( n13398 , n13397 , n8862 );
and ( n13399 , n8840 , n8851 );
or ( n13400 , n13398 , n13399 );
and ( n13401 , n13396 , n13400 );
and ( n13402 , n13390 , n13395 );
or ( n13403 , n13401 , n13402 );
and ( n13404 , n13388 , n13403 );
and ( n13405 , n13385 , n13387 );
or ( n13406 , n13404 , n13405 );
and ( n13407 , n13362 , n13406 );
and ( n13408 , n13359 , n13361 );
or ( n13409 , n13407 , n13408 );
xor ( n13410 , n13330 , n13409 );
xor ( n13411 , n13003 , n13089 );
xor ( n13412 , n13411 , n13187 );
and ( n13413 , n13410 , n13412 );
and ( n13414 , n13330 , n13409 );
or ( n13415 , n13413 , n13414 );
or ( n13416 , n13328 , n13415 );
not ( n13417 , n13416 );
not ( n13418 , n7405 );
not ( n13419 , n13289 );
or ( n13420 , n13418 , n13419 );
and ( n13421 , n493 , n8282 );
not ( n13422 , n493 );
and ( n13423 , n13422 , n9167 );
or ( n13424 , n13421 , n13423 );
nand ( n13425 , n13424 , n7371 );
nand ( n13426 , n13420 , n13425 );
xor ( n13427 , n13300 , n13301 );
and ( n13428 , n13427 , n13312 );
and ( n13429 , n13300 , n13301 );
or ( n13430 , n13428 , n13429 );
xor ( n13431 , n13426 , n13430 );
not ( n13432 , n7326 );
not ( n13433 , n12941 );
or ( n13434 , n13432 , n13433 );
and ( n13435 , n495 , n8479 );
not ( n13436 , n495 );
and ( n13437 , n13436 , n8475 );
or ( n13438 , n13435 , n13437 );
nand ( n13439 , n13438 , n6939 );
nand ( n13440 , n13434 , n13439 );
xor ( n13441 , n13431 , n13440 );
xor ( n13442 , n12943 , n12953 );
and ( n13443 , n13442 , n12999 );
and ( n13444 , n12943 , n12953 );
or ( n13445 , n13443 , n13444 );
xor ( n13446 , n13441 , n13445 );
not ( n13447 , n7415 );
not ( n13448 , n12948 );
or ( n13449 , n13447 , n13448 );
and ( n13450 , n497 , n9049 );
not ( n13451 , n497 );
and ( n13452 , n13451 , n9050 );
nor ( n13453 , n13450 , n13452 );
nand ( n13454 , n13453 , n7517 );
nand ( n13455 , n13449 , n13454 );
and ( n13456 , n491 , n8589 );
not ( n13457 , n491 );
and ( n13458 , n13457 , n7812 );
nor ( n13459 , n13456 , n13458 );
not ( n13460 , n13459 );
not ( n13461 , n6843 );
and ( n13462 , n13460 , n13461 );
and ( n13463 , n13308 , n6719 );
nor ( n13464 , n13462 , n13463 );
not ( n13465 , n6848 );
not ( n13466 , n489 );
not ( n13467 , n8843 );
or ( n13468 , n13466 , n13467 );
nand ( n13469 , n7511 , n4046 );
nand ( n13470 , n13468 , n13469 );
not ( n13471 , n13470 );
or ( n13472 , n13465 , n13471 );
nand ( n13473 , n13296 , n6867 );
nand ( n13474 , n13472 , n13473 );
nand ( n13475 , n7321 , n489 );
xor ( n13476 , n13474 , n13475 );
xor ( n13477 , n13464 , n13476 );
xor ( n13478 , n13455 , n13477 );
not ( n13479 , n7558 );
and ( n13480 , n499 , n13277 );
not ( n13481 , n499 );
and ( n13482 , n13481 , n13063 );
nor ( n13483 , n13480 , n13482 );
not ( n13484 , n13483 );
or ( n13485 , n13479 , n13484 );
and ( n13486 , n499 , n13179 );
not ( n13487 , n499 );
and ( n13488 , n13487 , n13084 );
or ( n13489 , n13486 , n13488 );
nand ( n13490 , n13489 , n7813 );
nand ( n13491 , n13485 , n13490 );
xor ( n13492 , n13478 , n13491 );
xor ( n13493 , n13446 , n13492 );
xor ( n13494 , n13195 , n13273 );
and ( n13495 , n13494 , n13326 );
and ( n13496 , n13195 , n13273 );
or ( n13497 , n13495 , n13496 );
xor ( n13498 , n13493 , n13497 );
xor ( n13499 , n13280 , n13314 );
and ( n13500 , n13499 , n13325 );
and ( n13501 , n13280 , n13314 );
or ( n13502 , n13500 , n13501 );
xor ( n13503 , n12870 , n12929 );
and ( n13504 , n13503 , n13000 );
and ( n13505 , n12870 , n12929 );
or ( n13506 , n13504 , n13505 );
xor ( n13507 , n13502 , n13506 );
xor ( n13508 , n13284 , n13293 );
and ( n13509 , n13508 , n13313 );
and ( n13510 , n13284 , n13293 );
or ( n13511 , n13509 , n13510 );
not ( n13512 , n7828 );
not ( n13513 , n501 );
not ( n13514 , n12737 );
not ( n13515 , n13514 );
or ( n13516 , n13513 , n13515 );
nand ( n13517 , n12737 , n8260 );
nand ( n13518 , n13516 , n13517 );
not ( n13519 , n13518 );
or ( n13520 , n13512 , n13519 );
nand ( n13521 , n13321 , n8594 );
nand ( n13522 , n13520 , n13521 );
xor ( n13523 , n13511 , n13522 );
not ( n13524 , n8306 );
not ( n13525 , n12866 );
or ( n13526 , n13524 , n13525 );
not ( n13527 , n12851 );
nor ( n13528 , n13527 , n12728 );
buf ( n13529 , n13528 );
nand ( n13530 , n12586 , n13529 );
not ( n13531 , n13530 );
not ( n13532 , n13531 );
not ( n13533 , n12601 );
or ( n13534 , n13532 , n13533 );
not ( n13535 , n12628 );
and ( n13536 , n13535 , n13529 );
not ( n13537 , n12851 );
or ( n13538 , n12730 , n13537 );
nand ( n13539 , n13538 , n12849 );
not ( n13540 , n13539 );
not ( n13541 , n13540 );
nor ( n13542 , n13536 , n13541 );
nand ( n13543 , n13534 , n13542 );
not ( n13544 , n13543 );
and ( n13545 , n12750 , n12606 );
nor ( n13546 , n13545 , n13530 );
not ( n13547 , n13546 );
not ( n13548 , n12758 );
not ( n13549 , n12825 );
or ( n13550 , n13548 , n13549 );
nand ( n13551 , n13550 , n12838 );
not ( n13552 , n12825 );
nand ( n13553 , n13552 , n12757 );
nand ( n13554 , n13551 , n13553 );
not ( n13555 , n13554 );
not ( n13556 , n12708 );
not ( n13557 , n12791 );
or ( n13558 , n13556 , n13557 );
not ( n13559 , n12711 );
not ( n13560 , n12788 );
or ( n13561 , n13559 , n13560 );
nand ( n13562 , n13561 , n12766 );
nand ( n13563 , n13558 , n13562 );
not ( n13564 , n13563 );
and ( n13565 , n528 , n457 );
not ( n13566 , n12778 );
not ( n13567 , n8337 );
or ( n13568 , n13566 , n13567 );
xor ( n13569 , n457 , n526 );
nand ( n13570 , n7908 , n13569 );
nand ( n13571 , n13568 , n13570 );
xor ( n13572 , n13565 , n13571 );
not ( n13573 , n12803 );
not ( n13574 , n8327 );
or ( n13575 , n13573 , n13574 );
nand ( n13576 , n7026 , n463 );
nand ( n13577 , n13575 , n13576 );
xor ( n13578 , n13572 , n13577 );
xor ( n13579 , n12805 , n12811 );
and ( n13580 , n13579 , n12814 );
and ( n13581 , n12805 , n12811 );
or ( n13582 , n13580 , n13581 );
xor ( n13583 , n13578 , n13582 );
not ( n13584 , n12774 );
not ( n13585 , n12780 );
or ( n13586 , n13584 , n13585 );
not ( n13587 , n12773 );
not ( n13588 , n12780 );
not ( n13589 , n13588 );
or ( n13590 , n13587 , n13589 );
nand ( n13591 , n13590 , n12787 );
nand ( n13592 , n13586 , n13591 );
not ( n13593 , n12785 );
not ( n13594 , n7585 );
or ( n13595 , n13593 , n13594 );
xor ( n13596 , n461 , n522 );
nand ( n13597 , n7475 , n13596 );
nand ( n13598 , n13595 , n13597 );
not ( n13599 , n13598 );
not ( n13600 , n12809 );
not ( n13601 , n7881 );
or ( n13602 , n13600 , n13601 );
xor ( n13603 , n459 , n524 );
nand ( n13604 , n7888 , n13603 );
nand ( n13605 , n13602 , n13604 );
not ( n13606 , n13605 );
and ( n13607 , n13599 , n13606 );
and ( n13608 , n13598 , n13605 );
nor ( n13609 , n13607 , n13608 );
not ( n13610 , n13609 );
and ( n13611 , n13592 , n13610 );
not ( n13612 , n13592 );
and ( n13613 , n13612 , n13609 );
nor ( n13614 , n13611 , n13613 );
xor ( n13615 , n13583 , n13614 );
xor ( n13616 , n13564 , n13615 );
nand ( n13617 , n12818 , n12799 );
not ( n13618 , n13617 );
not ( n13619 , n12793 );
or ( n13620 , n13618 , n13619 );
not ( n13621 , n12799 );
nand ( n13622 , n13621 , n12815 );
nand ( n13623 , n13620 , n13622 );
xor ( n13624 , n13616 , n13623 );
nand ( n13625 , n13555 , n13624 );
not ( n13626 , n13624 );
nand ( n13627 , n13626 , n13554 );
nand ( n13628 , n13625 , n13627 );
not ( n13629 , n13628 );
nand ( n13630 , n13544 , n13547 , n13629 );
or ( n13631 , n13543 , n13546 );
nand ( n13632 , n13631 , n13628 );
nand ( n13633 , n13630 , n13632 );
buf ( n13634 , n13633 );
and ( n13635 , n13634 , n8880 );
not ( n13636 , n13634 );
and ( n13637 , n13636 , n503 );
or ( n13638 , n13635 , n13637 );
nand ( n13639 , n13638 , n504 );
nand ( n13640 , n13526 , n13639 );
xor ( n13641 , n13523 , n13640 );
xor ( n13642 , n13507 , n13641 );
xor ( n13643 , n13498 , n13642 );
not ( n13644 , n13643 );
xor ( n13645 , n13001 , n13190 );
and ( n13646 , n13645 , n13327 );
and ( n13647 , n13001 , n13190 );
or ( n13648 , n13646 , n13647 );
not ( n13649 , n13648 );
nand ( n13650 , n13644 , n13649 );
not ( n13651 , n13650 );
nor ( n13652 , n13417 , n13651 );
not ( n13653 , n13652 );
not ( n13654 , n8306 );
and ( n13655 , n503 , n13060 );
not ( n13656 , n503 );
and ( n13657 , n13656 , n13275 );
nor ( n13658 , n13655 , n13657 );
not ( n13659 , n13658 );
or ( n13660 , n13654 , n13659 );
nand ( n13661 , n13182 , n504 );
nand ( n13662 , n13660 , n13661 );
xor ( n13663 , n9091 , n9102 );
and ( n13664 , n13663 , n9107 );
and ( n13665 , n9091 , n9102 );
or ( n13666 , n13664 , n13665 );
xor ( n13667 , n13366 , n13372 );
xor ( n13668 , n13667 , n13382 );
xor ( n13669 , n13666 , n13668 );
not ( n13670 , n8871 );
not ( n13671 , n8297 );
or ( n13672 , n13670 , n13671 );
not ( n13673 , n13351 );
not ( n13674 , n7828 );
or ( n13675 , n13673 , n13674 );
nand ( n13676 , n13672 , n13675 );
and ( n13677 , n13669 , n13676 );
and ( n13678 , n13666 , n13668 );
or ( n13679 , n13677 , n13678 );
xor ( n13680 , n13662 , n13679 );
xor ( n13681 , n13332 , n13345 );
xor ( n13682 , n13681 , n13356 );
and ( n13683 , n13680 , n13682 );
and ( n13684 , n13662 , n13679 );
or ( n13685 , n13683 , n13684 );
xor ( n13686 , n13138 , n13148 );
xor ( n13687 , n13686 , n13184 );
xor ( n13688 , n13685 , n13687 );
xor ( n13689 , n13359 , n13361 );
xor ( n13690 , n13689 , n13406 );
and ( n13691 , n13688 , n13690 );
and ( n13692 , n13685 , n13687 );
or ( n13693 , n13691 , n13692 );
not ( n13694 , n13693 );
xor ( n13695 , n13330 , n13409 );
xor ( n13696 , n13695 , n13412 );
not ( n13697 , n13696 );
and ( n13698 , n13694 , n13697 );
xor ( n13699 , n13685 , n13687 );
xor ( n13700 , n13699 , n13690 );
xor ( n13701 , n13385 , n13387 );
xor ( n13702 , n13701 , n13403 );
not ( n13703 , n504 );
not ( n13704 , n13658 );
or ( n13705 , n13703 , n13704 );
not ( n13706 , n9052 );
nand ( n13707 , n13706 , n8306 );
nand ( n13708 , n13705 , n13707 );
xor ( n13709 , n13390 , n13395 );
xor ( n13710 , n13709 , n13400 );
xor ( n13711 , n13708 , n13710 );
xor ( n13712 , n8863 , n8875 );
and ( n13713 , n13712 , n9054 );
and ( n13714 , n8863 , n8875 );
or ( n13715 , n13713 , n13714 );
and ( n13716 , n13711 , n13715 );
and ( n13717 , n13708 , n13710 );
or ( n13718 , n13716 , n13717 );
xor ( n13719 , n13702 , n13718 );
xor ( n13720 , n13662 , n13679 );
xor ( n13721 , n13720 , n13682 );
and ( n13722 , n13719 , n13721 );
and ( n13723 , n13702 , n13718 );
or ( n13724 , n13722 , n13723 );
nor ( n13725 , n13700 , n13724 );
nor ( n13726 , n13698 , n13725 );
not ( n13727 , n13726 );
xor ( n13728 , n13702 , n13718 );
xor ( n13729 , n13728 , n13721 );
xor ( n13730 , n13666 , n13668 );
xor ( n13731 , n13730 , n13676 );
xor ( n13732 , n9060 , n9108 );
and ( n13733 , n13732 , n9113 );
and ( n13734 , n9060 , n9108 );
or ( n13735 , n13733 , n13734 );
xor ( n13736 , n13731 , n13735 );
xor ( n13737 , n13708 , n13710 );
xor ( n13738 , n13737 , n13715 );
and ( n13739 , n13736 , n13738 );
and ( n13740 , n13731 , n13735 );
or ( n13741 , n13739 , n13740 );
nor ( n13742 , n13729 , n13741 );
xor ( n13743 , n13731 , n13735 );
xor ( n13744 , n13743 , n13738 );
xor ( n13745 , n8836 , n9055 );
and ( n13746 , n13745 , n9114 );
and ( n13747 , n8836 , n9055 );
or ( n13748 , n13746 , n13747 );
nor ( n13749 , n13744 , n13748 );
nor ( n13750 , n13742 , n13749 );
not ( n13751 , n13750 );
xor ( n13752 , n8832 , n9115 );
and ( n13753 , n13752 , n9905 );
and ( n13754 , n8832 , n9115 );
or ( n13755 , n13753 , n13754 );
not ( n13756 , n13755 );
or ( n13757 , n13751 , n13756 );
not ( n13758 , n13742 );
and ( n13759 , n13744 , n13748 );
and ( n13760 , n13758 , n13759 );
and ( n13761 , n13729 , n13741 );
nor ( n13762 , n13760 , n13761 );
nand ( n13763 , n13757 , n13762 );
not ( n13764 , n13763 );
or ( n13765 , n13727 , n13764 );
and ( n13766 , n13700 , n13724 );
not ( n13767 , n13766 );
not ( n13768 , n13693 );
not ( n13769 , n13696 );
nand ( n13770 , n13768 , n13769 );
not ( n13771 , n13770 );
or ( n13772 , n13767 , n13771 );
not ( n13773 , n13769 );
nand ( n13774 , n13773 , n13693 );
nand ( n13775 , n13772 , n13774 );
not ( n13776 , n13775 );
nand ( n13777 , n13765 , n13776 );
not ( n13778 , n13777 );
or ( n13779 , n13653 , n13778 );
and ( n13780 , n13328 , n13415 );
not ( n13781 , n13780 );
not ( n13782 , n13650 );
or ( n13783 , n13781 , n13782 );
buf ( n13784 , n13643 );
nand ( n13785 , n13784 , n13648 );
nand ( n13786 , n13783 , n13785 );
not ( n13787 , n13786 );
nand ( n13788 , n13779 , n13787 );
not ( n13789 , n504 );
not ( n13790 , n503 );
xor ( n13791 , n13578 , n13582 );
and ( n13792 , n13791 , n13614 );
and ( n13793 , n13578 , n13582 );
or ( n13794 , n13792 , n13793 );
not ( n13795 , n13794 );
and ( n13796 , n527 , n457 );
xor ( n13797 , n13796 , n13598 );
not ( n13798 , n13603 );
not ( n13799 , n7881 );
or ( n13800 , n13798 , n13799 );
xor ( n13801 , n523 , n459 );
nand ( n13802 , n7888 , n13801 );
nand ( n13803 , n13800 , n13802 );
xor ( n13804 , n13797 , n13803 );
not ( n13805 , n13605 );
nand ( n13806 , n13805 , n13598 );
not ( n13807 , n13806 );
not ( n13808 , n13592 );
or ( n13809 , n13807 , n13808 );
not ( n13810 , n13598 );
nand ( n13811 , n13810 , n13605 );
nand ( n13812 , n13809 , n13811 );
xor ( n13813 , n13804 , n13812 );
xor ( n13814 , n13565 , n13571 );
and ( n13815 , n13814 , n13577 );
and ( n13816 , n13565 , n13571 );
or ( n13817 , n13815 , n13816 );
not ( n13818 , n13569 );
not ( n13819 , n8337 );
or ( n13820 , n13818 , n13819 );
xor ( n13821 , n457 , n525 );
nand ( n13822 , n7908 , n13821 );
nand ( n13823 , n13820 , n13822 );
not ( n13824 , n13596 );
not ( n13825 , n8719 );
or ( n13826 , n13824 , n13825 );
xor ( n13827 , n521 , n461 );
nand ( n13828 , n7475 , n13827 );
nand ( n13829 , n13826 , n13828 );
xor ( n13830 , n13823 , n13829 );
not ( n13831 , n7026 );
not ( n13832 , n13831 );
not ( n13833 , n12314 );
or ( n13834 , n13832 , n13833 );
nand ( n13835 , n13834 , n463 );
xor ( n13836 , n13830 , n13835 );
xnor ( n13837 , n13817 , n13836 );
xor ( n13838 , n13813 , n13837 );
or ( n13839 , n13795 , n13838 );
nand ( n13840 , n13838 , n13795 );
nand ( n13841 , n13839 , n13840 );
not ( n13842 , n13615 );
nand ( n13843 , n13842 , n13564 );
nand ( n13844 , n13843 , n13623 );
nand ( n13845 , n13615 , n13563 );
and ( n13846 , n13844 , n13845 );
nor ( n13847 , n13841 , n13846 );
not ( n13848 , n13847 );
nand ( n13849 , n13841 , n13846 );
nand ( n13850 , n13848 , n13849 );
not ( n13851 , n13850 );
not ( n13852 , n13851 );
nand ( n13853 , n12616 , n12587 );
and ( n13854 , n13529 , n13625 );
not ( n13855 , n13854 );
or ( n13856 , n13853 , n13855 );
and ( n13857 , n13854 , n13535 );
not ( n13858 , n13625 );
not ( n13859 , n13539 );
or ( n13860 , n13858 , n13859 );
nand ( n13861 , n13860 , n13627 );
nor ( n13862 , n13857 , n13861 );
nand ( n13863 , n13856 , n13862 );
not ( n13864 , n13863 );
not ( n13865 , n13864 );
or ( n13866 , n13852 , n13865 );
nand ( n13867 , n13863 , n13850 );
nand ( n13868 , n13866 , n13867 );
not ( n13869 , n13868 );
not ( n13870 , n13869 );
or ( n13871 , n13790 , n13870 );
buf ( n13872 , n13868 );
nand ( n13873 , n13872 , n8880 );
nand ( n13874 , n13871 , n13873 );
not ( n13875 , n13874 );
or ( n13876 , n13789 , n13875 );
nand ( n13877 , n13638 , n8306 );
nand ( n13878 , n13876 , n13877 );
xor ( n13879 , n13455 , n13477 );
and ( n13880 , n13879 , n13491 );
and ( n13881 , n13455 , n13477 );
or ( n13882 , n13880 , n13881 );
xor ( n13883 , n13878 , n13882 );
xor ( n13884 , n13511 , n13522 );
and ( n13885 , n13884 , n13640 );
and ( n13886 , n13511 , n13522 );
or ( n13887 , n13885 , n13886 );
xor ( n13888 , n13883 , n13887 );
xor ( n13889 , n13502 , n13506 );
and ( n13890 , n13889 , n13641 );
and ( n13891 , n13502 , n13506 );
or ( n13892 , n13890 , n13891 );
xor ( n13893 , n13888 , n13892 );
not ( n13894 , n13475 );
and ( n13895 , n13474 , n13894 );
not ( n13896 , n6842 );
and ( n13897 , n8581 , n6892 );
not ( n13898 , n8581 );
and ( n13899 , n13898 , n491 );
or ( n13900 , n13897 , n13899 );
not ( n13901 , n13900 );
or ( n13902 , n13896 , n13901 );
not ( n13903 , n13459 );
nand ( n13904 , n13903 , n6719 );
nand ( n13905 , n13902 , n13904 );
xor ( n13906 , n13895 , n13905 );
and ( n13907 , n489 , n7301 );
not ( n13908 , n6848 );
not ( n13909 , n489 );
not ( n13910 , n7678 );
or ( n13911 , n13909 , n13910 );
nand ( n13912 , n7677 , n4046 );
nand ( n13913 , n13911 , n13912 );
not ( n13914 , n13913 );
or ( n13915 , n13908 , n13914 );
nand ( n13916 , n13470 , n6867 );
nand ( n13917 , n13915 , n13916 );
xor ( n13918 , n13907 , n13917 );
xor ( n13919 , n13906 , n13918 );
not ( n13920 , n7517 );
and ( n13921 , n497 , n13058 );
not ( n13922 , n497 );
and ( n13923 , n13922 , n13275 );
nor ( n13924 , n13921 , n13923 );
not ( n13925 , n13924 );
or ( n13926 , n13920 , n13925 );
nand ( n13927 , n13453 , n7415 );
nand ( n13928 , n13926 , n13927 );
xor ( n13929 , n13919 , n13928 );
xor ( n13930 , n13426 , n13430 );
and ( n13931 , n13930 , n13440 );
and ( n13932 , n13426 , n13430 );
or ( n13933 , n13931 , n13932 );
xor ( n13934 , n13929 , n13933 );
nor ( n13935 , n13464 , n13476 );
not ( n13936 , n7371 );
and ( n13937 , n493 , n8255 );
not ( n13938 , n493 );
and ( n13939 , n13938 , n12900 );
or ( n13940 , n13937 , n13939 );
not ( n13941 , n13940 );
or ( n13942 , n13936 , n13941 );
nand ( n13943 , n13424 , n7405 );
nand ( n13944 , n13942 , n13943 );
xor ( n13945 , n13935 , n13944 );
not ( n13946 , n6939 );
and ( n13947 , n495 , n8795 );
not ( n13948 , n495 );
and ( n13949 , n13948 , n8792 );
or ( n13950 , n13947 , n13949 );
not ( n13951 , n13950 );
or ( n13952 , n13946 , n13951 );
nand ( n13953 , n13438 , n7326 );
nand ( n13954 , n13952 , n13953 );
xor ( n13955 , n13945 , n13954 );
not ( n13956 , n7828 );
not ( n13957 , n12865 );
and ( n13958 , n501 , n13957 );
not ( n13959 , n501 );
and ( n13960 , n13959 , n12868 );
or ( n13961 , n13958 , n13960 );
not ( n13962 , n13961 );
or ( n13963 , n13956 , n13962 );
nand ( n13964 , n13518 , n8297 );
nand ( n13965 , n13963 , n13964 );
xor ( n13966 , n13955 , n13965 );
not ( n13967 , n7813 );
not ( n13968 , n13167 );
and ( n13969 , n499 , n13968 );
not ( n13970 , n499 );
not ( n13971 , n13968 );
and ( n13972 , n13970 , n13971 );
or ( n13973 , n13969 , n13972 );
not ( n13974 , n13973 );
or ( n13975 , n13967 , n13974 );
nand ( n13976 , n13489 , n7558 );
nand ( n13977 , n13975 , n13976 );
xor ( n13978 , n13966 , n13977 );
xor ( n13979 , n13934 , n13978 );
xor ( n13980 , n13441 , n13445 );
and ( n13981 , n13980 , n13492 );
and ( n13982 , n13441 , n13445 );
or ( n13983 , n13981 , n13982 );
xor ( n13984 , n13979 , n13983 );
xor ( n13985 , n13893 , n13984 );
xor ( n13986 , n13493 , n13497 );
and ( n13987 , n13986 , n13642 );
and ( n13988 , n13493 , n13497 );
or ( n13989 , n13987 , n13988 );
or ( n13990 , n13985 , n13989 );
and ( n13991 , n13985 , n13989 );
not ( n13992 , n13991 );
nand ( n13993 , n13990 , n13992 );
xnor ( n13994 , n13788 , n13993 );
nand ( n13995 , n13994 , n9907 );
nand ( n13996 , n12212 , n13995 );
not ( n13997 , n6598 );
nand ( n13998 , n6548 , n6601 );
not ( n13999 , n13998 );
or ( n14000 , n13997 , n13999 );
or ( n14001 , n13998 , n6598 );
nand ( n14002 , n14000 , n14001 );
nand ( n14003 , n454 , n14002 );
not ( n14004 , n9798 );
or ( n14005 , n9735 , n9743 );
nand ( n14006 , n14005 , n9800 );
not ( n14007 , n14006 );
or ( n14008 , n14004 , n14007 );
or ( n14009 , n14006 , n9798 );
nand ( n14010 , n14008 , n14009 );
nand ( n14011 , n14010 , n9907 );
nand ( n14012 , n14003 , n14011 );
not ( n14013 , n454 );
not ( n14014 , n11367 );
not ( n14015 , n10741 );
or ( n14016 , n14014 , n14015 );
not ( n14017 , n11933 );
nand ( n14018 , n14016 , n14017 );
buf ( n14019 , n11939 );
buf ( n14020 , n11663 );
nand ( n14021 , n14019 , n14020 );
xnor ( n14022 , n14018 , n14021 );
not ( n14023 , n14022 );
or ( n14024 , n14013 , n14023 );
not ( n14025 , n13780 );
nand ( n14026 , n13416 , n14025 );
xnor ( n14027 , n14026 , n13777 );
nand ( n14028 , n14027 , n9907 );
nand ( n14029 , n14024 , n14028 );
buf ( n14030 , n13755 );
not ( n14031 , n13749 );
not ( n14032 , n13759 );
nand ( n14033 , n14031 , n14032 );
xnor ( n14034 , n14030 , n14033 );
nand ( n14035 , n14034 , n9907 );
nand ( n14036 , n6509 , n6605 );
xnor ( n121587 , n6602 , n14036 );
nand ( n14037 , n121587 , n454 );
not ( n14038 , n9884 );
not ( n14039 , n9889 );
nand ( n14040 , n14038 , n14039 );
xnor ( n14041 , n14040 , n9861 );
nand ( n14042 , n14041 , n9907 );
xor ( n14043 , n9687 , n9689 );
xor ( n14044 , n14043 , n9807 );
nand ( n14045 , n14044 , n9907 );
or ( n14046 , n3300 , n3298 );
nand ( n14047 , n14046 , n547 );
and ( n14048 , n537 , n5578 );
xor ( n14049 , n14047 , n14048 );
and ( n14050 , n5614 , n537 );
xor ( n14051 , n14049 , n14050 );
not ( n14052 , n3300 );
not ( n14053 , n547 );
or ( n14054 , n12134 , n11635 );
not ( n14055 , n12129 );
and ( n14056 , n12135 , n14055 );
xor ( n14057 , n12150 , n12156 );
and ( n14058 , n14057 , n12166 );
and ( n14059 , n12150 , n12156 );
or ( n14060 , n14058 , n14059 );
and ( n14061 , n507 , n489 );
not ( n14062 , n3711 );
not ( n14063 , n5487 );
not ( n14064 , n14063 );
or ( n14065 , n14062 , n14064 );
nand ( n14066 , n14065 , n491 );
xor ( n14067 , n14061 , n14066 );
or ( n14068 , n12158 , n12164 );
and ( n14069 , n489 , n11803 );
not ( n14070 , n489 );
and ( n14071 , n14070 , n505 );
nor ( n14072 , n14069 , n14071 );
or ( n14073 , n12160 , n14072 );
nand ( n14074 , n14068 , n14073 );
xor ( n14075 , n14067 , n14074 );
xor ( n14076 , n14060 , n14075 );
not ( n14077 , n12156 );
xor ( n14078 , n14076 , n14077 );
xor ( n14079 , n12149 , n12167 );
and ( n14080 , n14079 , n12175 );
and ( n14081 , n12149 , n12167 );
or ( n14082 , n14080 , n14081 );
nor ( n14083 , n14078 , n14082 );
not ( n14084 , n14083 );
xor ( n14085 , n14060 , n14075 );
not ( n14086 , n12156 );
and ( n14087 , n14085 , n14086 );
and ( n14088 , n14060 , n14075 );
or ( n14089 , n14087 , n14088 );
or ( n14090 , n12158 , n14072 );
or ( n14091 , n12160 , n4046 );
nand ( n14092 , n14090 , n14091 );
nand ( n14093 , n506 , n489 );
xor ( n14094 , n14092 , n14093 );
xor ( n14095 , n14061 , n14066 );
and ( n14096 , n14095 , n14074 );
and ( n14097 , n14061 , n14066 );
or ( n14098 , n14096 , n14097 );
xor ( n14099 , n14094 , n14098 );
or ( n14100 , n14089 , n14099 );
and ( n14101 , n12177 , n14084 , n14100 );
not ( n14102 , n14101 );
nor ( n14103 , n14056 , n14102 );
nand ( n14104 , n14054 , n14103 );
and ( n14105 , n5449 , n11614 );
nand ( n14106 , n14105 , n12129 , n14101 );
or ( n14107 , n12178 , n14083 );
nand ( n14108 , n14078 , n14082 );
nand ( n14109 , n14107 , n14108 );
and ( n14110 , n14109 , n14100 );
nand ( n14111 , n14089 , n14099 );
not ( n14112 , n14111 );
nor ( n14113 , n14110 , n14112 );
not ( n14114 , n14113 );
xor ( n14115 , n14092 , n14093 );
and ( n14116 , n14115 , n14098 );
and ( n14117 , n14092 , n14093 );
or ( n14118 , n14116 , n14117 );
not ( n14119 , n14118 );
not ( n14120 , n14093 );
nand ( n14121 , n505 , n489 );
not ( n14122 , n14121 );
or ( n14123 , n4835 , n4838 );
nand ( n14124 , n14123 , n489 );
not ( n14125 , n14124 );
or ( n14126 , n14122 , n14125 );
or ( n14127 , n14124 , n14121 );
nand ( n14128 , n14126 , n14127 );
not ( n14129 , n14128 );
or ( n14130 , n14120 , n14129 );
or ( n14131 , n14128 , n14093 );
nand ( n14132 , n14130 , n14131 );
not ( n14133 , n14132 );
and ( n14134 , n14119 , n14133 );
and ( n14135 , n14118 , n14132 );
nor ( n14136 , n14134 , n14135 );
not ( n14137 , n14136 );
nor ( n14138 , n14114 , n14137 );
nand ( n14139 , n14104 , n14106 , n14138 );
nand ( n14140 , n14106 , n14104 , n14113 );
nand ( n14141 , n14140 , n14137 );
nand ( n14142 , n14139 , n14141 , n455 );
xor ( n14143 , n12079 , n12094 );
and ( n14144 , n14143 , n12099 );
and ( n14145 , n12079 , n12094 );
or ( n14146 , n14144 , n14145 );
not ( n14147 , n12093 );
not ( n14148 , n2200 );
not ( n14149 , n3572 );
or ( n14150 , n14148 , n14149 );
nand ( n14151 , n14150 , n491 );
not ( n14152 , n4056 );
not ( n14153 , n12084 );
or ( n14154 , n14152 , n14153 );
xor ( n14155 , n489 , n4076 );
nand ( n14156 , n14155 , n4547 );
nand ( n14157 , n14154 , n14156 );
xor ( n14158 , n14151 , n14157 );
and ( n14159 , n489 , n4093 );
xor ( n14160 , n14158 , n14159 );
xor ( n14161 , n14147 , n14160 );
xor ( n14162 , n12088 , n12089 );
and ( n14163 , n14162 , n12093 );
and ( n14164 , n12088 , n12089 );
or ( n14165 , n14163 , n14164 );
xor ( n14166 , n14161 , n14165 );
or ( n14167 , n14146 , n14166 );
not ( n14168 , n14167 );
xor ( n14169 , n14147 , n14160 );
and ( n14170 , n14169 , n14165 );
and ( n14171 , n14147 , n14160 );
or ( n14172 , n14170 , n14171 );
and ( n14173 , n14155 , n4553 );
and ( n14174 , n4547 , n489 );
nor ( n14175 , n14173 , n14174 );
not ( n14176 , n14175 );
and ( n14177 , n456 , n474 );
not ( n14178 , n456 );
and ( n14179 , n14178 , n458 );
or ( n14180 , n14177 , n14179 );
nand ( n14181 , n14180 , n489 );
xor ( n14182 , n14176 , n14181 );
xor ( n14183 , n14151 , n14157 );
and ( n14184 , n14183 , n14159 );
and ( n14185 , n14151 , n14157 );
or ( n14186 , n14184 , n14185 );
xor ( n14187 , n14182 , n14186 );
nor ( n14188 , n14172 , n14187 );
nor ( n14189 , n14168 , n14188 );
not ( n14190 , n14189 );
not ( n14191 , n10751 );
nor ( n14192 , n14191 , n11536 );
or ( n14193 , n11492 , n11530 );
nand ( n14194 , n12075 , n12101 );
nand ( n14195 , n14193 , n12067 , n14194 );
not ( n14196 , n14195 );
and ( n14197 , n14192 , n10456 , n14196 );
not ( n14198 , n14197 );
not ( n14199 , n5599 );
or ( n14200 , n14198 , n14199 );
not ( n14201 , n14192 );
not ( n14202 , n11144 );
or ( n14203 , n14201 , n14202 );
nand ( n14204 , n14203 , n11554 );
and ( n14205 , n14204 , n14196 );
and ( n14206 , n12114 , n12102 );
nor ( n14207 , n14206 , n12105 );
not ( n14208 , n14207 );
nor ( n14209 , n14205 , n14208 );
nand ( n14210 , n14200 , n14209 );
not ( n14211 , n14210 );
or ( n14212 , n14190 , n14211 );
nand ( n14213 , n14146 , n14166 );
not ( n14214 , n14213 );
not ( n14215 , n14188 );
and ( n14216 , n14214 , n14215 );
and ( n14217 , n14172 , n14187 );
nor ( n14218 , n14216 , n14217 );
nand ( n14219 , n14212 , n14218 );
xor ( n14220 , n14176 , n14181 );
and ( n14221 , n14220 , n14186 );
and ( n14222 , n14176 , n14181 );
or ( n14223 , n14221 , n14222 );
not ( n14224 , n14223 );
or ( n14225 , n4056 , n4547 );
nand ( n14226 , n14225 , n489 );
and ( n14227 , n489 , n4076 );
xor ( n14228 , n14226 , n14227 );
not ( n14229 , n14181 );
xor ( n14230 , n14228 , n14229 );
not ( n14231 , n14230 );
and ( n14232 , n14224 , n14231 );
and ( n14233 , n14223 , n14230 );
nor ( n14234 , n14232 , n14233 );
not ( n14235 , n14234 );
nor ( n14236 , n14235 , n455 );
and ( n14237 , n14219 , n14236 );
not ( n14238 , n14219 );
nor ( n14239 , n14234 , n455 );
and ( n14240 , n14238 , n14239 );
nor ( n14241 , n14237 , n14240 );
nand ( n14242 , n14142 , n14241 );
not ( n14243 , n14242 );
or ( n14244 , n14053 , n14243 );
nand ( n14245 , n14142 , n14241 );
not ( n14246 , n14245 );
nand ( n14247 , n14246 , n2369 );
nand ( n14248 , n14244 , n14247 );
not ( n14249 , n14248 );
or ( n14250 , n14052 , n14249 );
nand ( n14251 , n3298 , n547 );
nand ( n14252 , n14250 , n14251 );
not ( n14253 , n3955 );
not ( n14254 , n541 );
buf ( n14255 , n11640 );
not ( n14256 , n14255 );
not ( n14257 , n14256 );
or ( n14258 , n14254 , n14257 );
nand ( n14259 , n14255 , n3023 );
nand ( n14260 , n14258 , n14259 );
not ( n14261 , n14260 );
or ( n14262 , n14253 , n14261 );
not ( n14263 , n541 );
not ( n14264 , n11241 );
not ( n14265 , n14264 );
or ( n14266 , n14263 , n14265 );
nand ( n14267 , n11241 , n3023 );
nand ( n14268 , n14266 , n14267 );
nand ( n14269 , n14268 , n3288 );
nand ( n14270 , n14262 , n14269 );
xor ( n14271 , n14252 , n14270 );
not ( n14272 , n3017 );
not ( n14273 , n545 );
nand ( n14274 , n12129 , n12177 );
nor ( n14275 , n14274 , n14083 );
not ( n14276 , n14275 );
not ( n14277 , n11637 );
or ( n14278 , n14276 , n14277 );
not ( n14279 , n12177 );
not ( n14280 , n12134 );
or ( n14281 , n14279 , n14280 );
nand ( n14282 , n14281 , n12178 );
and ( n14283 , n14282 , n14084 );
not ( n14284 , n14108 );
nor ( n14285 , n14283 , n14284 );
nand ( n14286 , n14278 , n14285 );
nand ( n14287 , n14100 , n14111 );
and ( n14288 , n14286 , n14287 );
nor ( n14289 , n14288 , n5088 );
not ( n14290 , n14289 );
not ( n14291 , n14286 );
not ( n14292 , n14287 );
nand ( n14293 , n14291 , n14292 );
not ( n14294 , n14293 );
or ( n14295 , n14290 , n14294 );
not ( n14296 , n14213 );
nor ( n14297 , n14217 , n14188 , n14296 );
nor ( n14298 , n14297 , n14296 , n455 );
not ( n14299 , n14298 );
nand ( n14300 , n5599 , n14197 );
not ( n14301 , n14300 );
nor ( n14302 , n11545 , n14195 );
and ( n14303 , n11147 , n14302 );
not ( n14304 , n14196 );
not ( n14305 , n11553 );
or ( n14306 , n14304 , n14305 );
nand ( n14307 , n14306 , n14207 );
nor ( n14308 , n14303 , n14307 );
not ( n14309 , n14308 );
or ( n14310 , n14301 , n14309 );
nand ( n14311 , n14310 , n14167 );
not ( n14312 , n14311 );
or ( n14313 , n14299 , n14312 );
not ( n14314 , n455 );
xor ( n14315 , n14172 , n14187 );
nand ( n14316 , n14314 , n14315 );
or ( n14317 , n14297 , n14316 );
nand ( n14318 , n14313 , n14317 );
nor ( n14319 , n14311 , n14316 );
nor ( n14320 , n14318 , n14319 );
nand ( n14321 , n14295 , n14320 );
not ( n14322 , n14321 );
not ( n14323 , n14322 );
not ( n14324 , n14323 );
or ( n14325 , n14273 , n14324 );
not ( n14326 , n14323 );
nand ( n14327 , n14326 , n706 );
nand ( n14328 , n14325 , n14327 );
not ( n14329 , n14328 );
or ( n14330 , n14272 , n14329 );
not ( n14331 , n545 );
not ( n14332 , n716 );
nand ( n14333 , n14167 , n14213 );
xnor ( n14334 , n14210 , n14333 );
not ( n14335 , n14334 );
or ( n14336 , n14332 , n14335 );
not ( n14337 , n14274 );
not ( n14338 , n14337 );
not ( n14339 , n11637 );
or ( n14340 , n14338 , n14339 );
not ( n14341 , n14282 );
nand ( n14342 , n14340 , n14341 );
nand ( n14343 , n14084 , n14108 );
not ( n14344 , n14343 );
and ( n14345 , n14342 , n14344 );
not ( n14346 , n14342 );
and ( n14347 , n14346 , n14343 );
nor ( n14348 , n14345 , n14347 );
nand ( n14349 , n14348 , n455 );
nand ( n14350 , n14336 , n14349 );
not ( n14351 , n14350 );
not ( n14352 , n14351 );
or ( n14353 , n14331 , n14352 );
not ( n14354 , n14351 );
nand ( n14355 , n14354 , n706 );
nand ( n14356 , n14353 , n14355 );
nand ( n14357 , n14356 , n2376 );
nand ( n14358 , n14330 , n14357 );
and ( n14359 , n14271 , n14358 );
and ( n14360 , n14252 , n14270 );
or ( n14361 , n14359 , n14360 );
xor ( n14362 , n14051 , n14361 );
not ( n14363 , n3134 );
xor ( n14364 , n537 , n10438 );
not ( n14365 , n14364 );
or ( n14366 , n14363 , n14365 );
or ( n14367 , n10473 , n537 );
nand ( n14368 , n537 , n10473 );
nand ( n14369 , n14367 , n14368 );
nand ( n14370 , n14369 , n11729 );
nand ( n14371 , n14366 , n14370 );
not ( n14372 , n2376 );
not ( n14373 , n14328 );
or ( n14374 , n14372 , n14373 );
not ( n14375 , n545 );
not ( n14376 , n14246 );
not ( n14377 , n14376 );
or ( n14378 , n14375 , n14377 );
not ( n14379 , n14376 );
nand ( n14380 , n14379 , n706 );
nand ( n14381 , n14378 , n14380 );
nand ( n14382 , n14381 , n3017 );
nand ( n14383 , n14374 , n14382 );
xor ( n14384 , n14371 , n14383 );
not ( n14385 , n3955 );
not ( n14386 , n541 );
not ( n14387 , n11903 );
or ( n14388 , n14386 , n14387 );
nand ( n14389 , n11908 , n3023 );
nand ( n14390 , n14388 , n14389 );
not ( n14391 , n14390 );
or ( n14392 , n14385 , n14391 );
nand ( n14393 , n14260 , n3288 );
nand ( n14394 , n14392 , n14393 );
xor ( n14395 , n14384 , n14394 );
xor ( n14396 , n14362 , n14395 );
buf ( n14397 , n3026 );
not ( n14398 , n14397 );
not ( n14399 , n3069 );
not ( n14400 , n11241 );
or ( n14401 , n14399 , n14400 );
nand ( n14402 , n14264 , n539 );
nand ( n14403 , n14401 , n14402 );
not ( n14404 , n14403 );
or ( n14405 , n14398 , n14404 );
not ( n14406 , n539 );
not ( n14407 , n11478 );
not ( n14408 , n14407 );
or ( n14409 , n14406 , n14408 );
nand ( n14410 , n11478 , n3069 );
nand ( n14411 , n14409 , n14410 );
nand ( n14412 , n14411 , n3103 );
nand ( n14413 , n14405 , n14412 );
not ( n14414 , n714 );
not ( n14415 , n543 );
not ( n14416 , n12186 );
not ( n14417 , n14416 );
or ( n14418 , n14415 , n14417 );
not ( n14419 , n14416 );
nand ( n14420 , n14419 , n2123 );
nand ( n14421 , n14418 , n14420 );
not ( n14422 , n14421 );
or ( n14423 , n14414 , n14422 );
not ( n14424 , n543 );
not ( n14425 , n14351 );
or ( n14426 , n14424 , n14425 );
not ( n14427 , n14350 );
not ( n14428 , n14427 );
nand ( n14429 , n14428 , n2123 );
nand ( n14430 , n14426 , n14429 );
nand ( n14431 , n2362 , n14430 );
nand ( n14432 , n14423 , n14431 );
xor ( n14433 , n14413 , n14432 );
not ( n14434 , n11729 );
xor ( n14435 , n537 , n5578 );
not ( n14436 , n14435 );
or ( n14437 , n14434 , n14436 );
nand ( n14438 , n14369 , n3134 );
nand ( n14439 , n14437 , n14438 );
not ( n14440 , n3103 );
not ( n14441 , n539 );
not ( n14442 , n10439 );
or ( n14443 , n14441 , n14442 );
not ( n14444 , n11741 );
nand ( n14445 , n14444 , n3069 );
nand ( n14446 , n14443 , n14445 );
not ( n14447 , n14446 );
or ( n14448 , n14440 , n14447 );
nand ( n14449 , n14411 , n14397 );
nand ( n14450 , n14448 , n14449 );
xor ( n14451 , n14439 , n14450 );
not ( n14452 , n14050 );
and ( n14453 , n14451 , n14452 );
and ( n14454 , n14439 , n14450 );
or ( n14455 , n14453 , n14454 );
xor ( n14456 , n14433 , n14455 );
not ( n14457 , n2362 );
not ( n14458 , n14421 );
or ( n14459 , n14457 , n14458 );
not ( n14460 , n2123 );
not ( n14461 , n11908 );
or ( n14462 , n14460 , n14461 );
nand ( n14463 , n11903 , n543 );
nand ( n14464 , n14462 , n14463 );
nand ( n14465 , n14464 , n714 );
nand ( n14466 , n14459 , n14465 );
or ( n14467 , n4022 , n4020 );
nand ( n14468 , n14467 , n549 );
and ( n14469 , n5093 , n537 );
xor ( n14470 , n14468 , n14469 );
nand ( n14471 , n4638 , n537 );
not ( n14472 , n14471 );
and ( n14473 , n14470 , n14472 );
and ( n14474 , n14468 , n14469 );
or ( n14475 , n14473 , n14474 );
xor ( n14476 , n14466 , n14475 );
not ( n14477 , n3298 );
not ( n14478 , n14248 );
or ( n14479 , n14477 , n14478 );
not ( n14480 , n547 );
not ( n14481 , n14322 );
not ( n14482 , n14481 );
or ( n14483 , n14480 , n14482 );
nand ( n14484 , n2369 , n14322 );
nand ( n14485 , n14483 , n14484 );
nand ( n14486 , n14485 , n3300 );
nand ( n14487 , n14479 , n14486 );
not ( n14488 , n3955 );
not ( n14489 , n14268 );
or ( n14490 , n14488 , n14489 );
nand ( n14491 , n14407 , n541 );
not ( n14492 , n14491 );
not ( n14493 , n11475 );
nand ( n14494 , n14493 , n3023 );
not ( n14495 , n14494 );
or ( n14496 , n14492 , n14495 );
nand ( n14497 , n14496 , n3288 );
nand ( n14498 , n14490 , n14497 );
xor ( n14499 , n14487 , n14498 );
not ( n14500 , n2376 );
not ( n14501 , n706 );
not ( n14502 , n14419 );
or ( n14503 , n14501 , n14502 );
nand ( n14504 , n12187 , n545 );
nand ( n14505 , n14503 , n14504 );
not ( n14506 , n14505 );
or ( n14507 , n14500 , n14506 );
nand ( n14508 , n14356 , n3017 );
nand ( n14509 , n14507 , n14508 );
and ( n14510 , n14499 , n14509 );
and ( n14511 , n14487 , n14498 );
or ( n14512 , n14510 , n14511 );
and ( n14513 , n14476 , n14512 );
and ( n14514 , n14466 , n14475 );
or ( n14515 , n14513 , n14514 );
xor ( n14516 , n14456 , n14515 );
not ( n14517 , n3134 );
not ( n14518 , n14435 );
or ( n14519 , n14517 , n14518 );
buf ( n14520 , n5606 );
or ( n14521 , n14520 , n3177 );
nand ( n14522 , n14520 , n3177 );
nand ( n14523 , n14521 , n14522 );
nand ( n14524 , n14523 , n11729 );
nand ( n14525 , n14519 , n14524 );
not ( n14526 , n14397 );
not ( n14527 , n14446 );
or ( n14528 , n14526 , n14527 );
not ( n14529 , n539 );
not ( n14530 , n11447 );
or ( n14531 , n14529 , n14530 );
nand ( n14532 , n10472 , n3069 );
nand ( n14533 , n14531 , n14532 );
nand ( n14534 , n14533 , n3103 );
nand ( n14535 , n14528 , n14534 );
xor ( n14536 , n14525 , n14535 );
not ( n14537 , n2362 );
not ( n14538 , n14464 );
or ( n14539 , n14537 , n14538 );
not ( n14540 , n543 );
not ( n14541 , n12050 );
not ( n14542 , n14541 );
or ( n14543 , n14540 , n14542 );
nand ( n14544 , n11644 , n2123 );
nand ( n14545 , n14543 , n14544 );
nand ( n14546 , n14545 , n714 );
nand ( n14547 , n14539 , n14546 );
and ( n14548 , n14536 , n14547 );
and ( n14549 , n14525 , n14535 );
or ( n14550 , n14548 , n14549 );
xor ( n14551 , n14439 , n14450 );
xor ( n14552 , n14551 , n14452 );
xor ( n14553 , n14550 , n14552 );
xor ( n14554 , n14252 , n14270 );
xor ( n14555 , n14554 , n14358 );
and ( n14556 , n14553 , n14555 );
and ( n14557 , n14550 , n14552 );
or ( n14558 , n14556 , n14557 );
xor ( n14559 , n14516 , n14558 );
xor ( n14560 , n14396 , n14559 );
xor ( n14561 , n14466 , n14475 );
xor ( n14562 , n14561 , n14512 );
not ( n14563 , n11729 );
not ( n14564 , n5093 );
not ( n14565 , n3177 );
or ( n14566 , n14564 , n14565 );
nand ( n14567 , n10631 , n537 );
nand ( n14568 , n14566 , n14567 );
not ( n14569 , n14568 );
or ( n14570 , n14563 , n14569 );
nand ( n14571 , n14523 , n3186 );
nand ( n14572 , n14570 , n14571 );
xor ( n14573 , n14572 , n14471 );
not ( n14574 , n3103 );
not ( n14575 , n539 );
not ( n14576 , n10672 );
or ( n14577 , n14575 , n14576 );
nand ( n14578 , n5582 , n3069 );
nand ( n14579 , n14577 , n14578 );
not ( n14580 , n14579 );
or ( n14581 , n14574 , n14580 );
nand ( n14582 , n14533 , n14397 );
nand ( n14583 , n14581 , n14582 );
and ( n14584 , n14573 , n14583 );
and ( n14585 , n14572 , n14471 );
or ( n14586 , n14584 , n14585 );
xor ( n14587 , n14468 , n14469 );
xor ( n14588 , n14587 , n14472 );
xor ( n14589 , n14586 , n14588 );
xor ( n14590 , n14525 , n14535 );
xor ( n14591 , n14590 , n14547 );
and ( n14592 , n14589 , n14591 );
and ( n14593 , n14586 , n14588 );
or ( n14594 , n14592 , n14593 );
xor ( n14595 , n14562 , n14594 );
not ( n14596 , n4022 );
and ( n14597 , n14246 , n549 );
not ( n14598 , n14246 );
and ( n14599 , n14598 , n4013 );
nor ( n14600 , n14597 , n14599 );
not ( n14601 , n14600 );
or ( n14602 , n14596 , n14601 );
nand ( n14603 , n6220 , n549 );
nand ( n14604 , n14602 , n14603 );
not ( n14605 , n3300 );
not ( n14606 , n547 );
not ( n14607 , n14427 );
or ( n14608 , n14606 , n14607 );
nand ( n14609 , n14350 , n2369 );
nand ( n14610 , n14608 , n14609 );
not ( n14611 , n14610 );
or ( n14612 , n14605 , n14611 );
nand ( n14613 , n14485 , n3298 );
nand ( n14614 , n14612 , n14613 );
xor ( n14615 , n14604 , n14614 );
and ( n14616 , n11907 , n545 );
not ( n14617 , n11907 );
and ( n14618 , n14617 , n706 );
or ( n14619 , n14616 , n14618 );
nand ( n14620 , n14619 , n2376 );
nand ( n14621 , n14505 , n3017 );
nand ( n14622 , n14620 , n14621 );
and ( n14623 , n14615 , n14622 );
and ( n14624 , n14604 , n14614 );
or ( n14625 , n14623 , n14624 );
nand ( n14626 , n4342 , n537 );
not ( n14627 , n6050 );
not ( n14628 , n6157 );
nand ( n14629 , n14627 , n14628 );
nand ( n14630 , n14626 , n14629 );
not ( n14631 , n3288 );
not ( n14632 , n541 );
not ( n14633 , n10439 );
or ( n14634 , n14632 , n14633 );
nand ( n14635 , n14444 , n3023 );
nand ( n14636 , n14634 , n14635 );
not ( n14637 , n14636 );
or ( n14638 , n14631 , n14637 );
not ( n14639 , n14491 );
not ( n14640 , n14494 );
or ( n14641 , n14639 , n14640 );
nand ( n14642 , n14641 , n3955 );
nand ( n14643 , n14638 , n14642 );
xor ( n14644 , n14630 , n14643 );
not ( n14645 , n2362 );
not ( n14646 , n14545 );
or ( n14647 , n14645 , n14646 );
and ( n14648 , n11241 , n543 );
not ( n14649 , n11241 );
and ( n14650 , n14649 , n3212 );
nor ( n14651 , n14648 , n14650 );
nand ( n14652 , n14651 , n714 );
nand ( n14653 , n14647 , n14652 );
and ( n14654 , n14644 , n14653 );
and ( n14655 , n14630 , n14643 );
or ( n14656 , n14654 , n14655 );
xor ( n14657 , n14625 , n14656 );
xor ( n14658 , n14487 , n14498 );
xor ( n14659 , n14658 , n14509 );
and ( n14660 , n14657 , n14659 );
and ( n14661 , n14625 , n14656 );
or ( n14662 , n14660 , n14661 );
and ( n14663 , n14595 , n14662 );
and ( n14664 , n14562 , n14594 );
or ( n14665 , n14663 , n14664 );
xor ( n14666 , n14560 , n14665 );
not ( n14667 , n14666 );
xor ( n14668 , n14550 , n14552 );
xor ( n14669 , n14668 , n14555 );
xor ( n14670 , n14562 , n14594 );
xor ( n14671 , n14670 , n14662 );
xor ( n14672 , n14669 , n14671 );
not ( n14673 , n3134 );
not ( n14674 , n14568 );
or ( n14675 , n14673 , n14674 );
not ( n14676 , n537 );
not ( n14677 , n10995 );
or ( n14678 , n14676 , n14677 );
nand ( n14679 , n11387 , n3177 );
nand ( n14680 , n14678 , n14679 );
nand ( n14681 , n11729 , n14680 );
nand ( n14682 , n14675 , n14681 );
not ( n14683 , n11729 );
not ( n14684 , n537 );
not ( n14685 , n4339 );
or ( n14686 , n14684 , n14685 );
nand ( n14687 , n4342 , n3177 );
nand ( n14688 , n14686 , n14687 );
not ( n14689 , n14688 );
or ( n14690 , n14683 , n14689 );
nand ( n14691 , n14680 , n3186 );
nand ( n14692 , n14690 , n14691 );
nand ( n14693 , n4652 , n537 );
not ( n14694 , n14693 );
and ( n14695 , n14692 , n14694 );
xor ( n14696 , n14682 , n14695 );
not ( n14697 , n539 );
not ( n14698 , n5607 );
or ( n14699 , n14697 , n14698 );
nand ( n14700 , n5614 , n3069 );
nand ( n14701 , n14699 , n14700 );
not ( n14702 , n14701 );
not ( n14703 , n3103 );
or ( n14704 , n14702 , n14703 );
not ( n14705 , n14579 );
or ( n14706 , n14705 , n10609 );
nand ( n14707 , n14704 , n14706 );
and ( n14708 , n14696 , n14707 );
and ( n14709 , n14682 , n14695 );
or ( n14710 , n14708 , n14709 );
xor ( n14711 , n14572 , n14471 );
xor ( n14712 , n14711 , n14583 );
xor ( n14713 , n14710 , n14712 );
not ( n14714 , n14603 );
nand ( n14715 , n14376 , n14714 );
nor ( n14716 , n6533 , n4013 );
nand ( n14717 , n14481 , n14716 );
nor ( n14718 , n6563 , n549 );
nand ( n14719 , n14246 , n14718 );
nor ( n14720 , n6533 , n549 );
nand ( n14721 , n14322 , n14720 );
nand ( n14722 , n14715 , n14717 , n14719 , n14721 );
not ( n14723 , n2362 );
not ( n14724 , n14651 );
or ( n14725 , n14723 , n14724 );
not ( n14726 , n543 );
not ( n14727 , n11475 );
or ( n14728 , n14726 , n14727 );
nand ( n14729 , n11478 , n2123 );
nand ( n14730 , n14728 , n14729 );
nand ( n14731 , n14730 , n714 );
nand ( n14732 , n14725 , n14731 );
xor ( n14733 , n14722 , n14732 );
not ( n14734 , n3300 );
not ( n14735 , n2369 );
not ( n14736 , n14419 );
or ( n14737 , n14735 , n14736 );
nand ( n14738 , n547 , n12187 );
nand ( n14739 , n14737 , n14738 );
not ( n14740 , n14739 );
or ( n14741 , n14734 , n14740 );
nand ( n14742 , n14610 , n3298 );
nand ( n14743 , n14741 , n14742 );
and ( n14744 , n14733 , n14743 );
and ( n14745 , n14722 , n14732 );
or ( n14746 , n14744 , n14745 );
and ( n14747 , n14713 , n14746 );
and ( n14748 , n14710 , n14712 );
or ( n14749 , n14747 , n14748 );
xor ( n14750 , n14586 , n14588 );
xor ( n14751 , n14750 , n14591 );
xor ( n14752 , n14749 , n14751 );
xor ( n14753 , n14630 , n14643 );
xor ( n14754 , n14753 , n14653 );
or ( n14755 , n14626 , n14629 );
nand ( n14756 , n14755 , n14630 );
not ( n14757 , n3955 );
not ( n14758 , n14636 );
or ( n14759 , n14757 , n14758 );
not ( n14760 , n541 );
not ( n14761 , n10473 );
or ( n14762 , n14760 , n14761 );
nand ( n14763 , n10472 , n3023 );
nand ( n14764 , n14762 , n14763 );
nand ( n14765 , n14764 , n3288 );
nand ( n14766 , n14759 , n14765 );
xor ( n14767 , n14756 , n14766 );
not ( n14768 , n3017 );
not ( n14769 , n14619 );
or ( n14770 , n14768 , n14769 );
not ( n14771 , n545 );
not ( n14772 , n14541 );
or ( n14773 , n14771 , n14772 );
nand ( n14774 , n11644 , n706 );
nand ( n14775 , n14773 , n14774 );
nand ( n14776 , n14775 , n2376 );
nand ( n14777 , n14770 , n14776 );
and ( n14778 , n14767 , n14777 );
and ( n14779 , n14756 , n14766 );
or ( n14780 , n14778 , n14779 );
xor ( n14781 , n14754 , n14780 );
xor ( n14782 , n14604 , n14614 );
xor ( n14783 , n14782 , n14622 );
and ( n14784 , n14781 , n14783 );
and ( n14785 , n14754 , n14780 );
or ( n14786 , n14784 , n14785 );
and ( n14787 , n14752 , n14786 );
and ( n14788 , n14749 , n14751 );
or ( n14789 , n14787 , n14788 );
and ( n14790 , n14672 , n14789 );
and ( n14791 , n14669 , n14671 );
or ( n14792 , n14790 , n14791 );
not ( n14793 , n14792 );
nand ( n14794 , n14667 , n14793 );
not ( n14795 , n14794 );
xor ( n14796 , n11988 , n12002 );
and ( n14797 , n14796 , n12032 );
and ( n14798 , n11988 , n12002 );
or ( n14799 , n14797 , n14798 );
not ( n14800 , n3955 );
not ( n14801 , n541 );
not ( n14802 , n10631 );
or ( n14803 , n14801 , n14802 );
nand ( n14804 , n5093 , n3023 );
nand ( n14805 , n14803 , n14804 );
not ( n14806 , n14805 );
or ( n14807 , n14800 , n14806 );
not ( n14808 , n11952 );
not ( n14809 , n11954 );
or ( n14810 , n14808 , n14809 );
nand ( n14811 , n14810 , n3288 );
nand ( n14812 , n14807 , n14811 );
xor ( n14813 , n12013 , n12015 );
and ( n14814 , n14813 , n12031 );
and ( n14815 , n12013 , n12015 );
or ( n14816 , n14814 , n14815 );
xor ( n14817 , n14812 , n14816 );
not ( n14818 , n2362 );
not ( n14819 , n543 );
not ( n14820 , n5577 );
or ( n14821 , n14819 , n14820 );
nand ( n14822 , n5582 , n2123 );
nand ( n14823 , n14821 , n14822 );
not ( n14824 , n14823 );
or ( n14825 , n14818 , n14824 );
nand ( n14826 , n11965 , n714 );
nand ( n14827 , n14825 , n14826 );
xor ( n14828 , n14817 , n14827 );
xor ( n14829 , n14799 , n14828 );
xor ( n14830 , n12056 , n12060 );
and ( n14831 , n14830 , n12194 );
and ( n14832 , n12056 , n12060 );
or ( n14833 , n14831 , n14832 );
xor ( n14834 , n14829 , n14833 );
xor ( n14835 , n12043 , n12195 );
and ( n14836 , n14835 , n12200 );
and ( n14837 , n12043 , n12195 );
or ( n14838 , n14836 , n14837 );
xor ( n14839 , n14834 , n14838 );
not ( n14840 , n3298 );
and ( n14841 , n11241 , n2369 );
not ( n14842 , n11241 );
and ( n14843 , n14842 , n547 );
or ( n14844 , n14841 , n14843 );
not ( n14845 , n14844 );
or ( n14846 , n14840 , n14845 );
nand ( n14847 , n11993 , n3300 );
nand ( n14848 , n14846 , n14847 );
not ( n14849 , n537 );
nor ( n14850 , n14849 , n2356 );
nand ( n14851 , n12028 , n14850 );
not ( n14852 , n14851 );
not ( n14853 , n3103 );
not ( n14854 , n12008 );
or ( n14855 , n14853 , n14854 );
and ( n14856 , n4338 , n11419 );
not ( n14857 , n4338 );
and ( n14858 , n14857 , n11416 );
nor ( n14859 , n14856 , n14858 );
nand ( n14860 , n14855 , n14859 );
xor ( n14861 , n14852 , n14860 );
nand ( n14862 , n4784 , n537 );
not ( n14863 , n12026 );
not ( n14864 , n14863 );
not ( n14865 , n11729 );
not ( n14866 , n14865 );
and ( n14867 , n14864 , n14866 );
and ( n14868 , n3630 , n3177 );
not ( n14869 , n3630 );
and ( n14870 , n14869 , n537 );
or ( n14871 , n14868 , n14870 );
and ( n14872 , n14871 , n3186 );
nor ( n14873 , n14867 , n14872 );
xor ( n14874 , n14862 , n14873 );
xor ( n14875 , n14861 , n14874 );
xor ( n14876 , n14848 , n14875 );
xor ( n14877 , n11958 , n11967 );
and ( n14878 , n14877 , n11978 );
and ( n14879 , n11958 , n11967 );
or ( n14880 , n14878 , n14879 );
xor ( n14881 , n14876 , n14880 );
not ( n14882 , n3017 );
not ( n14883 , n545 );
not ( n14884 , n10439 );
or ( n14885 , n14883 , n14884 );
nand ( n14886 , n10438 , n706 );
nand ( n14887 , n14885 , n14886 );
not ( n14888 , n14887 );
or ( n14889 , n14882 , n14888 );
nand ( n14890 , n2376 , n11974 );
nand ( n14891 , n14889 , n14890 );
not ( n14892 , n6220 );
and ( n14893 , n11902 , n4013 );
not ( n14894 , n11902 );
and ( n14895 , n14894 , n549 );
or ( n14896 , n14893 , n14895 );
not ( n14897 , n14896 );
or ( n14898 , n14892 , n14897 );
nand ( n14899 , n12054 , n4022 );
nand ( n14900 , n14898 , n14899 );
xor ( n14901 , n14891 , n14900 );
not ( n14902 , n551 );
not ( n14903 , n14427 );
or ( n14904 , n14902 , n14903 );
nand ( n14905 , n14350 , n4018 );
nand ( n14906 , n14904 , n14905 );
not ( n14907 , n14906 );
not ( n14908 , n552 );
or ( n14909 , n14907 , n14908 );
not ( n14910 , n5618 );
nand ( n14911 , n14910 , n12192 );
nand ( n14912 , n14909 , n14911 );
xor ( n14913 , n14901 , n14912 );
xor ( n14914 , n14881 , n14913 );
xor ( n14915 , n11979 , n11983 );
and ( n14916 , n14915 , n12033 );
and ( n14917 , n11979 , n11983 );
or ( n14918 , n14916 , n14917 );
xor ( n14919 , n14914 , n14918 );
xor ( n14920 , n14839 , n14919 );
xor ( n14921 , n12034 , n12038 );
and ( n14922 , n14921 , n12201 );
and ( n14923 , n12034 , n12038 );
or ( n14924 , n14922 , n14923 );
nor ( n14925 , n14920 , n14924 );
nor ( n14926 , n12202 , n11948 );
nor ( n14927 , n14925 , n14926 );
not ( n14928 , n3288 );
not ( n14929 , n14805 );
or ( n14930 , n14928 , n14929 );
and ( n14931 , n3023 , n5607 );
not ( n14932 , n3023 );
and ( n14933 , n14932 , n5614 );
nor ( n14934 , n14931 , n14933 );
nand ( n14935 , n14934 , n3955 );
nand ( n14936 , n14930 , n14935 );
not ( n14937 , n714 );
not ( n14938 , n14823 );
or ( n14939 , n14937 , n14938 );
not ( n14940 , n543 );
not ( n14941 , n11055 );
or ( n14942 , n14940 , n14941 );
nand ( n14943 , n10472 , n2123 );
nand ( n14944 , n14942 , n14943 );
nand ( n14945 , n14944 , n2362 );
nand ( n14946 , n14939 , n14945 );
xor ( n14947 , n14936 , n14946 );
not ( n14948 , n2376 );
not ( n14949 , n14887 );
or ( n14950 , n14948 , n14949 );
and ( n14951 , n10949 , n545 );
not ( n14952 , n10949 );
and ( n14953 , n14952 , n706 );
nor ( n14954 , n14951 , n14953 );
nand ( n14955 , n14954 , n3017 );
nand ( n14956 , n14950 , n14955 );
xor ( n14957 , n14947 , n14956 );
xor ( n14958 , n14891 , n14900 );
and ( n14959 , n14958 , n14912 );
and ( n14960 , n14891 , n14900 );
or ( n14961 , n14959 , n14960 );
xor ( n14962 , n14957 , n14961 );
not ( n14963 , n3298 );
not ( n14964 , n547 );
not ( n14965 , n11641 );
or ( n14966 , n14964 , n14965 );
nand ( n14967 , n12050 , n2369 );
nand ( n14968 , n14966 , n14967 );
not ( n14969 , n14968 );
or ( n14970 , n14963 , n14969 );
nand ( n14971 , n14844 , n3300 );
nand ( n14972 , n14970 , n14971 );
not ( n14973 , n3103 );
and ( n14974 , n4338 , n3069 );
not ( n14975 , n4338 );
and ( n14976 , n14975 , n539 );
or ( n14977 , n14974 , n14976 );
not ( n14978 , n14977 );
or ( n14979 , n14973 , n14978 );
and ( n14980 , n4635 , n11416 );
not ( n14981 , n4635 );
and ( n14982 , n14981 , n11419 );
nor ( n14983 , n14980 , n14982 );
nand ( n14984 , n14979 , n14983 );
nor ( n14985 , n14873 , n14862 );
xor ( n14986 , n14984 , n14985 );
and ( n14987 , n4792 , n537 );
not ( n14988 , n3186 );
not ( n14989 , n537 );
not ( n14990 , n3943 );
or ( n122542 , n14989 , n14990 );
nand ( n14991 , n3946 , n3177 );
nand ( n14992 , n122542 , n14991 );
not ( n14993 , n14992 );
or ( n14994 , n14988 , n14993 );
nand ( n14995 , n14871 , n11729 );
nand ( n14996 , n14994 , n14995 );
xor ( n14997 , n14987 , n14996 );
xor ( n14998 , n14986 , n14997 );
xor ( n14999 , n14972 , n14998 );
xor ( n15000 , n14812 , n14816 );
and ( n15001 , n15000 , n14827 );
and ( n15002 , n14812 , n14816 );
or ( n15003 , n15001 , n15002 );
xor ( n15004 , n14999 , n15003 );
xor ( n15005 , n14962 , n15004 );
xor ( n15006 , n14848 , n14875 );
and ( n15007 , n15006 , n14880 );
and ( n15008 , n14848 , n14875 );
or ( n15009 , n15007 , n15008 );
xor ( n15010 , n14852 , n14860 );
and ( n15011 , n15010 , n14874 );
and ( n15012 , n14852 , n14860 );
or ( n15013 , n15011 , n15012 );
nand ( n15014 , n11908 , n14720 );
nand ( n15015 , n11907 , n14716 );
nand ( n15016 , n14416 , n14714 );
nand ( n15017 , n12186 , n14718 );
nand ( n15018 , n15014 , n15015 , n15016 , n15017 );
xor ( n15019 , n15013 , n15018 );
not ( n15020 , n552 );
nor ( n15021 , n14481 , n4018 );
nor ( n15022 , n14322 , n551 );
nor ( n15023 , n15021 , n15022 );
not ( n15024 , n15023 );
or ( n15025 , n15020 , n15024 );
nand ( n15026 , n14906 , n5619 );
nand ( n15027 , n15025 , n15026 );
xor ( n15028 , n15019 , n15027 );
xor ( n15029 , n15009 , n15028 );
xor ( n15030 , n14799 , n14828 );
and ( n15031 , n15030 , n14833 );
and ( n15032 , n14799 , n14828 );
or ( n15033 , n15031 , n15032 );
xor ( n15034 , n15029 , n15033 );
xor ( n15035 , n15005 , n15034 );
xor ( n15036 , n14881 , n14913 );
and ( n15037 , n15036 , n14918 );
and ( n15038 , n14881 , n14913 );
or ( n15039 , n15037 , n15038 );
and ( n15040 , n15035 , n15039 );
and ( n15041 , n15005 , n15034 );
or ( n15042 , n15040 , n15041 );
not ( n15043 , n15042 );
xor ( n15044 , n15013 , n15018 );
and ( n15045 , n15044 , n15027 );
and ( n15046 , n15013 , n15018 );
or ( n15047 , n15045 , n15046 );
not ( n15048 , n3955 );
and ( n15049 , n541 , n5579 );
not ( n15050 , n541 );
and ( n15051 , n15050 , n5578 );
or ( n15052 , n15049 , n15051 );
not ( n15053 , n15052 );
or ( n15054 , n15048 , n15053 );
nand ( n15055 , n14934 , n3288 );
nand ( n15056 , n15054 , n15055 );
xor ( n15057 , n14984 , n14985 );
and ( n15058 , n15057 , n14997 );
and ( n15059 , n14984 , n14985 );
or ( n15060 , n15058 , n15059 );
xor ( n15061 , n15056 , n15060 );
not ( n15062 , n2362 );
and ( n15063 , n10438 , n2123 );
not ( n15064 , n10438 );
and ( n122617 , n15064 , n543 );
or ( n15065 , n15063 , n122617 );
not ( n15066 , n15065 );
or ( n15067 , n15062 , n15066 );
nand ( n15068 , n14944 , n714 );
nand ( n15069 , n15067 , n15068 );
xor ( n15070 , n15061 , n15069 );
xor ( n15071 , n15047 , n15070 );
xor ( n15072 , n14972 , n14998 );
and ( n15073 , n15072 , n15003 );
and ( n15074 , n14972 , n14998 );
or ( n15075 , n15073 , n15074 );
xor ( n15076 , n15071 , n15075 );
xor ( n15077 , n15009 , n15028 );
and ( n15078 , n15077 , n15033 );
and ( n15079 , n15009 , n15028 );
or ( n15080 , n15078 , n15079 );
xor ( n15081 , n15076 , n15080 );
not ( n15082 , n3017 );
not ( n15083 , n545 );
not ( n15084 , n11241 );
not ( n15085 , n15084 );
or ( n15086 , n15083 , n15085 );
nand ( n15087 , n11241 , n706 );
nand ( n15088 , n15086 , n15087 );
not ( n15089 , n15088 );
or ( n15090 , n15082 , n15089 );
nand ( n15091 , n14954 , n2376 );
nand ( n15092 , n15090 , n15091 );
not ( n15093 , n552 );
and ( n15094 , n14246 , n4018 );
not ( n15095 , n14246 );
and ( n15096 , n15095 , n551 );
or ( n15097 , n15094 , n15096 );
not ( n15098 , n15097 );
or ( n15099 , n15093 , n15098 );
nor ( n15100 , n14481 , n4018 );
not ( n15101 , n15100 );
not ( n15102 , n15022 );
nand ( n15103 , n15101 , n15102 , n5619 );
nand ( n15104 , n15099 , n15103 );
xor ( n15105 , n15092 , n15104 );
not ( n15106 , n4022 );
not ( n15107 , n549 );
not ( n15108 , n12187 );
or ( n15109 , n15107 , n15108 );
nand ( n15110 , n12190 , n4013 );
nand ( n15111 , n15109 , n15110 );
not ( n15112 , n15111 );
or ( n15113 , n15106 , n15112 );
not ( n15114 , n549 );
not ( n15115 , n14351 );
or ( n15116 , n15114 , n15115 );
nand ( n15117 , n14428 , n4013 );
nand ( n15118 , n15116 , n15117 );
nand ( n15119 , n6220 , n15118 );
nand ( n15120 , n15113 , n15119 );
xor ( n15121 , n15105 , n15120 );
not ( n15122 , n3298 );
not ( n15123 , n547 );
not ( n15124 , n11907 );
or ( n15125 , n15123 , n15124 );
nand ( n15126 , n11908 , n2369 );
nand ( n15127 , n15125 , n15126 );
not ( n15128 , n15127 );
or ( n15129 , n15122 , n15128 );
not ( n15130 , n11996 );
nand ( n15131 , n15130 , n14968 );
nand ( n15132 , n15129 , n15131 );
and ( n15133 , n14987 , n14996 );
not ( n15134 , n3025 );
not ( n15135 , n10631 );
not ( n15136 , n539 );
or ( n15137 , n15135 , n15136 );
nand ( n15138 , n5093 , n3069 );
nand ( n15139 , n15137 , n15138 );
not ( n15140 , n15139 );
or ( n15141 , n15134 , n15140 );
and ( n15142 , n10995 , n4701 );
and ( n15143 , n4638 , n4699 );
nor ( n15144 , n15142 , n15143 );
nand ( n15145 , n15141 , n15144 );
xor ( n15146 , n15133 , n15145 );
not ( n15147 , n537 );
nor ( n15148 , n15147 , n6156 );
not ( n15149 , n3186 );
not ( n15150 , n14688 );
or ( n15151 , n15149 , n15150 );
nand ( n15152 , n14992 , n11729 );
nand ( n15153 , n15151 , n15152 );
xor ( n15154 , n15148 , n15153 );
xor ( n15155 , n15146 , n15154 );
xor ( n15156 , n15132 , n15155 );
xor ( n15157 , n14936 , n14946 );
and ( n15158 , n15157 , n14956 );
and ( n15159 , n14936 , n14946 );
or ( n15160 , n15158 , n15159 );
xor ( n15161 , n15156 , n15160 );
xor ( n15162 , n15121 , n15161 );
xor ( n15163 , n14957 , n14961 );
and ( n15164 , n15163 , n15004 );
and ( n15165 , n14957 , n14961 );
or ( n15166 , n15164 , n15165 );
xor ( n15167 , n15162 , n15166 );
xor ( n15168 , n15081 , n15167 );
not ( n15169 , n15168 );
nand ( n15170 , n15043 , n15169 );
and ( n15171 , n14927 , n15170 );
xor ( n15172 , n15076 , n15080 );
and ( n15173 , n15172 , n15167 );
and ( n15174 , n15076 , n15080 );
or ( n15175 , n15173 , n15174 );
not ( n15176 , n15175 );
xor ( n15177 , n15092 , n15104 );
and ( n15178 , n15177 , n15120 );
and ( n15179 , n15092 , n15104 );
or ( n15180 , n15178 , n15179 );
not ( n15181 , n3955 );
not ( n15182 , n14764 );
or ( n15183 , n15181 , n15182 );
nand ( n15184 , n15052 , n3288 );
nand ( n15185 , n15183 , n15184 );
not ( n15186 , n714 );
not ( n15187 , n15065 );
or ( n15188 , n15186 , n15187 );
nand ( n15189 , n14730 , n2362 );
nand ( n15190 , n15188 , n15189 );
xor ( n15191 , n15185 , n15190 );
not ( n15192 , n2376 );
not ( n15193 , n15088 );
or ( n15194 , n15192 , n15193 );
not ( n15195 , n10512 );
nand ( n15196 , n15195 , n14775 );
nand ( n15197 , n15194 , n15196 );
xor ( n15198 , n15191 , n15197 );
xor ( n15199 , n15180 , n15198 );
not ( n15200 , n5619 );
not ( n15201 , n15097 );
or ( n15202 , n15200 , n15201 );
nand ( n15203 , n15202 , n14628 );
not ( n15204 , n14323 );
not ( n15205 , n549 );
or ( n15206 , n15204 , n15205 );
nand ( n15207 , n14326 , n4013 );
nand ( n15208 , n15206 , n15207 );
not ( n15209 , n15208 );
not ( n15210 , n4020 );
or ( n15211 , n15209 , n15210 );
nand ( n15212 , n15118 , n4022 );
nand ( n15213 , n15211 , n15212 );
xor ( n15214 , n15203 , n15213 );
not ( n15215 , n3300 );
not ( n15216 , n15127 );
or ( n15217 , n15215 , n15216 );
nand ( n15218 , n14739 , n3298 );
nand ( n15219 , n15217 , n15218 );
xor ( n15220 , n15214 , n15219 );
xor ( n15221 , n15199 , n15220 );
xor ( n15222 , n15132 , n15155 );
and ( n15223 , n15222 , n15160 );
and ( n15224 , n15132 , n15155 );
or ( n15225 , n15223 , n15224 );
xor ( n15226 , n15133 , n15145 );
and ( n15227 , n15226 , n15154 );
and ( n15228 , n15133 , n15145 );
or ( n15229 , n15227 , n15228 );
xor ( n15230 , n15056 , n15060 );
and ( n15231 , n15230 , n15069 );
and ( n15232 , n15056 , n15060 );
or ( n15233 , n15231 , n15232 );
xor ( n15234 , n15229 , n15233 );
not ( n15235 , n3103 );
not ( n15236 , n15139 );
or ( n15237 , n15235 , n15236 );
nand ( n15238 , n14701 , n14397 );
nand ( n15239 , n15237 , n15238 );
and ( n15240 , n15148 , n15153 );
xor ( n15241 , n15239 , n15240 );
and ( n15242 , n14692 , n14694 );
not ( n15243 , n14692 );
and ( n15244 , n15243 , n14693 );
nor ( n15245 , n15242 , n15244 );
xor ( n15246 , n15241 , n15245 );
xor ( n15247 , n15234 , n15246 );
xor ( n15248 , n15225 , n15247 );
xor ( n15249 , n15047 , n15070 );
and ( n15250 , n15249 , n15075 );
and ( n15251 , n15047 , n15070 );
or ( n15252 , n15250 , n15251 );
xor ( n15253 , n15248 , n15252 );
xor ( n15254 , n15221 , n15253 );
xor ( n15255 , n15121 , n15161 );
and ( n15256 , n15255 , n15166 );
and ( n15257 , n15121 , n15161 );
or ( n15258 , n15256 , n15257 );
xor ( n15259 , n15254 , n15258 );
not ( n15260 , n15259 );
nand ( n15261 , n15176 , n15260 );
buf ( n15262 , n15261 );
xor ( n15263 , n15005 , n15034 );
xor ( n15264 , n15263 , n15039 );
xor ( n15265 , n14834 , n14838 );
and ( n15266 , n15265 , n14919 );
and ( n15267 , n14834 , n14838 );
or ( n15268 , n15266 , n15267 );
or ( n15269 , n15264 , n15268 );
nand ( n15270 , n15171 , n11943 , n15262 , n15269 );
not ( n15271 , n15260 );
nor ( n15272 , n15271 , n15175 );
nor ( n15273 , n15042 , n15168 );
nor ( n15274 , n15272 , n15273 );
not ( n15275 , n15264 );
not ( n15276 , n15268 );
and ( n15277 , n15275 , n15276 );
not ( n15278 , n12204 );
nand ( n15279 , n14920 , n14924 );
not ( n15280 , n15279 );
or ( n15281 , n15278 , n15280 );
not ( n15282 , n14920 );
not ( n15283 , n14924 );
nand ( n15284 , n15282 , n15283 );
nand ( n15285 , n15281 , n15284 );
nand ( n15286 , n15264 , n15268 );
and ( n15287 , n15285 , n15286 );
nor ( n15288 , n15277 , n15287 );
and ( n15289 , n15274 , n15288 );
not ( n15290 , n15261 );
nand ( n15291 , n15042 , n15168 );
not ( n15292 , n15291 );
not ( n15293 , n15292 );
or ( n15294 , n15290 , n15293 );
nand ( n15295 , n15271 , n15175 );
nand ( n15296 , n15294 , n15295 );
nor ( n15297 , n15289 , n15296 );
nand ( n15298 , n15270 , n15297 );
not ( n15299 , n15298 );
xor ( n15300 , n14754 , n14780 );
xor ( n15301 , n15300 , n14783 );
xor ( n15302 , n14710 , n14712 );
xor ( n15303 , n15302 , n14746 );
xor ( n15304 , n15239 , n15240 );
and ( n15305 , n15304 , n15245 );
and ( n15306 , n15239 , n15240 );
or ( n15307 , n15305 , n15306 );
xor ( n15308 , n14682 , n14695 );
xor ( n15309 , n15308 , n14707 );
xor ( n15310 , n15307 , n15309 );
xor ( n15311 , n14756 , n14766 );
xor ( n15312 , n15311 , n14777 );
and ( n15313 , n15310 , n15312 );
and ( n15314 , n15307 , n15309 );
or ( n15315 , n15313 , n15314 );
xor ( n15316 , n15303 , n15315 );
xor ( n15317 , n15185 , n15190 );
and ( n15318 , n15317 , n15197 );
and ( n15319 , n15185 , n15190 );
or ( n15320 , n15318 , n15319 );
xor ( n15321 , n15203 , n15213 );
and ( n15322 , n15321 , n15219 );
and ( n15323 , n15203 , n15213 );
or ( n15324 , n15322 , n15323 );
xor ( n15325 , n15320 , n15324 );
xor ( n15326 , n14722 , n14732 );
xor ( n15327 , n15326 , n14743 );
and ( n15328 , n15325 , n15327 );
and ( n15329 , n15320 , n15324 );
or ( n15330 , n15328 , n15329 );
xor ( n15331 , n15316 , n15330 );
xor ( n15332 , n15301 , n15331 );
xor ( n15333 , n15229 , n15233 );
and ( n15334 , n15333 , n15246 );
and ( n15335 , n15229 , n15233 );
or ( n15336 , n15334 , n15335 );
xor ( n15337 , n15307 , n15309 );
xor ( n15338 , n15337 , n15312 );
xor ( n15339 , n15336 , n15338 );
xor ( n15340 , n15180 , n15198 );
and ( n15341 , n15340 , n15220 );
and ( n15342 , n15180 , n15198 );
or ( n15343 , n15341 , n15342 );
and ( n15344 , n15339 , n15343 );
and ( n15345 , n15336 , n15338 );
or ( n15346 , n15344 , n15345 );
xor ( n15347 , n15332 , n15346 );
xor ( n15348 , n15320 , n15324 );
xor ( n15349 , n15348 , n15327 );
xor ( n15350 , n15336 , n15338 );
xor ( n15351 , n15350 , n15343 );
xor ( n15352 , n15349 , n15351 );
xor ( n15353 , n15225 , n15247 );
and ( n15354 , n15353 , n15252 );
and ( n15355 , n15225 , n15247 );
or ( n15356 , n15354 , n15355 );
and ( n15357 , n15352 , n15356 );
and ( n15358 , n15349 , n15351 );
or ( n15359 , n15357 , n15358 );
nor ( n15360 , n15347 , n15359 );
xor ( n15361 , n15349 , n15351 );
xor ( n15362 , n15361 , n15356 );
xor ( n15363 , n15221 , n15253 );
and ( n15364 , n15363 , n15258 );
and ( n15365 , n15221 , n15253 );
or ( n15366 , n15364 , n15365 );
nor ( n15367 , n15362 , n15366 );
nor ( n15368 , n15360 , n15367 );
xor ( n15369 , n14669 , n14671 );
xor ( n15370 , n15369 , n14789 );
xor ( n15371 , n14625 , n14656 );
xor ( n15372 , n15371 , n14659 );
xor ( n15373 , n14749 , n14751 );
xor ( n15374 , n15373 , n14786 );
xor ( n15375 , n15372 , n15374 );
xor ( n15376 , n15303 , n15315 );
and ( n15377 , n15376 , n15330 );
and ( n15378 , n15303 , n15315 );
or ( n15379 , n15377 , n15378 );
and ( n15380 , n15375 , n15379 );
and ( n15381 , n15372 , n15374 );
or ( n15382 , n15380 , n15381 );
nor ( n15383 , n15370 , n15382 );
xor ( n15384 , n15372 , n15374 );
xor ( n15385 , n15384 , n15379 );
xor ( n15386 , n15301 , n15331 );
and ( n15387 , n15386 , n15346 );
and ( n15388 , n15301 , n15331 );
or ( n15389 , n15387 , n15388 );
nor ( n15390 , n15385 , n15389 );
nor ( n15391 , n15383 , n15390 );
and ( n15392 , n15368 , n15391 );
not ( n15393 , n15392 );
or ( n15394 , n15299 , n15393 );
nor ( n15395 , n15347 , n15359 );
nand ( n15396 , n15362 , n15366 );
or ( n15397 , n15395 , n15396 );
nand ( n15398 , n15347 , n15359 );
nand ( n15399 , n15397 , n15398 );
nand ( n15400 , n15399 , n15391 );
not ( n15401 , n15385 );
not ( n15402 , n15389 );
nor ( n15403 , n15401 , n15402 );
not ( n15404 , n15383 );
nand ( n15405 , n15403 , n15404 );
buf ( n15406 , n15370 );
nand ( n15407 , n15406 , n15382 );
and ( n15408 , n15400 , n15405 , n15407 );
nand ( n15409 , n15394 , n15408 );
not ( n15410 , n15409 );
or ( n15411 , n14795 , n15410 );
nand ( n15412 , n14666 , n14792 );
buf ( n15413 , n15412 );
nand ( n15414 , n15411 , n15413 );
xor ( n15415 , n14396 , n14559 );
and ( n15416 , n15415 , n14665 );
and ( n15417 , n14396 , n14559 );
or ( n15418 , n15416 , n15417 );
not ( n15419 , n15418 );
xor ( n15420 , n14047 , n14048 );
and ( n15421 , n15420 , n14050 );
and ( n15422 , n14047 , n14048 );
or ( n15423 , n15421 , n15422 );
xor ( n15424 , n14371 , n14383 );
and ( n15425 , n15424 , n14394 );
and ( n15426 , n14371 , n14383 );
or ( n15427 , n15425 , n15426 );
xor ( n15428 , n15423 , n15427 );
not ( n15429 , n2362 );
not ( n15430 , n543 );
not ( n15431 , n14323 );
or ( n15432 , n15430 , n15431 );
nand ( n15433 , n14326 , n2123 );
nand ( n15434 , n15432 , n15433 );
not ( n15435 , n15434 );
or ( n15436 , n15429 , n15435 );
nand ( n15437 , n14430 , n714 );
nand ( n15438 , n15436 , n15437 );
not ( n15439 , n3955 );
not ( n15440 , n541 );
not ( n15441 , n12187 );
or ( n15442 , n15440 , n15441 );
nand ( n15443 , n12190 , n3023 );
nand ( n15444 , n15442 , n15443 );
not ( n15445 , n15444 );
or ( n15446 , n15439 , n15445 );
nand ( n15447 , n14390 , n3288 );
nand ( n15448 , n15446 , n15447 );
xor ( n15449 , n15438 , n15448 );
not ( n15450 , n10473 );
nand ( n15451 , n15450 , n537 );
xor ( n15452 , n15449 , n15451 );
xor ( n15453 , n15428 , n15452 );
not ( n15454 , n11729 );
not ( n15455 , n14364 );
or ( n15456 , n15454 , n15455 );
not ( n15457 , n537 );
not ( n15458 , n14407 );
or ( n15459 , n15457 , n15458 );
not ( n15460 , n11475 );
nand ( n15461 , n15460 , n3177 );
nand ( n15462 , n15459 , n15461 );
nand ( n15463 , n15462 , n3134 );
nand ( n15464 , n15456 , n15463 );
not ( n15465 , n2376 );
not ( n15466 , n14381 );
or ( n15467 , n15465 , n15466 );
nand ( n15468 , n15467 , n11265 );
xor ( n15469 , n15464 , n15468 );
not ( n15470 , n3103 );
not ( n15471 , n14403 );
or ( n15472 , n15470 , n15471 );
not ( n15473 , n539 );
not ( n15474 , n14256 );
or ( n15475 , n15473 , n15474 );
nand ( n15476 , n14255 , n3069 );
nand ( n15477 , n15475 , n15476 );
nand ( n15478 , n15477 , n14397 );
nand ( n15479 , n15472 , n15478 );
xor ( n15480 , n15469 , n15479 );
xor ( n15481 , n14413 , n14432 );
and ( n15482 , n15481 , n14455 );
and ( n15483 , n14413 , n14432 );
or ( n15484 , n15482 , n15483 );
xor ( n15485 , n15480 , n15484 );
xor ( n15486 , n14051 , n14361 );
and ( n15487 , n15486 , n14395 );
and ( n15488 , n14051 , n14361 );
or ( n15489 , n15487 , n15488 );
xor ( n15490 , n15485 , n15489 );
xor ( n15491 , n15453 , n15490 );
xor ( n15492 , n14456 , n14515 );
and ( n15493 , n15492 , n14558 );
and ( n15494 , n14456 , n14515 );
or ( n15495 , n15493 , n15494 );
xor ( n15496 , n15491 , n15495 );
not ( n15497 , n15496 );
nand ( n15498 , n15419 , n15497 );
nand ( n15499 , n15418 , n15496 );
nand ( n15500 , n15498 , n15499 );
not ( n15501 , n15500 );
and ( n15502 , n15414 , n15501 );
not ( n15503 , n15414 );
and ( n15504 , n15503 , n15500 );
nor ( n15505 , n15502 , n15504 );
nand ( n15506 , n15505 , n454 );
xor ( n15507 , n9733 , n9801 );
xor ( n15508 , n15507 , n9804 );
nand ( n15509 , n15508 , n9907 );
not ( n15510 , n13416 );
not ( n15511 , n13777 );
or ( n15512 , n15510 , n15511 );
nand ( n15513 , n15512 , n14025 );
buf ( n15514 , n13650 );
nand ( n15515 , n15514 , n13785 );
xnor ( n15516 , n15513 , n15515 );
nand ( n15517 , n9907 , n15516 );
and ( n15518 , n489 , n13634 );
not ( n15519 , n15518 );
not ( n15520 , n7326 );
not ( n15521 , n719 );
and ( n15522 , n457 , n525 );
not ( n15523 , n7881 );
xnor ( n15524 , n459 , n522 );
or ( n15525 , n15523 , n15524 );
not ( n15526 , n7888 );
not ( n15527 , n521 );
and ( n15528 , n459 , n15527 );
not ( n15529 , n459 );
and ( n15530 , n15529 , n521 );
nor ( n15531 , n15528 , n15530 );
or ( n15532 , n15526 , n15531 );
nand ( n15533 , n15525 , n15532 );
xor ( n15534 , n15522 , n15533 );
or ( n15535 , n7475 , n8719 );
nand ( n15536 , n15535 , n461 );
xor ( n15537 , n15534 , n15536 );
xnor ( n15538 , n457 , n524 );
or ( n15539 , n15538 , n8336 );
not ( n15540 , n7908 );
xnor ( n15541 , n457 , n523 );
or ( n15542 , n15540 , n15541 );
nand ( n15543 , n15539 , n15542 );
and ( n15544 , n8719 , n13827 );
and ( n15545 , n7475 , n461 );
nor ( n15546 , n15544 , n15545 );
not ( n15547 , n15546 );
xor ( n15548 , n15543 , n15547 );
and ( n15549 , n457 , n526 );
not ( n15550 , n13801 );
not ( n15551 , n7881 );
or ( n15552 , n15550 , n15551 );
not ( n15553 , n15524 );
nand ( n15554 , n15553 , n7888 );
nand ( n15555 , n15552 , n15554 );
xor ( n15556 , n15549 , n15555 );
not ( n15557 , n13821 );
not ( n15558 , n8337 );
or ( n15559 , n15557 , n15558 );
not ( n15560 , n15538 );
nand ( n15561 , n15560 , n7908 );
nand ( n15562 , n15559 , n15561 );
and ( n15563 , n15556 , n15562 );
and ( n15564 , n15549 , n15555 );
or ( n15565 , n15563 , n15564 );
xor ( n15566 , n15548 , n15565 );
xor ( n15567 , n15537 , n15566 );
xor ( n15568 , n15549 , n15555 );
xor ( n15569 , n15568 , n15562 );
xor ( n15570 , n15546 , n15569 );
xor ( n15571 , n13823 , n13829 );
and ( n15572 , n15571 , n13835 );
and ( n15573 , n13823 , n13829 );
or ( n15574 , n15572 , n15573 );
and ( n15575 , n15570 , n15574 );
and ( n15576 , n15546 , n15569 );
or ( n15577 , n15575 , n15576 );
and ( n15578 , n15567 , n15577 );
and ( n15579 , n15537 , n15566 );
or ( n15580 , n15578 , n15579 );
and ( n15581 , n524 , n457 );
xnor ( n15582 , n457 , n522 );
or ( n15583 , n15540 , n15582 );
not ( n15584 , n15541 );
nand ( n15585 , n15584 , n8337 );
nand ( n15586 , n15583 , n15585 );
xor ( n15587 , n15581 , n15586 );
not ( n15588 , n15523 );
not ( n15589 , n15531 );
and ( n15590 , n15588 , n15589 );
not ( n15591 , n459 );
nor ( n15592 , n15591 , n15526 );
nor ( n15593 , n15590 , n15592 );
xor ( n15594 , n15587 , n15593 );
xor ( n15595 , n15522 , n15533 );
and ( n15596 , n15595 , n15536 );
and ( n15597 , n15522 , n15533 );
or ( n15598 , n15596 , n15597 );
xor ( n15599 , n15543 , n15547 );
and ( n15600 , n15599 , n15565 );
and ( n15601 , n15543 , n15547 );
or ( n15602 , n15600 , n15601 );
xor ( n15603 , n15598 , n15602 );
xor ( n15604 , n15594 , n15603 );
or ( n15605 , n15580 , n15604 );
xor ( n15606 , n15581 , n15586 );
xor ( n15607 , n15606 , n15593 );
and ( n15608 , n15598 , n15607 );
xor ( n15609 , n15581 , n15586 );
xor ( n15610 , n15609 , n15593 );
and ( n15611 , n15602 , n15610 );
and ( n15612 , n15598 , n15602 );
or ( n15613 , n15608 , n15611 , n15612 );
xor ( n15614 , n15581 , n15586 );
and ( n15615 , n15614 , n15593 );
and ( n15616 , n15581 , n15586 );
or ( n15617 , n15615 , n15616 );
not ( n15618 , n15593 );
xor ( n15619 , n15617 , n15618 );
or ( n15620 , n7881 , n7888 );
nand ( n15621 , n15620 , n459 );
and ( n15622 , n523 , n457 );
xor ( n15623 , n15621 , n15622 );
or ( n15624 , n15582 , n8336 );
not ( n15625 , n457 );
and ( n15626 , n15625 , n521 );
and ( n15627 , n15527 , n457 );
nor ( n15628 , n15626 , n15627 );
or ( n15629 , n15540 , n15628 );
nand ( n15630 , n15624 , n15629 );
xor ( n15631 , n15623 , n15630 );
xor ( n15632 , n15619 , n15631 );
nor ( n15633 , n15613 , n15632 );
not ( n15634 , n15633 );
xor ( n15635 , n15617 , n15618 );
and ( n15636 , n15635 , n15631 );
and ( n15637 , n15617 , n15618 );
or ( n15638 , n15636 , n15637 );
or ( n15639 , n15628 , n8336 );
or ( n15640 , n15540 , n15625 );
nand ( n15641 , n15639 , n15640 );
nand ( n15642 , n522 , n457 );
xor ( n15643 , n15641 , n15642 );
xor ( n15644 , n15621 , n15622 );
and ( n15645 , n15644 , n15630 );
and ( n15646 , n15621 , n15622 );
or ( n15647 , n15645 , n15646 );
xor ( n15648 , n15643 , n15647 );
or ( n15649 , n15638 , n15648 );
and ( n15650 , n15605 , n15634 , n15649 );
not ( n15651 , n15650 );
xor ( n15652 , n15537 , n15566 );
xor ( n15653 , n15652 , n15577 );
not ( n15654 , n15653 );
xor ( n15655 , n13796 , n13598 );
and ( n15656 , n15655 , n13803 );
and ( n15657 , n13796 , n13598 );
or ( n15658 , n15656 , n15657 );
not ( n15659 , n15658 );
xor ( n15660 , n15546 , n15569 );
xor ( n15661 , n15660 , n15574 );
not ( n15662 , n15661 );
or ( n15663 , n15659 , n15662 );
not ( n15664 , n15658 );
not ( n15665 , n15664 );
not ( n15666 , n15661 );
not ( n15667 , n15666 );
or ( n15668 , n15665 , n15667 );
or ( n15669 , n13836 , n13804 );
nand ( n15670 , n15669 , n13817 );
nand ( n15671 , n13836 , n13804 );
and ( n15672 , n15670 , n15671 );
not ( n15673 , n15672 );
nand ( n15674 , n15668 , n15673 );
nand ( n15675 , n15663 , n15674 );
not ( n15676 , n15675 );
nand ( n15677 , n15654 , n15676 );
not ( n15678 , n15677 );
xor ( n15679 , n13837 , n13804 );
not ( n15680 , n13812 );
nand ( n15681 , n15679 , n15680 );
not ( n15682 , n15681 );
not ( n15683 , n13794 );
or ( n15684 , n15682 , n15683 );
or ( n15685 , n15679 , n15680 );
nand ( n15686 , n15684 , n15685 );
xor ( n15687 , n15658 , n15672 );
xnor ( n15688 , n15687 , n15661 );
nor ( n15689 , n15686 , n15688 );
nor ( n15690 , n15678 , n15689 );
not ( n15691 , n15690 );
not ( n15692 , n12627 );
nand ( n15693 , n13849 , n13625 );
nor ( n15694 , n15693 , n12728 , n13537 );
not ( n15695 , n15694 );
or ( n15696 , n15692 , n15695 );
not ( n15697 , n15693 );
not ( n15698 , n15697 );
not ( n15699 , n13539 );
or ( n15700 , n15698 , n15699 );
not ( n15701 , n13627 );
nand ( n15702 , n15701 , n13849 );
nand ( n15703 , n15700 , n15702 );
not ( n15704 , n15703 );
nand ( n15705 , n15696 , n15704 );
not ( n15706 , n15705 );
nand ( n15707 , n13528 , n12563 , n12584 , n15697 );
nor ( n15708 , n15707 , n12604 );
nand ( n15709 , n15708 , n9038 );
not ( n15710 , n15707 );
nand ( n15711 , n12611 , n9024 );
and ( n15712 , n15711 , n12599 );
and ( n15713 , n15710 , n15712 );
nor ( n15714 , n15713 , n13847 );
nand ( n15715 , n15706 , n15709 , n15714 );
not ( n15716 , n15715 );
or ( n15717 , n15691 , n15716 );
nand ( n15718 , n15688 , n15686 );
not ( n15719 , n15718 );
not ( n15720 , n15719 );
not ( n15721 , n15677 );
or ( n15722 , n15720 , n15721 );
nand ( n15723 , n15675 , n15653 );
nand ( n15724 , n15722 , n15723 );
not ( n15725 , n15724 );
nand ( n15726 , n15717 , n15725 );
not ( n15727 , n15726 );
or ( n15728 , n15651 , n15727 );
nand ( n15729 , n15580 , n15604 );
or ( n15730 , n15729 , n15633 );
nand ( n15731 , n15613 , n15632 );
nand ( n15732 , n15730 , n15731 );
and ( n15733 , n15732 , n15649 );
and ( n15734 , n15638 , n15648 );
nor ( n15735 , n15733 , n15734 );
nand ( n15736 , n15728 , n15735 );
not ( n15737 , n15642 );
nand ( n15738 , n521 , n457 );
not ( n15739 , n15738 );
or ( n15740 , n8337 , n7908 );
nand ( n15741 , n15740 , n457 );
not ( n15742 , n15741 );
or ( n15743 , n15739 , n15742 );
or ( n15744 , n15741 , n15738 );
nand ( n15745 , n15743 , n15744 );
not ( n15746 , n15745 );
or ( n15747 , n15737 , n15746 );
or ( n15748 , n15745 , n15642 );
nand ( n15749 , n15747 , n15748 );
not ( n15750 , n15749 );
xor ( n15751 , n15641 , n15642 );
and ( n15752 , n15751 , n15647 );
and ( n15753 , n15641 , n15642 );
or ( n15754 , n15752 , n15753 );
not ( n15755 , n15754 );
or ( n15756 , n15750 , n15755 );
or ( n15757 , n15754 , n15749 );
nand ( n15758 , n15756 , n15757 );
xnor ( n15759 , n15736 , n15758 );
not ( n15760 , n15759 );
not ( n15761 , n15760 );
not ( n15762 , n15761 );
or ( n15763 , n15521 , n15762 );
nand ( n15764 , n495 , n15760 );
nand ( n15765 , n15763 , n15764 );
not ( n15766 , n15765 );
or ( n15767 , n15520 , n15766 );
nand ( n15768 , n6939 , n495 );
nand ( n15769 , n15767 , n15768 );
xor ( n15770 , n15519 , n15769 );
or ( n15771 , n7415 , n7517 );
nand ( n15772 , n15771 , n497 );
and ( n15773 , n489 , n12868 );
xor ( n15774 , n15772 , n15773 );
not ( n15775 , n6842 );
not ( n15776 , n491 );
not ( n15777 , n15689 );
not ( n15778 , n15777 );
not ( n15779 , n15715 );
or ( n15780 , n15778 , n15779 );
nand ( n15781 , n15780 , n15718 );
nand ( n15782 , n15723 , n15677 );
and ( n15783 , n15781 , n15782 );
not ( n15784 , n15781 );
not ( n15785 , n15782 );
and ( n15786 , n15784 , n15785 );
nor ( n15787 , n15783 , n15786 );
not ( n15788 , n15787 );
not ( n15789 , n15788 );
not ( n15790 , n15789 );
or ( n15791 , n15776 , n15790 );
nand ( n15792 , n15788 , n6892 );
nand ( n15793 , n15791 , n15792 );
not ( n15794 , n15793 );
or ( n15795 , n15775 , n15794 );
not ( n15796 , n491 );
buf ( n15797 , n15715 );
nand ( n15798 , n15777 , n15718 );
not ( n15799 , n15798 );
and ( n15800 , n15797 , n15799 );
not ( n15801 , n15797 );
and ( n15802 , n15801 , n15798 );
nor ( n15803 , n15800 , n15802 );
not ( n15804 , n15803 );
not ( n15805 , n15804 );
or ( n15806 , n15796 , n15805 );
not ( n15807 , n15804 );
nand ( n15808 , n15807 , n6892 );
nand ( n15809 , n15806 , n15808 );
nand ( n15810 , n15809 , n6719 );
nand ( n15811 , n15795 , n15810 );
and ( n15812 , n15774 , n15811 );
and ( n15813 , n15772 , n15773 );
or ( n15814 , n15812 , n15813 );
and ( n15815 , n15770 , n15814 );
and ( n15816 , n15519 , n15769 );
or ( n15817 , n15815 , n15816 );
or ( n15818 , n7326 , n6939 );
nand ( n15819 , n15818 , n495 );
not ( n15820 , n6848 );
xor ( n15821 , n489 , n15788 );
not ( n15822 , n15821 );
or ( n15823 , n15820 , n15822 );
xor ( n15824 , n489 , n15807 );
nand ( n15825 , n15824 , n6867 );
nand ( n15826 , n15823 , n15825 );
xor ( n15827 , n15819 , n15826 );
not ( n15828 , n13869 );
and ( n15829 , n489 , n15828 );
xor ( n15830 , n15827 , n15829 );
not ( n15831 , n6719 );
not ( n15832 , n15793 );
or ( n15833 , n15831 , n15832 );
not ( n15834 , n491 );
nand ( n15835 , n15729 , n15605 );
and ( n15836 , n15726 , n15835 );
not ( n15837 , n15726 );
not ( n15838 , n15835 );
and ( n15839 , n15837 , n15838 );
nor ( n15840 , n15836 , n15839 );
buf ( n15841 , n15840 );
not ( n15842 , n15841 );
or ( n15843 , n15834 , n15842 );
not ( n15844 , n15840 );
nand ( n15845 , n15844 , n6892 );
nand ( n15846 , n15843 , n15845 );
nand ( n15847 , n15846 , n6842 );
nand ( n15848 , n15833 , n15847 );
not ( n15849 , n6848 );
not ( n15850 , n15824 );
or ( n15851 , n15849 , n15850 );
xor ( n15852 , n489 , n15828 );
nand ( n15853 , n15852 , n6867 );
nand ( n15854 , n15851 , n15853 );
xor ( n15855 , n15848 , n15854 );
not ( n15856 , n7371 );
not ( n15857 , n15634 );
not ( n15858 , n15724 );
not ( n15859 , n15605 );
or ( n15860 , n15858 , n15859 );
nand ( n15861 , n15860 , n15729 );
not ( n15862 , n15861 );
or ( n15863 , n15857 , n15862 );
nand ( n15864 , n15863 , n15731 );
not ( n15865 , n15734 );
nand ( n15866 , n15865 , n15649 );
nand ( n15867 , n15864 , n15866 );
or ( n15868 , n15634 , n15866 );
or ( n15869 , n15868 , n15864 );
not ( n15870 , n15866 );
nand ( n15871 , n15870 , n15731 );
not ( n15872 , n15871 );
nand ( n15873 , n15634 , n15861 );
nand ( n15874 , n15872 , n15873 );
not ( n15875 , n15874 );
and ( n15876 , n15777 , n15677 , n15605 );
and ( n15877 , n15876 , n15634 , n15866 );
nand ( n15878 , n15877 , n15797 );
not ( n15879 , n15878 );
or ( n15880 , n15875 , n15879 );
not ( n15881 , n15877 );
nand ( n15882 , n15881 , n15876 , n15797 );
nand ( n15883 , n15880 , n15882 );
nand ( n15884 , n15867 , n15869 , n15883 );
not ( n15885 , n15884 );
buf ( n15886 , n15885 );
not ( n15887 , n15886 );
and ( n15888 , n493 , n15887 );
not ( n15889 , n493 );
and ( n15890 , n15889 , n15886 );
nor ( n15891 , n15888 , n15890 );
not ( n15892 , n15891 );
or ( n15893 , n15856 , n15892 );
not ( n15894 , n15876 );
not ( n15895 , n15797 );
or ( n15896 , n15894 , n15895 );
not ( n15897 , n15861 );
nand ( n15898 , n15896 , n15897 );
nand ( n15899 , n15634 , n15731 );
xnor ( n15900 , n15898 , n15899 );
not ( n15901 , n15900 );
and ( n15902 , n493 , n15901 );
not ( n15903 , n493 );
not ( n15904 , n15901 );
and ( n15905 , n15903 , n15904 );
or ( n15906 , n15902 , n15905 );
nand ( n15907 , n15906 , n7405 );
nand ( n15908 , n15893 , n15907 );
and ( n15909 , n15855 , n15908 );
and ( n15910 , n15848 , n15854 );
or ( n15911 , n15909 , n15910 );
xor ( n15912 , n15830 , n15911 );
not ( n15913 , n6719 );
not ( n15914 , n15846 );
or ( n15915 , n15913 , n15914 );
not ( n15916 , n491 );
not ( n15917 , n15901 );
or ( n15918 , n15916 , n15917 );
nand ( n15919 , n15904 , n6892 );
nand ( n15920 , n15918 , n15919 );
nand ( n15921 , n15920 , n6842 );
nand ( n15922 , n15915 , n15921 );
not ( n15923 , n7371 );
and ( n15924 , n493 , n15761 );
not ( n15925 , n493 );
and ( n15926 , n15925 , n15760 );
nor ( n15927 , n15924 , n15926 );
not ( n15928 , n15927 );
or ( n15929 , n15923 , n15928 );
nand ( n15930 , n15891 , n7405 );
nand ( n15931 , n15929 , n15930 );
xor ( n15932 , n15922 , n15931 );
xor ( n15933 , n15932 , n15518 );
xor ( n15934 , n15912 , n15933 );
xor ( n15935 , n15817 , n15934 );
not ( n15936 , n6848 );
not ( n15937 , n15852 );
or ( n15938 , n15936 , n15937 );
xor ( n15939 , n489 , n13634 );
nand ( n15940 , n15939 , n6867 );
nand ( n15941 , n15938 , n15940 );
not ( n15942 , n7371 );
not ( n15943 , n15906 );
or ( n15944 , n15942 , n15943 );
not ( n15945 , n493 );
not ( n15946 , n15841 );
or ( n15947 , n15945 , n15946 );
not ( n15948 , n493 );
nand ( n15949 , n15948 , n15844 );
nand ( n15950 , n15947 , n15949 );
nand ( n15951 , n7405 , n15950 );
nand ( n15952 , n15944 , n15951 );
xor ( n15953 , n15941 , n15952 );
and ( n15954 , n495 , n15886 );
not ( n15955 , n495 );
not ( n15956 , n15885 );
and ( n15957 , n15955 , n15956 );
or ( n15958 , n15954 , n15957 );
not ( n15959 , n15958 );
not ( n15960 , n7326 );
or ( n15961 , n15959 , n15960 );
nand ( n15962 , n15765 , n6939 );
nand ( n15963 , n15961 , n15962 );
and ( n15964 , n15953 , n15963 );
and ( n15965 , n15941 , n15952 );
or ( n15966 , n15964 , n15965 );
xor ( n15967 , n15848 , n15854 );
xor ( n15968 , n15967 , n15908 );
xor ( n15969 , n15966 , n15968 );
not ( n15970 , n6867 );
xor ( n15971 , n489 , n12868 );
not ( n15972 , n15971 );
or ( n15973 , n15970 , n15972 );
nand ( n15974 , n15939 , n6848 );
nand ( n15975 , n15973 , n15974 );
and ( n15976 , n489 , n12737 );
not ( n15977 , n7405 );
and ( n15978 , n493 , n15789 );
not ( n15979 , n493 );
buf ( n15980 , n15787 );
not ( n15981 , n15980 );
and ( n15982 , n15979 , n15981 );
or ( n15983 , n15978 , n15982 );
not ( n15984 , n15983 );
or ( n15985 , n15977 , n15984 );
nand ( n15986 , n15950 , n7371 );
nand ( n15987 , n15985 , n15986 );
xor ( n15988 , n15976 , n15987 );
not ( n15989 , n6719 );
not ( n15990 , n491 );
not ( n15991 , n13851 );
not ( n15992 , n13864 );
or ( n15993 , n15991 , n15992 );
nand ( n15994 , n15993 , n13867 );
not ( n15995 , n15994 );
not ( n15996 , n15995 );
or ( n15997 , n15990 , n15996 );
nand ( n15998 , n13872 , n6892 );
nand ( n15999 , n15997 , n15998 );
not ( n16000 , n15999 );
or ( n16001 , n15989 , n16000 );
nand ( n16002 , n15809 , n6842 );
nand ( n16003 , n16001 , n16002 );
and ( n16004 , n15988 , n16003 );
and ( n16005 , n15976 , n15987 );
or ( n16006 , n16004 , n16005 );
xor ( n16007 , n15975 , n16006 );
xor ( n16008 , n15772 , n15773 );
xor ( n16009 , n16008 , n15811 );
and ( n16010 , n16007 , n16009 );
and ( n16011 , n15975 , n16006 );
or ( n16012 , n16010 , n16011 );
and ( n16013 , n15969 , n16012 );
and ( n16014 , n15966 , n15968 );
or ( n16015 , n16013 , n16014 );
xor ( n16016 , n15935 , n16015 );
not ( n16017 , n16016 );
xor ( n16018 , n15519 , n15769 );
xor ( n16019 , n16018 , n15814 );
xor ( n16020 , n15966 , n15968 );
xor ( n16021 , n16020 , n16012 );
xor ( n16022 , n16019 , n16021 );
not ( n16023 , n6939 );
not ( n16024 , n15958 );
or ( n16025 , n16023 , n16024 );
and ( n16026 , n495 , n15901 );
not ( n16027 , n495 );
and ( n16028 , n16027 , n15904 );
or ( n16029 , n16026 , n16028 );
nand ( n16030 , n16029 , n7326 );
nand ( n16031 , n16025 , n16030 );
not ( n16032 , n7415 );
and ( n16033 , n497 , n15761 );
not ( n16034 , n497 );
and ( n16035 , n16034 , n15760 );
nor ( n16036 , n16033 , n16035 );
not ( n16037 , n16036 );
or ( n16038 , n16032 , n16037 );
nand ( n16039 , n16038 , n13236 );
xor ( n16040 , n16031 , n16039 );
not ( n16041 , n15975 );
and ( n16042 , n16040 , n16041 );
and ( n16043 , n16031 , n16039 );
or ( n16044 , n16042 , n16043 );
xor ( n16045 , n15941 , n15952 );
xor ( n16046 , n16045 , n15963 );
xor ( n16047 , n16044 , n16046 );
xor ( n16048 , n15975 , n16006 );
xor ( n16049 , n16048 , n16009 );
and ( n16050 , n16047 , n16049 );
and ( n16051 , n16044 , n16046 );
or ( n16052 , n16050 , n16051 );
and ( n16053 , n16022 , n16052 );
and ( n16054 , n16019 , n16021 );
or ( n16055 , n16053 , n16054 );
not ( n16056 , n16055 );
and ( n16057 , n16017 , n16056 );
xor ( n16058 , n16019 , n16021 );
xor ( n16059 , n16058 , n16052 );
or ( n16060 , n7558 , n7813 );
nand ( n16061 , n16060 , n499 );
not ( n16062 , n6848 );
not ( n16063 , n15971 );
or ( n16064 , n16062 , n16063 );
xor ( n16065 , n489 , n12737 );
nand ( n16066 , n16065 , n6867 );
nand ( n16067 , n16064 , n16066 );
xor ( n16068 , n16061 , n16067 );
and ( n16069 , n13971 , n489 );
and ( n16070 , n16068 , n16069 );
and ( n16071 , n16061 , n16067 );
or ( n16072 , n16070 , n16071 );
not ( n16073 , n7371 );
not ( n16074 , n15983 );
or ( n16075 , n16073 , n16074 );
and ( n16076 , n493 , n15804 );
not ( n16077 , n493 );
and ( n16078 , n16077 , n15807 );
or ( n16079 , n16076 , n16078 );
nand ( n16080 , n16079 , n7405 );
nand ( n16081 , n16075 , n16080 );
not ( n16082 , n13080 );
nand ( n16083 , n16082 , n489 );
not ( n16084 , n16083 );
xor ( n16085 , n16081 , n16084 );
not ( n16086 , n6842 );
not ( n16087 , n15999 );
or ( n16088 , n16086 , n16087 );
not ( n16089 , n491 );
not ( n16090 , n13634 );
not ( n16091 , n16090 );
or ( n16092 , n16089 , n16091 );
nand ( n16093 , n13634 , n6892 );
nand ( n16094 , n16092 , n16093 );
nand ( n16095 , n16094 , n6719 );
nand ( n16096 , n16088 , n16095 );
and ( n16097 , n16085 , n16096 );
and ( n16098 , n16081 , n16084 );
or ( n16099 , n16097 , n16098 );
xor ( n16100 , n16072 , n16099 );
xor ( n16101 , n15976 , n15987 );
xor ( n16102 , n16101 , n16003 );
and ( n16103 , n16100 , n16102 );
and ( n16104 , n16072 , n16099 );
or ( n16105 , n16103 , n16104 );
xor ( n16106 , n16044 , n16046 );
xor ( n16107 , n16106 , n16049 );
xor ( n16108 , n16105 , n16107 );
xor ( n16109 , n16031 , n16039 );
xor ( n16110 , n16109 , n16041 );
not ( n16111 , n6939 );
not ( n16112 , n16029 );
or ( n16113 , n16111 , n16112 );
not ( n16114 , n495 );
not ( n16115 , n15841 );
or ( n16116 , n16114 , n16115 );
not ( n16117 , n495 );
nand ( n16118 , n16117 , n15844 );
nand ( n16119 , n16116 , n16118 );
nand ( n16120 , n16119 , n7326 );
nand ( n16121 , n16113 , n16120 );
not ( n16122 , n7517 );
not ( n16123 , n16036 );
or ( n16124 , n16122 , n16123 );
and ( n16125 , n497 , n15886 );
not ( n16126 , n497 );
and ( n16127 , n16126 , n15956 );
or ( n16128 , n16125 , n16127 );
nand ( n16129 , n16128 , n7415 );
nand ( n16130 , n16124 , n16129 );
xor ( n16131 , n16121 , n16130 );
not ( n16132 , n16094 );
not ( n16133 , n6842 );
or ( n16134 , n16132 , n16133 );
nand ( n16135 , n13957 , n491 );
not ( n16136 , n16135 );
nand ( n16137 , n12868 , n6892 );
not ( n16138 , n16137 );
or ( n16139 , n16136 , n16138 );
nand ( n16140 , n16139 , n6719 );
nand ( n16141 , n16134 , n16140 );
not ( n16142 , n6848 );
not ( n16143 , n16065 );
or ( n16144 , n16142 , n16143 );
not ( n16145 , n489 );
not ( n16146 , n13968 );
or ( n16147 , n16145 , n16146 );
nand ( n16148 , n13167 , n4046 );
nand ( n16149 , n16147 , n16148 );
nand ( n16150 , n16149 , n6867 );
nand ( n16151 , n16144 , n16150 );
xor ( n16152 , n16141 , n16151 );
not ( n16153 , n7326 );
and ( n16154 , n495 , n15789 );
not ( n16155 , n495 );
and ( n16156 , n16155 , n15981 );
or ( n16157 , n16154 , n16156 );
not ( n16158 , n16157 );
or ( n16159 , n16153 , n16158 );
nand ( n16160 , n16119 , n8841 );
nand ( n16161 , n16159 , n16160 );
and ( n16162 , n16152 , n16161 );
and ( n16163 , n16141 , n16151 );
or ( n16164 , n16162 , n16163 );
and ( n16165 , n16131 , n16164 );
and ( n16166 , n16121 , n16130 );
or ( n16167 , n16165 , n16166 );
xor ( n16168 , n16110 , n16167 );
xor ( n16169 , n16061 , n16067 );
xor ( n16170 , n16169 , n16069 );
xor ( n16171 , n16081 , n16084 );
xor ( n16172 , n16171 , n16096 );
xor ( n16173 , n16170 , n16172 );
not ( n16174 , n7371 );
not ( n16175 , n16079 );
or ( n16176 , n16174 , n16175 );
and ( n16177 , n493 , n15995 );
not ( n16178 , n493 );
and ( n16179 , n16178 , n13872 );
or ( n16180 , n16177 , n16179 );
nand ( n16181 , n16180 , n7405 );
nand ( n16182 , n16176 , n16181 );
xor ( n16183 , n16182 , n16083 );
not ( n16184 , n7517 );
not ( n16185 , n16128 );
or ( n16186 , n16184 , n16185 );
and ( n16187 , n497 , n15901 );
not ( n16188 , n497 );
and ( n16189 , n16188 , n15904 );
or ( n16190 , n16187 , n16189 );
nand ( n16191 , n16190 , n7415 );
nand ( n16192 , n16186 , n16191 );
and ( n16193 , n16183 , n16192 );
and ( n16194 , n16182 , n16083 );
or ( n16195 , n16193 , n16194 );
and ( n16196 , n16173 , n16195 );
and ( n16197 , n16170 , n16172 );
or ( n16198 , n16196 , n16197 );
and ( n16199 , n16168 , n16198 );
and ( n16200 , n16110 , n16167 );
or ( n16201 , n16199 , n16200 );
and ( n16202 , n16108 , n16201 );
and ( n16203 , n16105 , n16107 );
or ( n16204 , n16202 , n16203 );
nor ( n16205 , n16059 , n16204 );
nor ( n16206 , n16057 , n16205 );
not ( n16207 , n16206 );
xor ( n16208 , n16072 , n16099 );
xor ( n16209 , n16208 , n16102 );
xor ( n16210 , n16110 , n16167 );
xor ( n16211 , n16210 , n16198 );
xor ( n16212 , n16209 , n16211 );
or ( n16213 , n8297 , n7828 );
nand ( n16214 , n16213 , n501 );
and ( n16215 , n13060 , n489 );
xor ( n16216 , n16214 , n16215 );
nand ( n16217 , n9046 , n489 );
not ( n16218 , n16217 );
and ( n16219 , n16216 , n16218 );
and ( n16220 , n16214 , n16215 );
or ( n16221 , n16219 , n16220 );
not ( n16222 , n7558 );
not ( n16223 , n15759 );
and ( n16224 , n499 , n16223 );
not ( n16225 , n499 );
and ( n16226 , n16225 , n15759 );
or ( n16227 , n16224 , n16226 );
not ( n16228 , n16227 );
or ( n16229 , n16222 , n16228 );
nand ( n16230 , n16229 , n7818 );
xor ( n16231 , n16221 , n16230 );
not ( n16232 , n6842 );
nand ( n16233 , n16137 , n16135 );
not ( n16234 , n16233 );
or ( n16235 , n16232 , n16234 );
not ( n16236 , n491 );
not ( n16237 , n12737 );
not ( n16238 , n16237 );
or ( n16239 , n16236 , n16238 );
or ( n16240 , n16237 , n491 );
nand ( n16241 , n16239 , n16240 );
nand ( n16242 , n16241 , n6719 );
nand ( n16243 , n16235 , n16242 );
not ( n16244 , n6848 );
not ( n16245 , n16149 );
or ( n16246 , n16244 , n16245 );
not ( n16247 , n489 );
not ( n16248 , n13083 );
or ( n16249 , n16247 , n16248 );
nand ( n16250 , n13084 , n4046 );
nand ( n16251 , n16249 , n16250 );
nand ( n16252 , n16251 , n6867 );
nand ( n16253 , n16246 , n16252 );
xor ( n16254 , n16243 , n16253 );
not ( n16255 , n8841 );
not ( n16256 , n16157 );
or ( n16257 , n16255 , n16256 );
and ( n16258 , n495 , n15804 );
not ( n16259 , n495 );
and ( n16260 , n16259 , n15807 );
or ( n16261 , n16258 , n16260 );
nand ( n16262 , n16261 , n7326 );
nand ( n16263 , n16257 , n16262 );
and ( n16264 , n16254 , n16263 );
and ( n16265 , n16243 , n16253 );
or ( n16266 , n16264 , n16265 );
and ( n16267 , n16231 , n16266 );
and ( n16268 , n16221 , n16230 );
or ( n16269 , n16267 , n16268 );
xor ( n16270 , n16121 , n16130 );
xor ( n16271 , n16270 , n16164 );
xor ( n16272 , n16269 , n16271 );
xor ( n16273 , n16141 , n16151 );
xor ( n16274 , n16273 , n16161 );
not ( n16275 , n7371 );
not ( n16276 , n16180 );
or ( n16277 , n16275 , n16276 );
and ( n16278 , n493 , n16090 );
not ( n16279 , n493 );
and ( n16280 , n16279 , n13634 );
or ( n16281 , n16278 , n16280 );
nand ( n16282 , n16281 , n7405 );
nand ( n16283 , n16277 , n16282 );
not ( n16284 , n7415 );
and ( n16285 , n497 , n15841 );
not ( n16286 , n497 );
and ( n16287 , n16286 , n15844 );
or ( n16288 , n16285 , n16287 );
not ( n16289 , n16288 );
or ( n16290 , n16284 , n16289 );
nand ( n16291 , n16190 , n7517 );
nand ( n16292 , n16290 , n16291 );
xor ( n16293 , n16283 , n16292 );
not ( n16294 , n7558 );
and ( n16295 , n1665 , n15885 );
not ( n16296 , n1665 );
and ( n16297 , n16296 , n15956 );
nor ( n16298 , n16295 , n16297 );
not ( n16299 , n16298 );
or ( n16300 , n16294 , n16299 );
nand ( n16301 , n16227 , n7813 );
nand ( n16302 , n16300 , n16301 );
and ( n16303 , n16293 , n16302 );
and ( n16304 , n16283 , n16292 );
or ( n16305 , n16303 , n16304 );
xor ( n16306 , n16274 , n16305 );
xor ( n16307 , n16182 , n16083 );
xor ( n16308 , n16307 , n16192 );
and ( n16309 , n16306 , n16308 );
and ( n16310 , n16274 , n16305 );
or ( n16311 , n16309 , n16310 );
and ( n16312 , n16272 , n16311 );
and ( n16313 , n16269 , n16271 );
or ( n16314 , n16312 , n16313 );
xor ( n16315 , n16212 , n16314 );
xor ( n16316 , n16170 , n16172 );
xor ( n16317 , n16316 , n16195 );
xor ( n16318 , n16269 , n16271 );
xor ( n16319 , n16318 , n16311 );
xor ( n16320 , n16317 , n16319 );
not ( n16321 , n6867 );
not ( n16322 , n4046 );
not ( n16323 , n13058 );
or ( n16324 , n16322 , n16323 );
nand ( n16325 , n13275 , n489 );
nand ( n16326 , n16324 , n16325 );
not ( n16327 , n16326 );
or ( n16328 , n16321 , n16327 );
nand ( n16329 , n16251 , n6848 );
nand ( n16330 , n16328 , n16329 );
xor ( n16331 , n16330 , n16217 );
nand ( n16332 , n8792 , n489 );
nand ( n16333 , n8304 , n9625 );
nand ( n16334 , n16332 , n16333 );
and ( n16335 , n16331 , n16334 );
and ( n16336 , n16330 , n16217 );
or ( n16337 , n16335 , n16336 );
xor ( n16338 , n16214 , n16215 );
xor ( n16339 , n16338 , n16218 );
xor ( n16340 , n16337 , n16339 );
not ( n16341 , n7371 );
not ( n16342 , n16281 );
or ( n16343 , n16341 , n16342 );
not ( n16344 , n493 );
not ( n16345 , n12866 );
or ( n16346 , n16344 , n16345 );
not ( n16347 , n493 );
nand ( n16348 , n16347 , n12868 );
nand ( n16349 , n16346 , n16348 );
nand ( n16350 , n16349 , n7405 );
nand ( n16351 , n16343 , n16350 );
not ( n16352 , n6842 );
not ( n16353 , n16241 );
or ( n16354 , n16352 , n16353 );
not ( n16355 , n491 );
not ( n16356 , n13168 );
or ( n16357 , n16355 , n16356 );
nand ( n16358 , n13167 , n6892 );
nand ( n16359 , n16357 , n16358 );
nand ( n16360 , n16359 , n6719 );
nand ( n16361 , n16354 , n16360 );
xor ( n16362 , n16351 , n16361 );
not ( n16363 , n7517 );
not ( n16364 , n16288 );
or ( n16365 , n16363 , n16364 );
not ( n16366 , n497 );
not ( n16367 , n15980 );
or ( n16368 , n16366 , n16367 );
or ( n16369 , n15980 , n497 );
nand ( n16370 , n16368 , n16369 );
nand ( n16371 , n16370 , n7415 );
nand ( n16372 , n16365 , n16371 );
and ( n16373 , n16362 , n16372 );
and ( n16374 , n16351 , n16361 );
or ( n16375 , n16373 , n16374 );
and ( n16376 , n16340 , n16375 );
and ( n16377 , n16337 , n16339 );
or ( n16378 , n16376 , n16377 );
xor ( n16379 , n16221 , n16230 );
xor ( n16380 , n16379 , n16266 );
xor ( n16381 , n16378 , n16380 );
xor ( n16382 , n16243 , n16253 );
xor ( n16383 , n16382 , n16263 );
xor ( n16384 , n16283 , n16292 );
xor ( n16385 , n16384 , n16302 );
xor ( n16386 , n16383 , n16385 );
not ( n16387 , n7326 );
and ( n16388 , n495 , n15995 );
not ( n16389 , n495 );
and ( n16390 , n16389 , n15828 );
or ( n16391 , n16388 , n16390 );
not ( n16392 , n16391 );
or ( n16393 , n16387 , n16392 );
nand ( n16394 , n16261 , n8841 );
nand ( n16395 , n16393 , n16394 );
not ( n16396 , n7813 );
not ( n16397 , n16298 );
or ( n16398 , n16396 , n16397 );
and ( n16399 , n499 , n15901 );
not ( n16400 , n499 );
xnor ( n16401 , n15898 , n15899 );
and ( n16402 , n16400 , n16401 );
or ( n16403 , n16399 , n16402 );
nand ( n16404 , n16403 , n7558 );
nand ( n16405 , n16398 , n16404 );
xor ( n16406 , n16395 , n16405 );
not ( n16407 , n8594 );
not ( n16408 , n501 );
not ( n16409 , n16223 );
or ( n16410 , n16408 , n16409 );
nand ( n16411 , n15759 , n8260 );
nand ( n16412 , n16410 , n16411 );
not ( n16413 , n16412 );
or ( n16414 , n16407 , n16413 );
nand ( n16415 , n7828 , n501 );
nand ( n16416 , n16414 , n16415 );
and ( n16417 , n16406 , n16416 );
and ( n16418 , n16395 , n16405 );
or ( n16419 , n16417 , n16418 );
and ( n16420 , n16386 , n16419 );
and ( n16421 , n16383 , n16385 );
or ( n16422 , n16420 , n16421 );
and ( n16423 , n16381 , n16422 );
and ( n16424 , n16378 , n16380 );
or ( n16425 , n16423 , n16424 );
and ( n16426 , n16320 , n16425 );
and ( n16427 , n16317 , n16319 );
or ( n16428 , n16426 , n16427 );
or ( n16429 , n16315 , n16428 );
not ( n16430 , n16429 );
xor ( n16431 , n16274 , n16305 );
xor ( n16432 , n16431 , n16308 );
xor ( n16433 , n16378 , n16380 );
xor ( n16434 , n16433 , n16422 );
xor ( n16435 , n16432 , n16434 );
xor ( n16436 , n16337 , n16339 );
xor ( n16437 , n16436 , n16375 );
not ( n16438 , n6848 );
not ( n16439 , n16326 );
or ( n16440 , n16438 , n16439 );
not ( n16441 , n489 );
not ( n16442 , n9045 );
or ( n16443 , n16441 , n16442 );
nand ( n16444 , n9046 , n4046 );
nand ( n16445 , n16443 , n16444 );
nand ( n16446 , n16445 , n6867 );
nand ( n16447 , n16440 , n16446 );
not ( n16448 , n6867 );
not ( n16449 , n489 );
not ( n16450 , n8795 );
or ( n16451 , n16449 , n16450 );
nand ( n16452 , n8792 , n4046 );
nand ( n16453 , n16451 , n16452 );
not ( n16454 , n16453 );
or ( n16455 , n16448 , n16454 );
nand ( n16456 , n16445 , n6848 );
nand ( n16457 , n16455 , n16456 );
not ( n16458 , n16457 );
nand ( n16459 , n8869 , n489 );
nor ( n16460 , n16458 , n16459 );
xor ( n16461 , n16447 , n16460 );
or ( n16462 , n16332 , n16333 );
nand ( n16463 , n16462 , n16334 );
and ( n16464 , n16461 , n16463 );
and ( n16465 , n16447 , n16460 );
or ( n16466 , n16464 , n16465 );
xor ( n16467 , n16330 , n16217 );
xor ( n16468 , n16467 , n16334 );
xor ( n16469 , n16466 , n16468 );
xor ( n16470 , n16351 , n16361 );
xor ( n16471 , n16470 , n16372 );
and ( n16472 , n16469 , n16471 );
and ( n16473 , n16466 , n16468 );
or ( n16474 , n16472 , n16473 );
xor ( n16475 , n16437 , n16474 );
and ( n16476 , n493 , n13514 );
not ( n16477 , n493 );
and ( n16478 , n16477 , n12737 );
or ( n16479 , n16476 , n16478 );
not ( n16480 , n16479 );
not ( n16481 , n7405 );
or ( n16482 , n16480 , n16481 );
nand ( n16483 , n16349 , n7371 );
nand ( n16484 , n16482 , n16483 );
not ( n16485 , n6842 );
not ( n16486 , n16359 );
or ( n16487 , n16485 , n16486 );
not ( n16488 , n491 );
not ( n16489 , n13179 );
or ( n16490 , n16488 , n16489 );
nand ( n16491 , n13079 , n6892 );
nand ( n16492 , n16490 , n16491 );
nand ( n16493 , n16492 , n6719 );
nand ( n16494 , n16487 , n16493 );
xor ( n16495 , n16484 , n16494 );
not ( n16496 , n7517 );
not ( n16497 , n16370 );
or ( n16498 , n16496 , n16497 );
not ( n16499 , n9237 );
not ( n16500 , n15803 );
or ( n16501 , n16499 , n16500 );
or ( n16502 , n15803 , n9237 );
nand ( n16503 , n16501 , n16502 );
nand ( n16504 , n16503 , n7415 );
nand ( n16505 , n16498 , n16504 );
and ( n16506 , n16495 , n16505 );
and ( n16507 , n16484 , n16494 );
or ( n16508 , n16506 , n16507 );
not ( n16509 , n8841 );
not ( n16510 , n16391 );
or ( n16511 , n16509 , n16510 );
not ( n16512 , n13633 );
and ( n16513 , n495 , n16512 );
not ( n16514 , n495 );
and ( n16515 , n16514 , n13634 );
or ( n16516 , n16513 , n16515 );
nand ( n16517 , n16516 , n7326 );
nand ( n16518 , n16511 , n16517 );
not ( n16519 , n7558 );
not ( n16520 , n499 );
not ( n16521 , n15841 );
or ( n16522 , n16520 , n16521 );
not ( n16523 , n499 );
nand ( n16524 , n16523 , n15844 );
nand ( n16525 , n16522 , n16524 );
not ( n16526 , n16525 );
or ( n16527 , n16519 , n16526 );
nand ( n16528 , n16403 , n7813 );
nand ( n16529 , n16527 , n16528 );
xor ( n16530 , n16518 , n16529 );
nand ( n16531 , n15869 , n15867 , n15883 );
and ( n16532 , n501 , n16531 );
not ( n16533 , n501 );
and ( n16534 , n16533 , n15885 );
nor ( n16535 , n16532 , n16534 );
nand ( n16536 , n16535 , n8594 );
nand ( n16537 , n16412 , n7828 );
nand ( n16538 , n16536 , n16537 );
and ( n16539 , n16530 , n16538 );
and ( n16540 , n16518 , n16529 );
or ( n16541 , n16539 , n16540 );
xor ( n16542 , n16508 , n16541 );
xor ( n16543 , n16395 , n16405 );
xor ( n16544 , n16543 , n16416 );
and ( n16545 , n16542 , n16544 );
and ( n16546 , n16508 , n16541 );
or ( n16547 , n16545 , n16546 );
and ( n16548 , n16475 , n16547 );
and ( n16549 , n16437 , n16474 );
or ( n16550 , n16548 , n16549 );
xor ( n16551 , n16435 , n16550 );
xor ( n16552 , n16383 , n16385 );
xor ( n16553 , n16552 , n16419 );
not ( n16554 , n6719 );
and ( n16555 , n13058 , n6892 );
not ( n16556 , n13058 );
and ( n16557 , n16556 , n491 );
or ( n16558 , n16555 , n16557 );
not ( n16559 , n16558 );
or ( n16560 , n16554 , n16559 );
nand ( n16561 , n16492 , n6842 );
nand ( n16562 , n16560 , n16561 );
and ( n16563 , n16453 , n6848 );
not ( n16564 , n8478 );
not ( n16565 , n4046 );
or ( n16566 , n16564 , n16565 );
or ( n16567 , n8478 , n4046 );
nand ( n16568 , n16566 , n16567 );
not ( n16569 , n16568 );
nor ( n16570 , n16569 , n7355 );
nor ( n16571 , n16563 , n16570 );
nand ( n16572 , n8254 , n489 );
nor ( n16573 , n16571 , n16572 );
xor ( n16574 , n16562 , n16573 );
not ( n16575 , n16459 );
not ( n16576 , n16457 );
or ( n16577 , n16575 , n16576 );
or ( n16578 , n16457 , n16459 );
nand ( n16579 , n16577 , n16578 );
and ( n16580 , n16574 , n16579 );
and ( n16581 , n16562 , n16573 );
or ( n16582 , n16580 , n16581 );
xor ( n16583 , n16447 , n16460 );
xor ( n16584 , n16583 , n16463 );
xor ( n16585 , n16582 , n16584 );
not ( n16586 , n495 );
not ( n16587 , n13957 );
or ( n16588 , n16586 , n16587 );
or ( n16589 , n13957 , n495 );
nand ( n16590 , n16588 , n16589 );
not ( n16591 , n16590 );
not ( n16592 , n7326 );
or ( n16593 , n16591 , n16592 );
nand ( n16594 , n16516 , n8841 );
nand ( n16595 , n16593 , n16594 );
not ( n16596 , n7371 );
not ( n16597 , n16479 );
or ( n16598 , n16596 , n16597 );
and ( n16599 , n493 , n13168 );
not ( n16600 , n493 );
and ( n16601 , n16600 , n13167 );
or ( n16602 , n16599 , n16601 );
nand ( n16603 , n16602 , n7405 );
nand ( n16604 , n16598 , n16603 );
xor ( n16605 , n16595 , n16604 );
not ( n16606 , n7558 );
and ( n16607 , n499 , n15789 );
not ( n16608 , n499 );
and ( n16609 , n16608 , n15981 );
or ( n16610 , n16607 , n16609 );
not ( n16611 , n16610 );
or ( n16612 , n16606 , n16611 );
nand ( n16613 , n16525 , n7813 );
nand ( n16614 , n16612 , n16613 );
and ( n16615 , n16605 , n16614 );
and ( n16616 , n16595 , n16604 );
or ( n16617 , n16615 , n16616 );
and ( n16618 , n16585 , n16617 );
and ( n16619 , n16582 , n16584 );
or ( n16620 , n16618 , n16619 );
xor ( n16621 , n16466 , n16468 );
xor ( n16622 , n16621 , n16471 );
xor ( n16623 , n16620 , n16622 );
xor ( n16624 , n16484 , n16494 );
xor ( n16625 , n16624 , n16505 );
not ( n16626 , n7517 );
not ( n16627 , n16503 );
or ( n16628 , n16626 , n16627 );
and ( n16629 , n497 , n15995 );
not ( n16630 , n497 );
and ( n16631 , n16630 , n15828 );
or ( n16632 , n16629 , n16631 );
nand ( n16633 , n16632 , n7415 );
nand ( n16634 , n16628 , n16633 );
not ( n16635 , n8260 );
not ( n16636 , n16401 );
or ( n16637 , n16635 , n16636 );
or ( n16638 , n16401 , n8260 );
nand ( n16639 , n16637 , n16638 );
not ( n16640 , n16639 );
not ( n16641 , n8594 );
or ( n16642 , n16640 , n16641 );
nor ( n16643 , n13674 , n501 );
and ( n16644 , n16531 , n16643 );
nor ( n16645 , n16531 , n16415 );
nor ( n16646 , n16644 , n16645 );
nand ( n16647 , n16642 , n16646 );
xor ( n16648 , n16634 , n16647 );
and ( n16649 , n489 , n9167 );
not ( n16650 , n6848 );
not ( n16651 , n16568 );
or ( n16652 , n16650 , n16651 );
not ( n16653 , n489 );
not ( n16654 , n8258 );
or ( n16655 , n16653 , n16654 );
nand ( n16656 , n8253 , n4046 );
nand ( n16657 , n16655 , n16656 );
nand ( n16658 , n16657 , n6867 );
nand ( n16659 , n16652 , n16658 );
and ( n16660 , n16649 , n16659 );
not ( n16661 , n6892 );
not ( n16662 , n9049 );
or ( n16663 , n16661 , n16662 );
nand ( n16664 , n9045 , n491 );
nand ( n16665 , n16663 , n16664 );
not ( n16666 , n16665 );
not ( n16667 , n6719 );
or ( n16668 , n16666 , n16667 );
not ( n16669 , n16558 );
or ( n16670 , n16669 , n6843 );
nand ( n16671 , n16668 , n16670 );
xor ( n16672 , n16660 , n16671 );
and ( n16673 , n16453 , n6848 );
nor ( n16674 , n16673 , n16570 );
xor ( n16675 , n16674 , n16572 );
and ( n16676 , n16672 , n16675 );
and ( n16677 , n16660 , n16671 );
or ( n16678 , n16676 , n16677 );
and ( n16679 , n16648 , n16678 );
and ( n16680 , n16634 , n16647 );
or ( n16681 , n16679 , n16680 );
xor ( n16682 , n16625 , n16681 );
xor ( n16683 , n16518 , n16529 );
xor ( n16684 , n16683 , n16538 );
and ( n16685 , n16682 , n16684 );
and ( n16686 , n16625 , n16681 );
or ( n16687 , n16685 , n16686 );
and ( n16688 , n16623 , n16687 );
and ( n16689 , n16620 , n16622 );
or ( n16690 , n16688 , n16689 );
xor ( n16691 , n16553 , n16690 );
xor ( n16692 , n16437 , n16474 );
xor ( n16693 , n16692 , n16547 );
and ( n16694 , n16691 , n16693 );
and ( n16695 , n16553 , n16690 );
or ( n16696 , n16694 , n16695 );
nand ( n16697 , n16551 , n16696 );
xor ( n16698 , n16432 , n16434 );
and ( n16699 , n16698 , n16550 );
and ( n16700 , n16432 , n16434 );
or ( n16701 , n16699 , n16700 );
xor ( n16702 , n16317 , n16319 );
xor ( n16703 , n16702 , n16425 );
nor ( n16704 , n16701 , n16703 );
or ( n16705 , n16697 , n16704 );
nand ( n16706 , n16701 , n16703 );
nand ( n16707 , n16705 , n16706 );
not ( n16708 , n16707 );
or ( n16709 , n16430 , n16708 );
nand ( n16710 , n16315 , n16428 );
nand ( n16711 , n16709 , n16710 );
xor ( n16712 , n16209 , n16211 );
and ( n16713 , n16712 , n16314 );
and ( n16714 , n16209 , n16211 );
or ( n16715 , n16713 , n16714 );
xor ( n16716 , n16105 , n16107 );
xor ( n16717 , n16716 , n16201 );
nor ( n16718 , n16715 , n16717 );
not ( n16719 , n16718 );
and ( n16720 , n16711 , n16719 );
and ( n16721 , n16715 , n16717 );
nor ( n16722 , n16720 , n16721 );
and ( n16723 , n13652 , n13775 );
nor ( n16724 , n16723 , n13786 );
and ( n16725 , n13726 , n13416 );
nand ( n16726 , n16725 , n13763 , n15514 );
and ( n16727 , n16724 , n16726 );
xor ( n16728 , n13878 , n13882 );
and ( n16729 , n16728 , n13887 );
and ( n16730 , n13878 , n13882 );
or ( n16731 , n16729 , n16730 );
xor ( n16732 , n13934 , n13978 );
and ( n16733 , n16732 , n13983 );
and ( n16734 , n13934 , n13978 );
or ( n16735 , n16733 , n16734 );
xor ( n16736 , n16731 , n16735 );
xor ( n16737 , n13955 , n13965 );
and ( n16738 , n16737 , n13977 );
and ( n16739 , n13955 , n13965 );
or ( n16740 , n16738 , n16739 );
not ( n16741 , n8594 );
not ( n16742 , n13961 );
or ( n16743 , n16741 , n16742 );
not ( n16744 , n8260 );
not ( n16745 , n13634 );
or ( n16746 , n16744 , n16745 );
nand ( n16747 , n16512 , n501 );
nand ( n16748 , n16746 , n16747 );
nand ( n16749 , n16748 , n7828 );
nand ( n16750 , n16743 , n16749 );
not ( n16751 , n7558 );
not ( n16752 , n13973 );
or ( n16753 , n16751 , n16752 );
not ( n16754 , n499 );
not ( n16755 , n13514 );
or ( n16756 , n16754 , n16755 );
not ( n16757 , n499 );
nand ( n16758 , n16757 , n12737 );
nand ( n16759 , n16756 , n16758 );
nand ( n16760 , n16759 , n7813 );
nand ( n16761 , n16753 , n16760 );
xor ( n16762 , n16750 , n16761 );
not ( n16763 , n504 );
not ( n16764 , n503 );
not ( n16765 , n15804 );
or ( n16766 , n16764 , n16765 );
nand ( n16767 , n15807 , n8880 );
nand ( n16768 , n16766 , n16767 );
not ( n16769 , n16768 );
or ( n16770 , n16763 , n16769 );
nand ( n16771 , n13874 , n8306 );
nand ( n16772 , n16770 , n16771 );
xor ( n16773 , n16762 , n16772 );
xor ( n16774 , n16740 , n16773 );
not ( n16775 , n7405 );
not ( n16776 , n13940 );
or ( n16777 , n16775 , n16776 );
and ( n16778 , n493 , n8479 );
not ( n16779 , n493 );
and ( n16780 , n16779 , n8478 );
or ( n16781 , n16778 , n16780 );
nand ( n16782 , n16781 , n7371 );
nand ( n16783 , n16777 , n16782 );
not ( n16784 , n7326 );
not ( n16785 , n13950 );
or ( n16786 , n16784 , n16785 );
and ( n16787 , n495 , n9050 );
not ( n16788 , n495 );
and ( n16789 , n16788 , n9046 );
or ( n16790 , n16787 , n16789 );
nand ( n16791 , n16790 , n6939 );
nand ( n16792 , n16786 , n16791 );
xor ( n16793 , n16783 , n16792 );
xor ( n16794 , n13895 , n13905 );
and ( n16795 , n16794 , n13918 );
and ( n16796 , n13895 , n13905 );
or ( n16797 , n16795 , n16796 );
xor ( n16798 , n16793 , n16797 );
xor ( n16799 , n13919 , n13928 );
and ( n16800 , n16799 , n13933 );
and ( n16801 , n13919 , n13928 );
or ( n16802 , n16800 , n16801 );
xor ( n16803 , n16798 , n16802 );
not ( n16804 , n7415 );
not ( n16805 , n13924 );
or ( n16806 , n16804 , n16805 );
and ( n16807 , n497 , n13080 );
not ( n16808 , n497 );
and ( n16809 , n16808 , n16082 );
or ( n16810 , n16807 , n16809 );
nand ( n16811 , n16810 , n7517 );
nand ( n16812 , n16806 , n16811 );
not ( n16813 , n6842 );
not ( n16814 , n491 );
not ( n16815 , n8285 );
or ( n16816 , n16814 , n16815 );
nand ( n16817 , n9167 , n6892 );
nand ( n16818 , n16816 , n16817 );
not ( n16819 , n16818 );
or ( n16820 , n16813 , n16819 );
nand ( n16821 , n13900 , n6719 );
nand ( n16822 , n16820 , n16821 );
and ( n16823 , n13907 , n13917 );
xor ( n16824 , n16822 , n16823 );
and ( n16825 , n7511 , n489 );
not ( n16826 , n6867 );
not ( n16827 , n13913 );
or ( n16828 , n16826 , n16827 );
and ( n16829 , n7811 , n4046 );
not ( n16830 , n7811 );
and ( n16831 , n16830 , n489 );
or ( n16832 , n16829 , n16831 );
nand ( n16833 , n16832 , n6848 );
nand ( n16834 , n16828 , n16833 );
xor ( n16835 , n16825 , n16834 );
xor ( n16836 , n16824 , n16835 );
xor ( n16837 , n16812 , n16836 );
xor ( n16838 , n13935 , n13944 );
and ( n16839 , n16838 , n13954 );
and ( n16840 , n13935 , n13944 );
or ( n16841 , n16839 , n16840 );
xor ( n16842 , n16837 , n16841 );
xor ( n16843 , n16803 , n16842 );
xor ( n16844 , n16774 , n16843 );
xor ( n16845 , n16736 , n16844 );
xor ( n16846 , n13888 , n13892 );
and ( n16847 , n16846 , n13984 );
and ( n16848 , n13888 , n13892 );
or ( n16849 , n16847 , n16848 );
or ( n16850 , n16845 , n16849 );
nand ( n16851 , n16850 , n13990 );
nor ( n16852 , n16727 , n16851 );
not ( n16853 , n13991 );
not ( n16854 , n16850 );
or ( n16855 , n16853 , n16854 );
buf ( n16856 , n16845 );
nand ( n16857 , n16856 , n16849 );
nand ( n16858 , n16855 , n16857 );
or ( n16859 , n16852 , n16858 );
not ( n16860 , n7371 );
and ( n16861 , n493 , n8795 );
not ( n16862 , n493 );
and ( n16863 , n16862 , n8792 );
or ( n16864 , n16861 , n16863 );
not ( n16865 , n16864 );
or ( n16866 , n16860 , n16865 );
nand ( n16867 , n16781 , n7405 );
nand ( n16868 , n16866 , n16867 );
xor ( n16869 , n16822 , n16823 );
and ( n16870 , n16869 , n16835 );
and ( n16871 , n16822 , n16823 );
or ( n16872 , n16870 , n16871 );
xor ( n16873 , n16868 , n16872 );
and ( n16874 , n495 , n13063 );
not ( n16875 , n495 );
and ( n16876 , n16875 , n13277 );
or ( n16877 , n16874 , n16876 );
not ( n16878 , n16877 );
or ( n16879 , n16878 , n6938 );
nand ( n16880 , n16790 , n7326 );
nand ( n16881 , n16879 , n16880 );
xor ( n16882 , n16873 , n16881 );
xor ( n16883 , n16812 , n16836 );
and ( n16884 , n16883 , n16841 );
and ( n16885 , n16812 , n16836 );
or ( n16886 , n16884 , n16885 );
xor ( n16887 , n16882 , n16886 );
xor ( n16888 , n16750 , n16761 );
and ( n16889 , n16888 , n16772 );
and ( n16890 , n16750 , n16761 );
or ( n16891 , n16889 , n16890 );
and ( n16892 , n16887 , n16891 );
and ( n16893 , n16882 , n16886 );
or ( n16894 , n16892 , n16893 );
not ( n16895 , n7558 );
not ( n16896 , n16759 );
or ( n16897 , n16895 , n16896 );
not ( n16898 , n499 );
not ( n16899 , n12866 );
or ( n16900 , n16898 , n16899 );
not ( n16901 , n12859 );
not ( n16902 , n12864 );
or ( n16903 , n16901 , n16902 );
nand ( n16904 , n16903 , n1808 );
nand ( n16905 , n16900 , n16904 );
nand ( n16906 , n16905 , n7813 );
nand ( n16907 , n16897 , n16906 );
not ( n16908 , n16810 );
not ( n16909 , n7415 );
or ( n16910 , n16908 , n16909 );
not ( n16911 , n7411 );
and ( n16912 , n497 , n13168 );
not ( n16913 , n497 );
and ( n16914 , n16913 , n13167 );
or ( n16915 , n16912 , n16914 );
nand ( n16916 , n16911 , n16915 );
nand ( n16917 , n16910 , n16916 );
xor ( n16918 , n16907 , n16917 );
and ( n16919 , n16834 , n16825 );
or ( n16920 , n12900 , n12976 );
nand ( n16921 , n8254 , n12979 );
nand ( n16922 , n16818 , n6719 );
nand ( n16923 , n16920 , n16921 , n16922 );
xor ( n16924 , n16919 , n16923 );
and ( n16925 , n7677 , n489 );
not ( n16926 , n6848 );
not ( n16927 , n489 );
not ( n16928 , n9278 );
or ( n16929 , n16927 , n16928 );
nand ( n16930 , n8581 , n4046 );
nand ( n16931 , n16929 , n16930 );
not ( n16932 , n16931 );
or ( n16933 , n16926 , n16932 );
nand ( n16934 , n16832 , n6867 );
nand ( n16935 , n16933 , n16934 );
xor ( n16936 , n16925 , n16935 );
xor ( n16937 , n16924 , n16936 );
xor ( n16938 , n16918 , n16937 );
not ( n16939 , n7828 );
and ( n16940 , n501 , n13869 );
not ( n16941 , n501 );
and ( n16942 , n16941 , n15994 );
or ( n16943 , n16940 , n16942 );
not ( n16944 , n16943 );
or ( n16945 , n16939 , n16944 );
nand ( n16946 , n16748 , n8594 );
nand ( n16947 , n16945 , n16946 );
xor ( n16948 , n16783 , n16792 );
and ( n16949 , n16948 , n16797 );
and ( n16950 , n16783 , n16792 );
or ( n16951 , n16949 , n16950 );
xor ( n16952 , n16947 , n16951 );
not ( n16953 , n8306 );
not ( n16954 , n16768 );
or ( n16955 , n16953 , n16954 );
not ( n16956 , n503 );
not ( n16957 , n15789 );
or ( n16958 , n16956 , n16957 );
nand ( n16959 , n15788 , n8880 );
nand ( n16960 , n16958 , n16959 );
nand ( n16961 , n16960 , n504 );
nand ( n16962 , n16955 , n16961 );
xor ( n16963 , n16952 , n16962 );
xor ( n16964 , n16938 , n16963 );
xor ( n16965 , n16798 , n16802 );
and ( n16966 , n16965 , n16842 );
and ( n16967 , n16798 , n16802 );
or ( n16968 , n16966 , n16967 );
and ( n16969 , n16964 , n16968 );
and ( n16970 , n16938 , n16963 );
or ( n16971 , n16969 , n16970 );
xor ( n16972 , n16894 , n16971 );
not ( n16973 , n7558 );
not ( n16974 , n16905 );
or ( n16975 , n16973 , n16974 );
and ( n16976 , n499 , n13633 );
not ( n16977 , n499 );
and ( n16978 , n16977 , n16512 );
nor ( n16979 , n16976 , n16978 );
nand ( n16980 , n16979 , n7813 );
nand ( n16981 , n16975 , n16980 );
not ( n16982 , n7517 );
and ( n16983 , n497 , n13514 );
not ( n16984 , n497 );
and ( n16985 , n16984 , n12737 );
or ( n16986 , n16983 , n16985 );
not ( n16987 , n16986 );
or ( n16988 , n16982 , n16987 );
nand ( n16989 , n16915 , n7415 );
nand ( n16990 , n16988 , n16989 );
xor ( n16991 , n16981 , n16990 );
not ( n16992 , n6719 );
not ( n16993 , n491 );
not ( n16994 , n8258 );
or ( n16995 , n16993 , n16994 );
nand ( n16996 , n8254 , n6892 );
nand ( n16997 , n16995 , n16996 );
not ( n16998 , n16997 );
or ( n16999 , n16992 , n16998 );
not ( n17000 , n8478 );
nand ( n17001 , n17000 , n491 );
not ( n17002 , n17001 );
nand ( n17003 , n8478 , n6892 );
not ( n17004 , n17003 );
or ( n17005 , n17002 , n17004 );
nand ( n17006 , n17005 , n6842 );
nand ( n17007 , n16999 , n17006 );
and ( n17008 , n16935 , n16925 );
xor ( n17009 , n17007 , n17008 );
not ( n17010 , n8589 );
nand ( n17011 , n17010 , n489 );
not ( n17012 , n17011 );
xor ( n17013 , n489 , n9167 );
not ( n17014 , n17013 );
not ( n17015 , n6848 );
or ( n17016 , n17014 , n17015 );
nand ( n17017 , n6867 , n16931 );
nand ( n17018 , n17016 , n17017 );
not ( n17019 , n17018 );
or ( n17020 , n17012 , n17019 );
or ( n17021 , n17018 , n17011 );
nand ( n17022 , n17020 , n17021 );
xor ( n17023 , n17009 , n17022 );
xor ( n17024 , n16991 , n17023 );
not ( n17025 , n7828 );
and ( n17026 , n8260 , n15804 );
not ( n17027 , n8260 );
and ( n17028 , n17027 , n15807 );
nor ( n17029 , n17026 , n17028 );
not ( n17030 , n17029 );
or ( n17031 , n17025 , n17030 );
nand ( n17032 , n16943 , n8297 );
nand ( n17033 , n17031 , n17032 );
not ( n17034 , n8306 );
not ( n17035 , n16960 );
or ( n17036 , n17034 , n17035 );
and ( n17037 , n503 , n15841 );
not ( n17038 , n503 );
and ( n17039 , n17038 , n15844 );
nor ( n17040 , n17037 , n17039 );
not ( n17041 , n17040 );
nand ( n17042 , n17041 , n504 );
nand ( n17043 , n17036 , n17042 );
xor ( n17044 , n17033 , n17043 );
xor ( n17045 , n16868 , n16872 );
and ( n17046 , n17045 , n16881 );
and ( n17047 , n16868 , n16872 );
or ( n17048 , n17046 , n17047 );
xor ( n17049 , n17044 , n17048 );
xor ( n17050 , n17024 , n17049 );
not ( n17051 , n7405 );
not ( n17052 , n16864 );
or ( n17053 , n17051 , n17052 );
and ( n17054 , n493 , n9050 );
not ( n17055 , n493 );
and ( n17056 , n17055 , n9049 );
or ( n17057 , n17054 , n17056 );
nand ( n17058 , n17057 , n7371 );
nand ( n17059 , n17053 , n17058 );
xor ( n17060 , n16919 , n16923 );
and ( n17061 , n17060 , n16936 );
and ( n17062 , n16919 , n16923 );
or ( n17063 , n17061 , n17062 );
xor ( n17064 , n17059 , n17063 );
not ( n17065 , n7326 );
not ( n17066 , n16877 );
or ( n17067 , n17065 , n17066 );
and ( n17068 , n495 , n13179 );
not ( n17069 , n495 );
and ( n17070 , n17069 , n13084 );
or ( n17071 , n17068 , n17070 );
nand ( n17072 , n17071 , n8841 );
nand ( n17073 , n17067 , n17072 );
xor ( n17074 , n17064 , n17073 );
xor ( n17075 , n16907 , n16917 );
and ( n17076 , n17075 , n16937 );
and ( n17077 , n16907 , n16917 );
or ( n17078 , n17076 , n17077 );
xor ( n17079 , n17074 , n17078 );
xor ( n17080 , n16947 , n16951 );
and ( n17081 , n17080 , n16962 );
and ( n17082 , n16947 , n16951 );
or ( n17083 , n17081 , n17082 );
xor ( n17084 , n17079 , n17083 );
xor ( n17085 , n17050 , n17084 );
xor ( n17086 , n16972 , n17085 );
xor ( n17087 , n16882 , n16886 );
xor ( n17088 , n17087 , n16891 );
xor ( n17089 , n16938 , n16963 );
xor ( n17090 , n17089 , n16968 );
xor ( n17091 , n17088 , n17090 );
xor ( n17092 , n16740 , n16773 );
and ( n17093 , n17092 , n16843 );
and ( n17094 , n16740 , n16773 );
or ( n17095 , n17093 , n17094 );
and ( n17096 , n17091 , n17095 );
and ( n17097 , n17088 , n17090 );
or ( n17098 , n17096 , n17097 );
nor ( n17099 , n17086 , n17098 );
xor ( n17100 , n17088 , n17090 );
xor ( n17101 , n17100 , n17095 );
xor ( n17102 , n16731 , n16735 );
and ( n17103 , n17102 , n16844 );
and ( n17104 , n16731 , n16735 );
or ( n17105 , n17103 , n17104 );
nor ( n17106 , n17101 , n17105 );
nor ( n17107 , n17099 , n17106 );
nand ( n17108 , n16859 , n17107 );
not ( n17109 , n17099 );
and ( n17110 , n17101 , n17105 );
and ( n17111 , n17109 , n17110 );
and ( n17112 , n17086 , n17098 );
nor ( n17113 , n17111 , n17112 );
nand ( n17114 , n17108 , n17113 );
xor ( n17115 , n16508 , n16541 );
xor ( n17116 , n17115 , n16544 );
xor ( n17117 , n16620 , n16622 );
xor ( n17118 , n17117 , n16687 );
xor ( n17119 , n17116 , n17118 );
not ( n17120 , n8306 );
xor ( n17121 , n503 , n15759 );
not ( n17122 , n17121 );
or ( n17123 , n17120 , n17122 );
nand ( n17124 , n17123 , n9625 );
xor ( n17125 , n16562 , n16573 );
xor ( n17126 , n17125 , n16579 );
xor ( n17127 , n17124 , n17126 );
and ( n17128 , n16512 , n497 );
not ( n17129 , n16512 );
and ( n17130 , n17129 , n1009 );
or ( n17131 , n17128 , n17130 );
nand ( n17132 , n17131 , n7414 );
nand ( n17133 , n13228 , n13872 );
not ( n17134 , n13236 );
nand ( n17135 , n17134 , n13869 );
nand ( n17136 , n17132 , n17133 , n17135 );
not ( n17137 , n6719 );
and ( n17138 , n491 , n8795 );
not ( n17139 , n491 );
and ( n17140 , n17139 , n8792 );
or ( n17141 , n17138 , n17140 );
not ( n17142 , n17141 );
or ( n17143 , n17137 , n17142 );
and ( n17144 , n9049 , n12979 );
nor ( n17145 , n9046 , n12976 );
nor ( n17146 , n17144 , n17145 );
nand ( n17147 , n17143 , n17146 );
not ( n17148 , n6848 );
not ( n17149 , n16657 );
or ( n17150 , n17148 , n17149 );
nand ( n17151 , n17013 , n6867 );
nand ( n17152 , n17150 , n17151 );
not ( n17153 , n17152 );
not ( n17154 , n9278 );
nand ( n17155 , n17154 , n489 );
nor ( n17156 , n17153 , n17155 );
xor ( n17157 , n17147 , n17156 );
not ( n17158 , n16649 );
not ( n17159 , n17158 );
not ( n17160 , n16659 );
or ( n17161 , n17159 , n17160 );
or ( n17162 , n16659 , n17158 );
nand ( n17163 , n17161 , n17162 );
and ( n17164 , n17157 , n17163 );
and ( n17165 , n17147 , n17156 );
or ( n17166 , n17164 , n17165 );
xor ( n17167 , n17136 , n17166 );
not ( n17168 , n7813 );
not ( n17169 , n16610 );
or ( n17170 , n17168 , n17169 );
and ( n17171 , n499 , n15804 );
not ( n17172 , n499 );
and ( n17173 , n17172 , n15807 );
or ( n17174 , n17171 , n17173 );
nand ( n17175 , n17174 , n7558 );
nand ( n17176 , n17170 , n17175 );
and ( n17177 , n17167 , n17176 );
and ( n17178 , n17136 , n17166 );
or ( n17179 , n17177 , n17178 );
and ( n17180 , n17127 , n17179 );
and ( n17181 , n17124 , n17126 );
or ( n17182 , n17180 , n17181 );
xor ( n17183 , n16582 , n16584 );
xor ( n17184 , n17183 , n16617 );
xor ( n17185 , n17182 , n17184 );
xor ( n17186 , n16625 , n16681 );
xor ( n17187 , n17186 , n16684 );
and ( n17188 , n17185 , n17187 );
and ( n17189 , n17182 , n17184 );
or ( n17190 , n17188 , n17189 );
and ( n17191 , n17119 , n17190 );
and ( n17192 , n17116 , n17118 );
or ( n17193 , n17191 , n17192 );
not ( n17194 , n17193 );
xor ( n17195 , n16553 , n16690 );
xor ( n17196 , n17195 , n16693 );
not ( n17197 , n17196 );
nand ( n17198 , n17194 , n17197 );
xor ( n17199 , n16595 , n16604 );
xor ( n17200 , n17199 , n16614 );
not ( n17201 , n16590 );
not ( n17202 , n8841 );
or ( n17203 , n17201 , n17202 );
and ( n17204 , n12737 , n495 );
not ( n17205 , n12737 );
and ( n17206 , n17205 , n1554 );
nor ( n17207 , n17204 , n17206 );
nand ( n17208 , n17207 , n7326 );
nand ( n17209 , n17203 , n17208 );
not ( n17210 , n7371 );
not ( n17211 , n16602 );
or ( n17212 , n17210 , n17211 );
and ( n17213 , n493 , n13083 );
not ( n17214 , n493 );
and ( n17215 , n17214 , n13084 );
or ( n17216 , n17213 , n17215 );
nand ( n17217 , n17216 , n7405 );
nand ( n17218 , n17212 , n17217 );
xor ( n17219 , n17209 , n17218 );
not ( n17220 , n8594 );
not ( n17221 , n501 );
not ( n17222 , n15841 );
or ( n17223 , n17221 , n17222 );
or ( n17224 , n15841 , n501 );
nand ( n17225 , n17223 , n17224 );
not ( n17226 , n17225 );
or ( n17227 , n17220 , n17226 );
not ( n17228 , n15901 );
and ( n17229 , n17228 , n16643 );
not ( n17230 , n16415 );
and ( n17231 , n15901 , n17230 );
nor ( n17232 , n17229 , n17231 );
nand ( n17233 , n17227 , n17232 );
and ( n17234 , n17219 , n17233 );
and ( n17235 , n17209 , n17218 );
or ( n17236 , n17234 , n17235 );
xor ( n17237 , n17200 , n17236 );
not ( n17238 , n504 );
not ( n17239 , n17121 );
or ( n17240 , n17238 , n17239 );
not ( n17241 , n503 );
not ( n17242 , n15885 );
or ( n17243 , n17241 , n17242 );
nand ( n17244 , n16531 , n8880 );
nand ( n17245 , n17243 , n17244 );
nand ( n17246 , n17245 , n8306 );
nand ( n17247 , n17240 , n17246 );
not ( n17248 , n7371 );
not ( n17249 , n17216 );
or ( n17250 , n17248 , n17249 );
and ( n17251 , n493 , n13059 );
not ( n17252 , n493 );
and ( n17253 , n17252 , n13058 );
or ( n17254 , n17251 , n17253 );
nand ( n17255 , n17254 , n7405 );
nand ( n17256 , n17250 , n17255 );
not ( n17257 , n8841 );
not ( n17258 , n17207 );
or ( n17259 , n17257 , n17258 );
nor ( n17260 , n13221 , n495 );
and ( n17261 , n13167 , n17260 );
nand ( n17262 , n7326 , n495 );
nor ( n17263 , n13167 , n17262 );
nor ( n17264 , n17261 , n17263 );
nand ( n17265 , n17259 , n17264 );
xor ( n17266 , n17256 , n17265 );
not ( n17267 , n7415 );
and ( n17268 , n497 , n12866 );
not ( n17269 , n497 );
and ( n17270 , n17269 , n12868 );
or ( n17271 , n17268 , n17270 );
not ( n17272 , n17271 );
or ( n17273 , n17267 , n17272 );
nand ( n17274 , n17131 , n7517 );
nand ( n17275 , n17273 , n17274 );
and ( n17276 , n17266 , n17275 );
and ( n17277 , n17256 , n17265 );
or ( n17278 , n17276 , n17277 );
xor ( n17279 , n17247 , n17278 );
xor ( n17280 , n16660 , n16671 );
xor ( n17281 , n17280 , n16675 );
and ( n17282 , n17279 , n17281 );
and ( n17283 , n17247 , n17278 );
or ( n17284 , n17282 , n17283 );
and ( n17285 , n17237 , n17284 );
and ( n17286 , n17200 , n17236 );
or ( n17287 , n17285 , n17286 );
xor ( n17288 , n16634 , n16647 );
xor ( n17289 , n17288 , n16678 );
xor ( n17290 , n17124 , n17126 );
xor ( n17291 , n17290 , n17179 );
xor ( n17292 , n17289 , n17291 );
xor ( n17293 , n17209 , n17218 );
xor ( n17294 , n17293 , n17233 );
nor ( n17295 , n8296 , n8260 );
nand ( n17296 , n15789 , n17295 );
nand ( n17297 , n15841 , n17230 );
nand ( n17298 , n15844 , n16643 );
nand ( n17299 , n15788 , n9436 );
nand ( n17300 , n17296 , n17297 , n17298 , n17299 );
not ( n17301 , n17018 );
nor ( n17302 , n17301 , n17011 );
not ( n17303 , n6842 );
not ( n17304 , n17141 );
or ( n17305 , n17303 , n17304 );
not ( n17306 , n17003 );
not ( n17307 , n17001 );
or ( n17308 , n17306 , n17307 );
nand ( n17309 , n17308 , n6719 );
nand ( n17310 , n17305 , n17309 );
xor ( n17311 , n17302 , n17310 );
not ( n17312 , n17155 );
not ( n17313 , n17152 );
or ( n17314 , n17312 , n17313 );
or ( n17315 , n17152 , n17155 );
nand ( n17316 , n17314 , n17315 );
and ( n17317 , n17311 , n17316 );
and ( n17318 , n17302 , n17310 );
or ( n17319 , n17317 , n17318 );
xor ( n17320 , n17300 , n17319 );
and ( n17321 , n499 , n15995 );
not ( n17322 , n499 );
and ( n17323 , n17322 , n15828 );
or ( n17324 , n17321 , n17323 );
not ( n17325 , n17324 );
or ( n17326 , n17325 , n7557 );
not ( n17327 , n17174 );
or ( n17328 , n17327 , n7814 );
nand ( n17329 , n17326 , n17328 );
and ( n17330 , n17320 , n17329 );
and ( n17331 , n17300 , n17319 );
or ( n17332 , n17330 , n17331 );
xor ( n17333 , n17294 , n17332 );
xor ( n17334 , n17136 , n17166 );
xor ( n17335 , n17334 , n17176 );
and ( n17336 , n17333 , n17335 );
and ( n17337 , n17294 , n17332 );
or ( n17338 , n17336 , n17337 );
and ( n17339 , n17292 , n17338 );
and ( n17340 , n17289 , n17291 );
or ( n17341 , n17339 , n17340 );
xor ( n17342 , n17287 , n17341 );
xor ( n17343 , n17182 , n17184 );
xor ( n17344 , n17343 , n17187 );
xor ( n17345 , n17342 , n17344 );
not ( n17346 , n17345 );
xor ( n17347 , n17200 , n17236 );
xor ( n17348 , n17347 , n17284 );
xor ( n17349 , n17289 , n17291 );
xor ( n17350 , n17349 , n17338 );
xor ( n17351 , n17348 , n17350 );
not ( n17352 , n8306 );
not ( n17353 , n17228 );
not ( n17354 , n8880 );
or ( n17355 , n17353 , n17354 );
nand ( n17356 , n15901 , n503 );
nand ( n17357 , n17355 , n17356 );
not ( n17358 , n17357 );
or ( n17359 , n17352 , n17358 );
nand ( n17360 , n17245 , n504 );
nand ( n17361 , n17359 , n17360 );
xor ( n17362 , n17147 , n17156 );
xor ( n17363 , n17362 , n17163 );
xor ( n17364 , n17361 , n17363 );
xor ( n17365 , n17007 , n17008 );
and ( n17366 , n17365 , n17022 );
and ( n17367 , n17007 , n17008 );
or ( n17368 , n17366 , n17367 );
not ( n17369 , n7371 );
not ( n17370 , n17254 );
or ( n17371 , n17369 , n17370 );
nand ( n17372 , n17057 , n7405 );
nand ( n17373 , n17371 , n17372 );
xor ( n17374 , n17368 , n17373 );
not ( n17375 , n8841 );
and ( n17376 , n495 , n13167 );
not ( n17377 , n495 );
and ( n17378 , n17377 , n13968 );
nor ( n17379 , n17376 , n17378 );
not ( n17380 , n17379 );
or ( n17381 , n17375 , n17380 );
nand ( n17382 , n17071 , n7326 );
nand ( n17383 , n17381 , n17382 );
and ( n17384 , n17374 , n17383 );
and ( n17385 , n17368 , n17373 );
or ( n17386 , n17384 , n17385 );
and ( n17387 , n17364 , n17386 );
and ( n17388 , n17361 , n17363 );
or ( n17389 , n17387 , n17388 );
xor ( n17390 , n17247 , n17278 );
xor ( n17391 , n17390 , n17281 );
xor ( n17392 , n17389 , n17391 );
xor ( n17393 , n17256 , n17265 );
xor ( n17394 , n17393 , n17275 );
not ( n17395 , n7415 );
not ( n17396 , n16986 );
or ( n17397 , n17395 , n17396 );
nand ( n17398 , n17271 , n7517 );
nand ( n17399 , n17397 , n17398 );
not ( n17400 , n15788 );
not ( n17401 , n16415 );
and ( n17402 , n17400 , n17401 );
and ( n17403 , n15807 , n9436 );
nor ( n17404 , n17402 , n17403 );
and ( n17405 , n15804 , n17295 );
not ( n17406 , n16643 );
nor ( n17407 , n17406 , n15980 );
nor ( n17408 , n17405 , n17407 );
nand ( n17409 , n17404 , n17408 );
xor ( n17410 , n17399 , n17409 );
not ( n17411 , n504 );
not ( n17412 , n17357 );
or ( n17413 , n17411 , n17412 );
or ( n17414 , n17040 , n8304 );
nand ( n17415 , n17413 , n17414 );
and ( n17416 , n17410 , n17415 );
and ( n17417 , n17399 , n17409 );
or ( n17418 , n17416 , n17417 );
xor ( n17419 , n17394 , n17418 );
not ( n17420 , n7813 );
not ( n17421 , n17324 );
or ( n17422 , n17420 , n17421 );
nand ( n17423 , n16979 , n7558 );
nand ( n17424 , n17422 , n17423 );
xor ( n17425 , n17302 , n17310 );
xor ( n17426 , n17425 , n17316 );
xor ( n17427 , n17424 , n17426 );
xor ( n17428 , n17059 , n17063 );
and ( n17429 , n17428 , n17073 );
and ( n17430 , n17059 , n17063 );
or ( n17431 , n17429 , n17430 );
and ( n17432 , n17427 , n17431 );
and ( n17433 , n17424 , n17426 );
or ( n17434 , n17432 , n17433 );
and ( n17435 , n17419 , n17434 );
and ( n17436 , n17394 , n17418 );
or ( n17437 , n17435 , n17436 );
and ( n17438 , n17392 , n17437 );
and ( n17439 , n17389 , n17391 );
or ( n17440 , n17438 , n17439 );
and ( n17441 , n17351 , n17440 );
and ( n17442 , n17348 , n17350 );
or ( n17443 , n17441 , n17442 );
not ( n17444 , n17443 );
nand ( n17445 , n17346 , n17444 );
nand ( n17446 , n17198 , n17445 );
not ( n17447 , n17446 );
xor ( n17448 , n17116 , n17118 );
xor ( n17449 , n17448 , n17190 );
xor ( n17450 , n17287 , n17341 );
and ( n17451 , n17450 , n17344 );
and ( n17452 , n17287 , n17341 );
or ( n17453 , n17451 , n17452 );
nor ( n17454 , n17449 , n17453 );
xor ( n17455 , n17348 , n17350 );
xor ( n17456 , n17455 , n17440 );
xor ( n17457 , n17294 , n17332 );
xor ( n17458 , n17457 , n17335 );
xor ( n17459 , n17389 , n17391 );
xor ( n17460 , n17459 , n17437 );
xor ( n17461 , n17458 , n17460 );
xor ( n17462 , n17300 , n17319 );
xor ( n17463 , n17462 , n17329 );
xor ( n17464 , n17361 , n17363 );
xor ( n17465 , n17464 , n17386 );
xor ( n17466 , n17463 , n17465 );
xor ( n17467 , n16981 , n16990 );
and ( n17468 , n17467 , n17023 );
and ( n17469 , n16981 , n16990 );
or ( n17470 , n17468 , n17469 );
xor ( n17471 , n17368 , n17373 );
xor ( n17472 , n17471 , n17383 );
xor ( n17473 , n17470 , n17472 );
xor ( n17474 , n17424 , n17426 );
xor ( n17475 , n17474 , n17431 );
and ( n17476 , n17473 , n17475 );
and ( n17477 , n17470 , n17472 );
or ( n17478 , n17476 , n17477 );
and ( n17479 , n17466 , n17478 );
and ( n17480 , n17463 , n17465 );
or ( n17481 , n17479 , n17480 );
and ( n17482 , n17461 , n17481 );
and ( n17483 , n17458 , n17460 );
or ( n17484 , n17482 , n17483 );
nor ( n17485 , n17456 , n17484 );
nor ( n17486 , n17454 , n17485 );
xor ( n17487 , n17458 , n17460 );
xor ( n17488 , n17487 , n17481 );
not ( n17489 , n17488 );
xor ( n17490 , n17394 , n17418 );
xor ( n17491 , n17490 , n17434 );
xor ( n17492 , n17033 , n17043 );
and ( n17493 , n17492 , n17048 );
and ( n17494 , n17033 , n17043 );
or ( n17495 , n17493 , n17494 );
xor ( n17496 , n17399 , n17409 );
xor ( n17497 , n17496 , n17415 );
xor ( n17498 , n17495 , n17497 );
xor ( n17499 , n17074 , n17078 );
and ( n17500 , n17499 , n17083 );
and ( n17501 , n17074 , n17078 );
or ( n17502 , n17500 , n17501 );
and ( n17503 , n17498 , n17502 );
and ( n17504 , n17495 , n17497 );
or ( n17505 , n17503 , n17504 );
xor ( n17506 , n17491 , n17505 );
xor ( n17507 , n17463 , n17465 );
xor ( n17508 , n17507 , n17478 );
and ( n17509 , n17506 , n17508 );
and ( n17510 , n17491 , n17505 );
or ( n17511 , n17509 , n17510 );
not ( n17512 , n17511 );
nand ( n17513 , n17489 , n17512 );
xor ( n17514 , n17470 , n17472 );
xor ( n17515 , n17514 , n17475 );
xor ( n17516 , n17495 , n17497 );
xor ( n17517 , n17516 , n17502 );
xor ( n17518 , n17515 , n17517 );
xor ( n17519 , n17024 , n17049 );
and ( n17520 , n17519 , n17084 );
and ( n17521 , n17024 , n17049 );
or ( n17522 , n17520 , n17521 );
xor ( n17523 , n17518 , n17522 );
xor ( n17524 , n16894 , n16971 );
and ( n17525 , n17524 , n17085 );
and ( n17526 , n16894 , n16971 );
or ( n17527 , n17525 , n17526 );
nor ( n17528 , n17523 , n17527 );
xor ( n17529 , n17491 , n17505 );
xor ( n17530 , n17529 , n17508 );
xor ( n17531 , n17515 , n17517 );
and ( n17532 , n17531 , n17522 );
and ( n17533 , n17515 , n17517 );
or ( n17534 , n17532 , n17533 );
nor ( n17535 , n17530 , n17534 );
nor ( n17536 , n17528 , n17535 );
nand ( n17537 , n17513 , n17536 );
not ( n17538 , n17537 );
nand ( n17539 , n17114 , n17447 , n17486 , n17538 );
nand ( n17540 , n17449 , n17453 );
nand ( n17541 , n17345 , n17443 );
and ( n17542 , n17540 , n17541 );
not ( n17543 , n17542 );
and ( n17544 , n17456 , n17484 );
nand ( n17545 , n17544 , n17445 );
not ( n17546 , n17545 );
or ( n17547 , n17543 , n17546 );
nor ( n17548 , n17196 , n17193 );
nor ( n17549 , n17454 , n17548 );
nand ( n17550 , n17547 , n17549 );
nand ( n17551 , n17539 , n17550 );
nand ( n17552 , n17488 , n17511 );
nand ( n17553 , n17530 , n17534 );
and ( n17554 , n17552 , n17553 );
nand ( n17555 , n17523 , n17527 );
not ( n17556 , n17555 );
not ( n17557 , n17530 );
not ( n17558 , n17534 );
nand ( n17559 , n17557 , n17558 );
nand ( n17560 , n17556 , n17559 );
nand ( n17561 , n17554 , n17560 );
nor ( n17562 , n17548 , n17485 );
nand ( n17563 , n17561 , n17562 );
not ( n17564 , n17449 );
not ( n17565 , n17453 );
nand ( n17566 , n17564 , n17565 );
nand ( n17567 , n17566 , n17445 , n17513 );
or ( n17568 , n17563 , n17567 );
nand ( n17569 , n17196 , n17193 );
nand ( n17570 , n17568 , n17569 );
or ( n17571 , n17551 , n17570 );
nor ( n17572 , n16551 , n16696 );
nor ( n17573 , n16701 , n16703 );
nor ( n17574 , n17572 , n17573 );
nand ( n17575 , n17574 , n16429 );
nor ( n17576 , n17575 , n16718 );
nand ( n17577 , n17571 , n17576 );
nand ( n17578 , n16722 , n17577 );
not ( n17579 , n17578 );
or ( n17580 , n16207 , n17579 );
nor ( n17581 , n16055 , n16016 );
nand ( n17582 , n16204 , n16059 );
or ( n17583 , n17581 , n17582 );
nand ( n17584 , n16055 , n16016 );
nand ( n17585 , n17583 , n17584 );
buf ( n17586 , n17585 );
not ( n17587 , n17586 );
nand ( n17588 , n17580 , n17587 );
and ( n17589 , n489 , n15807 );
not ( n17590 , n6842 );
not ( n17591 , n491 );
not ( n17592 , n15886 );
or ( n17593 , n17591 , n17592 );
nand ( n17594 , n15887 , n6892 );
nand ( n17595 , n17593 , n17594 );
not ( n17596 , n17595 );
or ( n17597 , n17590 , n17596 );
nand ( n17598 , n15920 , n6719 );
nand ( n17599 , n17597 , n17598 );
xor ( n17600 , n17589 , n17599 );
not ( n17601 , n7405 );
not ( n17602 , n15927 );
or ( n17603 , n17601 , n17602 );
nand ( n17604 , n17603 , n13032 );
xor ( n17605 , n17600 , n17604 );
not ( n17606 , n489 );
not ( n17607 , n15841 );
or ( n17608 , n17606 , n17607 );
nand ( n17609 , n15844 , n4046 );
nand ( n17610 , n17608 , n17609 );
not ( n17611 , n17610 );
not ( n17612 , n17611 );
not ( n17613 , n6898 );
and ( n17614 , n17612 , n17613 );
and ( n17615 , n15821 , n6867 );
nor ( n17616 , n17614 , n17615 );
xor ( n17617 , n15819 , n15826 );
and ( n17618 , n17617 , n15829 );
and ( n17619 , n15819 , n15826 );
or ( n17620 , n17618 , n17619 );
xor ( n17621 , n17616 , n17620 );
xor ( n17622 , n15922 , n15931 );
and ( n17623 , n17622 , n15518 );
and ( n17624 , n15922 , n15931 );
or ( n17625 , n17623 , n17624 );
xor ( n17626 , n17621 , n17625 );
xor ( n17627 , n17605 , n17626 );
xor ( n17628 , n15830 , n15911 );
and ( n17629 , n17628 , n15933 );
and ( n17630 , n15830 , n15911 );
or ( n17631 , n17629 , n17630 );
xor ( n17632 , n17627 , n17631 );
xor ( n17633 , n15817 , n15934 );
and ( n17634 , n17633 , n16015 );
and ( n17635 , n15817 , n15934 );
or ( n17636 , n17634 , n17635 );
or ( n17637 , n17632 , n17636 );
nand ( n17638 , n17636 , n17632 );
nand ( n17639 , n17637 , n17638 );
not ( n17640 , n17639 );
and ( n17641 , n17588 , n17640 );
not ( n17642 , n17588 );
and ( n17643 , n17642 , n17639 );
nor ( n17644 , n17641 , n17643 );
nand ( n17645 , n17644 , n9907 );
not ( n17646 , n454 );
buf ( n17647 , n15170 );
buf ( n17648 , n15292 );
not ( n17649 , n17648 );
and ( n17650 , n17647 , n17649 );
not ( n17651 , n15269 );
not ( n17652 , n14927 );
nand ( n17653 , n11924 , n11942 );
not ( n17654 , n17653 );
or ( n17655 , n17652 , n17654 );
buf ( n17656 , n15285 );
nand ( n17657 , n17655 , n17656 );
not ( n17658 , n17657 );
or ( n17659 , n17651 , n17658 );
buf ( n17660 , n15286 );
nand ( n17661 , n17659 , n17660 );
xor ( n17662 , n17650 , n17661 );
not ( n17663 , n17662 );
or ( n17664 , n17646 , n17663 );
not ( n17665 , n17106 );
not ( n17666 , n17665 );
not ( n17667 , n16851 );
not ( n17668 , n17667 );
not ( n17669 , n13788 );
or ( n17670 , n17668 , n17669 );
not ( n17671 , n16858 );
nand ( n17672 , n17670 , n17671 );
not ( n17673 , n17672 );
or ( n17674 , n17666 , n17673 );
not ( n17675 , n17110 );
nand ( n17676 , n17674 , n17675 );
not ( n17677 , n17109 );
nor ( n17678 , n17677 , n17112 );
and ( n17679 , n17676 , n17678 );
not ( n17680 , n17676 );
not ( n17681 , n17678 );
and ( n17682 , n17680 , n17681 );
nor ( n17683 , n17679 , n17682 );
nand ( n17684 , n17683 , n9907 );
nand ( n17685 , n17664 , n17684 );
not ( n17686 , n456 );
not ( n17687 , n17449 );
nand ( n17688 , n17687 , n17565 );
not ( n17689 , n17688 );
not ( n17690 , n17345 );
and ( n17691 , n17690 , n17444 );
not ( n17692 , n17456 );
not ( n17693 , n17484 );
and ( n17694 , n17692 , n17693 );
nor ( n17695 , n17691 , n17694 );
not ( n17696 , n17695 );
not ( n17697 , n17114 );
and ( n17698 , n17513 , n17536 );
not ( n17699 , n17698 );
or ( n17700 , n17697 , n17699 );
nand ( n17701 , n17561 , n17513 );
nand ( n17702 , n17700 , n17701 );
not ( n17703 , n17702 );
or ( n17704 , n17696 , n17703 );
nand ( n17705 , n17541 , n17545 );
not ( n17706 , n17705 );
nand ( n17707 , n17704 , n17706 );
not ( n17708 , n17707 );
or ( n17709 , n17689 , n17708 );
buf ( n17710 , n17540 );
nand ( n17711 , n17709 , n17710 );
nand ( n17712 , n17569 , n17198 );
not ( n17713 , n17712 );
and ( n17714 , n17711 , n17713 );
not ( n17715 , n17711 );
and ( n17716 , n17715 , n17712 );
nor ( n17717 , n17714 , n17716 );
not ( n17718 , n17717 );
not ( n17719 , n9907 );
or ( n17720 , n17718 , n17719 );
nand ( n17721 , n17720 , n15506 );
and ( n17722 , n17721 , n472 );
not ( n17723 , n15270 );
not ( n17724 , n15297 );
or ( n17725 , n17723 , n17724 );
buf ( n17726 , n15368 );
nand ( n17727 , n17725 , n17726 );
not ( n17728 , n15399 );
nand ( n17729 , n17727 , n17728 );
not ( n17730 , n15385 );
nand ( n17731 , n17730 , n15402 );
not ( n17732 , n15403 );
nand ( n17733 , n17731 , n17732 );
not ( n17734 , n17733 );
nand ( n17735 , n17729 , n17734 );
not ( n17736 , n17735 );
and ( n17737 , n17727 , n17733 , n17728 );
not ( n17738 , n454 );
nor ( n17739 , n17737 , n17738 );
not ( n17740 , n17739 );
or ( n17741 , n17736 , n17740 );
not ( n17742 , n17484 );
nand ( n17743 , n17742 , n17692 );
not ( n17744 , n17544 );
nand ( n17745 , n17743 , n17744 );
not ( n17746 , n17745 );
and ( n17747 , n17702 , n17746 );
not ( n17748 , n17702 );
and ( n17749 , n17748 , n17745 );
nor ( n17750 , n17747 , n17749 );
nand ( n17751 , n9907 , n17750 );
nand ( n17752 , n17741 , n17751 );
and ( n17753 , n17752 , n470 );
not ( n17754 , n9907 );
not ( n17755 , n17743 );
not ( n17756 , n17702 );
or ( n17757 , n17755 , n17756 );
nand ( n17758 , n17757 , n17744 );
not ( n17759 , n17345 );
nand ( n17760 , n17759 , n17444 );
nand ( n17761 , n17760 , n17541 );
not ( n17762 , n17761 );
and ( n17763 , n17758 , n17762 );
not ( n17764 , n17758 );
and ( n17765 , n17764 , n17761 );
nor ( n17766 , n17763 , n17765 );
not ( n17767 , n17766 );
or ( n17768 , n17754 , n17767 );
not ( n17769 , n17729 );
nand ( n17770 , n15404 , n15407 );
buf ( n17771 , n17770 );
nand ( n17772 , n17769 , n17771 , n17732 );
not ( n17773 , n17770 );
nand ( n17774 , n17729 , n17731 , n17773 );
not ( n17775 , n17732 );
and ( n17776 , n17775 , n17773 );
not ( n17777 , n454 );
nor ( n17778 , n17776 , n17777 );
not ( n17779 , n17731 );
nand ( n17780 , n17779 , n17771 , n17732 );
nand ( n17781 , n17772 , n17774 , n17778 , n17780 );
nand ( n17782 , n17768 , n17781 );
nand ( n17783 , n17782 , n471 );
not ( n17784 , n17783 );
xor ( n17785 , n17753 , n17784 );
not ( n17786 , n454 );
not ( n17787 , n15392 );
not ( n17788 , n15298 );
or ( n17789 , n17787 , n17788 );
nand ( n17790 , n17789 , n15408 );
nand ( n17791 , n15413 , n14794 );
not ( n17792 , n17791 );
and ( n17793 , n17790 , n17792 );
not ( n17794 , n17790 );
and ( n17795 , n17794 , n17791 );
nor ( n17796 , n17793 , n17795 );
not ( n17797 , n17796 );
or ( n17798 , n17786 , n17797 );
nand ( n17799 , n17688 , n17540 );
not ( n17800 , n17799 );
not ( n17801 , n17707 );
or ( n17802 , n17800 , n17801 );
not ( n17803 , n17695 );
not ( n17804 , n17702 );
or ( n17805 , n17803 , n17804 );
nor ( n17806 , n17799 , n17705 );
nand ( n17807 , n17805 , n17806 );
nand ( n17808 , n17802 , n17807 );
nand ( n17809 , n17808 , n9907 );
nand ( n17810 , n17798 , n17809 );
and ( n17811 , n17810 , n472 );
and ( n17812 , n17785 , n17811 );
and ( n17813 , n17753 , n17784 );
or ( n17814 , n17812 , n17813 );
xor ( n17815 , n17722 , n17814 );
and ( n17816 , n17752 , n469 );
and ( n17817 , n17810 , n471 );
xor ( n17818 , n17816 , n17817 );
and ( n17819 , n17782 , n470 );
xor ( n17820 , n17818 , n17819 );
xor ( n17821 , n17815 , n17820 );
not ( n17822 , n454 );
not ( n17823 , n17559 );
nor ( n17824 , n17823 , n17528 );
not ( n17825 , n17824 );
buf ( n17826 , n17114 );
not ( n17827 , n17826 );
or ( n17828 , n17825 , n17827 );
buf ( n17829 , n17553 );
and ( n17830 , n17560 , n17829 );
nand ( n17831 , n17828 , n17830 );
nand ( n17832 , n17513 , n17552 );
xnor ( n17833 , n17831 , n17832 );
nand ( n17834 , n17822 , n17833 );
or ( n17835 , n15362 , n15366 );
not ( n17836 , n17835 );
buf ( n17837 , n15298 );
not ( n17838 , n17837 );
or ( n17839 , n17836 , n17838 );
buf ( n17840 , n15396 );
nand ( n17841 , n17839 , n17840 );
not ( n17842 , n15395 );
nand ( n17843 , n17842 , n15398 );
and ( n17844 , n17843 , n454 );
and ( n17845 , n17841 , n17844 );
not ( n17846 , n17841 );
not ( n17847 , n17843 );
and ( n17848 , n17847 , n454 );
and ( n17849 , n17846 , n17848 );
nor ( n17850 , n17845 , n17849 );
nand ( n17851 , n17834 , n17850 );
and ( n17852 , n17851 , n469 );
and ( n17853 , n17752 , n471 );
not ( n17854 , n17528 );
not ( n17855 , n17854 );
not ( n17856 , n17826 );
or ( n17857 , n17855 , n17856 );
nand ( n17858 , n17857 , n17555 );
nand ( n17859 , n17559 , n17829 );
xnor ( n17860 , n17858 , n17859 );
not ( n17861 , n17860 );
not ( n17862 , n9907 );
or ( n17863 , n17861 , n17862 );
not ( n17864 , n17837 );
nand ( n17865 , n17835 , n17840 );
buf ( n17866 , n17865 );
nand ( n17867 , n17864 , n17866 );
not ( n17868 , n17865 );
nand ( n17869 , n17837 , n17868 );
nand ( n17870 , n17867 , n17869 , n454 );
nand ( n17871 , n17863 , n17870 );
not ( n17872 , n17871 );
not ( n17873 , n469 );
nor ( n17874 , n17872 , n17873 );
xor ( n17875 , n17853 , n17874 );
not ( n17876 , n17782 );
not ( n17877 , n472 );
nor ( n17878 , n17876 , n17877 );
and ( n17879 , n17875 , n17878 );
and ( n17880 , n17853 , n17874 );
or ( n17881 , n17879 , n17880 );
xor ( n17882 , n17852 , n17881 );
xor ( n17883 , n17753 , n17784 );
xor ( n17884 , n17883 , n17811 );
and ( n17885 , n17882 , n17884 );
and ( n17886 , n17852 , n17881 );
or ( n17887 , n17885 , n17886 );
nor ( n17888 , n17821 , n17887 );
xor ( n17889 , n17852 , n17881 );
xor ( n17890 , n17889 , n17884 );
and ( n17891 , n17851 , n470 );
and ( n17892 , n17752 , n472 );
not ( n17893 , n9907 );
nor ( n17894 , n17556 , n17528 );
xor ( n17895 , n17894 , n17826 );
not ( n17896 , n17895 );
or ( n17897 , n17893 , n17896 );
not ( n17898 , n17649 );
nand ( n17899 , n17661 , n17647 );
not ( n17900 , n17899 );
or ( n17901 , n17898 , n17900 );
not ( n17902 , n17738 );
nand ( n17903 , n15262 , n15295 );
nand ( n17904 , n17902 , n17903 );
nand ( n17905 , n17901 , n17904 );
not ( n17906 , n17903 );
not ( n17907 , n17738 );
and ( n17908 , n17906 , n17907 );
nor ( n17909 , n17908 , n17648 );
nand ( n17910 , n17899 , n17909 );
nand ( n17911 , n17905 , n17910 );
nand ( n17912 , n17897 , n17911 );
and ( n17913 , n17912 , n469 );
xor ( n17914 , n17892 , n17913 );
and ( n17915 , n17871 , n470 );
and ( n17916 , n17914 , n17915 );
and ( n17917 , n17892 , n17913 );
or ( n17918 , n17916 , n17917 );
xor ( n17919 , n17891 , n17918 );
xor ( n17920 , n17853 , n17874 );
xor ( n17921 , n17920 , n17878 );
and ( n17922 , n17919 , n17921 );
and ( n17923 , n17891 , n17918 );
or ( n17924 , n17922 , n17923 );
nand ( n17925 , n17890 , n17924 );
or ( n17926 , n17888 , n17925 );
nand ( n17927 , n17821 , n17887 );
nand ( n17928 , n17926 , n17927 );
not ( n17929 , n17928 );
and ( n17930 , n17721 , n471 );
xor ( n17931 , n17816 , n17817 );
and ( n17932 , n17931 , n17819 );
and ( n17933 , n17816 , n17817 );
or ( n17934 , n17932 , n17933 );
xor ( n17935 , n17930 , n17934 );
and ( n17936 , n17810 , n470 );
and ( n17937 , n17782 , n469 );
xor ( n17938 , n17936 , n17937 );
not ( n17939 , n9907 );
not ( n17940 , n17572 );
nand ( n17941 , n17940 , n16697 );
not ( n17942 , n17941 );
not ( n17943 , n17570 );
nand ( n17944 , n17943 , n17539 , n17550 );
not ( n17945 , n17944 );
or ( n17946 , n17942 , n17945 );
or ( n17947 , n17944 , n17941 );
nand ( n17948 , n17946 , n17947 );
not ( n17949 , n17948 );
or ( n17950 , n17939 , n17949 );
nand ( n17951 , n14794 , n15498 );
not ( n17952 , n17951 );
not ( n17953 , n17952 );
not ( n17954 , n17790 );
or ( n17955 , n17953 , n17954 );
nor ( n17956 , n15418 , n15496 );
or ( n17957 , n17956 , n15412 );
nand ( n17958 , n17957 , n15499 );
not ( n17959 , n17958 );
nand ( n17960 , n17955 , n17959 );
not ( n17961 , n17960 );
xor ( n17962 , n15423 , n15427 );
and ( n17963 , n17962 , n15452 );
and ( n17964 , n15423 , n15427 );
or ( n17965 , n17963 , n17964 );
or ( n17966 , n2376 , n3017 );
nand ( n17967 , n17966 , n545 );
and ( n17968 , n537 , n10438 );
xor ( n17969 , n17967 , n17968 );
not ( n17970 , n543 );
buf ( n17971 , n14379 );
not ( n17972 , n17971 );
not ( n17973 , n17972 );
or ( n17974 , n17970 , n17973 );
nand ( n17975 , n17971 , n2123 );
nand ( n17976 , n17974 , n17975 );
not ( n17977 , n17976 );
not ( n17978 , n2362 );
or ( n17979 , n17977 , n17978 );
nand ( n17980 , n714 , n15434 );
nand ( n17981 , n17979 , n17980 );
xor ( n17982 , n17969 , n17981 );
not ( n17983 , n14397 );
not ( n17984 , n3069 );
not ( n17985 , n11903 );
not ( n17986 , n17985 );
or ( n17987 , n17984 , n17986 );
nand ( n17988 , n539 , n11903 );
nand ( n17989 , n17987 , n17988 );
not ( n17990 , n17989 );
or ( n17991 , n17983 , n17990 );
nand ( n17992 , n15477 , n3103 );
nand ( n17993 , n17991 , n17992 );
not ( n17994 , n11729 );
not ( n17995 , n15462 );
or ( n17996 , n17994 , n17995 );
not ( n17997 , n3177 );
not ( n17998 , n11241 );
or ( n17999 , n17997 , n17998 );
nand ( n18000 , n14264 , n537 );
nand ( n18001 , n17999 , n18000 );
nand ( n18002 , n18001 , n3133 );
nand ( n18003 , n17996 , n18002 );
xor ( n18004 , n17993 , n18003 );
not ( n18005 , n3288 );
not ( n18006 , n15444 );
or ( n18007 , n18005 , n18006 );
not ( n18008 , n541 );
not ( n18009 , n14351 );
or ( n18010 , n18008 , n18009 );
nand ( n18011 , n14354 , n3023 );
nand ( n18012 , n18010 , n18011 );
nand ( n18013 , n18012 , n3955 );
nand ( n18014 , n18007 , n18013 );
xor ( n18015 , n18004 , n18014 );
xor ( n18016 , n17982 , n18015 );
not ( n18017 , n15451 );
xor ( n18018 , n15464 , n15468 );
and ( n18019 , n18018 , n15479 );
and ( n18020 , n15464 , n15468 );
or ( n18021 , n18019 , n18020 );
xor ( n18022 , n18017 , n18021 );
xor ( n18023 , n15438 , n15448 );
and ( n18024 , n18023 , n15451 );
and ( n18025 , n15438 , n15448 );
or ( n18026 , n18024 , n18025 );
xor ( n18027 , n18022 , n18026 );
xor ( n18028 , n18016 , n18027 );
xor ( n18029 , n17965 , n18028 );
xor ( n18030 , n15480 , n15484 );
and ( n18031 , n18030 , n15489 );
and ( n18032 , n15480 , n15484 );
or ( n18033 , n18031 , n18032 );
xor ( n18034 , n18029 , n18033 );
xor ( n18035 , n15453 , n15490 );
and ( n18036 , n18035 , n15495 );
and ( n18037 , n15453 , n15490 );
or ( n18038 , n18036 , n18037 );
nor ( n18039 , n18034 , n18038 );
not ( n18040 , n18039 );
nand ( n18041 , n18038 , n18034 );
and ( n18042 , n18040 , n18041 );
not ( n18043 , n18042 );
nand ( n18044 , n17961 , n18043 );
nand ( n18045 , n17960 , n18042 );
nand ( n18046 , n18044 , n18045 , n454 );
nand ( n18047 , n17950 , n18046 );
and ( n18048 , n18047 , n472 );
xor ( n18049 , n17938 , n18048 );
xor ( n18050 , n17935 , n18049 );
not ( n18051 , n18050 );
xor ( n18052 , n17722 , n17814 );
and ( n18053 , n18052 , n17820 );
and ( n18054 , n17722 , n17814 );
or ( n18055 , n18053 , n18054 );
not ( n18056 , n18055 );
and ( n18057 , n18051 , n18056 );
not ( n18058 , n14397 );
not ( n18059 , n539 );
not ( n18060 , n14416 );
or ( n18061 , n18059 , n18060 );
nand ( n18062 , n14419 , n3069 );
nand ( n18063 , n18061 , n18062 );
not ( n18064 , n18063 );
or ( n18065 , n18058 , n18064 );
nand ( n18066 , n17989 , n3103 );
nand ( n18067 , n18065 , n18066 );
nand ( n18068 , n11478 , n537 );
xor ( n18069 , n18067 , n18068 );
xor ( n18070 , n17993 , n18003 );
and ( n18071 , n18070 , n18014 );
and ( n18072 , n17993 , n18003 );
or ( n18073 , n18071 , n18072 );
xor ( n18074 , n18069 , n18073 );
xor ( n18075 , n17967 , n17968 );
and ( n18076 , n18075 , n17981 );
and ( n18077 , n17967 , n17968 );
or ( n18078 , n18076 , n18077 );
not ( n18079 , n714 );
not ( n18080 , n17976 );
or ( n18081 , n18079 , n18080 );
nand ( n18082 , n2362 , n543 );
nand ( n18083 , n18081 , n18082 );
not ( n18084 , n3186 );
xor ( n18085 , n537 , n14255 );
not ( n18086 , n18085 );
or ( n18087 , n18084 , n18086 );
nand ( n18088 , n18001 , n11729 );
nand ( n18089 , n18087 , n18088 );
xor ( n18090 , n18083 , n18089 );
not ( n18091 , n3955 );
not ( n18092 , n541 );
not ( n18093 , n14323 );
or ( n18094 , n18092 , n18093 );
nand ( n18095 , n14326 , n3023 );
nand ( n18096 , n18094 , n18095 );
not ( n18097 , n18096 );
or ( n18098 , n18091 , n18097 );
nand ( n18099 , n18012 , n3288 );
nand ( n18100 , n18098 , n18099 );
xor ( n18101 , n18090 , n18100 );
xor ( n18102 , n18078 , n18101 );
xor ( n18103 , n18017 , n18021 );
and ( n18104 , n18103 , n18026 );
and ( n18105 , n18017 , n18021 );
or ( n18106 , n18104 , n18105 );
xor ( n18107 , n18102 , n18106 );
xor ( n18108 , n18074 , n18107 );
xor ( n18109 , n17982 , n18015 );
and ( n18110 , n18109 , n18027 );
and ( n18111 , n17982 , n18015 );
or ( n18112 , n18110 , n18111 );
xor ( n18113 , n18108 , n18112 );
xor ( n18114 , n17965 , n18028 );
and ( n18115 , n18114 , n18033 );
and ( n18116 , n17965 , n18028 );
or ( n18117 , n18115 , n18116 );
nand ( n18118 , n18113 , n18117 );
not ( n18119 , n18118 );
nor ( n18120 , n18117 , n18113 );
nor ( n18121 , n18119 , n18120 );
buf ( n18122 , n18041 );
and ( n18123 , n18121 , n18122 );
nand ( n18124 , n18123 , n17961 );
not ( n18125 , n18124 );
not ( n18126 , n18040 );
nor ( n18127 , n18126 , n18121 );
and ( n18128 , n17960 , n18127 );
not ( n18129 , n18122 );
nor ( n18130 , n18129 , n18040 );
not ( n18131 , n18130 );
not ( n18132 , n18121 );
or ( n18133 , n18131 , n18132 );
or ( n18134 , n18121 , n18122 );
nand ( n18135 , n18133 , n18134 );
nor ( n18136 , n18128 , n18135 );
not ( n18137 , n18136 );
or ( n18138 , n18125 , n18137 );
nand ( n18139 , n18138 , n454 );
not ( n18140 , n17940 );
not ( n18141 , n17944 );
or ( n18142 , n18140 , n18141 );
nand ( n18143 , n18142 , n16697 );
not ( n18144 , n18143 );
not ( n18145 , n17573 );
nand ( n18146 , n18145 , n16706 );
nand ( n18147 , n18144 , n18146 );
not ( n18148 , n18146 );
nand ( n18149 , n18148 , n18143 );
nand ( n18150 , n18147 , n18149 , n9907 );
nand ( n18151 , n18139 , n18150 );
and ( n18152 , n18151 , n472 );
xor ( n18153 , n17936 , n17937 );
and ( n18154 , n18153 , n18048 );
and ( n18155 , n17936 , n17937 );
or ( n18156 , n18154 , n18155 );
xor ( n18157 , n18152 , n18156 );
not ( n18158 , n17810 );
nor ( n18159 , n18158 , n17873 );
not ( n18160 , n9907 );
not ( n18161 , n17948 );
or ( n18162 , n18160 , n18161 );
nand ( n18163 , n18162 , n18046 );
and ( n18164 , n18163 , n471 );
xor ( n18165 , n18159 , n18164 );
and ( n18166 , n17721 , n470 );
xor ( n18167 , n18165 , n18166 );
xor ( n18168 , n18157 , n18167 );
not ( n18169 , n18168 );
xor ( n18170 , n17930 , n17934 );
and ( n18171 , n18170 , n18049 );
and ( n18172 , n17930 , n17934 );
or ( n18173 , n18171 , n18172 );
not ( n18174 , n18173 );
and ( n18175 , n18169 , n18174 );
nor ( n18176 , n18057 , n18175 );
not ( n18177 , n18176 );
or ( n18178 , n17929 , n18177 );
nand ( n18179 , n18050 , n18055 );
not ( n18180 , n18179 );
nand ( n18181 , n18168 , n18173 );
not ( n18182 , n18181 );
or ( n18183 , n18180 , n18182 );
not ( n18184 , n18168 );
nand ( n18185 , n18184 , n18174 );
nand ( n18186 , n18183 , n18185 );
nand ( n18187 , n18178 , n18186 );
not ( n18188 , n18187 );
and ( n18189 , n17912 , n472 );
not ( n18190 , n13990 );
not ( n18191 , n13788 );
or ( n18192 , n18190 , n18191 );
nand ( n18193 , n18192 , n13992 );
nand ( n18194 , n16850 , n16857 );
xnor ( n18195 , n18193 , n18194 );
not ( n18196 , n18195 );
not ( n18197 , n9907 );
or ( n18198 , n18196 , n18197 );
not ( n18199 , n12203 );
not ( n18200 , n11944 );
or ( n18201 , n18199 , n18200 );
not ( n18202 , n12205 );
not ( n18203 , n14925 );
and ( n18204 , n18203 , n15279 );
not ( n18205 , n18204 );
nor ( n18206 , n18202 , n18205 );
nand ( n18207 , n18201 , n18206 );
not ( n18208 , n18204 );
nand ( n18209 , n11944 , n18208 , n12203 );
not ( n18210 , n12205 );
nand ( n18211 , n18210 , n18208 );
nand ( n18212 , n18207 , n18209 , n18211 );
nand ( n18213 , n18212 , n454 );
nand ( n18214 , n18198 , n18213 );
and ( n18215 , n18214 , n470 );
and ( n18216 , n13996 , n469 );
xor ( n18217 , n18215 , n18216 );
and ( n18218 , n17685 , n472 );
and ( n18219 , n18217 , n18218 );
and ( n18220 , n18215 , n18216 );
or ( n18221 , n18219 , n18220 );
xor ( n18222 , n18189 , n18221 );
not ( n18223 , n18195 );
not ( n18224 , n9907 );
or ( n18225 , n18223 , n18224 );
nand ( n18226 , n18225 , n18213 );
and ( n18227 , n18226 , n469 );
and ( n18228 , n17685 , n471 );
xor ( n18229 , n18227 , n18228 );
not ( n18230 , n15286 );
nor ( n18231 , n15268 , n15264 );
nor ( n18232 , n18230 , n18231 );
xor ( n18233 , n17657 , n18232 );
nand ( n18234 , n18233 , n454 );
nand ( n18235 , n17665 , n17675 );
xnor ( n18236 , n18235 , n17672 );
nand ( n18237 , n9907 , n18236 );
nand ( n18238 , n18234 , n18237 );
and ( n18239 , n18238 , n470 );
xor ( n18240 , n18229 , n18239 );
xor ( n18241 , n18222 , n18240 );
not ( n18242 , n18241 );
and ( n18243 , n18238 , n471 );
not ( n18244 , n454 );
not ( n18245 , n14020 );
not ( n18246 , n14018 );
or ( n18247 , n18245 , n18246 );
nand ( n18248 , n18247 , n14019 );
nand ( n18249 , n11917 , n11921 );
nand ( n18250 , n11923 , n18249 );
not ( n18251 , n18250 );
and ( n18252 , n18248 , n18251 );
not ( n18253 , n18248 );
and ( n18254 , n18253 , n18250 );
nor ( n18255 , n18252 , n18254 );
not ( n18256 , n18255 );
or ( n18257 , n18244 , n18256 );
nand ( n18258 , n18257 , n15517 );
and ( n18259 , n18258 , n469 );
and ( n18260 , n18226 , n471 );
xor ( n18261 , n18259 , n18260 );
and ( n18262 , n13996 , n470 );
and ( n18263 , n18261 , n18262 );
and ( n18264 , n18259 , n18260 );
or ( n18265 , n18263 , n18264 );
xor ( n18266 , n18243 , n18265 );
xor ( n18267 , n18215 , n18216 );
xor ( n18268 , n18267 , n18218 );
and ( n18269 , n18266 , n18268 );
and ( n18270 , n18243 , n18265 );
or ( n18271 , n18269 , n18270 );
not ( n18272 , n18271 );
nand ( n18273 , n18242 , n18272 );
and ( n18274 , n18238 , n472 );
and ( n18275 , n14029 , n469 );
and ( n18276 , n18258 , n470 );
xor ( n18277 , n18275 , n18276 );
and ( n18278 , n18214 , n472 );
and ( n18279 , n18277 , n18278 );
and ( n18280 , n18275 , n18276 );
or ( n18281 , n18279 , n18280 );
xor ( n18282 , n18274 , n18281 );
xor ( n18283 , n18259 , n18260 );
xor ( n18284 , n18283 , n18262 );
and ( n18285 , n18282 , n18284 );
and ( n18286 , n18274 , n18281 );
or ( n18287 , n18285 , n18286 );
xor ( n18288 , n18243 , n18265 );
xor ( n18289 , n18288 , n18268 );
nor ( n18290 , n18287 , n18289 );
xor ( n18291 , n18274 , n18281 );
xor ( n18292 , n18291 , n18284 );
and ( n18293 , n13996 , n471 );
not ( n18294 , n454 );
not ( n18295 , n11359 );
nand ( n18296 , n18295 , n11932 );
not ( n18297 , n18296 );
not ( n18298 , n11366 );
not ( n18299 , n18298 );
not ( n18300 , n10741 );
or ( n18301 , n18299 , n18300 );
buf ( n18302 , n11930 );
nand ( n18303 , n18301 , n18302 );
not ( n18304 , n18303 );
or ( n18305 , n18297 , n18304 );
or ( n18306 , n18303 , n18296 );
nand ( n18307 , n18305 , n18306 );
not ( n18308 , n18307 );
or ( n18309 , n18294 , n18308 );
nand ( n18310 , n13770 , n13774 );
not ( n18311 , n18310 );
not ( n18312 , n13725 );
not ( n18313 , n18312 );
not ( n18314 , n13763 );
or ( n18315 , n18313 , n18314 );
not ( n18316 , n13766 );
nand ( n18317 , n18315 , n18316 );
not ( n18318 , n18317 );
or ( n18319 , n18311 , n18318 );
or ( n18320 , n18317 , n18310 );
nand ( n18321 , n18319 , n18320 );
nand ( n18322 , n18321 , n9907 );
nand ( n18323 , n18309 , n18322 );
and ( n18324 , n18323 , n469 );
and ( n18325 , n14029 , n470 );
xor ( n18326 , n18324 , n18325 );
and ( n18327 , n18258 , n471 );
and ( n18328 , n18326 , n18327 );
and ( n18329 , n18324 , n18325 );
or ( n18330 , n18328 , n18329 );
xor ( n18331 , n18293 , n18330 );
xor ( n18332 , n18275 , n18276 );
xor ( n18333 , n18332 , n18278 );
and ( n18334 , n18331 , n18333 );
and ( n18335 , n18293 , n18330 );
or ( n18336 , n18334 , n18335 );
nand ( n18337 , n18292 , n18336 );
or ( n18338 , n18290 , n18337 );
nand ( n18339 , n18289 , n18287 );
nand ( n18340 , n18338 , n18339 );
and ( n18341 , n17912 , n471 );
xor ( n18342 , n18227 , n18228 );
and ( n18343 , n18342 , n18239 );
and ( n18344 , n18227 , n18228 );
or ( n18345 , n18343 , n18344 );
xor ( n18346 , n18341 , n18345 );
and ( n18347 , n17685 , n470 );
and ( n18348 , n18234 , n18237 );
nor ( n18349 , n18348 , n7074 );
xor ( n18350 , n18347 , n18349 );
and ( n18351 , n17871 , n472 );
xor ( n18352 , n18350 , n18351 );
xor ( n18353 , n18346 , n18352 );
not ( n18354 , n18353 );
xor ( n18355 , n18189 , n18221 );
and ( n18356 , n18355 , n18240 );
and ( n18357 , n18189 , n18221 );
or ( n18358 , n18356 , n18357 );
not ( n18359 , n18358 );
nand ( n18360 , n18354 , n18359 );
nand ( n18361 , n18273 , n18340 , n18360 );
not ( n18362 , n18353 );
and ( n18363 , n18362 , n18359 );
nand ( n18364 , n18241 , n18271 );
nor ( n18365 , n18363 , n18364 );
and ( n18366 , n18353 , n18358 );
nor ( n18367 , n18365 , n18366 );
nand ( n18368 , n18361 , n18367 );
xor ( n18369 , n17891 , n17918 );
xor ( n18370 , n18369 , n17921 );
not ( n18371 , n18370 );
and ( n18372 , n17851 , n471 );
and ( n18373 , n17685 , n469 );
and ( n18374 , n17871 , n471 );
xor ( n18375 , n18373 , n18374 );
and ( n18376 , n17912 , n470 );
and ( n18377 , n18375 , n18376 );
and ( n18378 , n18373 , n18374 );
or ( n18379 , n18377 , n18378 );
xor ( n18380 , n18372 , n18379 );
xor ( n18381 , n17892 , n17913 );
xor ( n18382 , n18381 , n17915 );
and ( n18383 , n18380 , n18382 );
and ( n18384 , n18372 , n18379 );
or ( n18385 , n18383 , n18384 );
not ( n18386 , n18385 );
nand ( n18387 , n18371 , n18386 );
and ( n18388 , n17834 , n17850 );
nor ( n18389 , n18388 , n6725 );
xor ( n18390 , n18347 , n18349 );
and ( n18391 , n18390 , n18351 );
and ( n18392 , n18347 , n18349 );
or ( n18393 , n18391 , n18392 );
xor ( n18394 , n18389 , n18393 );
xor ( n18395 , n18373 , n18374 );
xor ( n18396 , n18395 , n18376 );
xor ( n18397 , n18394 , n18396 );
not ( n18398 , n18397 );
xor ( n18399 , n18341 , n18345 );
and ( n18400 , n18399 , n18352 );
and ( n18401 , n18341 , n18345 );
or ( n18402 , n18400 , n18401 );
not ( n18403 , n18402 );
nand ( n18404 , n18398 , n18403 );
xor ( n18405 , n18372 , n18379 );
xor ( n18406 , n18405 , n18382 );
not ( n18407 , n18406 );
xor ( n18408 , n18389 , n18393 );
and ( n18409 , n18408 , n18396 );
and ( n18410 , n18389 , n18393 );
or ( n18411 , n18409 , n18410 );
not ( n18412 , n18411 );
nand ( n18413 , n18407 , n18412 );
nand ( n18414 , n18404 , n18413 );
not ( n18415 , n18414 );
nand ( n18416 , n18368 , n18387 , n18415 );
not ( n18417 , n18416 );
nor ( n18418 , n17821 , n17887 );
nor ( n18419 , n17890 , n17924 );
nor ( n18420 , n18418 , n18419 );
nand ( n18421 , n18176 , n18420 );
not ( n18422 , n18421 );
nand ( n18423 , n18417 , n18422 );
buf ( n18424 , n18271 );
nor ( n18425 , n18424 , n18241 );
nor ( n18426 , n18358 , n18353 );
nor ( n18427 , n18425 , n18426 );
not ( n18428 , n18289 );
not ( n18429 , n18287 );
and ( n18430 , n18428 , n18429 );
nor ( n18431 , n18292 , n18336 );
nor ( n18432 , n18430 , n18431 );
nand ( n18433 , n18427 , n18432 );
not ( n18434 , n18433 );
nand ( n18435 , n18434 , n18415 );
and ( n18436 , n13996 , n472 );
and ( n18437 , n18323 , n470 );
not ( n18438 , n454 );
nand ( n18439 , n18298 , n18302 );
xnor ( n18440 , n10741 , n18439 );
not ( n18441 , n18440 );
or ( n18442 , n18438 , n18441 );
nand ( n18443 , n18312 , n18316 );
xnor ( n18444 , n13763 , n18443 );
nand ( n18445 , n18444 , n9907 );
nand ( n18446 , n18442 , n18445 );
and ( n18447 , n18446 , n469 );
xor ( n18448 , n18437 , n18447 );
and ( n18449 , n14029 , n471 );
and ( n18450 , n18448 , n18449 );
and ( n18451 , n18437 , n18447 );
or ( n18452 , n18450 , n18451 );
xor ( n18453 , n18436 , n18452 );
xor ( n18454 , n18324 , n18325 );
xor ( n18455 , n18454 , n18327 );
xor ( n18456 , n18453 , n18455 );
not ( n18457 , n18456 );
and ( n18458 , n18258 , n472 );
not ( n18459 , n14031 );
not ( n18460 , n14030 );
or ( n18461 , n18459 , n18460 );
nand ( n18462 , n18461 , n14032 );
not ( n18463 , n13758 );
nor ( n18464 , n18463 , n13761 );
xor ( n18465 , n18462 , n18464 );
not ( n18466 , n18465 );
not ( n18467 , n9907 );
or ( n18468 , n18466 , n18467 );
or ( n18469 , n10723 , n10718 );
buf ( n18470 , n10732 );
nand ( n18471 , n18469 , n18470 );
not ( n18472 , n10739 );
nand ( n18473 , n18472 , n10736 );
not ( n18474 , n10737 );
nand ( n18475 , n18471 , n18473 , n18474 );
not ( n18476 , n18473 );
and ( n18477 , n18476 , n10737 );
nor ( n18478 , n18477 , n17777 );
nand ( n18479 , n18476 , n18470 , n18469 );
nand ( n18480 , n18475 , n18478 , n18479 );
nand ( n18481 , n18468 , n18480 );
and ( n18482 , n18481 , n469 );
and ( n18483 , n18323 , n471 );
xor ( n18484 , n18482 , n18483 );
and ( n18485 , n18446 , n470 );
and ( n18486 , n18484 , n18485 );
and ( n18487 , n18482 , n18483 );
or ( n18488 , n18486 , n18487 );
xor ( n18489 , n18458 , n18488 );
xor ( n18490 , n18437 , n18447 );
xor ( n18491 , n18490 , n18449 );
and ( n18492 , n18489 , n18491 );
and ( n18493 , n18458 , n18488 );
or ( n18494 , n18492 , n18493 );
not ( n18495 , n18494 );
nand ( n18496 , n18457 , n18495 );
not ( n18497 , n18496 );
xor ( n18498 , n18293 , n18330 );
xor ( n18499 , n18498 , n18333 );
xor ( n18500 , n18436 , n18452 );
and ( n18501 , n18500 , n18455 );
and ( n18502 , n18436 , n18452 );
or ( n18503 , n18501 , n18502 );
nor ( n18504 , n18499 , n18503 );
nor ( n18505 , n18497 , n18504 );
not ( n18506 , n18505 );
xor ( n18507 , n18458 , n18488 );
xor ( n18508 , n18507 , n18491 );
and ( n18509 , n14029 , n472 );
and ( n18510 , n18481 , n470 );
not ( n18511 , n454 );
nand ( n18512 , n18469 , n18474 );
xnor ( n18513 , n18470 , n18512 );
not ( n18514 , n18513 );
or ( n18515 , n18511 , n18514 );
nand ( n18516 , n18515 , n14035 );
and ( n18517 , n18516 , n469 );
xor ( n18518 , n18510 , n18517 );
and ( n18519 , n18323 , n472 );
and ( n18520 , n18518 , n18519 );
and ( n18521 , n18510 , n18517 );
or ( n18522 , n18520 , n18521 );
xor ( n18523 , n18509 , n18522 );
xor ( n18524 , n18482 , n18483 );
xor ( n18525 , n18524 , n18485 );
and ( n18526 , n18523 , n18525 );
and ( n18527 , n18509 , n18522 );
or ( n18528 , n18526 , n18527 );
nor ( n18529 , n18508 , n18528 );
xor ( n18530 , n18509 , n18522 );
xor ( n18531 , n18530 , n18525 );
and ( n18532 , n18446 , n471 );
and ( n18533 , n9909 , n469 );
and ( n18534 , n18481 , n471 );
xor ( n18535 , n18533 , n18534 );
and ( n18536 , n18516 , n470 );
and ( n18537 , n18535 , n18536 );
and ( n18538 , n18533 , n18534 );
or ( n18539 , n18537 , n18538 );
xor ( n18540 , n18532 , n18539 );
xor ( n18541 , n18510 , n18517 );
xor ( n18542 , n18541 , n18519 );
and ( n18543 , n18540 , n18542 );
and ( n18544 , n18532 , n18539 );
or ( n18545 , n18543 , n18544 );
nor ( n18546 , n18531 , n18545 );
nor ( n18547 , n18529 , n18546 );
not ( n18548 , n18547 );
and ( n18549 , n18516 , n471 );
not ( n18550 , n454 );
buf ( n18551 , n6135 );
nand ( n18552 , n6042 , n18551 );
not ( n18553 , n18552 );
not ( n18554 , n6701 );
not ( n18555 , n9923 );
or ( n18556 , n18554 , n18555 );
nand ( n18557 , n18556 , n6133 );
not ( n18558 , n18557 );
or ( n18559 , n18553 , n18558 );
or ( n18560 , n18557 , n18552 );
nand ( n18561 , n18559 , n18560 );
not ( n18562 , n18561 );
or ( n18563 , n18550 , n18562 );
not ( n18564 , n9931 );
not ( n18565 , n9934 );
or ( n18566 , n18564 , n18565 );
nand ( n18567 , n18566 , n9932 );
not ( n18568 , n9899 );
nand ( n18569 , n18568 , n9896 );
xnor ( n18570 , n18567 , n18569 );
nand ( n18571 , n18570 , n9907 );
nand ( n18572 , n18563 , n18571 );
and ( n18573 , n18572 , n469 );
and ( n18574 , n9909 , n471 );
xor ( n18575 , n18573 , n18574 );
and ( n18576 , n9920 , n470 );
and ( n18577 , n18575 , n18576 );
and ( n18578 , n18573 , n18574 );
or ( n18579 , n18577 , n18578 );
xor ( n18580 , n18549 , n18579 );
and ( n18581 , n9909 , n470 );
and ( n18582 , n9920 , n469 );
xor ( n18583 , n18581 , n18582 );
and ( n18584 , n18481 , n472 );
xor ( n18585 , n18583 , n18584 );
xor ( n18586 , n18580 , n18585 );
and ( n18587 , n18516 , n472 );
and ( n18588 , n9937 , n469 );
and ( n18589 , n18572 , n470 );
xor ( n18590 , n18588 , n18589 );
and ( n18591 , n9909 , n472 );
and ( n18592 , n18590 , n18591 );
and ( n18593 , n18588 , n18589 );
or ( n18594 , n18592 , n18593 );
xor ( n18595 , n18587 , n18594 );
xor ( n18596 , n18573 , n18574 );
xor ( n18597 , n18596 , n18576 );
and ( n18598 , n18595 , n18597 );
and ( n18599 , n18587 , n18594 );
or ( n18600 , n18598 , n18599 );
nor ( n18601 , n18586 , n18600 );
xor ( n18602 , n18587 , n18594 );
xor ( n18603 , n18602 , n18597 );
and ( n18604 , n9920 , n471 );
not ( n18605 , n454 );
and ( n18606 , n6138 , n6199 );
not ( n18607 , n6138 );
and ( n18608 , n18607 , n6200 );
nor ( n18609 , n18606 , n18608 );
not ( n18610 , n18609 );
not ( n18611 , n6696 );
not ( n18612 , n18611 );
or ( n18613 , n18610 , n18612 );
not ( n18614 , n6699 );
not ( n18615 , n6201 );
or ( n18616 , n18614 , n18615 );
not ( n18617 , n18611 );
nand ( n18618 , n18616 , n18617 );
nand ( n18619 , n18613 , n18618 );
not ( n18620 , n18619 );
or ( n18621 , n18605 , n18620 );
not ( n18622 , n14038 );
not ( n18623 , n9861 );
or ( n18624 , n18622 , n18623 );
nand ( n18625 , n18624 , n14039 );
not ( n18626 , n18625 );
not ( n18627 , n9891 );
nand ( n18628 , n18627 , n9888 );
not ( n18629 , n18628 );
or ( n18630 , n18626 , n18629 );
or ( n18631 , n18628 , n18625 );
nand ( n18632 , n18630 , n18631 );
nand ( n18633 , n18632 , n9907 );
nand ( n18634 , n18621 , n18633 );
and ( n18635 , n18634 , n469 );
and ( n18636 , n9937 , n470 );
xor ( n18637 , n18635 , n18636 );
and ( n18638 , n18572 , n471 );
and ( n18639 , n18637 , n18638 );
and ( n18640 , n18635 , n18636 );
or ( n18641 , n18639 , n18640 );
xor ( n18642 , n18604 , n18641 );
xor ( n18643 , n18588 , n18589 );
xor ( n18644 , n18643 , n18591 );
and ( n18645 , n18642 , n18644 );
and ( n18646 , n18604 , n18641 );
or ( n18647 , n18645 , n18646 );
nor ( n18648 , n18603 , n18647 );
nor ( n18649 , n18601 , n18648 );
not ( n18650 , n18649 );
and ( n18651 , n18572 , n472 );
not ( n18652 , n9953 );
nor ( n18653 , n18652 , n17873 );
not ( n18654 , n454 );
buf ( n18655 , n6690 );
nand ( n18656 , n18655 , n6695 );
not ( n18657 , n18656 );
not ( n18658 , n6687 );
not ( n18659 , n9944 );
or ( n18660 , n18658 , n18659 );
nand ( n18661 , n18660 , n9945 );
not ( n18662 , n18661 );
or ( n18663 , n18657 , n18662 );
or ( n18664 , n18661 , n18656 );
nand ( n18665 , n18663 , n18664 );
not ( n18666 , n18665 );
or ( n18667 , n18654 , n18666 );
nand ( n18668 , n18667 , n14042 );
not ( n18669 , n18668 );
nor ( n18670 , n18669 , n7742 );
xor ( n18671 , n18653 , n18670 );
and ( n18672 , n18634 , n471 );
and ( n18673 , n18671 , n18672 );
and ( n18674 , n18653 , n18670 );
or ( n18675 , n18673 , n18674 );
xor ( n18676 , n18651 , n18675 );
and ( n18677 , n18668 , n469 );
and ( n18678 , n18634 , n470 );
xor ( n18679 , n18677 , n18678 );
and ( n18680 , n9937 , n471 );
xor ( n18681 , n18679 , n18680 );
xor ( n18682 , n18676 , n18681 );
and ( n18683 , n9937 , n472 );
and ( n18684 , n9971 , n469 );
and ( n18685 , n9953 , n470 );
xor ( n18686 , n18684 , n18685 );
and ( n18687 , n18668 , n471 );
and ( n18688 , n18686 , n18687 );
and ( n18689 , n18684 , n18685 );
or ( n18690 , n18688 , n18689 );
xor ( n18691 , n18683 , n18690 );
xor ( n18692 , n18653 , n18670 );
xor ( n18693 , n18692 , n18672 );
and ( n18694 , n18691 , n18693 );
and ( n18695 , n18683 , n18690 );
or ( n18696 , n18694 , n18695 );
or ( n18697 , n18682 , n18696 );
and ( n18698 , n9920 , n472 );
xor ( n18699 , n18677 , n18678 );
and ( n18700 , n18699 , n18680 );
and ( n18701 , n18677 , n18678 );
or ( n18702 , n18700 , n18701 );
xor ( n18703 , n18698 , n18702 );
xor ( n18704 , n18635 , n18636 );
xor ( n18705 , n18704 , n18638 );
xor ( n18706 , n18703 , n18705 );
xor ( n18707 , n18651 , n18675 );
and ( n18708 , n18707 , n18681 );
and ( n18709 , n18651 , n18675 );
or ( n18710 , n18708 , n18709 );
nor ( n18711 , n18706 , n18710 );
not ( n18712 , n18711 );
nand ( n18713 , n18697 , n18712 );
xor ( n18714 , n18604 , n18641 );
xor ( n18715 , n18714 , n18644 );
xor ( n18716 , n18698 , n18702 );
and ( n18717 , n18716 , n18705 );
and ( n18718 , n18698 , n18702 );
or ( n18719 , n18717 , n18718 );
nor ( n18720 , n18715 , n18719 );
nor ( n18721 , n18713 , n18720 );
not ( n18722 , n18721 );
and ( n18723 , n18634 , n472 );
and ( n18724 , n9987 , n469 );
and ( n18725 , n9971 , n470 );
xor ( n18726 , n18724 , n18725 );
and ( n18727 , n9953 , n471 );
and ( n18728 , n18726 , n18727 );
and ( n18729 , n18724 , n18725 );
or ( n18730 , n18728 , n18729 );
xor ( n18731 , n18723 , n18730 );
xor ( n18732 , n18684 , n18685 );
xor ( n18733 , n18732 , n18687 );
and ( n18734 , n18731 , n18733 );
and ( n18735 , n18723 , n18730 );
or ( n18736 , n18734 , n18735 );
xor ( n18737 , n18683 , n18690 );
xor ( n18738 , n18737 , n18693 );
xor ( n18739 , n18736 , n18738 );
and ( n18740 , n10008 , n469 );
and ( n18741 , n9987 , n470 );
xor ( n18742 , n18740 , n18741 );
and ( n18743 , n9971 , n471 );
and ( n18744 , n18742 , n18743 );
and ( n18745 , n18740 , n18741 );
or ( n18746 , n18744 , n18745 );
and ( n18747 , n18668 , n472 );
xor ( n18748 , n18746 , n18747 );
xor ( n18749 , n18724 , n18725 );
xor ( n18750 , n18749 , n18727 );
and ( n18751 , n18748 , n18750 );
and ( n18752 , n18746 , n18747 );
or ( n18753 , n18751 , n18752 );
xor ( n18754 , n18723 , n18730 );
xor ( n18755 , n18754 , n18733 );
xor ( n18756 , n18753 , n18755 );
xor ( n18757 , n18746 , n18747 );
xor ( n18758 , n18757 , n18750 );
and ( n18759 , n9953 , n472 );
and ( n18760 , n10028 , n469 );
and ( n18761 , n10008 , n470 );
xor ( n18762 , n18760 , n18761 );
and ( n18763 , n9987 , n471 );
and ( n18764 , n18762 , n18763 );
and ( n18765 , n18760 , n18761 );
or ( n18766 , n18764 , n18765 );
xor ( n18767 , n18759 , n18766 );
xor ( n18768 , n18740 , n18741 );
xor ( n18769 , n18768 , n18743 );
and ( n18770 , n18767 , n18769 );
and ( n18771 , n18759 , n18766 );
or ( n18772 , n18770 , n18771 );
or ( n18773 , n18758 , n18772 );
not ( n18774 , n18773 );
xor ( n18775 , n18759 , n18766 );
xor ( n18776 , n18775 , n18769 );
and ( n18777 , n9971 , n472 );
not ( n18778 , n454 );
not ( n18779 , n6608 );
nand ( n18780 , n18779 , n6477 );
not ( n18781 , n6606 );
and ( n18782 , n18780 , n18781 );
not ( n18783 , n18780 );
and ( n18784 , n18783 , n6606 );
nor ( n18785 , n18782 , n18784 );
not ( n18786 , n18785 );
or ( n18787 , n18778 , n18786 );
nand ( n18788 , n18787 , n14045 );
and ( n18789 , n18788 , n469 );
and ( n18790 , n10028 , n470 );
xor ( n18791 , n18789 , n18790 );
and ( n18792 , n10008 , n471 );
and ( n18793 , n18791 , n18792 );
and ( n18794 , n18789 , n18790 );
or ( n18795 , n18793 , n18794 );
xor ( n18796 , n18777 , n18795 );
xor ( n18797 , n18760 , n18761 );
xor ( n18798 , n18797 , n18763 );
and ( n18799 , n18796 , n18798 );
and ( n18800 , n18777 , n18795 );
or ( n18801 , n18799 , n18800 );
or ( n18802 , n18776 , n18801 );
not ( n18803 , n18802 );
xor ( n18804 , n18777 , n18795 );
xor ( n18805 , n18804 , n18798 );
nand ( n18806 , n14037 , n15509 );
and ( n18807 , n18806 , n469 );
and ( n18808 , n18788 , n470 );
xor ( n18809 , n18807 , n18808 );
nand ( n18810 , n470 , n18806 );
nand ( n18811 , n469 , n14012 );
nor ( n18812 , n18810 , n18811 );
and ( n18813 , n18809 , n18812 );
and ( n18814 , n18807 , n18808 );
or ( n18815 , n18813 , n18814 );
and ( n18816 , n9987 , n472 );
xor ( n18817 , n18815 , n18816 );
and ( n18818 , n10028 , n471 );
and ( n18819 , n18788 , n471 );
not ( n18820 , n18810 );
not ( n18821 , n18811 );
not ( n18822 , n18821 );
or ( n18823 , n18820 , n18822 );
nand ( n18824 , n470 , n18806 , n18811 );
nand ( n18825 , n18823 , n18824 );
xor ( n18826 , n18819 , n18825 );
nand ( n18827 , n14012 , n470 );
not ( n18828 , n18827 );
not ( n18829 , n18828 );
not ( n18830 , n15509 );
not ( n18831 , n14037 );
or ( n18832 , n18830 , n18831 );
nand ( n18833 , n18832 , n471 );
nor ( n18834 , n18829 , n18833 );
and ( n18835 , n18826 , n18834 );
and ( n18836 , n18819 , n18825 );
or ( n18837 , n18835 , n18836 );
xor ( n18838 , n18818 , n18837 );
and ( n18839 , n10008 , n472 );
and ( n18840 , n18838 , n18839 );
and ( n18841 , n18818 , n18837 );
or ( n18842 , n18840 , n18841 );
and ( n18843 , n18817 , n18842 );
and ( n18844 , n18815 , n18816 );
or ( n18845 , n18843 , n18844 );
or ( n18846 , n18805 , n18845 );
not ( n18847 , n18846 );
xor ( n18848 , n18815 , n18816 );
xor ( n18849 , n18848 , n18842 );
xor ( n18850 , n18789 , n18790 );
xor ( n18851 , n18850 , n18792 );
nor ( n18852 , n18849 , n18851 );
xor ( n18853 , n18818 , n18837 );
xor ( n18854 , n18853 , n18839 );
xor ( n18855 , n18807 , n18808 );
xor ( n18856 , n18855 , n18812 );
xor ( n18857 , n18854 , n18856 );
not ( n18858 , n10028 );
nor ( n18859 , n18858 , n17877 );
xor ( n18860 , n18819 , n18825 );
xor ( n18861 , n18860 , n18834 );
xor ( n18862 , n18859 , n18861 );
nand ( n18863 , n472 , n14012 );
or ( n18864 , n18833 , n18863 );
and ( n18865 , n18788 , n472 );
not ( n18866 , n18865 );
and ( n18867 , n18864 , n18866 );
and ( n18868 , n18833 , n18828 );
not ( n18869 , n18833 );
and ( n18870 , n18869 , n18827 );
nor ( n18871 , n18868 , n18870 );
or ( n18872 , n18867 , n18871 );
or ( n18873 , n18866 , n18864 );
nand ( n18874 , n18872 , n18873 );
and ( n18875 , n18862 , n18874 );
and ( n18876 , n18859 , n18861 );
or ( n18877 , n18875 , n18876 );
and ( n18878 , n18857 , n18877 );
and ( n18879 , n18854 , n18856 );
nor ( n18880 , n18878 , n18879 );
or ( n18881 , n18852 , n18880 );
nand ( n18882 , n18849 , n18851 );
nand ( n18883 , n18881 , n18882 );
not ( n18884 , n18883 );
or ( n18885 , n18847 , n18884 );
nand ( n18886 , n18805 , n18845 );
nand ( n18887 , n18885 , n18886 );
not ( n18888 , n18887 );
or ( n18889 , n18803 , n18888 );
nand ( n18890 , n18776 , n18801 );
nand ( n18891 , n18889 , n18890 );
not ( n18892 , n18891 );
or ( n18893 , n18774 , n18892 );
nand ( n18894 , n18758 , n18772 );
nand ( n18895 , n18893 , n18894 );
and ( n18896 , n18756 , n18895 );
and ( n18897 , n18753 , n18755 );
or ( n18898 , n18896 , n18897 );
and ( n18899 , n18739 , n18898 );
and ( n18900 , n18736 , n18738 );
or ( n18901 , n18899 , n18900 );
not ( n18902 , n18901 );
or ( n18903 , n18722 , n18902 );
not ( n18904 , n18720 );
nand ( n18905 , n18682 , n18696 );
or ( n18906 , n18711 , n18905 );
nand ( n18907 , n18706 , n18710 );
nand ( n18908 , n18906 , n18907 );
and ( n18909 , n18904 , n18908 );
and ( n18910 , n18715 , n18719 );
nor ( n18911 , n18909 , n18910 );
nand ( n18912 , n18903 , n18911 );
not ( n18913 , n18912 );
or ( n18914 , n18650 , n18913 );
not ( n18915 , n18601 );
nand ( n18916 , n18647 , n18603 );
not ( n18917 , n18916 );
and ( n18918 , n18915 , n18917 );
and ( n18919 , n18586 , n18600 );
nor ( n18920 , n18918 , n18919 );
nand ( n18921 , n18914 , n18920 );
not ( n18922 , n18921 );
xor ( n18923 , n18532 , n18539 );
xor ( n18924 , n18923 , n18542 );
and ( n18925 , n18446 , n472 );
xor ( n18926 , n18581 , n18582 );
and ( n18927 , n18926 , n18584 );
and ( n18928 , n18581 , n18582 );
or ( n18929 , n18927 , n18928 );
xor ( n18930 , n18925 , n18929 );
xor ( n18931 , n18533 , n18534 );
xor ( n18932 , n18931 , n18536 );
and ( n18933 , n18930 , n18932 );
and ( n18934 , n18925 , n18929 );
or ( n18935 , n18933 , n18934 );
nor ( n18936 , n18924 , n18935 );
xor ( n18937 , n18925 , n18929 );
xor ( n18938 , n18937 , n18932 );
xor ( n18939 , n18549 , n18579 );
and ( n18940 , n18939 , n18585 );
and ( n18941 , n18549 , n18579 );
or ( n18942 , n18940 , n18941 );
nor ( n18943 , n18938 , n18942 );
nor ( n18944 , n18936 , n18943 );
not ( n18945 , n18944 );
or ( n18946 , n18922 , n18945 );
not ( n18947 , n18936 );
nand ( n18948 , n18938 , n18942 );
not ( n18949 , n18948 );
and ( n18950 , n18947 , n18949 );
and ( n18951 , n18924 , n18935 );
nor ( n18952 , n18950 , n18951 );
nand ( n18953 , n18946 , n18952 );
not ( n18954 , n18953 );
or ( n18955 , n18548 , n18954 );
not ( n18956 , n18529 );
nand ( n18957 , n18531 , n18545 );
not ( n18958 , n18957 );
and ( n18959 , n18956 , n18958 );
and ( n18960 , n18508 , n18528 );
nor ( n18961 , n18959 , n18960 );
nand ( n18962 , n18955 , n18961 );
not ( n18963 , n18962 );
or ( n18964 , n18506 , n18963 );
not ( n18965 , n18504 );
nand ( n18966 , n18456 , n18494 );
not ( n18967 , n18966 );
and ( n18968 , n18965 , n18967 );
and ( n18969 , n18499 , n18503 );
nor ( n18970 , n18968 , n18969 );
nand ( n18971 , n18964 , n18970 );
nand ( n18972 , n18387 , n18971 );
nor ( n18973 , n18435 , n18972 );
nand ( n18974 , n18973 , n18422 );
not ( n18975 , n18387 );
not ( n18976 , n18397 );
nor ( n18977 , n18976 , n18403 );
not ( n18978 , n18977 );
not ( n18979 , n18413 );
or ( n18980 , n18978 , n18979 );
buf ( n18981 , n18406 );
nand ( n18982 , n18981 , n18411 );
nand ( n18983 , n18980 , n18982 );
not ( n18984 , n18983 );
or ( n18985 , n18975 , n18984 );
buf ( n18986 , n18385 );
nand ( n18987 , n18370 , n18986 );
nand ( n18988 , n18985 , n18987 );
nand ( n18989 , n18422 , n18988 );
nand ( n18990 , n18188 , n18423 , n18974 , n18989 );
buf ( n18991 , n18990 );
not ( n18992 , n18991 );
not ( n18993 , n17575 );
not ( n18994 , n18993 );
not ( n18995 , n17944 );
or ( n18996 , n18994 , n18995 );
not ( n18997 , n16711 );
nand ( n18998 , n18996 , n18997 );
not ( n18999 , n16719 );
nor ( n19000 , n18999 , n16721 );
xor ( n19001 , n18998 , n19000 );
not ( n19002 , n19001 );
not ( n19003 , n9907 );
or ( n19004 , n19002 , n19003 );
nor ( n19005 , n18113 , n18117 );
nor ( n19006 , n19005 , n18039 );
not ( n19007 , n19006 );
nor ( n19008 , n19007 , n17951 );
xor ( n19009 , n18067 , n18068 );
and ( n19010 , n19009 , n18073 );
and ( n19011 , n18067 , n18068 );
or ( n19012 , n19010 , n19011 );
xor ( n19013 , n18083 , n18089 );
and ( n19014 , n19013 , n18100 );
and ( n19015 , n18083 , n18089 );
or ( n19016 , n19014 , n19015 );
or ( n19017 , n714 , n2362 );
nand ( n19018 , n19017 , n543 );
not ( n19019 , n3955 );
xor ( n19020 , n541 , n17971 );
not ( n19021 , n19020 );
or ( n19022 , n19019 , n19021 );
nand ( n19023 , n18096 , n3288 );
nand ( n19024 , n19022 , n19023 );
xor ( n19025 , n19018 , n19024 );
not ( n19026 , n3186 );
xor ( n19027 , n537 , n17985 );
not ( n19028 , n19027 );
or ( n19029 , n19026 , n19028 );
nand ( n19030 , n18085 , n11729 );
nand ( n19031 , n19029 , n19030 );
xor ( n19032 , n19025 , n19031 );
xor ( n19033 , n19016 , n19032 );
nor ( n19034 , n3177 , n14264 );
not ( n19035 , n3103 );
not ( n19036 , n18063 );
or ( n19037 , n19035 , n19036 );
not ( n19038 , n539 );
not ( n19039 , n14351 );
or ( n19040 , n19038 , n19039 );
nand ( n19041 , n14354 , n3069 );
nand ( n19042 , n19040 , n19041 );
nand ( n19043 , n19042 , n14397 );
nand ( n19044 , n19037 , n19043 );
xor ( n19045 , n19034 , n19044 );
not ( n19046 , n18068 );
xor ( n19047 , n19045 , n19046 );
xor ( n19048 , n19033 , n19047 );
xor ( n19049 , n19012 , n19048 );
xor ( n19050 , n18078 , n18101 );
and ( n19051 , n19050 , n18106 );
and ( n19052 , n18078 , n18101 );
or ( n19053 , n19051 , n19052 );
xor ( n19054 , n19049 , n19053 );
not ( n19055 , n19054 );
xor ( n19056 , n18074 , n18107 );
and ( n19057 , n19056 , n18112 );
and ( n19058 , n18074 , n18107 );
or ( n19059 , n19057 , n19058 );
not ( n19060 , n19059 );
nand ( n19061 , n19055 , n19060 );
nand ( n19062 , n19008 , n19061 );
not ( n19063 , n19062 );
not ( n19064 , n19063 );
not ( n19065 , n17790 );
or ( n19066 , n19064 , n19065 );
or ( n19067 , n18120 , n18041 );
nand ( n19068 , n19067 , n18118 );
nand ( n19069 , n19068 , n19061 );
nor ( n19070 , n18039 , n19005 );
nand ( n19071 , n19061 , n19070 , n17958 );
nand ( n19072 , n19054 , n19059 );
nand ( n19073 , n19069 , n19071 , n19072 );
not ( n19074 , n19073 );
nand ( n19075 , n19066 , n19074 );
buf ( n19076 , n19075 );
xor ( n19077 , n19012 , n19048 );
and ( n19078 , n19077 , n19053 );
and ( n19079 , n19012 , n19048 );
or ( n19080 , n19078 , n19079 );
and ( n19081 , n537 , n14255 );
not ( n19082 , n14397 );
and ( n19083 , n539 , n14326 );
not ( n19084 , n539 );
and ( n19085 , n19084 , n14323 );
nor ( n19086 , n19083 , n19085 );
not ( n19087 , n19086 );
or ( n19088 , n19082 , n19087 );
nand ( n19089 , n3103 , n19042 );
nand ( n19090 , n19088 , n19089 );
xor ( n19091 , n19081 , n19090 );
not ( n19092 , n11729 );
not ( n19093 , n19027 );
or ( n19094 , n19092 , n19093 );
xor ( n19095 , n14419 , n537 );
nand ( n19096 , n19095 , n3186 );
nand ( n19097 , n19094 , n19096 );
xor ( n19098 , n19091 , n19097 );
not ( n19099 , n11032 );
not ( n19100 , n3023 );
and ( n19101 , n19099 , n19100 );
and ( n19102 , n19020 , n3288 );
nor ( n19103 , n19101 , n19102 );
xor ( n19104 , n19018 , n19024 );
and ( n19105 , n19104 , n19031 );
and ( n19106 , n19018 , n19024 );
or ( n19107 , n19105 , n19106 );
xor ( n19108 , n19103 , n19107 );
xor ( n19109 , n19034 , n19044 );
and ( n19110 , n19109 , n19046 );
and ( n19111 , n19034 , n19044 );
or ( n19112 , n19110 , n19111 );
xor ( n19113 , n19108 , n19112 );
xor ( n19114 , n19098 , n19113 );
xor ( n19115 , n19016 , n19032 );
and ( n19116 , n19115 , n19047 );
and ( n19117 , n19016 , n19032 );
or ( n19118 , n19116 , n19117 );
xor ( n19119 , n19114 , n19118 );
or ( n19120 , n19080 , n19119 );
nand ( n19121 , n19119 , n19080 );
nand ( n19122 , n19120 , n19121 );
not ( n19123 , n19122 );
and ( n19124 , n19076 , n19123 );
not ( n19125 , n19076 );
and ( n19126 , n19125 , n19122 );
nor ( n19127 , n19124 , n19126 );
nand ( n19128 , n19127 , n454 );
nand ( n19129 , n19004 , n19128 );
and ( n19130 , n19129 , n472 );
and ( n19131 , n18163 , n470 );
not ( n19132 , n17721 );
nor ( n19133 , n19132 , n17873 );
xor ( n19134 , n19131 , n19133 );
not ( n19135 , n9907 );
nand ( n19136 , n16429 , n16710 );
not ( n19137 , n19136 );
not ( n19138 , n17574 );
not ( n19139 , n17944 );
or ( n19140 , n19138 , n19139 );
not ( n19141 , n16707 );
nand ( n19142 , n19140 , n19141 );
not ( n19143 , n19142 );
or ( n19144 , n19137 , n19143 );
or ( n19145 , n19136 , n19142 );
nand ( n19146 , n19144 , n19145 );
not ( n19147 , n19146 );
or ( n19148 , n19135 , n19147 );
not ( n19149 , n19008 );
not ( n19150 , n15409 );
or ( n19151 , n19149 , n19150 );
not ( n19152 , n19070 );
not ( n19153 , n17958 );
or ( n19154 , n19152 , n19153 );
not ( n19155 , n19068 );
nand ( n19156 , n19154 , n19155 );
not ( n19157 , n19156 );
nand ( n19158 , n19151 , n19157 );
nand ( n19159 , n19061 , n19072 );
not ( n19160 , n19159 );
and ( n19161 , n19158 , n19160 );
not ( n19162 , n19158 );
and ( n19163 , n19162 , n19159 );
nor ( n19164 , n19161 , n19163 );
nand ( n19165 , n19164 , n454 );
nand ( n19166 , n19148 , n19165 );
and ( n19167 , n19166 , n472 );
and ( n19168 , n19134 , n19167 );
and ( n19169 , n19131 , n19133 );
or ( n19170 , n19168 , n19169 );
xor ( n19171 , n19130 , n19170 );
and ( n19172 , n18047 , n469 );
and ( n19173 , n19166 , n471 );
xor ( n19174 , n19172 , n19173 );
nand ( n19175 , n18139 , n18150 );
and ( n19176 , n19175 , n470 );
xor ( n19177 , n19174 , n19176 );
xor ( n19178 , n19171 , n19177 );
not ( n19179 , n19178 );
not ( n19180 , n19179 );
and ( n19181 , n18151 , n471 );
xor ( n19182 , n18159 , n18164 );
and ( n19183 , n19182 , n18166 );
and ( n19184 , n18159 , n18164 );
or ( n19185 , n19183 , n19184 );
xor ( n19186 , n19181 , n19185 );
xor ( n19187 , n19131 , n19133 );
xor ( n19188 , n19187 , n19167 );
and ( n19189 , n19186 , n19188 );
and ( n19190 , n19181 , n19185 );
or ( n19191 , n19189 , n19190 );
nor ( n19192 , n19180 , n19191 );
not ( n19193 , n19192 );
nand ( n19194 , n19178 , n19191 );
buf ( n19195 , n19194 );
nand ( n19196 , n19193 , n19195 );
xor ( n19197 , n19181 , n19185 );
xor ( n19198 , n19197 , n19188 );
xor ( n19199 , n18152 , n18156 );
and ( n19200 , n19199 , n18167 );
and ( n19201 , n18152 , n18156 );
or ( n19202 , n19200 , n19201 );
nand ( n19203 , n19198 , n19202 );
not ( n19204 , n19203 );
nor ( n19205 , n19196 , n19204 );
nand ( n19206 , n18992 , n19205 );
or ( n19207 , n19198 , n19202 );
and ( n19208 , n19196 , n19207 );
nand ( n19209 , n18991 , n19208 );
not ( n19210 , n19196 );
not ( n19211 , n19207 );
nand ( n19212 , n19211 , n19203 );
not ( n19213 , n19212 );
and ( n19214 , n19210 , n19213 );
and ( n19215 , n19196 , n19204 );
nor ( n19216 , n19214 , n19215 );
and ( n19217 , n19206 , n19209 , n19216 );
and ( n19218 , n716 , n17686 );
nor ( n19219 , n19218 , n454 );
buf ( n19220 , n19219 );
not ( n19221 , n19220 );
or ( n19222 , n19217 , n19221 );
nor ( n19223 , n527 , n543 );
nor ( n19224 , n528 , n544 );
nor ( n19225 , n19223 , n19224 );
not ( n19226 , n19225 );
nand ( n19227 , n536 , n552 );
nand ( n19228 , n535 , n551 );
nand ( n19229 , n19227 , n19228 );
or ( n19230 , n535 , n551 );
nor ( n19231 , n534 , n550 );
not ( n19232 , n19231 );
nand ( n19233 , n19229 , n19230 , n19232 );
not ( n19234 , n19233 );
nand ( n19235 , n534 , n550 );
nand ( n19236 , n533 , n549 );
and ( n19237 , n19235 , n19236 );
not ( n19238 , n19237 );
or ( n19239 , n19234 , n19238 );
or ( n19240 , n531 , n547 );
or ( n19241 , n532 , n548 );
nand ( n19242 , n19240 , n19241 );
or ( n19243 , n529 , n545 );
nor ( n19244 , n533 , n549 );
not ( n19245 , n19244 );
nor ( n19246 , n530 , n546 );
not ( n19247 , n19246 );
nand ( n19248 , n19243 , n19245 , n19247 );
nor ( n19249 , n19242 , n19248 );
nand ( n19250 , n19239 , n19249 );
nand ( n19251 , n530 , n546 );
nand ( n19252 , n529 , n545 );
nand ( n19253 , n531 , n547 );
and ( n19254 , n19251 , n19252 , n19253 );
not ( n19255 , n19254 );
nand ( n19256 , n532 , n548 );
not ( n19257 , n19256 );
nand ( n19258 , n19257 , n19240 );
not ( n19259 , n19258 );
or ( n19260 , n19255 , n19259 );
not ( n19261 , n19247 );
not ( n19262 , n19243 );
or ( n19263 , n19261 , n19262 );
nand ( n19264 , n19263 , n19252 );
nand ( n19265 , n19260 , n19264 );
nand ( n19266 , n19250 , n19265 );
not ( n19267 , n19266 );
or ( n19268 , n19226 , n19267 );
nand ( n19269 , n528 , n544 );
or ( n19270 , n19223 , n19269 );
nand ( n19271 , n527 , n543 );
nand ( n19272 , n19270 , n19271 );
not ( n19273 , n19272 );
nand ( n19274 , n19268 , n19273 );
nor ( n19275 , n526 , n542 );
not ( n19276 , n19275 );
nand ( n19277 , n526 , n542 );
nand ( n19278 , n19276 , n19277 );
not ( n19279 , n19278 );
and ( n19280 , n19274 , n19279 );
not ( n19281 , n19274 );
and ( n19282 , n19281 , n19278 );
nor ( n19283 , n19280 , n19282 );
not ( n19284 , n19224 );
not ( n19285 , n19284 );
not ( n19286 , n19266 );
or ( n19287 , n19285 , n19286 );
nand ( n19288 , n19287 , n19269 );
not ( n19289 , n19271 );
nor ( n19290 , n19289 , n19223 );
xor ( n19291 , n19288 , n19290 );
xor ( n19292 , n19283 , n19291 );
not ( n19293 , n19292 );
and ( n19294 , n19225 , n19276 );
not ( n19295 , n19294 );
nand ( n19296 , n19250 , n19265 );
not ( n19297 , n19296 );
or ( n19298 , n19295 , n19297 );
and ( n19299 , n19272 , n19276 );
not ( n19300 , n19277 );
nor ( n19301 , n19299 , n19300 );
nand ( n19302 , n19298 , n19301 );
nor ( n19303 , n525 , n541 );
and ( n19304 , n525 , n541 );
nor ( n19305 , n19303 , n19304 );
not ( n19306 , n19305 );
and ( n19307 , n19302 , n19306 );
not ( n19308 , n19302 );
and ( n19309 , n19308 , n19305 );
nor ( n19310 , n19307 , n19309 );
not ( n19311 , n19310 );
and ( n19312 , n19283 , n19311 );
not ( n19313 , n19283 );
and ( n19314 , n19313 , n19310 );
nor ( n19315 , n19312 , n19314 );
and ( n19316 , n19293 , n19315 );
not ( n19317 , n19316 );
not ( n19318 , n19311 );
not ( n19319 , n19318 );
not ( n19320 , n703 );
and ( n19321 , n691 , n19320 );
not ( n19322 , n691 );
and ( n19323 , n19322 , n703 );
nor ( n19324 , n19321 , n19323 );
not ( n19325 , n19324 );
buf ( n19326 , n19325 );
not ( n19327 , n19326 );
not ( n19328 , n19327 );
not ( n19329 , n988 );
not ( n19330 , n19329 );
and ( n19331 , n703 , n19330 );
not ( n19332 , n703 );
and ( n19333 , n19332 , n19329 );
or ( n19334 , n19331 , n19333 );
nand ( n19335 , n19324 , n19334 );
not ( n19336 , n19335 );
not ( n19337 , n19336 );
not ( n19338 , n19337 );
or ( n19339 , n19328 , n19338 );
buf ( n19340 , n19329 );
nand ( n19341 , n19339 , n19340 );
not ( n19342 , n14180 );
not ( n19343 , n19342 );
not ( n19344 , n10146 );
or ( n19345 , n19343 , n19344 );
nand ( n19346 , n2547 , n14180 );
nand ( n19347 , n19345 , n19346 );
not ( n19348 , n19347 );
not ( n19349 , n19348 );
not ( n19350 , n3592 );
buf ( n19351 , n19350 );
nand ( n19352 , n496 , n512 );
not ( n19353 , n19352 );
nor ( n19354 , n496 , n512 );
nor ( n19355 , n19353 , n19354 );
nor ( n19356 , n503 , n519 );
not ( n19357 , n19356 );
not ( n19358 , n503 );
not ( n19359 , n519 );
or ( n19360 , n19358 , n19359 );
nand ( n19361 , n504 , n520 );
nand ( n19362 , n19360 , n19361 );
nor ( n19363 , n502 , n518 );
not ( n19364 , n19363 );
nand ( n19365 , n19357 , n19362 , n19364 );
nand ( n19366 , n502 , n518 );
nand ( n19367 , n501 , n517 );
nand ( n19368 , n19365 , n19366 , n19367 );
not ( n19369 , n19368 );
nor ( n19370 , n498 , n514 );
nor ( n19371 , n497 , n513 );
nor ( n19372 , n19370 , n19371 );
nor ( n19373 , n501 , n517 );
not ( n19374 , n19373 );
nor ( n19375 , n499 , n515 );
not ( n19376 , n19375 );
not ( n19377 , n500 );
nand ( n19378 , n19377 , n1836 );
and ( n19379 , n19372 , n19374 , n19376 , n19378 );
not ( n19380 , n19379 );
or ( n19381 , n19369 , n19380 );
nand ( n19382 , n500 , n516 );
not ( n19383 , n19382 );
nand ( n19384 , n19376 , n19383 );
not ( n19385 , n19384 );
nand ( n19386 , n498 , n514 );
nand ( n19387 , n497 , n513 );
nand ( n19388 , n499 , n515 );
and ( n19389 , n19386 , n19387 , n19388 );
not ( n19390 , n19389 );
or ( n19391 , n19385 , n19390 );
or ( n19392 , n19371 , n19370 );
nand ( n19393 , n19392 , n19387 );
nand ( n19394 , n19391 , n19393 );
nand ( n19395 , n19381 , n19394 );
buf ( n19396 , n19395 );
xor ( n19397 , n19355 , n19396 );
not ( n19398 , n19397 );
not ( n19399 , n19398 );
xor ( n19400 , n19351 , n19399 );
not ( n19401 , n19400 );
or ( n19402 , n19349 , n19401 );
nand ( n19403 , n19376 , n19378 );
nor ( n19404 , n19403 , n19370 );
not ( n19405 , n19404 );
nor ( n19406 , n501 , n517 );
not ( n19407 , n19406 );
nand ( n19408 , n19357 , n19407 , n19364 );
not ( n19409 , n19362 );
or ( n19410 , n19408 , n19409 );
not ( n19411 , n19373 );
not ( n19412 , n19366 );
and ( n19413 , n19411 , n19412 );
not ( n19414 , n19367 );
nor ( n19415 , n19413 , n19414 );
nand ( n19416 , n19410 , n19415 );
not ( n19417 , n19416 );
or ( n19418 , n19405 , n19417 );
not ( n19419 , n19383 );
not ( n19420 , n19376 );
or ( n19421 , n19419 , n19420 );
nand ( n19422 , n19421 , n19388 );
not ( n19423 , n19370 );
and ( n19424 , n19422 , n19423 );
not ( n19425 , n19386 );
nor ( n19426 , n19424 , n19425 );
nand ( n19427 , n19418 , n19426 );
not ( n19428 , n19387 );
nor ( n19429 , n19428 , n19371 );
and ( n19430 , n19427 , n19429 );
not ( n19431 , n19427 );
not ( n19432 , n19429 );
and ( n19433 , n19431 , n19432 );
nor ( n19434 , n19430 , n19433 );
not ( n19435 , n19434 );
not ( n19436 , n19435 );
xor ( n19437 , n19351 , n19436 );
and ( n19438 , n19350 , n14180 );
not ( n19439 , n19350 );
and ( n19440 , n19439 , n19342 );
nor ( n19441 , n19438 , n19440 );
nand ( n19442 , n19347 , n19441 );
not ( n19443 , n19442 );
nand ( n19444 , n19437 , n19443 );
nand ( n19445 , n19402 , n19444 );
xor ( n19446 , n19341 , n19445 );
not ( n19447 , n19403 );
not ( n19448 , n19447 );
not ( n19449 , n19416 );
or ( n19450 , n19448 , n19449 );
not ( n19451 , n19422 );
nand ( n19452 , n19450 , n19451 );
not ( n19453 , n19386 );
nor ( n19454 , n19453 , n19370 );
and ( n19455 , n19452 , n19454 );
not ( n19456 , n19452 );
not ( n19457 , n19454 );
and ( n19458 , n19456 , n19457 );
nor ( n19459 , n19455 , n19458 );
not ( n19460 , n19459 );
not ( n19461 , n19460 );
and ( n19462 , n19461 , n19351 );
and ( n19463 , n19446 , n19462 );
and ( n19464 , n19341 , n19445 );
or ( n19465 , n19463 , n19464 );
not ( n19466 , n778 );
not ( n19467 , n19330 );
or ( n19468 , n19466 , n19467 );
not ( n19469 , n777 );
nand ( n19470 , n19469 , n19329 );
nand ( n19471 , n19468 , n19470 );
not ( n19472 , n19471 );
not ( n19473 , n778 );
buf ( n19474 , n873 );
not ( n19475 , n19474 );
not ( n19476 , n19475 );
or ( n19477 , n19473 , n19476 );
nand ( n19478 , n19469 , n19474 );
nand ( n19479 , n19477 , n19478 );
and ( n19480 , n19472 , n19479 );
buf ( n19481 , n19480 );
not ( n19482 , n19481 );
buf ( n19483 , n19474 );
not ( n19484 , n19483 );
nor ( n19485 , n491 , n507 );
nor ( n19486 , n492 , n508 );
nor ( n19487 , n19485 , n19486 );
nor ( n19488 , n490 , n506 );
not ( n19489 , n19488 );
and ( n19490 , n19487 , n19489 );
not ( n19491 , n19490 );
not ( n19492 , n493 );
not ( n19493 , n509 );
and ( n19494 , n19492 , n19493 );
nor ( n19495 , n494 , n510 );
nor ( n19496 , n19494 , n19495 );
nor ( n19497 , n495 , n511 );
nor ( n19498 , n19497 , n19354 );
nand ( n19499 , n19496 , n19498 );
nor ( n19500 , n19491 , n19499 );
not ( n19501 , n19500 );
not ( n19502 , n19396 );
or ( n19503 , n19501 , n19502 );
nor ( n19504 , n495 , n511 );
nand ( n19505 , n496 , n512 );
or ( n19506 , n19504 , n19505 );
nand ( n19507 , n495 , n511 );
nand ( n19508 , n19506 , n19507 );
not ( n19509 , n19508 );
nor ( n19510 , n493 , n509 );
nor ( n19511 , n19510 , n19495 );
not ( n19512 , n19511 );
or ( n19513 , n19509 , n19512 );
not ( n19514 , n19510 );
nand ( n19515 , n494 , n510 );
not ( n19516 , n19515 );
and ( n19517 , n19514 , n19516 );
and ( n19518 , n493 , n509 );
nor ( n19519 , n19517 , n19518 );
nand ( n19520 , n19513 , n19519 );
and ( n19521 , n19490 , n19520 );
not ( n19522 , n19489 );
nand ( n19523 , n492 , n508 );
not ( n19524 , n19523 );
not ( n19525 , n19524 );
not ( n19526 , n19485 );
not ( n19527 , n19526 );
or ( n19528 , n19525 , n19527 );
nand ( n19529 , n491 , n507 );
nand ( n19530 , n19528 , n19529 );
not ( n19531 , n19530 );
or ( n19532 , n19522 , n19531 );
nand ( n19533 , n490 , n506 );
nand ( n19534 , n19532 , n19533 );
nor ( n19535 , n19521 , n19534 );
nand ( n19536 , n19503 , n19535 );
nand ( n19537 , n489 , n505 );
not ( n19538 , n19537 );
nor ( n19539 , n489 , n505 );
nor ( n19540 , n19538 , n19539 );
and ( n19541 , n19536 , n19540 );
not ( n19542 , n19536 );
not ( n19543 , n19540 );
and ( n19544 , n19542 , n19543 );
nor ( n19545 , n19541 , n19544 );
not ( n19546 , n19545 );
not ( n19547 , n19546 );
or ( n19548 , n19484 , n19547 );
not ( n19549 , n19483 );
nand ( n19550 , n19549 , n19545 );
nand ( n19551 , n19548 , n19550 );
not ( n19552 , n19551 );
or ( n19553 , n19482 , n19552 );
not ( n19554 , n19486 );
and ( n19555 , n19526 , n19554 );
nor ( n19556 , n19488 , n19539 );
and ( n19557 , n19555 , n19556 );
not ( n19558 , n19557 );
nor ( n19559 , n19558 , n19499 );
not ( n19560 , n19559 );
not ( n19561 , n19396 );
or ( n19562 , n19560 , n19561 );
and ( n19563 , n19557 , n19520 );
not ( n19564 , n19556 );
not ( n19565 , n19530 );
or ( n19566 , n19564 , n19565 );
or ( n19567 , n19533 , n19539 );
nand ( n19568 , n19567 , n19537 );
not ( n19569 , n19568 );
nand ( n19570 , n19566 , n19569 );
nor ( n19571 , n19563 , n19570 );
nand ( n19572 , n19562 , n19571 );
not ( n19573 , n19483 );
and ( n19574 , n19572 , n19573 );
not ( n19575 , n19572 );
and ( n19576 , n19575 , n19483 );
or ( n19577 , n19574 , n19576 );
not ( n19578 , n19472 );
nand ( n19579 , n19577 , n19578 );
nand ( n19580 , n19553 , n19579 );
and ( n19581 , n2948 , n4971 );
not ( n19582 , n2948 );
and ( n19583 , n19582 , n951 );
nor ( n19584 , n19581 , n19583 );
not ( n19585 , n19584 );
not ( n19586 , n19585 );
buf ( n19587 , n1036 );
buf ( n19588 , n19587 );
not ( n19589 , n19588 );
not ( n19590 , n19499 );
not ( n19591 , n19590 );
not ( n19592 , n19396 );
or ( n19593 , n19591 , n19592 );
not ( n19594 , n19520 );
nand ( n19595 , n19593 , n19594 );
nor ( n19596 , n19486 , n19524 );
and ( n19597 , n19595 , n19596 );
not ( n19598 , n19595 );
not ( n19599 , n19596 );
and ( n19600 , n19598 , n19599 );
nor ( n19601 , n19597 , n19600 );
not ( n19602 , n19601 );
not ( n19603 , n19602 );
or ( n19604 , n19589 , n19603 );
buf ( n19605 , n19601 );
not ( n19606 , n19588 );
nand ( n19607 , n19605 , n19606 );
nand ( n19608 , n19604 , n19607 );
not ( n19609 , n19608 );
or ( n19610 , n19586 , n19609 );
not ( n19611 , n19495 );
and ( n19612 , n19498 , n19611 );
not ( n19613 , n19612 );
not ( n19614 , n19395 );
or ( n19615 , n19613 , n19614 );
not ( n19616 , n19611 );
not ( n19617 , n19508 );
or ( n19618 , n19616 , n19617 );
nand ( n19619 , n494 , n510 );
nand ( n19620 , n19618 , n19619 );
not ( n19621 , n19620 );
nand ( n19622 , n19615 , n19621 );
nand ( n19623 , n493 , n509 );
not ( n19624 , n19623 );
nor ( n19625 , n19624 , n19510 );
xor ( n19626 , n19622 , n19625 );
buf ( n19627 , n19626 );
not ( n19628 , n19627 );
and ( n19629 , n19606 , n19628 );
not ( n19630 , n19606 );
and ( n19631 , n19630 , n19627 );
nor ( n19632 , n19629 , n19631 );
not ( n19633 , n19584 );
not ( n19634 , n2948 );
not ( n19635 , n19634 );
not ( n19636 , n19587 );
not ( n19637 , n19636 );
or ( n19638 , n19635 , n19637 );
buf ( n19639 , n2948 );
nand ( n19640 , n19587 , n19639 );
nand ( n19641 , n19638 , n19640 );
nor ( n19642 , n19633 , n19641 );
buf ( n19643 , n19642 );
nand ( n19644 , n19632 , n19643 );
nand ( n19645 , n19610 , n19644 );
xor ( n19646 , n19580 , n19645 );
buf ( n19647 , n2177 );
not ( n19648 , n19647 );
and ( n19649 , n10146 , n19648 );
not ( n19650 , n10146 );
and ( n19651 , n19650 , n19647 );
or ( n19652 , n19649 , n19651 );
xor ( n19653 , n19647 , n19587 );
nor ( n19654 , n19652 , n19653 );
buf ( n19655 , n19654 );
not ( n19656 , n19655 );
not ( n19657 , n10146 );
not ( n19658 , n19657 );
not ( n19659 , n19354 );
not ( n19660 , n19659 );
not ( n19661 , n19395 );
or ( n19662 , n19660 , n19661 );
nand ( n19663 , n19662 , n19352 );
not ( n19664 , n19507 );
nor ( n19665 , n19664 , n19497 );
xor ( n19666 , n19663 , n19665 );
not ( n19667 , n19666 );
not ( n19668 , n19667 );
or ( n19669 , n19658 , n19668 );
nand ( n19670 , n19666 , n10146 );
nand ( n19671 , n19669 , n19670 );
not ( n19672 , n19671 );
or ( n19673 , n19656 , n19672 );
not ( n19674 , n19657 );
not ( n19675 , n19498 );
not ( n19676 , n19395 );
or ( n19677 , n19675 , n19676 );
not ( n19678 , n19508 );
nand ( n19679 , n19677 , n19678 );
not ( n19680 , n19619 );
nor ( n19681 , n19680 , n19495 );
xor ( n19682 , n19679 , n19681 );
not ( n19683 , n19682 );
not ( n19684 , n19683 );
or ( n19685 , n19674 , n19684 );
not ( n19686 , n19683 );
not ( n19687 , n19657 );
nand ( n19688 , n19686 , n19687 );
nand ( n19689 , n19685 , n19688 );
buf ( n19690 , n19653 );
nand ( n19691 , n19689 , n19690 );
nand ( n19692 , n19673 , n19691 );
and ( n19693 , n19646 , n19692 );
and ( n19694 , n19580 , n19645 );
or ( n19695 , n19693 , n19694 );
xor ( n19696 , n19465 , n19695 );
not ( n19697 , n19348 );
xor ( n19698 , n19351 , n19666 );
not ( n19699 , n19698 );
or ( n19700 , n19697 , n19699 );
nand ( n19701 , n19400 , n19443 );
nand ( n19702 , n19700 , n19701 );
not ( n19703 , n19585 );
nor ( n19704 , n19499 , n19486 );
not ( n19705 , n19704 );
not ( n19706 , n19396 );
or ( n19707 , n19705 , n19706 );
not ( n19708 , n19554 );
not ( n19709 , n19520 );
or ( n19710 , n19708 , n19709 );
nand ( n19711 , n19710 , n19523 );
not ( n19712 , n19711 );
nand ( n19713 , n19707 , n19712 );
nand ( n19714 , n19526 , n19529 );
not ( n19715 , n19714 );
and ( n19716 , n19713 , n19715 );
not ( n19717 , n19713 );
and ( n19718 , n19717 , n19714 );
nor ( n19719 , n19716 , n19718 );
not ( n19720 , n19719 );
not ( n19721 , n19720 );
and ( n19722 , n19588 , n19721 );
not ( n19723 , n19588 );
and ( n19724 , n19723 , n19720 );
nor ( n19725 , n19722 , n19724 );
not ( n19726 , n19725 );
or ( n19727 , n19703 , n19726 );
nand ( n19728 , n19608 , n19643 );
nand ( n19729 , n19727 , n19728 );
xor ( n19730 , n19702 , n19729 );
not ( n19731 , n19577 );
not ( n19732 , n19731 );
not ( n19733 , n19481 );
not ( n19734 , n19733 );
and ( n19735 , n19732 , n19734 );
and ( n19736 , n19578 , n19483 );
nor ( n19737 , n19735 , n19736 );
xor ( n19738 , n19730 , n19737 );
xor ( n19739 , n19696 , n19738 );
and ( n19740 , n19351 , n19436 );
xnor ( n19741 , n697 , n19483 );
not ( n19742 , n19741 );
not ( n19743 , n19742 );
not ( n19744 , n11107 );
not ( n19745 , n19744 );
buf ( n19746 , n19545 );
not ( n19747 , n19746 );
not ( n19748 , n19747 );
or ( n19749 , n19745 , n19748 );
nand ( n19750 , n19746 , n11107 );
nand ( n19751 , n19749 , n19750 );
not ( n19752 , n19751 );
or ( n19753 , n19743 , n19752 );
not ( n19754 , n19744 );
nand ( n19755 , n19489 , n19533 );
not ( n19756 , n19755 );
not ( n19757 , n19756 );
not ( n19758 , n19555 );
nor ( n19759 , n19758 , n19499 );
not ( n19760 , n19759 );
not ( n19761 , n19396 );
or ( n19762 , n19760 , n19761 );
and ( n19763 , n19555 , n19520 );
nor ( n19764 , n19763 , n19530 );
nand ( n19765 , n19762 , n19764 );
not ( n19766 , n19765 );
not ( n19767 , n19766 );
or ( n19768 , n19757 , n19767 );
nand ( n19769 , n19765 , n19755 );
nand ( n19770 , n19768 , n19769 );
not ( n19771 , n19770 );
not ( n19772 , n19771 );
or ( n19773 , n19754 , n19772 );
buf ( n19774 , n19770 );
nand ( n19775 , n19774 , n11107 );
nand ( n19776 , n19773 , n19775 );
not ( n19777 , n697 );
not ( n19778 , n11107 );
or ( n19779 , n19777 , n19778 );
not ( n19780 , n697 );
nand ( n19781 , n11108 , n19780 );
nand ( n19782 , n19779 , n19781 );
and ( n19783 , n19741 , n19782 );
buf ( n19784 , n19783 );
nand ( n19785 , n19776 , n19784 );
nand ( n19786 , n19753 , n19785 );
xor ( n19787 , n19740 , n19786 );
not ( n19788 , n19690 );
not ( n19789 , n19657 );
not ( n19790 , n19628 );
or ( n19791 , n19789 , n19790 );
nand ( n19792 , n19627 , n19687 );
nand ( n19793 , n19791 , n19792 );
not ( n19794 , n19793 );
or ( n19795 , n19788 , n19794 );
nand ( n19796 , n19689 , n19655 );
nand ( n19797 , n19795 , n19796 );
xor ( n19798 , n19787 , n19797 );
not ( n19799 , n19784 );
and ( n19800 , n19744 , n19721 );
not ( n19801 , n19744 );
and ( n19802 , n19801 , n19720 );
nor ( n19803 , n19800 , n19802 );
not ( n19804 , n19803 );
or ( n19805 , n19799 , n19804 );
nand ( n19806 , n19776 , n19742 );
nand ( n19807 , n19805 , n19806 );
xor ( n19808 , n19340 , n19572 );
not ( n19809 , n19337 );
and ( n19810 , n19808 , n19809 );
and ( n19811 , n19326 , n19340 );
nor ( n19812 , n19810 , n19811 );
not ( n19813 , n19812 );
xor ( n19814 , n19807 , n19813 );
not ( n19815 , n19351 );
not ( n19816 , n19460 );
or ( n19817 , n19815 , n19816 );
not ( n19818 , n19351 );
nand ( n19819 , n19461 , n19818 );
nand ( n19820 , n19817 , n19819 );
not ( n19821 , n19820 );
not ( n19822 , n19443 );
or ( n19823 , n19821 , n19822 );
not ( n19824 , n19348 );
not ( n19825 , n19824 );
nand ( n19826 , n19825 , n19437 );
nand ( n19827 , n19823 , n19826 );
nand ( n19828 , n19365 , n19366 );
not ( n19829 , n19828 );
not ( n19830 , n19378 );
nor ( n19831 , n19406 , n19830 );
not ( n19832 , n19831 );
or ( n19833 , n19829 , n19832 );
or ( n19834 , n19830 , n19367 );
nand ( n19835 , n19834 , n19382 );
not ( n19836 , n19835 );
nand ( n19837 , n19833 , n19836 );
nand ( n19838 , n19376 , n19388 );
not ( n19839 , n19838 );
and ( n19840 , n19837 , n19839 );
not ( n19841 , n19837 );
and ( n19842 , n19841 , n19838 );
nor ( n19843 , n19840 , n19842 );
buf ( n19844 , n19843 );
and ( n19845 , n19351 , n19844 );
xor ( n19846 , n19827 , n19845 );
not ( n19847 , n19481 );
not ( n19848 , n19483 );
not ( n19849 , n19771 );
or ( n19850 , n19848 , n19849 );
nand ( n19851 , n19774 , n19573 );
nand ( n19852 , n19850 , n19851 );
not ( n19853 , n19852 );
or ( n19854 , n19847 , n19853 );
nand ( n19855 , n19551 , n19578 );
nand ( n19856 , n19854 , n19855 );
and ( n19857 , n19846 , n19856 );
and ( n19858 , n19827 , n19845 );
or ( n19859 , n19857 , n19858 );
and ( n19860 , n19814 , n19859 );
and ( n19861 , n19807 , n19813 );
or ( n19862 , n19860 , n19861 );
xor ( n19863 , n19798 , n19862 );
not ( n19864 , n19643 );
and ( n19865 , n19682 , n19588 );
not ( n19866 , n19682 );
and ( n19867 , n19866 , n19606 );
nor ( n19868 , n19865 , n19867 );
not ( n19869 , n19868 );
or ( n19870 , n19864 , n19869 );
nand ( n19871 , n19632 , n19585 );
nand ( n19872 , n19870 , n19871 );
not ( n19873 , n691 );
nor ( n19874 , n19873 , n685 );
buf ( n19875 , n19874 );
buf ( n19876 , n685 );
or ( n19877 , n19875 , n19876 );
buf ( n19878 , n691 );
nand ( n19879 , n19877 , n19878 );
not ( n19880 , n19879 );
nor ( n19881 , n19383 , n19830 );
not ( n19882 , n19881 );
not ( n19883 , n19416 );
not ( n19884 , n19883 );
or ( n19885 , n19882 , n19884 );
not ( n19886 , n19881 );
nand ( n19887 , n19886 , n19416 );
nand ( n19888 , n19885 , n19887 );
not ( n19889 , n19888 );
not ( n19890 , n19889 );
nand ( n19891 , n19890 , n19351 );
nand ( n19892 , n19880 , n19891 );
xor ( n19893 , n19872 , n19892 );
not ( n19894 , n19657 );
not ( n19895 , n19398 );
or ( n19896 , n19894 , n19895 );
nand ( n19897 , n19399 , n10146 );
nand ( n19898 , n19896 , n19897 );
not ( n19899 , n19898 );
not ( n19900 , n19655 );
or ( n19901 , n19899 , n19900 );
not ( n19902 , n19671 );
not ( n19903 , n19690 );
or ( n19904 , n19902 , n19903 );
nand ( n19905 , n19901 , n19904 );
and ( n19906 , n19893 , n19905 );
and ( n19907 , n19872 , n19892 );
or ( n19908 , n19906 , n19907 );
xor ( n19909 , n19341 , n19445 );
xor ( n19910 , n19909 , n19462 );
xor ( n19911 , n19908 , n19910 );
xor ( n19912 , n19580 , n19645 );
xor ( n19913 , n19912 , n19692 );
and ( n19914 , n19911 , n19913 );
and ( n19915 , n19908 , n19910 );
or ( n19916 , n19914 , n19915 );
xor ( n19917 , n19863 , n19916 );
xor ( n19918 , n19739 , n19917 );
xor ( n19919 , n19807 , n19813 );
xor ( n19920 , n19919 , n19859 );
not ( n19921 , n19742 );
not ( n19922 , n19803 );
or ( n19923 , n19921 , n19922 );
not ( n19924 , n19744 );
not ( n19925 , n19602 );
or ( n19926 , n19924 , n19925 );
nand ( n19927 , n19605 , n11107 );
nand ( n19928 , n19926 , n19927 );
nand ( n19929 , n19928 , n19784 );
nand ( n19930 , n19923 , n19929 );
xor ( n19931 , n19930 , n19812 );
not ( n19932 , n19809 );
xor ( n19933 , n19340 , n19545 );
not ( n19934 , n19933 );
or ( n19935 , n19932 , n19934 );
nand ( n19936 , n19808 , n19326 );
nand ( n19937 , n19935 , n19936 );
not ( n19938 , n19643 );
not ( n19939 , n19588 );
not ( n19940 , n19667 );
or ( n19941 , n19939 , n19940 );
nand ( n19942 , n19666 , n19606 );
nand ( n19943 , n19941 , n19942 );
not ( n19944 , n19943 );
or ( n19945 , n19938 , n19944 );
nand ( n19946 , n19868 , n19585 );
nand ( n19947 , n19945 , n19946 );
xor ( n19948 , n19937 , n19947 );
not ( n19949 , n19578 );
not ( n19950 , n19852 );
or ( n19951 , n19949 , n19950 );
not ( n19952 , n19483 );
not ( n19953 , n19720 );
or ( n19954 , n19952 , n19953 );
nand ( n19955 , n19719 , n19573 );
nand ( n19956 , n19954 , n19955 );
nand ( n19957 , n19956 , n19481 );
nand ( n19958 , n19951 , n19957 );
and ( n19959 , n19948 , n19958 );
and ( n19960 , n19937 , n19947 );
or ( n19961 , n19959 , n19960 );
and ( n19962 , n19931 , n19961 );
and ( n19963 , n19930 , n19812 );
or ( n19964 , n19962 , n19963 );
xor ( n19965 , n19920 , n19964 );
xor ( n19966 , n19908 , n19910 );
xor ( n19967 , n19966 , n19913 );
and ( n19968 , n19965 , n19967 );
and ( n19969 , n19920 , n19964 );
or ( n19970 , n19968 , n19969 );
and ( n19971 , n19918 , n19970 );
and ( n19972 , n19739 , n19917 );
or ( n19973 , n19971 , n19972 );
xor ( n19974 , n19465 , n19695 );
and ( n19975 , n19974 , n19738 );
and ( n19976 , n19465 , n19695 );
or ( n19977 , n19975 , n19976 );
xor ( n19978 , n19702 , n19729 );
and ( n19979 , n19978 , n19737 );
and ( n19980 , n19702 , n19729 );
or ( n19981 , n19979 , n19980 );
not ( n19982 , n19655 );
not ( n19983 , n19793 );
or ( n19984 , n19982 , n19983 );
not ( n19985 , n19657 );
not ( n19986 , n19602 );
or ( n19987 , n19985 , n19986 );
not ( n19988 , n19602 );
nand ( n19989 , n19988 , n19687 );
nand ( n19990 , n19987 , n19989 );
nand ( n19991 , n19990 , n19690 );
nand ( n19992 , n19984 , n19991 );
not ( n19993 , n19443 );
not ( n19994 , n19698 );
or ( n19995 , n19993 , n19994 );
xor ( n19996 , n19351 , n19686 );
nand ( n19997 , n19996 , n19348 );
nand ( n19998 , n19995 , n19997 );
xor ( n19999 , n19992 , n19998 );
not ( n20000 , n19643 );
not ( n20001 , n19725 );
or ( n20002 , n20000 , n20001 );
xnor ( n20003 , n19606 , n19774 );
nand ( n20004 , n20003 , n19585 );
nand ( n20005 , n20002 , n20004 );
xor ( n20006 , n19999 , n20005 );
xor ( n20007 , n19981 , n20006 );
not ( n20008 , n19737 );
xor ( n20009 , n19740 , n19786 );
and ( n20010 , n20009 , n19797 );
and ( n20011 , n19740 , n19786 );
or ( n20012 , n20010 , n20011 );
xor ( n20013 , n20008 , n20012 );
not ( n20014 , n19472 );
not ( n20015 , n19733 );
or ( n20016 , n20014 , n20015 );
nand ( n20017 , n20016 , n19483 );
and ( n20018 , n19351 , n19399 );
xor ( n20019 , n20017 , n20018 );
not ( n20020 , n19784 );
not ( n20021 , n19751 );
or ( n20022 , n20020 , n20021 );
not ( n20023 , n19572 );
and ( n20024 , n11107 , n20023 );
not ( n20025 , n11107 );
and ( n20026 , n20025 , n19572 );
nor ( n20027 , n20024 , n20026 );
nand ( n20028 , n20027 , n19742 );
nand ( n20029 , n20022 , n20028 );
xor ( n20030 , n20019 , n20029 );
xor ( n20031 , n20013 , n20030 );
xor ( n20032 , n20007 , n20031 );
xor ( n20033 , n19977 , n20032 );
xor ( n20034 , n19798 , n19862 );
and ( n20035 , n20034 , n19916 );
and ( n20036 , n19798 , n19862 );
or ( n20037 , n20035 , n20036 );
xor ( n20038 , n20033 , n20037 );
nand ( n20039 , n19973 , n20038 );
not ( n20040 , n20039 );
nor ( n20041 , n20038 , n19973 );
nor ( n20042 , n20040 , n20041 );
xor ( n20043 , n19739 , n19917 );
xor ( n20044 , n20043 , n19970 );
not ( n20045 , n20044 );
not ( n20046 , n19655 );
not ( n20047 , n19657 );
not ( n20048 , n19435 );
or ( n20049 , n20047 , n20048 );
nand ( n20050 , n19436 , n10146 );
nand ( n20051 , n20049 , n20050 );
not ( n20052 , n20051 );
or ( n20053 , n20046 , n20052 );
nand ( n20054 , n19898 , n19690 );
nand ( n20055 , n20053 , n20054 );
not ( n20056 , n19443 );
xor ( n20057 , n19351 , n19844 );
not ( n20058 , n20057 );
or ( n20059 , n20056 , n20058 );
nand ( n20060 , n19820 , n19348 );
nand ( n20061 , n20059 , n20060 );
xor ( n20062 , n20055 , n20061 );
not ( n20063 , n19742 );
not ( n20064 , n19928 );
or ( n20065 , n20063 , n20064 );
and ( n20066 , n11108 , n19627 );
not ( n20067 , n11108 );
and ( n20068 , n20067 , n19628 );
nor ( n20069 , n20066 , n20068 );
nand ( n20070 , n20069 , n19784 );
nand ( n20071 , n20065 , n20070 );
and ( n20072 , n20062 , n20071 );
and ( n20073 , n20055 , n20061 );
or ( n20074 , n20072 , n20073 );
xor ( n20075 , n19827 , n19845 );
xor ( n20076 , n20075 , n19856 );
xor ( n20077 , n20074 , n20076 );
xor ( n20078 , n19872 , n19892 );
xor ( n20079 , n20078 , n19905 );
and ( n20080 , n20077 , n20079 );
and ( n20081 , n20074 , n20076 );
or ( n20082 , n20080 , n20081 );
xor ( n20083 , n19920 , n19964 );
xor ( n20084 , n20083 , n19967 );
xor ( n20085 , n20082 , n20084 );
not ( n20086 , n19879 );
not ( n20087 , n19891 );
not ( n20088 , n20087 );
or ( n20089 , n20086 , n20088 );
nand ( n20090 , n20089 , n19892 );
and ( n20091 , n19407 , n19367 );
xor ( n20092 , n20091 , n19828 );
and ( n20093 , n19351 , n20092 );
not ( n20094 , n19875 );
not ( n20095 , n19878 );
and ( n20096 , n19572 , n20095 );
not ( n20097 , n19572 );
and ( n20098 , n20097 , n19878 );
or ( n20099 , n20096 , n20098 );
not ( n20100 , n20099 );
or ( n20101 , n20094 , n20100 );
nand ( n20102 , n19878 , n19876 );
nand ( n20103 , n20101 , n20102 );
and ( n20104 , n20093 , n20103 );
xor ( n20105 , n20090 , n20104 );
not ( n20106 , n19348 );
not ( n20107 , n19351 );
buf ( n20108 , n19888 );
not ( n20109 , n20108 );
not ( n20110 , n20109 );
or ( n20111 , n20107 , n20110 );
nand ( n20112 , n20108 , n19818 );
nand ( n20113 , n20111 , n20112 );
not ( n20114 , n20113 );
or ( n20115 , n20106 , n20114 );
xor ( n20116 , n19351 , n20092 );
nand ( n20117 , n20116 , n19443 );
nand ( n20118 , n20115 , n20117 );
not ( n20119 , n20118 );
not ( n20120 , n19361 );
not ( n20121 , n20120 );
not ( n20122 , n19357 );
or ( n20123 , n20121 , n20122 );
nand ( n20124 , n503 , n519 );
nand ( n20125 , n20123 , n20124 );
and ( n20126 , n19364 , n19366 );
xor ( n20127 , n20125 , n20126 );
nand ( n20128 , n20127 , n19351 );
nor ( n20129 , n20119 , n20128 );
not ( n20130 , n19690 );
not ( n20131 , n20051 );
or ( n20132 , n20130 , n20131 );
not ( n20133 , n19657 );
not ( n20134 , n19460 );
or ( n20135 , n20133 , n20134 );
nand ( n20136 , n19461 , n19687 );
nand ( n20137 , n20135 , n20136 );
nand ( n20138 , n20137 , n19655 );
nand ( n20139 , n20132 , n20138 );
xor ( n20140 , n20129 , n20139 );
not ( n20141 , n19348 );
not ( n20142 , n20057 );
or ( n20143 , n20141 , n20142 );
nand ( n20144 , n20113 , n19443 );
nand ( n20145 , n20143 , n20144 );
and ( n20146 , n20140 , n20145 );
and ( n20147 , n20129 , n20139 );
or ( n20148 , n20146 , n20147 );
and ( n20149 , n20105 , n20148 );
and ( n20150 , n20090 , n20104 );
or ( n20151 , n20149 , n20150 );
xor ( n20152 , n19930 , n19812 );
xor ( n20153 , n20152 , n19961 );
xor ( n20154 , n20151 , n20153 );
not ( n20155 , n19784 );
not ( n20156 , n19744 );
not ( n20157 , n19683 );
or ( n20158 , n20156 , n20157 );
nand ( n20159 , n19682 , n11107 );
nand ( n20160 , n20158 , n20159 );
not ( n20161 , n20160 );
or ( n20162 , n20155 , n20161 );
nand ( n20163 , n20069 , n19742 );
nand ( n20164 , n20162 , n20163 );
not ( n20165 , n19326 );
not ( n20166 , n19933 );
or ( n20167 , n20165 , n20166 );
not ( n20168 , n19755 );
not ( n20169 , n19340 );
not ( n20170 , n20169 );
or ( n20171 , n20168 , n20170 );
or ( n20172 , n20169 , n19755 );
nand ( n20173 , n20171 , n20172 );
and ( n20174 , n20173 , n19766 );
not ( n20175 , n20173 );
and ( n20176 , n20175 , n19765 );
nor ( n20177 , n20174 , n20176 );
nand ( n20178 , n20177 , n19809 );
nand ( n20179 , n20167 , n20178 );
xor ( n20180 , n20164 , n20179 );
not ( n20181 , n19643 );
not ( n20182 , n19588 );
not ( n20183 , n19398 );
or ( n20184 , n20182 , n20183 );
nand ( n20185 , n19399 , n19606 );
nand ( n20186 , n20184 , n20185 );
not ( n20187 , n20186 );
or ( n20188 , n20181 , n20187 );
not ( n20189 , n19943 );
or ( n20190 , n20189 , n19584 );
nand ( n20191 , n20188 , n20190 );
and ( n20192 , n20180 , n20191 );
and ( n20193 , n20164 , n20179 );
or ( n20194 , n20192 , n20193 );
xor ( n20195 , n20055 , n20061 );
xor ( n20196 , n20195 , n20071 );
xor ( n20197 , n20194 , n20196 );
xor ( n20198 , n19937 , n19947 );
xor ( n20199 , n20198 , n19958 );
and ( n20200 , n20197 , n20199 );
and ( n20201 , n20194 , n20196 );
or ( n20202 , n20200 , n20201 );
and ( n20203 , n20154 , n20202 );
and ( n20204 , n20151 , n20153 );
or ( n20205 , n20203 , n20204 );
and ( n20206 , n20085 , n20205 );
and ( n20207 , n20082 , n20084 );
or ( n20208 , n20206 , n20207 );
not ( n20209 , n20208 );
and ( n20210 , n20045 , n20209 );
xor ( n20211 , n20082 , n20084 );
xor ( n20212 , n20211 , n20205 );
xor ( n20213 , n20074 , n20076 );
xor ( n20214 , n20213 , n20079 );
xor ( n20215 , n20151 , n20153 );
xor ( n20216 , n20215 , n20202 );
xor ( n20217 , n20214 , n20216 );
not ( n20218 , n19481 );
and ( n20219 , n19602 , n19483 );
not ( n20220 , n19602 );
and ( n20221 , n20220 , n19573 );
or ( n20222 , n20219 , n20221 );
not ( n20223 , n20222 );
or ( n20224 , n20218 , n20223 );
nand ( n20225 , n19956 , n19578 );
nand ( n20226 , n20224 , n20225 );
xor ( n20227 , n20093 , n20103 );
xor ( n20228 , n20226 , n20227 );
not ( n20229 , n20128 );
and ( n20230 , n20118 , n20229 );
not ( n20231 , n20118 );
and ( n20232 , n20231 , n20128 );
nor ( n20233 , n20230 , n20232 );
not ( n20234 , n19585 );
not ( n20235 , n20186 );
or ( n20236 , n20234 , n20235 );
not ( n20237 , n19588 );
not ( n20238 , n19435 );
or ( n20239 , n20237 , n20238 );
nand ( n20240 , n19436 , n19606 );
nand ( n20241 , n20239 , n20240 );
nand ( n20242 , n20241 , n19643 );
nand ( n20243 , n20236 , n20242 );
and ( n20244 , n20233 , n20243 );
and ( n20245 , n20228 , n20244 );
and ( n20246 , n20226 , n20227 );
or ( n20247 , n20245 , n20246 );
xor ( n20248 , n20090 , n20104 );
xor ( n20249 , n20248 , n20148 );
xor ( n20250 , n20247 , n20249 );
not ( n20251 , n19655 );
and ( n20252 , n19657 , n19844 );
not ( n20253 , n19657 );
not ( n20254 , n19844 );
and ( n20255 , n20253 , n20254 );
nor ( n20256 , n20252 , n20255 );
not ( n20257 , n20256 );
or ( n20258 , n20251 , n20257 );
nand ( n20259 , n20137 , n19690 );
nand ( n20260 , n20258 , n20259 );
not ( n20261 , n19784 );
and ( n20262 , n19744 , n19666 );
not ( n20263 , n19744 );
and ( n20264 , n20263 , n19667 );
nor ( n20265 , n20262 , n20264 );
not ( n20266 , n20265 );
or ( n20267 , n20261 , n20266 );
nand ( n20268 , n20160 , n19742 );
nand ( n20269 , n20267 , n20268 );
xor ( n20270 , n20260 , n20269 );
and ( n20271 , n20095 , n19546 );
not ( n20272 , n20095 );
and ( n20273 , n20272 , n19545 );
or ( n20274 , n20271 , n20273 );
not ( n20275 , n19875 );
or ( n20276 , n20274 , n20275 );
not ( n20277 , n20099 );
not ( n20278 , n19876 );
or ( n20279 , n20277 , n20278 );
nand ( n20280 , n20276 , n20279 );
and ( n20281 , n20270 , n20280 );
and ( n20282 , n20260 , n20269 );
or ( n20283 , n20281 , n20282 );
xor ( n20284 , n20129 , n20139 );
xor ( n20285 , n20284 , n20145 );
xor ( n20286 , n20283 , n20285 );
xor ( n20287 , n20164 , n20179 );
xor ( n20288 , n20287 , n20191 );
and ( n20289 , n20286 , n20288 );
and ( n20290 , n20283 , n20285 );
or ( n20291 , n20289 , n20290 );
and ( n20292 , n20250 , n20291 );
and ( n20293 , n20247 , n20249 );
or ( n20294 , n20292 , n20293 );
and ( n20295 , n20217 , n20294 );
and ( n20296 , n20214 , n20216 );
or ( n20297 , n20295 , n20296 );
nor ( n20298 , n20212 , n20297 );
nor ( n20299 , n20210 , n20298 );
not ( n20300 , n20299 );
xor ( n20301 , n20214 , n20216 );
xor ( n20302 , n20301 , n20294 );
xor ( n20303 , n20194 , n20196 );
xor ( n20304 , n20303 , n20199 );
xor ( n20305 , n20226 , n20227 );
xor ( n20306 , n20305 , n20244 );
not ( n20307 , n19809 );
not ( n20308 , n19340 );
not ( n20309 , n19720 );
or ( n20310 , n20308 , n20309 );
nand ( n20311 , n19719 , n20169 );
nand ( n20312 , n20310 , n20311 );
not ( n20313 , n20312 );
or ( n20314 , n20307 , n20313 );
nand ( n20315 , n20177 , n19326 );
nand ( n20316 , n20314 , n20315 );
not ( n20317 , n19481 );
not ( n20318 , n19483 );
not ( n20319 , n19628 );
or ( n20320 , n20318 , n20319 );
nand ( n20321 , n19627 , n19573 );
nand ( n20322 , n20320 , n20321 );
not ( n20323 , n20322 );
or ( n20324 , n20317 , n20323 );
nand ( n20325 , n20222 , n19578 );
nand ( n20326 , n20324 , n20325 );
xor ( n20327 , n20316 , n20326 );
not ( n20328 , n19351 );
buf ( n20329 , n20127 );
not ( n20330 , n20329 );
not ( n20331 , n20330 );
or ( n20332 , n20328 , n20331 );
not ( n20333 , n19350 );
nand ( n20334 , n20333 , n20329 );
nand ( n20335 , n20332 , n20334 );
nand ( n20336 , n20335 , n19443 );
nand ( n20337 , n20116 , n19348 );
nand ( n20338 , n20336 , n20337 );
and ( n20339 , n19357 , n20124 );
and ( n20340 , n20339 , n20120 );
not ( n20341 , n20339 );
not ( n20342 , n20120 );
and ( n20343 , n20341 , n20342 );
nor ( n20344 , n20340 , n20343 );
buf ( n20345 , n20344 );
and ( n20346 , n19350 , n20345 );
xor ( n20347 , n20338 , n20346 );
not ( n20348 , n19690 );
not ( n20349 , n20256 );
or ( n20350 , n20348 , n20349 );
not ( n20351 , n19657 );
not ( n20352 , n20109 );
or ( n20353 , n20351 , n20352 );
not ( n20354 , n19657 );
nand ( n20355 , n20354 , n20108 );
nand ( n20356 , n20353 , n20355 );
nand ( n20357 , n20356 , n19655 );
nand ( n20358 , n20350 , n20357 );
and ( n20359 , n20347 , n20358 );
and ( n20360 , n20338 , n20346 );
or ( n20361 , n20359 , n20360 );
and ( n20362 , n20327 , n20361 );
and ( n20363 , n20316 , n20326 );
or ( n20364 , n20362 , n20363 );
xor ( n20365 , n20306 , n20364 );
xor ( n20366 , n20233 , n20243 );
not ( n20367 , n19585 );
not ( n20368 , n20241 );
or ( n20369 , n20367 , n20368 );
not ( n20370 , n19588 );
not ( n20371 , n19460 );
or ( n20372 , n20370 , n20371 );
nand ( n20373 , n19459 , n19606 );
nand ( n20374 , n20372 , n20373 );
nand ( n20375 , n20374 , n19643 );
nand ( n20376 , n20369 , n20375 );
not ( n20377 , n19744 );
not ( n20378 , n19398 );
or ( n20379 , n20377 , n20378 );
nand ( n20380 , n19399 , n11107 );
nand ( n20381 , n20379 , n20380 );
not ( n20382 , n20381 );
not ( n20383 , n19784 );
or ( n20384 , n20382 , n20383 );
not ( n20385 , n20265 );
not ( n20386 , n19742 );
or ( n20387 , n20385 , n20386 );
nand ( n20388 , n20384 , n20387 );
xor ( n20389 , n20376 , n20388 );
and ( n20390 , n20095 , n19771 );
not ( n20391 , n20095 );
and ( n20392 , n20391 , n19774 );
or ( n20393 , n20390 , n20392 );
or ( n20394 , n20393 , n20275 );
or ( n20395 , n20274 , n20278 );
nand ( n20396 , n20394 , n20395 );
and ( n20397 , n20389 , n20396 );
and ( n20398 , n20376 , n20388 );
or ( n20399 , n20397 , n20398 );
xor ( n20400 , n20366 , n20399 );
not ( n20401 , n19809 );
and ( n20402 , n19601 , n20169 );
not ( n20403 , n19601 );
and ( n20404 , n20403 , n19340 );
or ( n20405 , n20402 , n20404 );
not ( n20406 , n20405 );
or ( n20407 , n20401 , n20406 );
nand ( n20408 , n20312 , n19326 );
nand ( n20409 , n20407 , n20408 );
xor ( n20410 , n504 , n520 );
buf ( n20411 , n20410 );
and ( n20412 , n20411 , n19351 );
not ( n20413 , n19443 );
xor ( n20414 , n19350 , n20345 );
not ( n20415 , n20414 );
or ( n20416 , n20413 , n20415 );
nand ( n20417 , n20335 , n19348 );
nand ( n20418 , n20416 , n20417 );
xor ( n20419 , n20412 , n20418 );
not ( n20420 , n19442 );
not ( n20421 , n20411 );
and ( n20422 , n19350 , n20421 );
not ( n20423 , n19350 );
not ( n20424 , n20410 );
not ( n20425 , n20424 );
and ( n20426 , n20423 , n20425 );
nor ( n20427 , n20422 , n20426 );
not ( n20428 , n20427 );
and ( n20429 , n20420 , n20428 );
and ( n20430 , n20414 , n19348 );
nor ( n20431 , n20429 , n20430 );
not ( n20432 , n19342 );
not ( n20433 , n10146 );
or ( n20434 , n20432 , n20433 );
nand ( n20435 , n20434 , n20411 );
nand ( n20436 , n19351 , n19346 , n20435 );
nor ( n20437 , n20431 , n20436 );
and ( n20438 , n20419 , n20437 );
and ( n20439 , n20412 , n20418 );
or ( n20440 , n20438 , n20439 );
xor ( n20441 , n20409 , n20440 );
not ( n20442 , n19481 );
not ( n20443 , n19483 );
not ( n20444 , n19683 );
or ( n20445 , n20443 , n20444 );
nand ( n20446 , n19686 , n19573 );
nand ( n20447 , n20445 , n20446 );
not ( n20448 , n20447 );
or ( n20449 , n20442 , n20448 );
nand ( n20450 , n20322 , n19578 );
nand ( n20451 , n20449 , n20450 );
and ( n20452 , n20441 , n20451 );
and ( n20453 , n20409 , n20440 );
or ( n20454 , n20452 , n20453 );
and ( n20455 , n20400 , n20454 );
and ( n20456 , n20366 , n20399 );
or ( n20457 , n20455 , n20456 );
and ( n20458 , n20365 , n20457 );
and ( n20459 , n20306 , n20364 );
or ( n20460 , n20458 , n20459 );
xor ( n20461 , n20304 , n20460 );
xor ( n20462 , n20247 , n20249 );
xor ( n20463 , n20462 , n20291 );
and ( n20464 , n20461 , n20463 );
and ( n20465 , n20304 , n20460 );
or ( n20466 , n20464 , n20465 );
nor ( n20467 , n20302 , n20466 );
xor ( n20468 , n20283 , n20285 );
xor ( n20469 , n20468 , n20288 );
xor ( n20470 , n20306 , n20364 );
xor ( n20471 , n20470 , n20457 );
xor ( n20472 , n20469 , n20471 );
xor ( n20473 , n20260 , n20269 );
xor ( n20474 , n20473 , n20280 );
xor ( n20475 , n20316 , n20326 );
xor ( n20476 , n20475 , n20361 );
xor ( n20477 , n20474 , n20476 );
not ( n20478 , n19690 );
not ( n20479 , n20356 );
or ( n20480 , n20478 , n20479 );
not ( n20481 , n19657 );
not ( n20482 , n20092 );
not ( n20483 , n20482 );
or ( n20484 , n20481 , n20483 );
nand ( n20485 , n20092 , n19687 );
nand ( n20486 , n20484 , n20485 );
nand ( n20487 , n20486 , n19655 );
nand ( n20488 , n20480 , n20487 );
not ( n20489 , n19643 );
and ( n20490 , n19588 , n19844 );
not ( n20491 , n19588 );
and ( n20492 , n20491 , n20254 );
nor ( n20493 , n20490 , n20492 );
not ( n20494 , n20493 );
or ( n20495 , n20489 , n20494 );
nand ( n20496 , n20374 , n19585 );
nand ( n20497 , n20495 , n20496 );
xor ( n20498 , n20488 , n20497 );
not ( n20499 , n19784 );
not ( n20500 , n11108 );
not ( n20501 , n19435 );
or ( n20502 , n20500 , n20501 );
nand ( n20503 , n19436 , n11107 );
nand ( n20504 , n20502 , n20503 );
not ( n20505 , n20504 );
or ( n20506 , n20499 , n20505 );
nand ( n20507 , n20381 , n19742 );
nand ( n20508 , n20506 , n20507 );
and ( n20509 , n20498 , n20508 );
and ( n20510 , n20488 , n20497 );
or ( n20511 , n20509 , n20510 );
xor ( n20512 , n20338 , n20346 );
xor ( n20513 , n20512 , n20358 );
xor ( n20514 , n20511 , n20513 );
xor ( n20515 , n20412 , n20418 );
xor ( n20516 , n20515 , n20437 );
not ( n20517 , n19809 );
not ( n20518 , n19340 );
not ( n20519 , n19628 );
or ( n20520 , n20518 , n20519 );
nand ( n20521 , n19627 , n20169 );
nand ( n20522 , n20520 , n20521 );
not ( n20523 , n20522 );
or ( n20524 , n20517 , n20523 );
nand ( n20525 , n20405 , n19326 );
nand ( n20526 , n20524 , n20525 );
xor ( n20527 , n20516 , n20526 );
not ( n20528 , n19878 );
not ( n20529 , n19720 );
or ( n20530 , n20528 , n20529 );
nand ( n20531 , n19719 , n20095 );
nand ( n20532 , n20530 , n20531 );
not ( n20533 , n20532 );
not ( n20534 , n19875 );
or ( n20535 , n20533 , n20534 );
or ( n20536 , n20393 , n20278 );
nand ( n20537 , n20535 , n20536 );
and ( n20538 , n20527 , n20537 );
and ( n20539 , n20516 , n20526 );
or ( n20540 , n20538 , n20539 );
and ( n20541 , n20514 , n20540 );
and ( n20542 , n20511 , n20513 );
or ( n20543 , n20541 , n20542 );
and ( n20544 , n20477 , n20543 );
and ( n20545 , n20474 , n20476 );
or ( n20546 , n20544 , n20545 );
and ( n20547 , n20472 , n20546 );
and ( n20548 , n20469 , n20471 );
or ( n20549 , n20547 , n20548 );
xor ( n20550 , n20304 , n20460 );
xor ( n20551 , n20550 , n20463 );
nand ( n20552 , n20549 , n20551 );
or ( n20553 , n20467 , n20552 );
nand ( n20554 , n20302 , n20466 );
nand ( n20555 , n20553 , n20554 );
not ( n20556 , n20555 );
or ( n20557 , n20300 , n20556 );
not ( n20558 , n20044 );
not ( n20559 , n20208 );
nand ( n20560 , n20558 , n20559 );
and ( n20561 , n20212 , n20297 );
and ( n20562 , n20560 , n20561 );
nor ( n20563 , n20558 , n20559 );
nor ( n20564 , n20562 , n20563 );
nand ( n20565 , n20557 , n20564 );
not ( n20566 , n20565 );
not ( n20567 , n19741 );
not ( n20568 , n20567 );
not ( n20569 , n11108 );
not ( n20570 , n20345 );
not ( n20571 , n20570 );
or ( n20572 , n20569 , n20571 );
nand ( n20573 , n20345 , n11107 );
nand ( n20574 , n20572 , n20573 );
not ( n20575 , n20574 );
or ( n20576 , n20568 , n20575 );
nor ( n20577 , n20411 , n697 , n19483 , n11107 );
and ( n20578 , n19483 , n11107 , n20411 , n697 );
nor ( n20579 , n20577 , n20578 );
nand ( n20580 , n20576 , n20579 );
not ( n20581 , n19483 );
nand ( n20582 , n20581 , n19780 );
and ( n20583 , n20582 , n20425 );
not ( n20584 , n697 );
not ( n20585 , n19483 );
or ( n20586 , n20584 , n20585 );
nand ( n20587 , n20586 , n11108 );
nor ( n20588 , n20583 , n20587 );
and ( n20589 , n20580 , n20588 );
not ( n20590 , n19809 );
not ( n20591 , n19330 );
and ( n20592 , n20591 , n20254 );
not ( n20593 , n20591 );
and ( n20594 , n20593 , n19844 );
or ( n20595 , n20592 , n20594 );
not ( n20596 , n20595 );
or ( n20597 , n20590 , n20596 );
xor ( n20598 , n19340 , n19459 );
nand ( n20599 , n20598 , n19326 );
nand ( n20600 , n20597 , n20599 );
xor ( n20601 , n20589 , n20600 );
not ( n20602 , n19876 );
xor ( n20603 , n19878 , n19397 );
not ( n20604 , n20603 );
or ( n20605 , n20602 , n20604 );
and ( n20606 , n20095 , n19435 );
not ( n20607 , n20095 );
and ( n20608 , n20607 , n19434 );
nor ( n20609 , n20606 , n20608 );
nand ( n20610 , n20609 , n19875 );
nand ( n20611 , n20605 , n20610 );
and ( n20612 , n20601 , n20611 );
and ( n20613 , n20589 , n20600 );
or ( n20614 , n20612 , n20613 );
not ( n20615 , n19742 );
not ( n20616 , n19744 );
not ( n20617 , n20482 );
or ( n20618 , n20616 , n20617 );
nand ( n20619 , n20092 , n11107 );
nand ( n20620 , n20618 , n20619 );
not ( n20621 , n20620 );
or ( n20622 , n20615 , n20621 );
not ( n20623 , n19744 );
not ( n20624 , n20127 );
not ( n20625 , n20624 );
or ( n20626 , n20623 , n20625 );
nand ( n20627 , n20329 , n11107 );
nand ( n20628 , n20626 , n20627 );
nand ( n20629 , n20628 , n19783 );
nand ( n20630 , n20622 , n20629 );
not ( n20631 , n11108 );
nand ( n20632 , n20631 , n19634 );
and ( n20633 , n20632 , n20411 );
not ( n20634 , n19639 );
not ( n20635 , n19744 );
or ( n20636 , n20634 , n20635 );
nand ( n20637 , n20636 , n19588 );
nor ( n20638 , n20633 , n20637 );
not ( n20639 , n19585 );
not ( n20640 , n19588 );
not ( n20641 , n20570 );
or ( n20642 , n20640 , n20641 );
nand ( n20643 , n20345 , n19606 );
nand ( n20644 , n20642 , n20643 );
not ( n20645 , n20644 );
or ( n20646 , n20639 , n20645 );
not ( n20647 , n20411 );
not ( n20648 , n19636 );
or ( n20649 , n20647 , n20648 );
nand ( n20650 , n20424 , n19588 );
nand ( n20651 , n20649 , n20650 );
nand ( n20652 , n19642 , n20651 );
nand ( n20653 , n20646 , n20652 );
xor ( n20654 , n20638 , n20653 );
xor ( n20655 , n20630 , n20654 );
not ( n20656 , n19326 );
not ( n20657 , n19330 );
not ( n20658 , n19434 );
or ( n20659 , n20657 , n20658 );
not ( n20660 , n19340 );
or ( n20661 , n19434 , n20660 );
nand ( n20662 , n20659 , n20661 );
not ( n20663 , n20662 );
or ( n20664 , n20656 , n20663 );
nand ( n20665 , n20598 , n19336 );
nand ( n20666 , n20664 , n20665 );
xor ( n20667 , n20655 , n20666 );
xor ( n20668 , n20614 , n20667 );
not ( n20669 , n19578 );
not ( n20670 , n19483 );
not ( n20671 , n20254 );
or ( n20672 , n20670 , n20671 );
nand ( n20673 , n19844 , n19573 );
nand ( n20674 , n20672 , n20673 );
not ( n20675 , n20674 );
or ( n20676 , n20669 , n20675 );
not ( n20677 , n19483 );
not ( n20678 , n19889 );
or ( n20679 , n20677 , n20678 );
nand ( n20680 , n19888 , n19573 );
nand ( n20681 , n20679 , n20680 );
nand ( n20682 , n20681 , n19481 );
nand ( n20683 , n20676 , n20682 );
nor ( n20684 , n19584 , n20421 );
not ( n20685 , n19742 );
not ( n20686 , n20628 );
or ( n20687 , n20685 , n20686 );
nand ( n20688 , n20574 , n19783 );
nand ( n20689 , n20687 , n20688 );
xor ( n20690 , n20684 , n20689 );
not ( n20691 , n19578 );
not ( n20692 , n20681 );
or ( n20693 , n20691 , n20692 );
not ( n20694 , n19483 );
not ( n20695 , n20482 );
or ( n20696 , n20694 , n20695 );
nand ( n20697 , n20092 , n19573 );
nand ( n20698 , n20696 , n20697 );
nand ( n20699 , n20698 , n19480 );
nand ( n20700 , n20693 , n20699 );
and ( n20701 , n20690 , n20700 );
and ( n20702 , n20684 , n20689 );
or ( n20703 , n20701 , n20702 );
xor ( n20704 , n20683 , n20703 );
not ( n20705 , n19876 );
not ( n20706 , n19878 );
not ( n20707 , n19667 );
or ( n20708 , n20706 , n20707 );
nand ( n20709 , n19666 , n20095 );
nand ( n20710 , n20708 , n20709 );
not ( n20711 , n20710 );
or ( n20712 , n20705 , n20711 );
nand ( n20713 , n20603 , n19875 );
nand ( n20714 , n20712 , n20713 );
xor ( n20715 , n20704 , n20714 );
xor ( n20716 , n20668 , n20715 );
xor ( n20717 , n20684 , n20689 );
xor ( n20718 , n20717 , n20700 );
not ( n20719 , n19578 );
not ( n20720 , n20698 );
or ( n20721 , n20719 , n20720 );
not ( n20722 , n19483 );
not ( n20723 , n20330 );
or ( n20724 , n20722 , n20723 );
not ( n20725 , n19483 );
nand ( n20726 , n20329 , n20725 );
nand ( n20727 , n20724 , n20726 );
nand ( n20728 , n20727 , n19480 );
nand ( n20729 , n20721 , n20728 );
xor ( n20730 , n20580 , n20588 );
xor ( n20731 , n20729 , n20730 );
not ( n20732 , n19326 );
not ( n20733 , n20595 );
or ( n20734 , n20732 , n20733 );
not ( n20735 , n19340 );
not ( n20736 , n19889 );
or ( n20737 , n20735 , n20736 );
nand ( n20738 , n20108 , n20660 );
nand ( n20739 , n20737 , n20738 );
nand ( n20740 , n20739 , n19809 );
nand ( n20741 , n20734 , n20740 );
and ( n20742 , n20731 , n20741 );
and ( n20743 , n20729 , n20730 );
or ( n20744 , n20742 , n20743 );
xor ( n20745 , n20718 , n20744 );
xor ( n20746 , n20589 , n20600 );
xor ( n20747 , n20746 , n20611 );
and ( n20748 , n20745 , n20747 );
and ( n20749 , n20718 , n20744 );
or ( n20750 , n20748 , n20749 );
or ( n20751 , n20716 , n20750 );
not ( n20752 , n20751 );
xor ( n20753 , n20718 , n20744 );
xor ( n20754 , n20753 , n20747 );
not ( n20755 , n19876 );
not ( n20756 , n20609 );
or ( n20757 , n20755 , n20756 );
and ( n20758 , n19878 , n19460 );
not ( n20759 , n19878 );
and ( n20760 , n20759 , n19459 );
or ( n20761 , n20758 , n20760 );
nand ( n20762 , n20761 , n19875 );
nand ( n20763 , n20757 , n20762 );
and ( n20764 , n20567 , n20425 );
not ( n20765 , n20345 );
nand ( n20766 , n19329 , n777 );
nor ( n20767 , n20766 , n19483 );
not ( n20768 , n20767 );
or ( n20769 , n20765 , n20768 );
not ( n20770 , n20345 );
not ( n20771 , n19329 );
nand ( n20772 , n20771 , n19469 );
nor ( n20773 , n20772 , n20725 );
nand ( n20774 , n20770 , n20773 , n19479 );
nand ( n20775 , n20769 , n20774 );
not ( n20776 , n20775 );
nand ( n20777 , n20727 , n19471 );
nand ( n20778 , n20776 , n20777 , C1 );
xor ( n20779 , n20764 , n20778 );
not ( n20780 , n20425 );
not ( n20781 , n19475 );
or ( n20782 , n20780 , n20781 );
nand ( n20783 , n19474 , n20424 );
nand ( n20784 , n20782 , n20783 );
and ( n20785 , n19479 , n20784 );
not ( n20786 , n20785 );
not ( n20787 , n19472 );
or ( n20788 , n20786 , n20787 );
xor ( n20789 , n19483 , n20345 );
nand ( n20790 , n20789 , n19471 );
nand ( n20791 , n20788 , n20790 );
not ( n20792 , n19475 );
nand ( n20793 , n20772 , n20411 );
nand ( n20794 , n20792 , n20766 , n20793 );
not ( n20795 , n20794 );
and ( n20796 , n20791 , n20795 );
and ( n20797 , n20779 , n20796 );
and ( n20798 , n20764 , n20778 );
or ( n20799 , n20797 , n20798 );
xor ( n20800 , n20763 , n20799 );
xor ( n20801 , n20729 , n20730 );
xor ( n20802 , n20801 , n20741 );
and ( n20803 , n20800 , n20802 );
and ( n20804 , n20763 , n20799 );
or ( n20805 , n20803 , n20804 );
or ( n20806 , n20754 , n20805 );
not ( n20807 , n19326 );
not ( n20808 , n20739 );
or ( n20809 , n20807 , n20808 );
and ( n20810 , n19340 , n20482 );
not ( n20811 , n19340 );
and ( n20812 , n20811 , n20092 );
or ( n20813 , n20810 , n20812 );
nand ( n20814 , n20813 , n19809 );
nand ( n20815 , n20809 , n20814 );
not ( n20816 , n19876 );
not ( n20817 , n20761 );
or ( n20818 , n20816 , n20817 );
not ( n20819 , n19878 );
not ( n20820 , n20254 );
or ( n20821 , n20819 , n20820 );
nand ( n20822 , n19844 , n20095 );
nand ( n20823 , n20821 , n20822 );
nand ( n20824 , n20823 , n19875 );
nand ( n20825 , n20818 , n20824 );
xor ( n20826 , n20815 , n20825 );
xor ( n20827 , n20764 , n20778 );
xor ( n20828 , n20827 , n20796 );
xor ( n20829 , n20826 , n20828 );
not ( n20830 , n20829 );
not ( n20831 , n19326 );
not ( n20832 , n20813 );
or ( n20833 , n20831 , n20832 );
not ( n20834 , n19340 );
not ( n20835 , n20624 );
or ( n20836 , n20834 , n20835 );
not ( n20837 , n20591 );
not ( n20838 , n20624 );
nand ( n20839 , n20837 , n20838 );
nand ( n20840 , n20836 , n20839 );
nand ( n20841 , n20840 , n19336 );
nand ( n20842 , n20833 , n20841 );
not ( n20843 , n20790 );
not ( n20844 , n20795 );
and ( n20845 , n20843 , n20844 );
nor ( n20846 , n20794 , n20784 );
not ( n20847 , n20846 );
not ( n20848 , n20790 );
or ( n20849 , n20847 , n20848 );
nand ( n20850 , n20794 , n20785 , n19472 );
nand ( n20851 , n20849 , n20850 );
nor ( n20852 , n20845 , n20851 );
not ( n20853 , n19471 );
nand ( n20854 , n20853 , n19479 );
nand ( n20855 , n20854 , n20790 , n20795 );
nand ( n20856 , n20852 , n20855 );
xor ( n20857 , n20842 , n20856 );
not ( n20858 , n19876 );
not ( n20859 , n20823 );
or ( n20860 , n20858 , n20859 );
and ( n20861 , n19878 , n19889 );
not ( n20862 , n19878 );
and ( n20863 , n20862 , n20108 );
or ( n20864 , n20861 , n20863 );
nand ( n20865 , n20864 , n19875 );
nand ( n20866 , n20860 , n20865 );
and ( n20867 , n20857 , n20866 );
and ( n20868 , n20842 , n20856 );
or ( n20869 , n20867 , n20868 );
not ( n20870 , n20869 );
nand ( n20871 , n20830 , n20870 );
not ( n20872 , n20871 );
not ( n20873 , n19876 );
not ( n20874 , n20864 );
or ( n20875 , n20873 , n20874 );
not ( n20876 , n19878 );
not ( n20877 , n20482 );
or ( n20878 , n20876 , n20877 );
nand ( n20879 , n20092 , n20095 );
nand ( n20880 , n20878 , n20879 );
nand ( n20881 , n20880 , n19875 );
nand ( n20882 , n20875 , n20881 );
and ( n20883 , n19471 , n20425 );
not ( n20884 , n19325 );
not ( n20885 , n20840 );
or ( n20886 , n20884 , n20885 );
not ( n20887 , n19340 );
not ( n20888 , n20570 );
or ( n20889 , n20887 , n20888 );
nand ( n20890 , n20345 , n20660 );
nand ( n20891 , n20889 , n20890 );
nand ( n20892 , n20891 , n19336 );
nand ( n20893 , n20886 , n20892 );
xor ( n20894 , n20883 , n20893 );
not ( n20895 , n19335 );
and ( n20896 , n20424 , n19340 );
not ( n20897 , n20424 );
and ( n20898 , n20897 , n19330 );
nor ( n20899 , n20896 , n20898 );
not ( n20900 , n20899 );
and ( n20901 , n20895 , n20900 );
and ( n20902 , n20891 , n19325 );
nor ( n20903 , n20901 , n20902 );
not ( n20904 , n703 );
buf ( n20905 , n691 );
not ( n20906 , n20905 );
or ( n20907 , n20904 , n20906 );
nand ( n20908 , n20907 , n20591 );
not ( n20909 , n20908 );
or ( n20910 , n19878 , n703 );
nand ( n20911 , n20910 , n20411 );
nand ( n20912 , n20909 , n20911 );
nor ( n20913 , n20903 , n20912 );
xor ( n20914 , n20894 , n20913 );
xor ( n20915 , n20882 , n20914 );
not ( n20916 , n19874 );
xor ( n20917 , n20905 , n20345 );
not ( n20918 , n20917 );
or ( n20919 , n20916 , n20918 );
and ( n20920 , n20905 , n20329 );
not ( n20921 , n20905 );
and ( n20922 , n20921 , n20624 );
nor ( n20923 , n20920 , n20922 );
nand ( n20924 , n20923 , n19876 );
nand ( n20925 , n20919 , n20924 );
not ( n20926 , n20925 );
nand ( n20927 , n19326 , n20425 );
nand ( n20928 , n20926 , n20927 );
not ( n20929 , n20425 );
not ( n20930 , n19874 );
not ( n20931 , n20930 );
and ( n20932 , n20929 , n20931 );
and ( n20933 , n20917 , n19876 );
nor ( n20934 , n20932 , n20933 );
nand ( n20935 , n20425 , n19876 );
nand ( n20936 , n20935 , n19878 );
nor ( n20937 , n20934 , n20936 );
buf ( n20938 , n20937 );
and ( n20939 , n20928 , n20938 );
not ( n20940 , n20927 );
nand ( n20941 , n20940 , n20925 );
not ( n20942 , n20941 );
nor ( n20943 , n20939 , n20942 );
xor ( n20944 , n20912 , n20903 );
not ( n20945 , n19876 );
not ( n20946 , n20880 );
or ( n20947 , n20945 , n20946 );
nand ( n20948 , n20923 , n19875 );
nand ( n20949 , n20947 , n20948 );
nor ( n20950 , n20944 , n20949 );
or ( n20951 , n20943 , n20950 );
nand ( n20952 , n20944 , n20949 );
nand ( n20953 , n20951 , n20952 );
and ( n20954 , n20915 , n20953 );
and ( n20955 , n20882 , n20914 );
or ( n20956 , n20954 , n20955 );
not ( n20957 , n20956 );
xor ( n20958 , n20842 , n20856 );
xor ( n20959 , n20958 , n20866 );
not ( n20960 , n20959 );
xor ( n20961 , n20883 , n20893 );
and ( n20962 , n20961 , n20913 );
and ( n20963 , n20883 , n20893 );
or ( n20964 , n20962 , n20963 );
not ( n20965 , n20964 );
nand ( n20966 , n20960 , n20965 );
not ( n20967 , n20966 );
or ( n20968 , n20957 , n20967 );
buf ( n20969 , n20959 );
nand ( n20970 , n20969 , n20964 );
nand ( n20971 , n20968 , n20970 );
not ( n20972 , n20971 );
or ( n20973 , n20872 , n20972 );
nand ( n20974 , n20829 , n20869 );
nand ( n20975 , n20973 , n20974 );
xor ( n20976 , n20763 , n20799 );
xor ( n20977 , n20976 , n20802 );
xor ( n20978 , n20815 , n20825 );
and ( n20979 , n20978 , n20828 );
and ( n20980 , n20815 , n20825 );
or ( n20981 , n20979 , n20980 );
or ( n20982 , n20977 , n20981 );
nand ( n20983 , n20806 , n20975 , n20982 );
and ( n20984 , n20977 , n20981 );
nand ( n20985 , n20806 , n20984 );
buf ( n20986 , n20754 );
nand ( n20987 , n20986 , n20805 );
nand ( n20988 , n20983 , n20985 , n20987 );
not ( n20989 , n20988 );
or ( n20990 , n20752 , n20989 );
nand ( n20991 , n20716 , n20750 );
nand ( n20992 , n20990 , n20991 );
not ( n20993 , n20992 );
not ( n20994 , n19578 );
not ( n20995 , n19483 );
not ( n20996 , n19435 );
or ( n20997 , n20995 , n20996 );
nand ( n20998 , n19436 , n19573 );
nand ( n20999 , n20997 , n20998 );
not ( n21000 , n20999 );
or ( n21001 , n20994 , n21000 );
and ( n21002 , n19460 , n19483 );
not ( n21003 , n19460 );
and ( n21004 , n21003 , n19573 );
or ( n21005 , n21002 , n21004 );
nand ( n21006 , n21005 , n19481 );
nand ( n21007 , n21001 , n21006 );
and ( n21008 , n19653 , n20411 );
not ( n21009 , n19585 );
not ( n21010 , n19588 );
not ( n21011 , n20624 );
or ( n21012 , n21010 , n21011 );
nand ( n21013 , n20329 , n19606 );
nand ( n21014 , n21012 , n21013 );
not ( n21015 , n21014 );
or ( n21016 , n21009 , n21015 );
nand ( n21017 , n20644 , n19642 );
nand ( n21018 , n21016 , n21017 );
xor ( n21019 , n21008 , n21018 );
not ( n21020 , n19742 );
not ( n21021 , n19744 );
not ( n21022 , n19889 );
or ( n21023 , n21021 , n21022 );
not ( n21024 , n11108 );
nand ( n21025 , n21024 , n19888 );
nand ( n21026 , n21023 , n21025 );
not ( n21027 , n21026 );
or ( n21028 , n21020 , n21027 );
nand ( n21029 , n20620 , n19783 );
nand ( n21030 , n21028 , n21029 );
and ( n21031 , n21019 , n21030 );
and ( n21032 , n21008 , n21018 );
or ( n21033 , n21031 , n21032 );
xor ( n21034 , n21007 , n21033 );
not ( n21035 , n19326 );
not ( n21036 , n19340 );
not ( n21037 , n19667 );
or ( n21038 , n21036 , n21037 );
nand ( n21039 , n19666 , n20169 );
nand ( n21040 , n21038 , n21039 );
not ( n21041 , n21040 );
or ( n21042 , n21035 , n21041 );
and ( n21043 , n19397 , n20660 );
not ( n21044 , n19397 );
and ( n21045 , n21044 , n19340 );
or ( n21046 , n21043 , n21045 );
nand ( n21047 , n21046 , n19809 );
nand ( n21048 , n21042 , n21047 );
xor ( n21049 , n21034 , n21048 );
xor ( n21050 , n21008 , n21018 );
xor ( n21051 , n21050 , n21030 );
not ( n21052 , n19875 );
not ( n21053 , n20710 );
or ( n21054 , n21052 , n21053 );
not ( n21055 , n19878 );
not ( n21056 , n19683 );
or ( n21057 , n21055 , n21056 );
nand ( n21058 , n19682 , n20095 );
nand ( n21059 , n21057 , n21058 );
nand ( n21060 , n21059 , n19876 );
nand ( n21061 , n21054 , n21060 );
xor ( n21062 , n21051 , n21061 );
xor ( n21063 , n20630 , n20654 );
and ( n21064 , n21063 , n20666 );
and ( n21065 , n20630 , n20654 );
or ( n21066 , n21064 , n21065 );
and ( n21067 , n21062 , n21066 );
and ( n21068 , n21051 , n21061 );
or ( n21069 , n21067 , n21068 );
xor ( n21070 , n21049 , n21069 );
not ( n21071 , n19876 );
not ( n21072 , n19878 );
not ( n21073 , n19628 );
or ( n21074 , n21072 , n21073 );
nand ( n21075 , n19627 , n20095 );
nand ( n21076 , n21074 , n21075 );
not ( n21077 , n21076 );
or ( n21078 , n21071 , n21077 );
nand ( n21079 , n21059 , n19875 );
nand ( n21080 , n21078 , n21079 );
not ( n21081 , n19585 );
not ( n21082 , n19588 );
not ( n21083 , n20482 );
or ( n21084 , n21082 , n21083 );
nand ( n21085 , n20092 , n19606 );
nand ( n21086 , n21084 , n21085 );
not ( n21087 , n21086 );
or ( n21088 , n21081 , n21087 );
nand ( n21089 , n21014 , n19643 );
nand ( n21090 , n21088 , n21089 );
nand ( n21091 , n19636 , n19648 );
and ( n21092 , n21091 , n20411 );
not ( n21093 , n19647 );
not ( n21094 , n19588 );
or ( n21095 , n21093 , n21094 );
nand ( n21096 , n21095 , n19657 );
nor ( n21097 , n21092 , n21096 );
not ( n21098 , n19653 );
not ( n21099 , n19657 );
not ( n21100 , n20570 );
or ( n21101 , n21099 , n21100 );
nand ( n21102 , n20345 , n10146 );
nand ( n21103 , n21101 , n21102 );
not ( n21104 , n21103 );
or ( n21105 , n21098 , n21104 );
not ( n21106 , n20411 );
not ( n21107 , n10146 );
or ( n21108 , n21106 , n21107 );
nand ( n21109 , n20424 , n19657 );
nand ( n21110 , n21108 , n21109 );
nand ( n21111 , n19654 , n21110 );
nand ( n21112 , n21105 , n21111 );
xor ( n21113 , n21097 , n21112 );
xor ( n21114 , n21090 , n21113 );
not ( n21115 , n19742 );
not ( n21116 , n19744 );
not ( n21117 , n20254 );
or ( n21118 , n21116 , n21117 );
nand ( n21119 , n19844 , n11107 );
nand ( n21120 , n21118 , n21119 );
not ( n21121 , n21120 );
or ( n21122 , n21115 , n21121 );
nand ( n21123 , n21026 , n19784 );
nand ( n21124 , n21122 , n21123 );
xor ( n21125 , n21114 , n21124 );
xor ( n21126 , n21080 , n21125 );
and ( n21127 , n20638 , n20653 );
not ( n21128 , n19326 );
not ( n21129 , n21046 );
or ( n21130 , n21128 , n21129 );
nand ( n21131 , n20662 , n19809 );
nand ( n21132 , n21130 , n21131 );
xor ( n21133 , n21127 , n21132 );
not ( n21134 , n19481 );
not ( n21135 , n20674 );
or ( n21136 , n21134 , n21135 );
nand ( n21137 , n21005 , n19578 );
nand ( n21138 , n21136 , n21137 );
and ( n21139 , n21133 , n21138 );
and ( n21140 , n21127 , n21132 );
or ( n21141 , n21139 , n21140 );
xor ( n21142 , n21126 , n21141 );
xor ( n21143 , n21070 , n21142 );
not ( n21144 , n21143 );
xor ( n21145 , n21127 , n21132 );
xor ( n21146 , n21145 , n21138 );
xor ( n21147 , n20683 , n20703 );
and ( n21148 , n21147 , n20714 );
and ( n21149 , n20683 , n20703 );
or ( n21150 , n21148 , n21149 );
xor ( n21151 , n21146 , n21150 );
xor ( n21152 , n21051 , n21061 );
xor ( n21153 , n21152 , n21066 );
and ( n21154 , n21151 , n21153 );
and ( n21155 , n21146 , n21150 );
or ( n21156 , n21154 , n21155 );
not ( n21157 , n21156 );
and ( n21158 , n21144 , n21157 );
xor ( n21159 , n21146 , n21150 );
xor ( n21160 , n21159 , n21153 );
xor ( n21161 , n20614 , n20667 );
and ( n21162 , n21161 , n20715 );
and ( n21163 , n20614 , n20667 );
or ( n21164 , n21162 , n21163 );
nor ( n21165 , n21160 , n21164 );
nor ( n21166 , n21158 , n21165 );
not ( n21167 , n21166 );
or ( n21168 , n20993 , n21167 );
not ( n21169 , n21143 );
not ( n21170 , n21156 );
nand ( n21171 , n21169 , n21170 );
and ( n21172 , n21160 , n21164 );
and ( n21173 , n21171 , n21172 );
not ( n21174 , n21143 );
nor ( n21175 , n21174 , n21170 );
nor ( n21176 , n21173 , n21175 );
nand ( n21177 , n21168 , n21176 );
not ( n21178 , n19875 );
not ( n21179 , n19878 );
not ( n21180 , n19602 );
or ( n21181 , n21179 , n21180 );
nand ( n21182 , n19601 , n20095 );
nand ( n21183 , n21181 , n21182 );
not ( n21184 , n21183 );
or ( n21185 , n21178 , n21184 );
nand ( n21186 , n20532 , n19876 );
nand ( n21187 , n21185 , n21186 );
not ( n21188 , n19578 );
not ( n21189 , n19483 );
not ( n21190 , n19667 );
or ( n21191 , n21189 , n21190 );
nand ( n21192 , n19666 , n19573 );
nand ( n21193 , n21191 , n21192 );
not ( n21194 , n21193 );
or ( n21195 , n21188 , n21194 );
not ( n21196 , n19483 );
not ( n21197 , n19398 );
or ( n21198 , n21196 , n21197 );
nand ( n21199 , n19397 , n19573 );
nand ( n21200 , n21198 , n21199 );
nand ( n21201 , n21200 , n19481 );
nand ( n21202 , n21195 , n21201 );
xor ( n21203 , n21187 , n21202 );
not ( n21204 , n19690 );
not ( n21205 , n20486 );
or ( n21206 , n21204 , n21205 );
and ( n21207 , n19657 , n20624 );
not ( n21208 , n19657 );
and ( n21209 , n21208 , n20127 );
or ( n21210 , n21207 , n21209 );
nand ( n21211 , n21210 , n19655 );
nand ( n21212 , n21206 , n21211 );
xor ( n21213 , n20431 , n20436 );
xor ( n21214 , n21212 , n21213 );
not ( n21215 , n19585 );
not ( n21216 , n20493 );
or ( n21217 , n21215 , n21216 );
not ( n21218 , n19588 );
not ( n21219 , n19889 );
or ( n21220 , n21218 , n21219 );
nand ( n21221 , n19890 , n19606 );
nand ( n21222 , n21220 , n21221 );
nand ( n21223 , n21222 , n19643 );
nand ( n21224 , n21217 , n21223 );
xor ( n21225 , n21214 , n21224 );
xor ( n21226 , n21203 , n21225 );
xor ( n21227 , n21090 , n21113 );
and ( n21228 , n21227 , n21124 );
and ( n21229 , n21090 , n21113 );
or ( n21230 , n21228 , n21229 );
not ( n21231 , n19585 );
not ( n21232 , n21222 );
or ( n21233 , n21231 , n21232 );
nand ( n21234 , n21086 , n19643 );
nand ( n21235 , n21233 , n21234 );
not ( n21236 , n19481 );
not ( n21237 , n20999 );
or ( n21238 , n21236 , n21237 );
nand ( n21239 , n21200 , n19578 );
nand ( n21240 , n21238 , n21239 );
xor ( n21241 , n21235 , n21240 );
not ( n21242 , n19742 );
and ( n21243 , n19460 , n19744 );
not ( n21244 , n19460 );
and ( n21245 , n21244 , n11107 );
or ( n21246 , n21243 , n21245 );
not ( n21247 , n21246 );
or ( n21248 , n21242 , n21247 );
nand ( n21249 , n21120 , n19784 );
nand ( n21250 , n21248 , n21249 );
xor ( n21251 , n21241 , n21250 );
xor ( n21252 , n21230 , n21251 );
xor ( n21253 , n21007 , n21033 );
and ( n21254 , n21253 , n21048 );
and ( n21255 , n21007 , n21033 );
or ( n21256 , n21254 , n21255 );
and ( n21257 , n21252 , n21256 );
and ( n21258 , n21230 , n21251 );
or ( n21259 , n21257 , n21258 );
xor ( n21260 , n21226 , n21259 );
xor ( n21261 , n21235 , n21240 );
and ( n21262 , n21261 , n21250 );
and ( n21263 , n21235 , n21240 );
or ( n21264 , n21262 , n21263 );
not ( n21265 , n19326 );
not ( n21266 , n19340 );
not ( n21267 , n19683 );
or ( n21268 , n21266 , n21267 );
nand ( n21269 , n19682 , n20169 );
nand ( n21270 , n21268 , n21269 );
not ( n21271 , n21270 );
or ( n21272 , n21265 , n21271 );
nand ( n21273 , n21040 , n19809 );
nand ( n21274 , n21272 , n21273 );
and ( n21275 , n19348 , n20425 );
not ( n21276 , n19690 );
not ( n21277 , n21210 );
or ( n21278 , n21276 , n21277 );
nand ( n21279 , n21103 , n19655 );
nand ( n21280 , n21278 , n21279 );
xor ( n21281 , n21275 , n21280 );
and ( n21282 , n21097 , n21112 );
xor ( n21283 , n21281 , n21282 );
xor ( n21284 , n21274 , n21283 );
not ( n21285 , n19876 );
not ( n21286 , n21183 );
or ( n21287 , n21285 , n21286 );
nand ( n21288 , n21076 , n19875 );
nand ( n21289 , n21287 , n21288 );
and ( n21290 , n21284 , n21289 );
and ( n21291 , n21274 , n21283 );
or ( n21292 , n21290 , n21291 );
xor ( n21293 , n21264 , n21292 );
not ( n21294 , n19742 );
not ( n21295 , n20504 );
or ( n21296 , n21294 , n21295 );
nand ( n21297 , n21246 , n19784 );
nand ( n21298 , n21296 , n21297 );
not ( n21299 , n19326 );
not ( n21300 , n20522 );
or ( n21301 , n21299 , n21300 );
nand ( n21302 , n21270 , n19809 );
nand ( n21303 , n21301 , n21302 );
xor ( n21304 , n21298 , n21303 );
xor ( n21305 , n21275 , n21280 );
and ( n21306 , n21305 , n21282 );
and ( n21307 , n21275 , n21280 );
or ( n21308 , n21306 , n21307 );
xor ( n21309 , n21304 , n21308 );
xor ( n21310 , n21293 , n21309 );
xor ( n21311 , n21260 , n21310 );
not ( n21312 , n21311 );
xor ( n21313 , n21274 , n21283 );
xor ( n21314 , n21313 , n21289 );
xor ( n21315 , n21080 , n21125 );
and ( n21316 , n21315 , n21141 );
and ( n21317 , n21080 , n21125 );
or ( n21318 , n21316 , n21317 );
xor ( n21319 , n21314 , n21318 );
xor ( n21320 , n21230 , n21251 );
xor ( n21321 , n21320 , n21256 );
and ( n21322 , n21319 , n21321 );
and ( n21323 , n21314 , n21318 );
or ( n21324 , n21322 , n21323 );
not ( n21325 , n21324 );
nand ( n21326 , n21312 , n21325 );
xor ( n21327 , n21314 , n21318 );
xor ( n21328 , n21327 , n21321 );
xor ( n21329 , n21049 , n21069 );
and ( n21330 , n21329 , n21142 );
and ( n21331 , n21049 , n21069 );
or ( n21332 , n21330 , n21331 );
or ( n21333 , n21328 , n21332 );
nand ( n21334 , n21177 , n21326 , n21333 );
not ( n21335 , n21311 );
nand ( n21336 , n21335 , n21325 );
and ( n21337 , n21328 , n21332 );
nand ( n21338 , n21336 , n21337 );
nand ( n21339 , n21311 , n21324 );
nand ( n21340 , n21334 , n21338 , n21339 );
not ( n21341 , n21340 );
not ( n21342 , n19481 );
not ( n21343 , n21193 );
or ( n21344 , n21342 , n21343 );
nand ( n21345 , n20447 , n19578 );
nand ( n21346 , n21344 , n21345 );
xor ( n21347 , n21212 , n21213 );
and ( n21348 , n21347 , n21224 );
and ( n21349 , n21212 , n21213 );
or ( n21350 , n21348 , n21349 );
xor ( n21351 , n21346 , n21350 );
xor ( n21352 , n20488 , n20497 );
xor ( n21353 , n21352 , n20508 );
xor ( n21354 , n21351 , n21353 );
xor ( n21355 , n21264 , n21292 );
and ( n21356 , n21355 , n21309 );
and ( n21357 , n21264 , n21292 );
or ( n21358 , n21356 , n21357 );
xor ( n21359 , n21354 , n21358 );
xor ( n21360 , n21298 , n21303 );
and ( n21361 , n21360 , n21308 );
and ( n21362 , n21298 , n21303 );
or ( n21363 , n21361 , n21362 );
xor ( n21364 , n20516 , n20526 );
xor ( n21365 , n21364 , n20537 );
xor ( n21366 , n21363 , n21365 );
xor ( n21367 , n21187 , n21202 );
and ( n21368 , n21367 , n21225 );
and ( n21369 , n21187 , n21202 );
or ( n21370 , n21368 , n21369 );
xor ( n21371 , n21366 , n21370 );
xor ( n21372 , n21359 , n21371 );
not ( n21373 , n21372 );
xor ( n21374 , n21226 , n21259 );
and ( n21375 , n21374 , n21310 );
and ( n21376 , n21226 , n21259 );
or ( n21377 , n21375 , n21376 );
not ( n21378 , n21377 );
and ( n21379 , n21373 , n21378 );
xor ( n21380 , n21346 , n21350 );
and ( n21381 , n21380 , n21353 );
and ( n21382 , n21346 , n21350 );
or ( n21383 , n21381 , n21382 );
xor ( n21384 , n21363 , n21365 );
and ( n21385 , n21384 , n21370 );
and ( n21386 , n21363 , n21365 );
or ( n21387 , n21385 , n21386 );
xor ( n21388 , n21383 , n21387 );
xor ( n21389 , n20409 , n20440 );
xor ( n21390 , n21389 , n20451 );
xor ( n21391 , n20376 , n20388 );
xor ( n21392 , n21391 , n20396 );
xor ( n21393 , n21390 , n21392 );
xor ( n21394 , n20511 , n20513 );
xor ( n21395 , n21394 , n20540 );
xor ( n21396 , n21393 , n21395 );
xor ( n21397 , n21388 , n21396 );
xor ( n21398 , n21354 , n21358 );
and ( n21399 , n21398 , n21371 );
and ( n21400 , n21354 , n21358 );
or ( n21401 , n21399 , n21400 );
nor ( n21402 , n21397 , n21401 );
nor ( n21403 , n21379 , n21402 );
not ( n21404 , n21403 );
or ( n21405 , n21341 , n21404 );
not ( n21406 , n21402 );
nand ( n21407 , n21372 , n21377 );
not ( n21408 , n21407 );
and ( n21409 , n21406 , n21408 );
nand ( n21410 , n21397 , n21401 );
not ( n21411 , n21410 );
nor ( n21412 , n21409 , n21411 );
nand ( n21413 , n21405 , n21412 );
nor ( n21414 , n20466 , n20302 );
nor ( n21415 , n20549 , n20551 );
nor ( n21416 , n21414 , n21415 );
xor ( n21417 , n20469 , n20471 );
xor ( n21418 , n21417 , n20546 );
not ( n21419 , n21418 );
xor ( n21420 , n20366 , n20399 );
xor ( n21421 , n21420 , n20454 );
xor ( n21422 , n20474 , n20476 );
xor ( n21423 , n21422 , n20543 );
xor ( n21424 , n21421 , n21423 );
xor ( n21425 , n21390 , n21392 );
and ( n21426 , n21425 , n21395 );
and ( n21427 , n21390 , n21392 );
or ( n21428 , n21426 , n21427 );
and ( n21429 , n21424 , n21428 );
and ( n21430 , n21421 , n21423 );
or ( n21431 , n21429 , n21430 );
not ( n21432 , n21431 );
and ( n21433 , n21419 , n21432 );
xor ( n21434 , n21421 , n21423 );
xor ( n21435 , n21434 , n21428 );
xor ( n21436 , n21383 , n21387 );
and ( n21437 , n21436 , n21396 );
and ( n21438 , n21383 , n21387 );
or ( n21439 , n21437 , n21438 );
nor ( n21440 , n21435 , n21439 );
nor ( n21441 , n21433 , n21440 );
nand ( n21442 , n21413 , n21416 , n20299 , n21441 );
and ( n21443 , n21435 , n21439 );
not ( n21444 , n21443 );
not ( n21445 , n21418 );
not ( n21446 , n21431 );
nand ( n21447 , n21445 , n21446 );
not ( n21448 , n21447 );
or ( n21449 , n21444 , n21448 );
nand ( n21450 , n21418 , n21431 );
nand ( n21451 , n21449 , n21450 );
nand ( n21452 , n20299 , n21416 , n21451 );
nand ( n21453 , n20566 , n21442 , n21452 );
buf ( n21454 , n21453 );
xor ( n21455 , n20042 , n21454 );
buf ( n21456 , n21455 );
and ( n21457 , n19319 , n21456 );
not ( n21458 , n19319 );
not ( n21459 , n21456 );
and ( n21460 , n21458 , n21459 );
nor ( n21461 , n21457 , n21460 );
not ( n21462 , n21461 );
or ( n21463 , n19317 , n21462 );
not ( n21464 , n20041 );
not ( n21465 , n21464 );
not ( n21466 , n21454 );
or ( n21467 , n21465 , n21466 );
nand ( n21468 , n21467 , n20039 );
not ( n21469 , n19690 );
not ( n21470 , n19657 );
not ( n21471 , n19720 );
or ( n21472 , n21470 , n21471 );
or ( n21473 , n19720 , n19657 );
nand ( n21474 , n21472 , n21473 );
not ( n21475 , n21474 );
or ( n21476 , n21469 , n21475 );
not ( n21477 , n19990 );
not ( n21478 , n19655 );
or ( n21479 , n21477 , n21478 );
nand ( n21480 , n21476 , n21479 );
not ( n21481 , n20027 );
not ( n21482 , n19784 );
or ( n21483 , n21481 , n21482 );
or ( n21484 , n20386 , n11107 );
nand ( n21485 , n21483 , n21484 );
not ( n21486 , n21485 );
xor ( n21487 , n21480 , n21486 );
xor ( n21488 , n19992 , n19998 );
and ( n21489 , n21488 , n20005 );
and ( n21490 , n19992 , n19998 );
or ( n21491 , n21489 , n21490 );
xor ( n21492 , n21487 , n21491 );
xor ( n21493 , n20017 , n20018 );
and ( n21494 , n21493 , n20029 );
and ( n21495 , n20017 , n20018 );
or ( n21496 , n21494 , n21495 );
not ( n21497 , n19643 );
not ( n21498 , n20003 );
or ( n21499 , n21497 , n21498 );
not ( n21500 , n19588 );
not ( n21501 , n19747 );
or ( n21502 , n21500 , n21501 );
nand ( n21503 , n19746 , n19606 );
nand ( n21504 , n21502 , n21503 );
nand ( n21505 , n21504 , n19585 );
nand ( n21506 , n21499 , n21505 );
not ( n21507 , n19348 );
xor ( n21508 , n19351 , n19627 );
not ( n21509 , n21508 );
or ( n21510 , n21507 , n21509 );
nand ( n21511 , n19996 , n19443 );
nand ( n21512 , n21510 , n21511 );
xor ( n21513 , n21506 , n21512 );
and ( n21514 , n19351 , n19666 );
xor ( n21515 , n21513 , n21514 );
xor ( n21516 , n21496 , n21515 );
xor ( n21517 , n20008 , n20012 );
and ( n21518 , n21517 , n20030 );
and ( n21519 , n20008 , n20012 );
or ( n21520 , n21518 , n21519 );
xor ( n21521 , n21516 , n21520 );
xor ( n21522 , n21492 , n21521 );
xor ( n21523 , n19981 , n20006 );
and ( n21524 , n21523 , n20031 );
and ( n21525 , n19981 , n20006 );
or ( n21526 , n21524 , n21525 );
xor ( n21527 , n21522 , n21526 );
not ( n21528 , n21527 );
xor ( n21529 , n19977 , n20032 );
and ( n21530 , n21529 , n20037 );
and ( n21531 , n19977 , n20032 );
or ( n21532 , n21530 , n21531 );
not ( n21533 , n21532 );
nor ( n21534 , n21528 , n21533 );
not ( n21535 , n21534 );
nand ( n21536 , n21528 , n21533 );
nand ( n21537 , n21535 , n21536 );
not ( n21538 , n21537 );
and ( n21539 , n21468 , n21538 );
not ( n21540 , n21468 );
and ( n21541 , n21540 , n21537 );
nor ( n21542 , n21539 , n21541 );
buf ( n21543 , n21542 );
and ( n21544 , n19319 , n21543 );
not ( n21545 , n19319 );
not ( n21546 , n21543 );
and ( n21547 , n21545 , n21546 );
nor ( n21548 , n21544 , n21547 );
buf ( n21549 , n19292 );
nand ( n21550 , n21548 , n21549 );
nand ( n21551 , n21463 , n21550 );
nor ( n21552 , n19303 , n19275 );
nand ( n21553 , n21552 , n19225 );
not ( n21554 , n21553 );
not ( n21555 , n21554 );
not ( n21556 , n19296 );
or ( n21557 , n21555 , n21556 );
not ( n21558 , n19272 );
not ( n21559 , n21552 );
or ( n21560 , n21558 , n21559 );
not ( n21561 , n19303 );
not ( n21562 , n19277 );
and ( n21563 , n21561 , n21562 );
nor ( n21564 , n21563 , n19304 );
nand ( n21565 , n21560 , n21564 );
not ( n21566 , n21565 );
nand ( n21567 , n21557 , n21566 );
nor ( n21568 , n524 , n540 );
not ( n21569 , n21568 );
nand ( n21570 , n524 , n540 );
and ( n21571 , n21569 , n21570 );
xor ( n21572 , n21567 , n21571 );
and ( n21573 , n21572 , n19310 );
not ( n21574 , n21572 );
and ( n21575 , n21574 , n19311 );
nor ( n21576 , n21573 , n21575 );
not ( n21577 , n21576 );
not ( n21578 , n21577 );
nor ( n21579 , n21553 , n21568 );
not ( n21580 , n21579 );
not ( n21581 , n19266 );
or ( n21582 , n21580 , n21581 );
not ( n21583 , n21569 );
not ( n21584 , n21565 );
or ( n21585 , n21583 , n21584 );
nand ( n21586 , n21585 , n21570 );
not ( n21587 , n21586 );
nand ( n21588 , n21582 , n21587 );
nor ( n21589 , n523 , n539 );
not ( n21590 , n21589 );
nand ( n21591 , n523 , n539 );
nand ( n21592 , n21590 , n21591 );
xnor ( n21593 , n21588 , n21592 );
not ( n21594 , n21593 );
not ( n21595 , n21594 );
not ( n21596 , n21595 );
not ( n21597 , n20298 );
not ( n21598 , n21597 );
not ( n21599 , n21416 );
not ( n21600 , n21441 );
not ( n21601 , n21403 );
not ( n21602 , n21340 );
or ( n21603 , n21601 , n21602 );
nand ( n21604 , n21603 , n21412 );
not ( n21605 , n21604 );
or ( n21606 , n21600 , n21605 );
not ( n21607 , n21451 );
nand ( n21608 , n21606 , n21607 );
not ( n21609 , n21608 );
or ( n21610 , n21599 , n21609 );
not ( n21611 , n20555 );
nand ( n21612 , n21610 , n21611 );
not ( n21613 , n21612 );
or ( n21614 , n21598 , n21613 );
not ( n21615 , n20561 );
nand ( n21616 , n21614 , n21615 );
not ( n21617 , n20563 );
nand ( n21618 , n21617 , n20560 );
xnor ( n21619 , n21616 , n21618 );
not ( n21620 , n21619 );
not ( n21621 , n21620 );
or ( n21622 , n21596 , n21621 );
not ( n21623 , n21595 );
nand ( n21624 , n21619 , n21623 );
nand ( n21625 , n21622 , n21624 );
not ( n21626 , n21625 );
or ( n21627 , n21578 , n21626 );
not ( n21628 , n21595 );
nand ( n21629 , n21597 , n21615 );
not ( n21630 , n21629 );
not ( n21631 , n21630 );
not ( n21632 , n21612 );
not ( n21633 , n21632 );
or ( n21634 , n21631 , n21633 );
nand ( n21635 , n21612 , n21629 );
nand ( n21636 , n21634 , n21635 );
not ( n21637 , n21636 );
not ( n21638 , n21637 );
or ( n21639 , n21628 , n21638 );
nand ( n21640 , n21636 , n21623 );
nand ( n21641 , n21639 , n21640 );
not ( n21642 , n21572 );
and ( n21643 , n21594 , n21642 );
and ( n21644 , n21593 , n21572 );
nor ( n21645 , n21643 , n21644 );
and ( n21646 , n21576 , n21645 );
nand ( n21647 , n21641 , n21646 );
nand ( n21648 , n21627 , n21647 );
xor ( n21649 , n21551 , n21648 );
not ( n21650 , n19291 );
not ( n21651 , n21650 );
and ( n21652 , n19284 , n19269 );
and ( n21653 , n21652 , n19296 );
not ( n21654 , n21652 );
not ( n21655 , n19296 );
and ( n21656 , n21654 , n21655 );
or ( n21657 , n21653 , n21656 );
not ( n21658 , n21657 );
or ( n21659 , n21651 , n21658 );
or ( n21660 , n21650 , n21657 );
nand ( n21661 , n21659 , n21660 );
not ( n21662 , n21657 );
nand ( n21663 , n19243 , n19252 );
not ( n21664 , n21663 );
nor ( n21665 , n19242 , n19246 );
not ( n21666 , n21665 );
nor ( n21667 , n19231 , n19244 );
not ( n21668 , n21667 );
not ( n21669 , n19227 );
not ( n21670 , n21669 );
not ( n21671 , n19230 );
or ( n21672 , n21670 , n21671 );
nand ( n21673 , n21672 , n19228 );
not ( n21674 , n21673 );
or ( n21675 , n21668 , n21674 );
not ( n21676 , n19236 );
nor ( n21677 , n19235 , n19244 );
nor ( n21678 , n21676 , n21677 );
nand ( n21679 , n21675 , n21678 );
not ( n21680 , n21679 );
or ( n21681 , n21666 , n21680 );
not ( n21682 , n19247 );
nand ( n21683 , n19258 , n19253 );
not ( n21684 , n21683 );
or ( n21685 , n21682 , n21684 );
nand ( n21686 , n21685 , n19251 );
not ( n21687 , n21686 );
nand ( n21688 , n21681 , n21687 );
not ( n21689 , n21688 );
or ( n21690 , n21664 , n21689 );
or ( n21691 , n21688 , n21663 );
nand ( n21692 , n21690 , n21691 );
not ( n21693 , n21692 );
or ( n21694 , n21662 , n21693 );
or ( n21695 , n21692 , n21657 );
nand ( n21696 , n21694 , n21695 );
nor ( n21697 , n21661 , n21696 );
buf ( n21698 , n21697 );
not ( n21699 , n21698 );
xor ( n21700 , n21492 , n21521 );
and ( n21701 , n21700 , n21526 );
and ( n21702 , n21492 , n21521 );
or ( n21703 , n21701 , n21702 );
xor ( n21704 , n21480 , n21486 );
and ( n21705 , n21704 , n21491 );
and ( n21706 , n21480 , n21486 );
or ( n21707 , n21705 , n21706 );
xor ( n21708 , n21506 , n21512 );
and ( n21709 , n21708 , n21514 );
and ( n21710 , n21506 , n21512 );
or ( n21711 , n21709 , n21710 );
not ( n21712 , n20386 );
not ( n21713 , n21482 );
or ( n21714 , n21712 , n21713 );
nand ( n21715 , n21714 , n19744 );
not ( n21716 , n19643 );
not ( n21717 , n21504 );
or ( n21718 , n21716 , n21717 );
and ( n21719 , n19588 , n19572 );
not ( n21720 , n19588 );
and ( n21721 , n21720 , n20023 );
nor ( n21722 , n21719 , n21721 );
nand ( n21723 , n21722 , n19585 );
nand ( n21724 , n21718 , n21723 );
xor ( n21725 , n21715 , n21724 );
not ( n21726 , n19443 );
not ( n21727 , n21508 );
or ( n21728 , n21726 , n21727 );
xor ( n21729 , n19351 , n19988 );
not ( n21730 , n21729 );
or ( n21731 , n21730 , n19824 );
nand ( n21732 , n21728 , n21731 );
xor ( n21733 , n21725 , n21732 );
xor ( n21734 , n21711 , n21733 );
and ( n21735 , n19351 , n19686 );
not ( n21736 , n19690 );
not ( n21737 , n19657 );
not ( n21738 , n19774 );
not ( n21739 , n21738 );
or ( n21740 , n21737 , n21739 );
nand ( n21741 , n19774 , n19687 );
nand ( n21742 , n21740 , n21741 );
not ( n21743 , n21742 );
or ( n21744 , n21736 , n21743 );
nand ( n21745 , n21474 , n19655 );
nand ( n21746 , n21744 , n21745 );
xor ( n21747 , n21735 , n21746 );
xor ( n21748 , n21747 , n21485 );
xor ( n21749 , n21734 , n21748 );
xor ( n21750 , n21707 , n21749 );
xor ( n21751 , n21496 , n21515 );
and ( n21752 , n21751 , n21520 );
and ( n21753 , n21496 , n21515 );
or ( n21754 , n21752 , n21753 );
xor ( n21755 , n21750 , n21754 );
nor ( n21756 , n21703 , n21755 );
not ( n21757 , n21756 );
nand ( n21758 , n21703 , n21755 );
and ( n21759 , n21757 , n21758 );
not ( n21760 , n21536 );
nor ( n21761 , n21760 , n20041 );
not ( n21762 , n21761 );
not ( n21763 , n21453 );
or ( n21764 , n21762 , n21763 );
and ( n21765 , n20040 , n21536 );
nor ( n21766 , n21765 , n21534 );
nand ( n21767 , n21764 , n21766 );
xor ( n21768 , n21759 , n21767 );
not ( n21769 , n21768 );
and ( n21770 , n21651 , n21769 );
not ( n21771 , n21651 );
and ( n21772 , n21771 , n21768 );
or ( n21773 , n21770 , n21772 );
not ( n21774 , n21773 );
or ( n21775 , n21699 , n21774 );
not ( n21776 , n21651 );
xor ( n21777 , n21707 , n21749 );
and ( n21778 , n21777 , n21754 );
and ( n21779 , n21707 , n21749 );
or ( n21780 , n21778 , n21779 );
and ( n21781 , n19351 , n19627 );
not ( n21782 , n19655 );
not ( n21783 , n21742 );
or ( n21784 , n21782 , n21783 );
not ( n21785 , n19657 );
not ( n21786 , n19747 );
or ( n21787 , n21785 , n21786 );
nand ( n21788 , n19746 , n19687 );
nand ( n21789 , n21787 , n21788 );
nand ( n21790 , n21789 , n19690 );
nand ( n21791 , n21784 , n21790 );
xor ( n21792 , n21781 , n21791 );
not ( n21793 , n19443 );
not ( n21794 , n21729 );
or ( n21795 , n21793 , n21794 );
xor ( n21796 , n19351 , n19721 );
nand ( n21797 , n21796 , n19348 );
nand ( n21798 , n21795 , n21797 );
xor ( n21799 , n21792 , n21798 );
and ( n21800 , n21722 , n19643 );
and ( n21801 , n19585 , n19588 );
nor ( n21802 , n21800 , n21801 );
xor ( n21803 , n21715 , n21724 );
and ( n21804 , n21803 , n21732 );
and ( n21805 , n21715 , n21724 );
or ( n21806 , n21804 , n21805 );
xor ( n21807 , n21802 , n21806 );
xor ( n21808 , n21735 , n21746 );
and ( n21809 , n21808 , n21485 );
and ( n21810 , n21735 , n21746 );
or ( n21811 , n21809 , n21810 );
xor ( n21812 , n21807 , n21811 );
xor ( n21813 , n21799 , n21812 );
xor ( n21814 , n21711 , n21733 );
and ( n21815 , n21814 , n21748 );
and ( n21816 , n21711 , n21733 );
or ( n21817 , n21815 , n21816 );
xor ( n21818 , n21813 , n21817 );
or ( n21819 , n21780 , n21818 );
not ( n21820 , n21819 );
not ( n21821 , n21820 );
nand ( n21822 , n21780 , n21818 );
nand ( n21823 , n21821 , n21822 );
not ( n21824 , n21757 );
not ( n21825 , n21767 );
or ( n21826 , n21824 , n21825 );
nand ( n21827 , n21826 , n21758 );
or ( n21828 , n21823 , n21827 );
nand ( n21829 , n21827 , n21823 );
nand ( n21830 , n21828 , n21829 );
not ( n21831 , n21830 );
not ( n21832 , n21831 );
or ( n21833 , n21776 , n21832 );
not ( n21834 , n21651 );
nand ( n21835 , n21830 , n21834 );
nand ( n21836 , n21833 , n21835 );
buf ( n21837 , n21696 );
nand ( n21838 , n21836 , n21837 );
nand ( n21839 , n21775 , n21838 );
xor ( n21840 , n21649 , n21839 );
and ( n21841 , n19232 , n19235 );
xor ( n21842 , n21841 , n21673 );
and ( n21843 , n19230 , n19228 );
xnor ( n21844 , n21843 , n19227 );
xnor ( n21845 , n21842 , n21844 );
not ( n21846 , n21845 );
not ( n21847 , n21846 );
nand ( n21848 , n19233 , n19235 );
and ( n21849 , n19245 , n19236 );
xor ( n21850 , n21848 , n21849 );
buf ( n21851 , n21850 );
not ( n21852 , n21851 );
not ( n21853 , n21852 );
nor ( n21854 , n19747 , n19818 );
and ( n21855 , n20023 , n19351 );
and ( n21856 , n19572 , n19818 );
nor ( n21857 , n21855 , n21856 );
not ( n21858 , n21857 );
and ( n21859 , n21858 , n19443 );
and ( n21860 , n19348 , n19351 );
nor ( n21861 , n21859 , n21860 );
xor ( n21862 , n21854 , n21861 );
not ( n21863 , n19903 );
not ( n21864 , n21478 );
or ( n21865 , n21863 , n21864 );
nand ( n21866 , n21865 , n19657 );
and ( n21867 , n19747 , n19351 );
and ( n21868 , n19746 , n19818 );
nor ( n21869 , n21867 , n21868 );
or ( n21870 , n21869 , n19442 );
or ( n21871 , n21857 , n19824 );
nand ( n21872 , n21870 , n21871 );
xor ( n21873 , n21866 , n21872 );
nor ( n21874 , n21738 , n19818 );
and ( n21875 , n21873 , n21874 );
and ( n21876 , n21866 , n21872 );
or ( n21877 , n21875 , n21876 );
and ( n21878 , n21862 , n21877 );
and ( n21879 , n21854 , n21861 );
or ( n21880 , n21878 , n21879 );
not ( n21881 , n21880 );
not ( n21882 , n21881 );
or ( n21883 , n19443 , n19348 );
nand ( n21884 , n21883 , n19351 );
nor ( n21885 , n20023 , n19818 );
xor ( n21886 , n21884 , n21885 );
not ( n21887 , n21861 );
xor ( n21888 , n21886 , n21887 );
not ( n21889 , n21888 );
not ( n21890 , n21889 );
and ( n21891 , n21882 , n21890 );
and ( n21892 , n21881 , n21889 );
nor ( n21893 , n21891 , n21892 );
not ( n21894 , n21893 );
or ( n21895 , n19643 , n19585 );
nand ( n21896 , n21895 , n19588 );
not ( n21897 , n19690 );
or ( n21898 , n19572 , n19687 );
or ( n21899 , n20023 , n19657 );
nand ( n21900 , n21898 , n21899 );
not ( n21901 , n21900 );
or ( n21902 , n21897 , n21901 );
nand ( n21903 , n21789 , n19655 );
nand ( n21904 , n21902 , n21903 );
xor ( n21905 , n21896 , n21904 );
and ( n21906 , n19351 , n19988 );
and ( n21907 , n21905 , n21906 );
and ( n21908 , n21896 , n21904 );
or ( n21909 , n21907 , n21908 );
not ( n21910 , n19443 );
and ( n21911 , n19818 , n19774 );
not ( n21912 , n19818 );
and ( n21913 , n21912 , n21738 );
or ( n21914 , n21911 , n21913 );
not ( n21915 , n21914 );
or ( n21916 , n21910 , n21915 );
or ( n21917 , n21869 , n19824 );
nand ( n21918 , n21916 , n21917 );
and ( n21919 , n19351 , n19721 );
xor ( n21920 , n21918 , n21919 );
and ( n21921 , n21900 , n19655 );
and ( n21922 , n19690 , n19657 );
nor ( n21923 , n21921 , n21922 );
xor ( n21924 , n21920 , n21923 );
xor ( n21925 , n21909 , n21924 );
not ( n21926 , n19443 );
not ( n21927 , n21796 );
or ( n21928 , n21926 , n21927 );
not ( n21929 , n21914 );
or ( n21930 , n21929 , n19824 );
nand ( n21931 , n21928 , n21930 );
not ( n21932 , n21802 );
xor ( n21933 , n21931 , n21932 );
xor ( n21934 , n21781 , n21791 );
and ( n21935 , n21934 , n21798 );
and ( n21936 , n21781 , n21791 );
or ( n21937 , n21935 , n21936 );
and ( n21938 , n21933 , n21937 );
and ( n21939 , n21931 , n21932 );
or ( n21940 , n21938 , n21939 );
and ( n21941 , n21925 , n21940 );
and ( n21942 , n21909 , n21924 );
or ( n21943 , n21941 , n21942 );
not ( n21944 , n21923 );
xor ( n21945 , n21866 , n21872 );
xor ( n21946 , n21945 , n21874 );
xor ( n21947 , n21944 , n21946 );
xor ( n21948 , n21918 , n21919 );
and ( n21949 , n21948 , n21923 );
and ( n21950 , n21918 , n21919 );
or ( n21951 , n21949 , n21950 );
xor ( n21952 , n21947 , n21951 );
nor ( n21953 , n21943 , n21952 );
xor ( n21954 , n21944 , n21946 );
and ( n21955 , n21954 , n21951 );
and ( n21956 , n21944 , n21946 );
or ( n21957 , n21955 , n21956 );
xor ( n21958 , n21854 , n21861 );
xor ( n21959 , n21958 , n21877 );
nor ( n21960 , n21957 , n21959 );
or ( n21961 , n21953 , n21960 );
not ( n21962 , n21961 );
xor ( n21963 , n21799 , n21812 );
and ( n21964 , n21963 , n21817 );
and ( n21965 , n21799 , n21812 );
or ( n21966 , n21964 , n21965 );
xor ( n21967 , n21896 , n21904 );
xor ( n21968 , n21967 , n21906 );
xor ( n21969 , n21931 , n21932 );
xor ( n21970 , n21969 , n21937 );
xor ( n21971 , n21968 , n21970 );
xor ( n21972 , n21802 , n21806 );
and ( n21973 , n21972 , n21811 );
and ( n21974 , n21802 , n21806 );
or ( n21975 , n21973 , n21974 );
xor ( n21976 , n21971 , n21975 );
nor ( n21977 , n21966 , n21976 );
xor ( n21978 , n21968 , n21970 );
and ( n21979 , n21978 , n21975 );
and ( n21980 , n21968 , n21970 );
or ( n21981 , n21979 , n21980 );
xor ( n21982 , n21909 , n21924 );
xor ( n21983 , n21982 , n21940 );
nor ( n21984 , n21981 , n21983 );
nor ( n21985 , n21977 , n21984 );
nand ( n21986 , n21819 , n21985 );
not ( n21987 , n21986 );
not ( n21988 , n21987 );
or ( n21989 , n21766 , n21756 );
nand ( n21990 , n21989 , n21758 );
not ( n21991 , n21990 );
or ( n21992 , n21988 , n21991 );
or ( n21993 , n21822 , n21977 );
nand ( n21994 , n21966 , n21976 );
nand ( n21995 , n21993 , n21994 );
not ( n21996 , n21984 );
and ( n21997 , n21995 , n21996 );
and ( n21998 , n21981 , n21983 );
nor ( n21999 , n21997 , n21998 );
nand ( n22000 , n21992 , n21999 );
nand ( n22001 , n21962 , n22000 );
nor ( n22002 , n21756 , n21986 );
nand ( n22003 , n21761 , n22002 );
nor ( n22004 , n22003 , n21961 );
nand ( n22005 , n21454 , n22004 );
nand ( n22006 , n21943 , n21952 );
not ( n22007 , n22006 );
not ( n22008 , n21960 );
and ( n22009 , n22007 , n22008 );
and ( n22010 , n21957 , n21959 );
nor ( n22011 , n22009 , n22010 );
nand ( n22012 , n22001 , n22005 , n22011 );
not ( n22013 , n22012 );
not ( n22014 , n22013 );
or ( n22015 , n21894 , n22014 );
not ( n22016 , n21893 );
nand ( n22017 , n22016 , n22012 );
nand ( n22018 , n22015 , n22017 );
and ( n22019 , n21853 , n22018 );
not ( n22020 , n21853 );
not ( n22021 , n22018 );
and ( n22022 , n22020 , n22021 );
nor ( n22023 , n22019 , n22022 );
not ( n22024 , n22023 );
or ( n22025 , n21847 , n22024 );
nor ( n22026 , n21960 , n22010 );
not ( n22027 , n22026 );
nor ( n22028 , n22003 , n21953 );
nand ( n22029 , n21453 , n22028 );
not ( n22030 , n21953 );
nand ( n22031 , n22000 , n22030 );
nand ( n22032 , n22029 , n22031 , n22006 );
not ( n22033 , n22032 );
not ( n22034 , n22033 );
or ( n22035 , n22027 , n22034 );
not ( n22036 , n22026 );
nand ( n22037 , n22036 , n22032 );
nand ( n22038 , n22035 , n22037 );
and ( n22039 , n21853 , n22038 );
not ( n22040 , n21853 );
not ( n22041 , n22038 );
and ( n22042 , n22040 , n22041 );
nor ( n22043 , n22039 , n22042 );
and ( n22044 , n21842 , n21851 );
not ( n22045 , n21842 );
not ( n22046 , n21851 );
and ( n22047 , n22045 , n22046 );
nor ( n22048 , n22044 , n22047 );
nand ( n22049 , n21845 , n22048 );
not ( n22050 , n22049 );
buf ( n22051 , n22050 );
nand ( n22052 , n22043 , n22051 );
nand ( n22053 , n22025 , n22052 );
nand ( n22054 , n19241 , n19256 );
not ( n22055 , n21679 );
xor ( n22056 , n22054 , n22055 );
and ( n22057 , n21850 , n22056 );
not ( n22058 , n21850 );
not ( n22059 , n22056 );
and ( n22060 , n22058 , n22059 );
or ( n22061 , n22057 , n22060 );
not ( n22062 , n22061 );
not ( n22063 , n22062 );
not ( n22064 , n19241 );
not ( n22065 , n21679 );
or ( n22066 , n22064 , n22065 );
nand ( n22067 , n22066 , n19256 );
nand ( n22068 , n19240 , n19253 );
xnor ( n22069 , n22067 , n22068 );
not ( n22070 , n22069 );
not ( n22071 , n22070 );
not ( n22072 , n22003 );
not ( n22073 , n22072 );
not ( n22074 , n21454 );
or ( n22075 , n22073 , n22074 );
not ( n22076 , n22000 );
nand ( n22077 , n22075 , n22076 );
nand ( n22078 , n22030 , n22006 );
and ( n22079 , n22077 , n22078 );
not ( n22080 , n22077 );
not ( n22081 , n22078 );
and ( n22082 , n22080 , n22081 );
or ( n22083 , n22079 , n22082 );
and ( n22084 , n22071 , n22083 );
not ( n22085 , n22071 );
not ( n22086 , n22083 );
and ( n22087 , n22085 , n22086 );
nor ( n22088 , n22084 , n22087 );
not ( n22089 , n22088 );
or ( n22090 , n22063 , n22089 );
nor ( n22091 , n21998 , n21984 );
not ( n22092 , n22091 );
nor ( n22093 , n21756 , n21820 );
not ( n22094 , n22093 );
nor ( n22095 , n22094 , n21977 );
not ( n22096 , n22095 );
not ( n22097 , n21767 );
or ( n22098 , n22096 , n22097 );
or ( n22099 , n21758 , n21820 );
nand ( n22100 , n22099 , n21822 );
not ( n22101 , n21977 );
and ( n22102 , n22100 , n22101 );
not ( n22103 , n21994 );
nor ( n22104 , n22102 , n22103 );
nand ( n22105 , n22098 , n22104 );
not ( n22106 , n22105 );
not ( n22107 , n22106 );
or ( n22108 , n22092 , n22107 );
not ( n22109 , n22091 );
nand ( n22110 , n22109 , n22105 );
nand ( n22111 , n22108 , n22110 );
and ( n22112 , n22071 , n22111 );
not ( n22113 , n22071 );
not ( n22114 , n22111 );
and ( n22115 , n22113 , n22114 );
nor ( n22116 , n22112 , n22115 );
and ( n22117 , n22070 , n22059 );
and ( n22118 , n22069 , n22056 );
nor ( n22119 , n22117 , n22118 );
and ( n22120 , n22119 , n22061 );
buf ( n22121 , n22120 );
nand ( n22122 , n22116 , n22121 );
nand ( n22123 , n22090 , n22122 );
xor ( n22124 , n22053 , n22123 );
and ( n22125 , n19247 , n19251 );
not ( n22126 , n19242 );
not ( n22127 , n22126 );
not ( n22128 , n21679 );
or ( n22129 , n22127 , n22128 );
not ( n22130 , n21683 );
nand ( n22131 , n22129 , n22130 );
xor ( n22132 , n22125 , n22131 );
xor ( n22133 , n22132 , n22069 );
buf ( n22134 , n22133 );
not ( n22135 , n22134 );
not ( n22136 , n21692 );
not ( n22137 , n22136 );
nand ( n22138 , n22101 , n21994 );
not ( n22139 , n22138 );
not ( n22140 , n22139 );
not ( n22141 , n22093 );
not ( n22142 , n21767 );
or ( n22143 , n22141 , n22142 );
not ( n22144 , n22100 );
nand ( n22145 , n22143 , n22144 );
not ( n22146 , n22145 );
not ( n22147 , n22146 );
or ( n22148 , n22140 , n22147 );
nand ( n22149 , n22145 , n22138 );
nand ( n22150 , n22148 , n22149 );
and ( n22151 , n22137 , n22150 );
not ( n22152 , n22137 );
not ( n22153 , n22150 );
and ( n22154 , n22152 , n22153 );
nor ( n22155 , n22151 , n22154 );
not ( n22156 , n22155 );
or ( n22157 , n22135 , n22156 );
and ( n22158 , n22137 , n21830 );
not ( n22159 , n22137 );
and ( n22160 , n22159 , n21831 );
nor ( n22161 , n22158 , n22160 );
buf ( n22162 , n21692 );
xor ( n22163 , n22132 , n22162 );
not ( n22164 , n22163 );
nor ( n22165 , n22164 , n22133 );
buf ( n22166 , n22165 );
nand ( n22167 , n22161 , n22166 );
nand ( n22168 , n22157 , n22167 );
and ( n22169 , n22124 , n22168 );
and ( n22170 , n22053 , n22123 );
or ( n22171 , n22169 , n22170 );
xor ( n22172 , n21840 , n22171 );
not ( n22173 , n22051 );
not ( n22174 , n22023 );
or ( n22175 , n22173 , n22174 );
nand ( n22176 , n21846 , n21853 );
nand ( n22177 , n22175 , n22176 );
buf ( n22178 , n21844 );
not ( n22179 , n22178 );
not ( n22180 , n22179 );
not ( n22181 , n19296 );
nor ( n22182 , n21589 , n21568 );
nor ( n22183 , n522 , n538 );
nor ( n22184 , n521 , n537 );
nor ( n22185 , n22183 , n22184 );
and ( n22186 , n22182 , n22185 );
and ( n22187 , n21554 , n22186 );
not ( n22188 , n22187 );
or ( n22189 , n22181 , n22188 );
and ( n22190 , n21565 , n22186 );
not ( n22191 , n22185 );
not ( n22192 , n21570 );
not ( n22193 , n22192 );
not ( n22194 , n21590 );
or ( n22195 , n22193 , n22194 );
nand ( n22196 , n22195 , n21591 );
not ( n22197 , n22196 );
or ( n22198 , n22191 , n22197 );
not ( n22199 , n22184 );
nand ( n22200 , n522 , n538 );
not ( n22201 , n22200 );
and ( n22202 , n22199 , n22201 );
and ( n22203 , n521 , n537 );
nor ( n22204 , n22202 , n22203 );
nand ( n22205 , n22198 , n22204 );
nor ( n22206 , n22190 , n22205 );
nand ( n22207 , n22189 , n22206 );
not ( n22208 , n22183 );
and ( n22209 , n22182 , n22208 );
not ( n22210 , n22209 );
nor ( n22211 , n22210 , n21553 );
not ( n22212 , n22211 );
not ( n22213 , n19266 );
or ( n22214 , n22212 , n22213 );
and ( n22215 , n22209 , n21565 );
not ( n22216 , n22208 );
not ( n22217 , n22196 );
or ( n22218 , n22216 , n22217 );
nand ( n22219 , n22218 , n22200 );
nor ( n22220 , n22215 , n22219 );
nand ( n22221 , n22214 , n22220 );
nor ( n22222 , n22203 , n22184 );
xor ( n22223 , n22221 , n22222 );
xnor ( n22224 , n22207 , n22223 );
not ( n22225 , n22224 );
not ( n22226 , n22225 );
not ( n22227 , n21440 );
not ( n22228 , n21443 );
nand ( n22229 , n22227 , n22228 );
xnor ( n22230 , n21413 , n22229 );
buf ( n22231 , n22230 );
not ( n22232 , n22231 );
or ( n22233 , n22226 , n22232 );
not ( n22234 , n21402 );
and ( n22235 , n22234 , n21410 );
or ( n22236 , n21372 , n21377 );
not ( n22237 , n22236 );
not ( n22238 , n21340 );
or ( n22239 , n22237 , n22238 );
nand ( n22240 , n22239 , n21407 );
xor ( n22241 , n22235 , n22240 );
nand ( n22242 , n22224 , n22207 );
not ( n22243 , n22242 );
nand ( n22244 , n22241 , n22243 );
nand ( n22245 , n22233 , n22244 );
not ( n22246 , n22245 );
or ( n22247 , n22180 , n22246 );
not ( n22248 , n22245 );
nand ( n22249 , n22248 , n22178 );
nand ( n22250 , n22247 , n22249 );
and ( n22251 , n21554 , n22182 );
not ( n22252 , n22251 );
not ( n22253 , n19296 );
or ( n22254 , n22252 , n22253 );
and ( n22255 , n21565 , n22182 );
nor ( n22256 , n22255 , n22196 );
nand ( n22257 , n22254 , n22256 );
nand ( n22258 , n22208 , n22200 );
xnor ( n22259 , n22257 , n22258 );
and ( n22260 , n22259 , n21594 );
not ( n22261 , n22259 );
and ( n22262 , n22261 , n21593 );
nor ( n22263 , n22260 , n22262 );
not ( n22264 , n22263 );
not ( n22265 , n22264 );
not ( n22266 , n22265 );
not ( n22267 , n22266 );
buf ( n22268 , n22223 );
not ( n22269 , n22268 );
not ( n22270 , n21415 );
nand ( n22271 , n22270 , n20552 );
xnor ( n22272 , n22271 , n21608 );
buf ( n22273 , n22272 );
not ( n22274 , n22273 );
not ( n22275 , n22274 );
or ( n22276 , n22269 , n22275 );
not ( n22277 , n22268 );
nand ( n22278 , n22273 , n22277 );
nand ( n22279 , n22276 , n22278 );
not ( n22280 , n22279 );
or ( n22281 , n22267 , n22280 );
not ( n22282 , n22268 );
nand ( n22283 , n21447 , n21450 );
not ( n22284 , n22227 );
not ( n22285 , n21604 );
or ( n22286 , n22284 , n22285 );
nand ( n22287 , n22286 , n22228 );
xnor ( n22288 , n22283 , n22287 );
not ( n22289 , n22288 );
not ( n22290 , n22289 );
or ( n22291 , n22282 , n22290 );
nand ( n22292 , n22288 , n22277 );
nand ( n22293 , n22291 , n22292 );
not ( n22294 , n22223 );
not ( n22295 , n22259 );
and ( n22296 , n22294 , n22295 );
and ( n22297 , n22223 , n22259 );
nor ( n22298 , n22296 , n22297 );
and ( n22299 , n22263 , n22298 );
nand ( n22300 , n22293 , n22299 );
nand ( n22301 , n22281 , n22300 );
xor ( n22302 , n22250 , n22301 );
not ( n22303 , n21577 );
not ( n22304 , n21641 );
or ( n22305 , n22303 , n22304 );
not ( n22306 , n21414 );
nand ( n22307 , n22306 , n20554 );
not ( n22308 , n22270 );
not ( n22309 , n21608 );
or ( n22310 , n22308 , n22309 );
nand ( n22311 , n22310 , n20552 );
or ( n22312 , n22307 , n22311 );
nand ( n22313 , n22311 , n22307 );
nand ( n22314 , n22312 , n22313 );
and ( n22315 , n21595 , n22314 );
not ( n22316 , n21595 );
not ( n22317 , n22314 );
and ( n22318 , n22316 , n22317 );
nor ( n22319 , n22315 , n22318 );
nand ( n22320 , n22319 , n21646 );
nand ( n22321 , n22305 , n22320 );
and ( n22322 , n22302 , n22321 );
and ( n22323 , n22250 , n22301 );
or ( n22324 , n22322 , n22323 );
xor ( n22325 , n22177 , n22324 );
not ( n22326 , n22121 );
not ( n22327 , n22088 );
or ( n22328 , n22326 , n22327 );
not ( n22329 , n22071 );
not ( n22330 , n22041 );
or ( n22331 , n22329 , n22330 );
nand ( n22332 , n22070 , n22038 );
nand ( n22333 , n22331 , n22332 );
nand ( n22334 , n22062 , n22333 );
nand ( n22335 , n22328 , n22334 );
xor ( n22336 , n22325 , n22335 );
and ( n22337 , n22172 , n22336 );
and ( n22338 , n21840 , n22171 );
or ( n22339 , n22337 , n22338 );
or ( n22340 , n22051 , n21846 );
nand ( n22341 , n22340 , n21853 );
not ( n22342 , n22243 );
not ( n22343 , n22288 );
or ( n22344 , n22342 , n22343 );
nand ( n22345 , n22273 , n22225 );
nand ( n22346 , n22344 , n22345 );
xor ( n22347 , n22341 , n22346 );
not ( n22348 , n22266 );
not ( n22349 , n22268 );
not ( n22350 , n21637 );
or ( n22351 , n22349 , n22350 );
nand ( n22352 , n21636 , n22277 );
nand ( n22353 , n22351 , n22352 );
not ( n22354 , n22353 );
or ( n22355 , n22348 , n22354 );
not ( n22356 , n22268 );
not ( n22357 , n22317 );
or ( n22358 , n22356 , n22357 );
nand ( n22359 , n22314 , n22277 );
nand ( n22360 , n22358 , n22359 );
nand ( n22361 , n22360 , n22299 );
nand ( n22362 , n22355 , n22361 );
xor ( n22363 , n22347 , n22362 );
nand ( n22364 , n22288 , n22225 );
nand ( n22365 , n22231 , n22243 );
and ( n22366 , n22364 , n22365 );
xor ( n22367 , n22249 , n22366 );
not ( n22368 , n22266 );
not ( n22369 , n22360 );
or ( n22370 , n22368 , n22369 );
nand ( n22371 , n22279 , n22299 );
nand ( n22372 , n22370 , n22371 );
and ( n22373 , n22367 , n22372 );
and ( n22374 , n22249 , n22366 );
or ( n22375 , n22373 , n22374 );
not ( n22376 , n22366 );
not ( n22377 , n21549 );
and ( n22378 , n19319 , n21768 );
not ( n22379 , n19319 );
and ( n22380 , n22379 , n21769 );
nor ( n22381 , n22378 , n22380 );
not ( n22382 , n22381 );
or ( n22383 , n22377 , n22382 );
nand ( n22384 , n21548 , n19316 );
nand ( n22385 , n22383 , n22384 );
xor ( n22386 , n22376 , n22385 );
not ( n22387 , n21577 );
and ( n22388 , n21595 , n21456 );
not ( n22389 , n21595 );
and ( n22390 , n22389 , n21459 );
nor ( n22391 , n22388 , n22390 );
not ( n22392 , n22391 );
or ( n22393 , n22387 , n22392 );
nand ( n22394 , n21625 , n21646 );
nand ( n22395 , n22393 , n22394 );
xor ( n22396 , n22386 , n22395 );
xor ( n22397 , n22375 , n22396 );
xor ( n22398 , n22363 , n22397 );
not ( n22399 , n22134 );
and ( n22400 , n22137 , n22111 );
not ( n22401 , n22137 );
and ( n22402 , n22401 , n22114 );
nor ( n22403 , n22400 , n22402 );
not ( n22404 , n22403 );
or ( n22405 , n22399 , n22404 );
nand ( n22406 , n22155 , n22166 );
nand ( n22407 , n22405 , n22406 );
not ( n22408 , n22407 );
not ( n22409 , n22225 );
not ( n22410 , n22241 );
or ( n22411 , n22409 , n22410 );
nand ( n22412 , n22236 , n21407 );
and ( n22413 , n21340 , n22412 );
not ( n22414 , n21340 );
not ( n22415 , n22412 );
and ( n22416 , n22414 , n22415 );
or ( n22417 , n22413 , n22416 );
not ( n22418 , n22417 );
or ( n22419 , n22418 , n22242 );
nand ( n22420 , n22411 , n22419 );
not ( n22421 , n22266 );
not ( n22422 , n22293 );
or ( n22423 , n22421 , n22422 );
and ( n22424 , n22268 , n22231 );
not ( n22425 , n22268 );
not ( n22426 , n22231 );
and ( n22427 , n22425 , n22426 );
nor ( n22428 , n22424 , n22427 );
nand ( n22429 , n22428 , n22299 );
nand ( n22430 , n22423 , n22429 );
and ( n22431 , n22420 , n22430 );
not ( n22432 , n19319 );
not ( n22433 , n21620 );
or ( n22434 , n22432 , n22433 );
nand ( n22435 , n21619 , n19318 );
nand ( n22436 , n22434 , n22435 );
not ( n22437 , n22436 );
not ( n22438 , n19316 );
or ( n22439 , n22437 , n22438 );
nand ( n22440 , n21461 , n21549 );
nand ( n22441 , n22439 , n22440 );
xor ( n22442 , n22431 , n22441 );
not ( n22443 , n21837 );
not ( n22444 , n21773 );
or ( n22445 , n22443 , n22444 );
not ( n22446 , n21651 );
not ( n22447 , n21546 );
or ( n22448 , n22446 , n22447 );
nand ( n22449 , n21543 , n21834 );
nand ( n22450 , n22448 , n22449 );
nand ( n22451 , n22450 , n21698 );
nand ( n22452 , n22445 , n22451 );
and ( n22453 , n22442 , n22452 );
and ( n22454 , n22431 , n22441 );
or ( n22455 , n22453 , n22454 );
not ( n22456 , n22455 );
or ( n22457 , n22408 , n22456 );
or ( n22458 , n22455 , n22407 );
xor ( n22459 , n22249 , n22366 );
xor ( n22460 , n22459 , n22372 );
nand ( n22461 , n22458 , n22460 );
nand ( n22462 , n22457 , n22461 );
xor ( n22463 , n22398 , n22462 );
xor ( n22464 , n21551 , n21648 );
and ( n22465 , n22464 , n21839 );
and ( n22466 , n21551 , n21648 );
or ( n22467 , n22465 , n22466 );
xor ( n22468 , n22177 , n22324 );
and ( n22469 , n22468 , n22335 );
and ( n22470 , n22177 , n22324 );
or ( n22471 , n22469 , n22470 );
xor ( n22472 , n22467 , n22471 );
not ( n22473 , n22121 );
not ( n22474 , n22333 );
or ( n22475 , n22473 , n22474 );
and ( n22476 , n22071 , n22018 );
not ( n22477 , n22071 );
and ( n22478 , n22477 , n22021 );
nor ( n22479 , n22476 , n22478 );
nand ( n22480 , n22479 , n22062 );
nand ( n22481 , n22475 , n22480 );
not ( n22482 , n21698 );
not ( n22483 , n21836 );
or ( n22484 , n22482 , n22483 );
not ( n22485 , n21651 );
not ( n22486 , n22153 );
or ( n22487 , n22485 , n22486 );
nand ( n22488 , n22150 , n21834 );
nand ( n22489 , n22487 , n22488 );
nand ( n22490 , n22489 , n21837 );
nand ( n22491 , n22484 , n22490 );
xor ( n22492 , n22481 , n22491 );
not ( n22493 , n22134 );
not ( n22494 , n22137 );
not ( n22495 , n22086 );
or ( n22496 , n22494 , n22495 );
nand ( n22497 , n22083 , n22136 );
nand ( n22498 , n22496 , n22497 );
not ( n22499 , n22498 );
or ( n22500 , n22493 , n22499 );
nand ( n22501 , n22403 , n22166 );
nand ( n22502 , n22500 , n22501 );
xor ( n22503 , n22492 , n22502 );
xor ( n22504 , n22472 , n22503 );
xor ( n22505 , n22463 , n22504 );
xor ( n22506 , n22339 , n22505 );
not ( n22507 , n22455 );
xnor ( n22508 , n22407 , n22460 );
not ( n22509 , n22508 );
and ( n22510 , n22507 , n22509 );
and ( n22511 , n22455 , n22508 );
nor ( n22512 , n22510 , n22511 );
not ( n22513 , n22512 );
not ( n22514 , n22513 );
xor ( n22515 , n21840 , n22171 );
xor ( n22516 , n22515 , n22336 );
not ( n22517 , n22516 );
or ( n22518 , n22514 , n22517 );
or ( n22519 , n22516 , n22513 );
xor ( n22520 , n22250 , n22301 );
xor ( n22521 , n22520 , n22321 );
not ( n22522 , n22243 );
not ( n22523 , n21333 );
not ( n22524 , n21177 );
or ( n22525 , n22523 , n22524 );
not ( n22526 , n21337 );
nand ( n22527 , n22525 , n22526 );
not ( n22528 , n22527 );
not ( n22529 , n22528 );
nand ( n22530 , n21336 , n21339 );
not ( n22531 , n22530 );
not ( n22532 , n22531 );
or ( n22533 , n22529 , n22532 );
nand ( n22534 , n22530 , n22527 );
nand ( n22535 , n22533 , n22534 );
not ( n22536 , n22535 );
or ( n22537 , n22522 , n22536 );
nand ( n22538 , n22417 , n22225 );
nand ( n22539 , n22537 , n22538 );
not ( n22540 , n22266 );
not ( n22541 , n22428 );
or ( n22542 , n22540 , n22541 );
not ( n22543 , n22268 );
not ( n22544 , n22241 );
not ( n22545 , n22544 );
or ( n22546 , n22543 , n22545 );
nand ( n22547 , n22241 , n22277 );
nand ( n22548 , n22546 , n22547 );
nand ( n22549 , n22548 , n22299 );
nand ( n22550 , n22542 , n22549 );
and ( n22551 , n22539 , n22550 );
not ( n22552 , n21577 );
not ( n22553 , n22319 );
or ( n22554 , n22552 , n22553 );
and ( n22555 , n21595 , n22273 );
not ( n22556 , n21595 );
and ( n22557 , n22556 , n22274 );
nor ( n22558 , n22555 , n22557 );
nand ( n22559 , n22558 , n21646 );
nand ( n22560 , n22554 , n22559 );
xor ( n22561 , n22551 , n22560 );
xor ( n22562 , n22420 , n22430 );
and ( n22563 , n22561 , n22562 );
and ( n22564 , n22551 , n22560 );
or ( n22565 , n22563 , n22564 );
xor ( n22566 , n22521 , n22565 );
not ( n22567 , n19319 );
not ( n22568 , n21637 );
or ( n22569 , n22567 , n22568 );
nand ( n22570 , n21636 , n19318 );
nand ( n22571 , n22569 , n22570 );
not ( n22572 , n22571 );
not ( n22573 , n19316 );
nor ( n22574 , n22572 , n22573 );
and ( n22575 , n22436 , n21549 );
nor ( n22576 , n22574 , n22575 );
not ( n22577 , n22576 );
not ( n22578 , n22577 );
not ( n22579 , n21837 );
not ( n22580 , n22450 );
or ( n22581 , n22579 , n22580 );
and ( n22582 , n21651 , n21456 );
not ( n22583 , n21651 );
and ( n22584 , n22583 , n21459 );
nor ( n22585 , n22582 , n22584 );
nand ( n22586 , n22585 , n21698 );
nand ( n22587 , n22581 , n22586 );
not ( n22588 , n22587 );
or ( n22589 , n22578 , n22588 );
not ( n22590 , n22576 );
not ( n22591 , n22587 );
not ( n22592 , n22591 );
or ( n22593 , n22590 , n22592 );
xor ( n22594 , n22539 , n22550 );
not ( n22595 , n21646 );
not ( n22596 , n21595 );
not ( n22597 , n22289 );
or ( n22598 , n22596 , n22597 );
nand ( n22599 , n22288 , n21623 );
nand ( n22600 , n22598 , n22599 );
not ( n22601 , n22600 );
or ( n22602 , n22595 , n22601 );
nand ( n22603 , n22558 , n21577 );
nand ( n22604 , n22602 , n22603 );
xor ( n22605 , n22594 , n22604 );
not ( n22606 , n22225 );
not ( n22607 , n22535 );
or ( n22608 , n22606 , n22607 );
nand ( n22609 , n21333 , n22526 );
xnor ( n22610 , n22609 , n21177 );
buf ( n22611 , n22610 );
not ( n22612 , n22611 );
or ( n22613 , n22612 , n22242 );
nand ( n22614 , n22608 , n22613 );
nand ( n22615 , n22548 , n22266 );
not ( n22616 , n22268 );
not ( n22617 , n22418 );
or ( n22618 , n22616 , n22617 );
nand ( n22619 , n22417 , n22277 );
nand ( n22620 , n22618 , n22619 );
nand ( n22621 , n22620 , n22299 );
nand ( n22622 , n22615 , n22621 );
and ( n22623 , n22614 , n22622 );
and ( n22624 , n22605 , n22623 );
and ( n22625 , n22594 , n22604 );
or ( n22626 , n22624 , n22625 );
nand ( n22627 , n22593 , n22626 );
nand ( n22628 , n22589 , n22627 );
and ( n22629 , n22566 , n22628 );
and ( n22630 , n22521 , n22565 );
or ( n22631 , n22629 , n22630 );
nand ( n22632 , n22519 , n22631 );
nand ( n22633 , n22518 , n22632 );
xnor ( n22634 , n22506 , n22633 );
xor ( n22635 , n22631 , n22512 );
xor ( n22636 , n22516 , n22635 );
xor ( n22637 , n22431 , n22441 );
xor ( n22638 , n22637 , n22452 );
xor ( n22639 , n22053 , n22123 );
xor ( n22640 , n22639 , n22168 );
xor ( n22641 , n22638 , n22640 );
xor ( n22642 , n536 , n552 );
not ( n22643 , n22642 );
nand ( n22644 , n21844 , n22643 );
not ( n22645 , n22644 );
not ( n22646 , n22645 );
and ( n22647 , n22179 , n22021 );
not ( n22648 , n22179 );
and ( n22649 , n22648 , n22018 );
nor ( n22650 , n22647 , n22649 );
not ( n22651 , n22650 );
or ( n22652 , n22646 , n22651 );
nand ( n22653 , n22178 , n22642 );
nand ( n22654 , n22652 , n22653 );
not ( n22655 , n22134 );
not ( n22656 , n22161 );
or ( n22657 , n22655 , n22656 );
not ( n22658 , n22137 );
not ( n22659 , n21769 );
or ( n22660 , n22658 , n22659 );
nand ( n22661 , n21768 , n22136 );
nand ( n22662 , n22660 , n22661 );
nand ( n22663 , n22662 , n22166 );
nand ( n22664 , n22657 , n22663 );
nor ( n22665 , n22654 , n22664 );
not ( n22666 , n22043 );
not ( n22667 , n22666 );
not ( n22668 , n21845 );
and ( n22669 , n22667 , n22668 );
and ( n22670 , n21852 , n22086 );
not ( n22671 , n21852 );
and ( n22672 , n22671 , n22083 );
or ( n22673 , n22670 , n22672 );
not ( n22674 , n22673 );
and ( n22675 , n22674 , n22051 );
nor ( n22676 , n22669 , n22675 );
or ( n22677 , n22665 , n22676 );
nand ( n22678 , n22654 , n22664 );
nand ( n22679 , n22677 , n22678 );
and ( n22680 , n22641 , n22679 );
and ( n22681 , n22638 , n22640 );
or ( n22682 , n22680 , n22681 );
not ( n22683 , n22682 );
nand ( n22684 , n22636 , n22683 );
not ( n22685 , n22121 );
not ( n22686 , n22071 );
not ( n130240 , n22153 );
or ( n22687 , n22686 , n130240 );
nand ( n22688 , n22150 , n22070 );
nand ( n22689 , n22687 , n22688 );
not ( n22690 , n22689 );
or ( n22691 , n22685 , n22690 );
nand ( n22692 , n22116 , n22062 );
nand ( n22693 , n22691 , n22692 );
xor ( n22694 , n22551 , n22560 );
xor ( n22695 , n22694 , n22562 );
xor ( n22696 , n22693 , n22695 );
not ( n22697 , n19316 );
not ( n22698 , n19319 );
not ( n22699 , n22317 );
or ( n22700 , n22698 , n22699 );
nand ( n22701 , n22314 , n19318 );
nand ( n22702 , n22700 , n22701 );
not ( n22703 , n22702 );
or ( n22704 , n22697 , n22703 );
nand ( n22705 , n22571 , n21549 );
nand ( n22706 , n22704 , n22705 );
not ( n22707 , n21698 );
and ( n22708 , n21651 , n21619 );
not ( n22709 , n21651 );
and ( n22710 , n22709 , n21620 );
nor ( n22711 , n22708 , n22710 );
not ( n22712 , n22711 );
or ( n22713 , n22707 , n22712 );
nand ( n22714 , n22585 , n21837 );
nand ( n22715 , n22713 , n22714 );
xor ( n22716 , n22706 , n22715 );
not ( n22717 , n22225 );
not ( n22718 , n22611 );
or ( n22719 , n22717 , n22718 );
not ( n22720 , n21165 );
not ( n22721 , n22720 );
not ( n22722 , n20992 );
or ( n22723 , n22721 , n22722 );
not ( n22724 , n21172 );
nand ( n22725 , n22723 , n22724 );
not ( n22726 , n21170 );
not ( n22727 , n21169 );
or ( n22728 , n22726 , n22727 );
not ( n22729 , n21175 );
nand ( n22730 , n22728 , n22729 );
not ( n22731 , n22730 );
and ( n22732 , n22725 , n22731 );
not ( n22733 , n22725 );
and ( n22734 , n22733 , n22730 );
nor ( n22735 , n22732 , n22734 );
not ( n22736 , n22735 );
not ( n22737 , n22736 );
nand ( n22738 , n22737 , n22243 );
nand ( n22739 , n22719 , n22738 );
not ( n22740 , n22299 );
not ( n22741 , n22268 );
not ( n22742 , n22535 );
not ( n22743 , n22742 );
or ( n22744 , n22741 , n22743 );
nand ( n22745 , n22535 , n22277 );
nand ( n22746 , n22744 , n22745 );
not ( n22747 , n22746 );
or ( n22748 , n22740 , n22747 );
nand ( n22749 , n22620 , n22266 );
nand ( n22750 , n22748 , n22749 );
and ( n22751 , n22739 , n22750 );
xor ( n22752 , n22614 , n22622 );
xor ( n22753 , n22751 , n22752 );
not ( n22754 , n21577 );
not ( n22755 , n22600 );
or ( n22756 , n22754 , n22755 );
and ( n22757 , n21623 , n22426 );
not ( n22758 , n21623 );
and ( n22759 , n22758 , n22231 );
or ( n22760 , n22757 , n22759 );
not ( n22761 , n22760 );
nand ( n22762 , n22761 , n21646 );
nand ( n22763 , n22756 , n22762 );
and ( n22764 , n22753 , n22763 );
and ( n22765 , n22751 , n22752 );
or ( n22766 , n22764 , n22765 );
and ( n22767 , n22716 , n22766 );
and ( n22768 , n22706 , n22715 );
or ( n22769 , n22767 , n22768 );
and ( n22770 , n22696 , n22769 );
and ( n22771 , n22693 , n22695 );
or ( n22772 , n22770 , n22771 );
xor ( n22773 , n22521 , n22565 );
xor ( n22774 , n22773 , n22628 );
xor ( n22775 , n22772 , n22774 );
xor ( n22776 , n22638 , n22640 );
xor ( n22777 , n22776 , n22679 );
and ( n22778 , n22775 , n22777 );
and ( n22779 , n22772 , n22774 );
or ( n22780 , n22778 , n22779 );
and ( n22781 , n22684 , n22780 );
not ( n22782 , n22636 );
and ( n22783 , n22782 , n22682 );
nor ( n22784 , n22781 , n22783 );
nor ( n22785 , n22634 , n22784 );
not ( n22786 , n22785 );
nand ( n22787 , n22634 , n22784 );
nand ( n22788 , n22786 , n22787 );
xor ( n22789 , n22706 , n22715 );
xor ( n22790 , n22789 , n22766 );
not ( n22791 , n22166 );
not ( n22792 , n22136 );
not ( n22793 , n21456 );
or ( n22794 , n22792 , n22793 );
nand ( n22795 , n21459 , n22137 );
nand ( n22796 , n22794 , n22795 );
not ( n22797 , n22796 );
or ( n22798 , n22791 , n22797 );
not ( n22799 , n22136 );
not ( n22800 , n21543 );
or ( n22801 , n22799 , n22800 );
nand ( n22802 , n21546 , n22137 );
nand ( n22803 , n22801 , n22802 );
nand ( n22804 , n22803 , n22134 );
nand ( n22805 , n22798 , n22804 );
not ( n22806 , n22642 );
not ( n22807 , n22178 );
not ( n22808 , n22041 );
or ( n22809 , n22807 , n22808 );
nand ( n22810 , n22038 , n22179 );
nand ( n22811 , n22809 , n22810 );
not ( n22812 , n22811 );
or ( n22813 , n22806 , n22812 );
not ( n22814 , n22178 );
not ( n22815 , n22086 );
or ( n22816 , n22814 , n22815 );
nand ( n22817 , n22083 , n22179 );
nand ( n22818 , n22816 , n22817 );
nand ( n22819 , n22818 , n22645 );
nand ( n22820 , n22813 , n22819 );
xor ( n22821 , n22805 , n22820 );
not ( n22822 , n21853 );
not ( n22823 , n22153 );
or ( n22824 , n22822 , n22823 );
nand ( n22825 , n22150 , n21852 );
nand ( n22826 , n22824 , n22825 );
not ( n22827 , n22826 );
not ( n22828 , n22051 );
or ( n22829 , n22827 , n22828 );
and ( n22830 , n21852 , n22111 );
not ( n22831 , n21852 );
and ( n22832 , n22831 , n22114 );
nor ( n22833 , n22830 , n22832 );
or ( n22834 , n22833 , n21845 );
nand ( n22835 , n22829 , n22834 );
and ( n22836 , n22821 , n22835 );
and ( n22837 , n22805 , n22820 );
or ( n22838 , n22836 , n22837 );
xor ( n22839 , n22790 , n22838 );
xor ( n22840 , n22751 , n22752 );
xor ( n22841 , n22840 , n22763 );
and ( n22842 , n22070 , n21830 );
not ( n22843 , n22070 );
and ( n22844 , n22843 , n21831 );
nor ( n22845 , n22842 , n22844 );
or ( n22846 , n22845 , n22061 );
not ( n22847 , n22071 );
not ( n22848 , n21769 );
or ( n22849 , n22847 , n22848 );
nand ( n22850 , n21768 , n22070 );
nand ( n22851 , n22849 , n22850 );
nand ( n22852 , n22851 , n22121 );
nand ( n22853 , n22846 , n22852 );
xor ( n22854 , n22841 , n22853 );
and ( n22855 , n19318 , n22288 );
not ( n22856 , n19318 );
and ( n22857 , n22856 , n22289 );
nor ( n22858 , n22855 , n22857 );
or ( n22859 , n22858 , n22573 );
and ( n22860 , n19318 , n22273 );
not ( n22861 , n19318 );
and ( n22862 , n22861 , n22274 );
nor ( n22863 , n22860 , n22862 );
not ( n22864 , n21549 );
or ( n22865 , n22863 , n22864 );
nand ( n22866 , n22859 , n22865 );
and ( n22867 , n21834 , n22317 );
not ( n22868 , n21834 );
and ( n22869 , n22868 , n22314 );
or ( n22870 , n22867 , n22869 );
not ( n22871 , n21698 );
or ( n22872 , n22870 , n22871 );
and ( n22873 , n21834 , n21637 );
not ( n22874 , n21834 );
and ( n22875 , n22874 , n21636 );
or ( n22876 , n22873 , n22875 );
not ( n22877 , n21837 );
or ( n22878 , n22876 , n22877 );
nand ( n22879 , n22872 , n22878 );
xor ( n22880 , n22866 , n22879 );
not ( n22881 , n22225 );
nand ( n22882 , n22720 , n22724 );
xnor ( n22883 , n20992 , n22882 );
buf ( n22884 , n22883 );
not ( n22885 , n22884 );
or ( n22886 , n22881 , n22885 );
buf ( n22887 , n20988 );
nand ( n22888 , n20751 , n20991 );
or ( n22889 , n22887 , n22888 );
nand ( n22890 , n22888 , n22887 );
nand ( n22891 , n22889 , n22890 );
not ( n22892 , n22891 );
or ( n22893 , n22892 , n22242 );
nand ( n22894 , n22886 , n22893 );
not ( n22895 , n22264 );
not ( n22896 , n22268 );
not ( n22897 , n22612 );
or ( n22898 , n22896 , n22897 );
nand ( n22899 , n22611 , n22277 );
nand ( n22900 , n22898 , n22899 );
not ( n22901 , n22900 );
or ( n22902 , n22895 , n22901 );
not ( n22903 , n22268 );
not ( n22904 , n22736 );
or ( n22905 , n22903 , n22904 );
nand ( n22906 , n22737 , n22277 );
nand ( n22907 , n22905 , n22906 );
nand ( n22908 , n22907 , n22299 );
nand ( n22909 , n22902 , n22908 );
and ( n22910 , n22894 , n22909 );
not ( n22911 , n21595 );
not ( n22912 , n22418 );
or ( n22913 , n22911 , n22912 );
nand ( n22914 , n22417 , n21623 );
nand ( n22915 , n22913 , n22914 );
not ( n22916 , n22915 );
not ( n22917 , n21646 );
or ( n22918 , n22916 , n22917 );
and ( n22919 , n21623 , n22544 );
not ( n22920 , n21623 );
and ( n22921 , n22920 , n22241 );
or ( n22922 , n22919 , n22921 );
or ( n22923 , n22922 , n21576 );
nand ( n22924 , n22918 , n22923 );
xor ( n22925 , n22910 , n22924 );
not ( n22926 , n22884 );
not ( n22927 , n22926 );
not ( n22928 , n22242 );
and ( n22929 , n22927 , n22928 );
and ( n22930 , n22737 , n22225 );
nor ( n22931 , n22929 , n22930 );
and ( n22932 , n22746 , n22266 );
not ( n22933 , n22900 );
not ( n22934 , n22299 );
nor ( n22935 , n22933 , n22934 );
nor ( n22936 , n22932 , n22935 );
xor ( n22937 , n22931 , n22936 );
and ( n22938 , n22925 , n22937 );
and ( n22939 , n22910 , n22924 );
or ( n22940 , n22938 , n22939 );
and ( n22941 , n22880 , n22940 );
and ( n22942 , n22866 , n22879 );
or ( n22943 , n22941 , n22942 );
and ( n22944 , n22854 , n22943 );
and ( n22945 , n22841 , n22853 );
or ( n22946 , n22944 , n22945 );
xor ( n22947 , n22839 , n22946 );
xor ( n22948 , n22805 , n22820 );
xor ( n22949 , n22948 , n22835 );
xor ( n22950 , n22841 , n22853 );
xor ( n22951 , n22950 , n22943 );
xor ( n22952 , n22949 , n22951 );
xor ( n22953 , n22866 , n22879 );
xor ( n22954 , n22953 , n22940 );
xor ( n22955 , n22910 , n22924 );
xor ( n22956 , n22955 , n22937 );
not ( n22957 , n22121 );
not ( n22958 , n22071 );
not ( n22959 , n21459 );
or ( n22960 , n22958 , n22959 );
nand ( n22961 , n21456 , n22070 );
nand ( n22962 , n22960 , n22961 );
not ( n22963 , n22962 );
or ( n22964 , n22957 , n22963 );
not ( n22965 , n22071 );
not ( n22966 , n21546 );
or ( n22967 , n22965 , n22966 );
nand ( n22968 , n21543 , n22070 );
nand ( n22969 , n22967 , n22968 );
nand ( n22970 , n22969 , n22062 );
nand ( n22971 , n22964 , n22970 );
xor ( n22972 , n22956 , n22971 );
not ( n22973 , n22134 );
buf ( n22974 , n21619 );
and ( n22975 , n22137 , n22974 );
not ( n22976 , n22137 );
and ( n22977 , n22976 , n21620 );
nor ( n22978 , n22975 , n22977 );
not ( n22979 , n22978 );
or ( n22980 , n22973 , n22979 );
not ( n22981 , n22137 );
not ( n22982 , n21637 );
or ( n22983 , n22981 , n22982 );
nand ( n22984 , n21636 , n22136 );
nand ( n22985 , n22983 , n22984 );
nand ( n22986 , n22985 , n22166 );
nand ( n22987 , n22980 , n22986 );
and ( n22988 , n22972 , n22987 );
and ( n22989 , n22956 , n22971 );
or ( n22990 , n22988 , n22989 );
xor ( n22991 , n22954 , n22990 );
not ( n22992 , n21549 );
not ( n22993 , n19319 );
not ( n22994 , n22426 );
or ( n22995 , n22993 , n22994 );
nand ( n22996 , n22231 , n19318 );
nand ( n22997 , n22995 , n22996 );
not ( n22998 , n22997 );
or ( n22999 , n22992 , n22998 );
and ( n23000 , n19319 , n22241 );
not ( n23001 , n19319 );
and ( n23002 , n23001 , n22544 );
nor ( n23003 , n23000 , n23002 );
nand ( n23004 , n23003 , n19316 );
nand ( n23005 , n22999 , n23004 );
not ( n23006 , n21698 );
and ( n23007 , n21651 , n22288 );
not ( n23008 , n21651 );
and ( n23009 , n23008 , n22289 );
nor ( n23010 , n23007 , n23009 );
not ( n23011 , n23010 );
or ( n23012 , n23006 , n23011 );
and ( n23013 , n21651 , n22273 );
not ( n23014 , n21651 );
and ( n23015 , n23014 , n22274 );
nor ( n23016 , n23013 , n23015 );
nand ( n23017 , n23016 , n21837 );
nand ( n23018 , n23012 , n23017 );
xor ( n23019 , n23005 , n23018 );
not ( n23020 , n22264 );
and ( n23021 , n22268 , n22884 );
not ( n23022 , n22268 );
and ( n23023 , n23022 , n22926 );
nor ( n23024 , n23021 , n23023 );
not ( n23025 , n23024 );
or ( n23026 , n23020 , n23025 );
not ( n23027 , n22892 );
and ( n23028 , n22277 , n23027 );
not ( n23029 , n22277 );
and ( n23030 , n23029 , n22892 );
nor ( n23031 , n23028 , n23030 );
not ( n23032 , n23031 );
nand ( n23033 , n23032 , n22299 );
nand ( n23034 , n23026 , n23033 );
not ( n23035 , n23034 );
not ( n23036 , n20975 );
not ( n23037 , n23036 );
not ( n23038 , n20984 );
nand ( n23039 , n23038 , n20982 );
not ( n23040 , n23039 );
not ( n23041 , n23040 );
or ( n23042 , n23037 , n23041 );
nand ( n23043 , n23039 , n20975 );
nand ( n23044 , n23042 , n23043 );
not ( n23045 , n23044 );
not ( n23046 , n23045 );
and ( n23047 , n23046 , n22243 );
nand ( n23048 , n20806 , n20987 );
not ( n23049 , n20982 );
not ( n23050 , n20975 );
or ( n23051 , n23049 , n23050 );
nand ( n23052 , n23051 , n23038 );
or ( n23053 , n23048 , n23052 );
nand ( n23054 , n23052 , n23048 );
nand ( n23055 , n23053 , n23054 );
not ( n23056 , n23055 );
not ( n23057 , n23056 );
and ( n23058 , n23057 , n22225 );
nor ( n23059 , n23047 , n23058 );
nor ( n23060 , n23035 , n23059 );
not ( n23061 , n21577 );
and ( n23062 , n21595 , n22535 );
not ( n23063 , n21595 );
and ( n23064 , n23063 , n22742 );
nor ( n23065 , n23062 , n23064 );
not ( n23066 , n23065 );
or ( n23067 , n23061 , n23066 );
and ( n23068 , n21595 , n22611 );
not ( n23069 , n21595 );
and ( n23070 , n23069 , n22612 );
nor ( n23071 , n23068 , n23070 );
nand ( n23072 , n23071 , n21646 );
nand ( n23073 , n23067 , n23072 );
xor ( n23074 , n23060 , n23073 );
not ( n23075 , n22225 );
not ( n23076 , n23027 );
or ( n23077 , n23075 , n23076 );
or ( n23078 , n23056 , n22242 );
nand ( n23079 , n23077 , n23078 );
not ( n23080 , n22264 );
not ( n23081 , n22907 );
or ( n23082 , n23080 , n23081 );
nand ( n23083 , n23024 , n22299 );
nand ( n23084 , n23082 , n23083 );
xor ( n23085 , n23079 , n23084 );
and ( n23086 , n23074 , n23085 );
and ( n23087 , n23060 , n23073 );
or ( n23088 , n23086 , n23087 );
and ( n23089 , n23019 , n23088 );
and ( n23090 , n23005 , n23018 );
or ( n23091 , n23089 , n23090 );
not ( n23092 , n21646 );
not ( n23093 , n23065 );
or ( n23094 , n23092 , n23093 );
nand ( n23095 , n22915 , n21577 );
nand ( n23096 , n23094 , n23095 );
and ( n23097 , n23079 , n23084 );
xor ( n23098 , n23096 , n23097 );
xor ( n23099 , n22894 , n22909 );
and ( n23100 , n23098 , n23099 );
and ( n23101 , n23096 , n23097 );
or ( n23102 , n23100 , n23101 );
not ( n23103 , n21549 );
not ( n23104 , n22858 );
not ( n23105 , n23104 );
or ( n23106 , n23103 , n23105 );
nand ( n23107 , n22997 , n19316 );
nand ( n23108 , n23106 , n23107 );
xor ( n23109 , n23102 , n23108 );
not ( n23110 , n21698 );
not ( n23111 , n23016 );
or ( n23112 , n23110 , n23111 );
not ( n23113 , n22870 );
nand ( n23114 , n23113 , n21837 );
nand ( n23115 , n23112 , n23114 );
xor ( n23116 , n23109 , n23115 );
xor ( n23117 , n23091 , n23116 );
not ( n23118 , n22051 );
not ( n23119 , n21853 );
not ( n23120 , n21769 );
or ( n23121 , n23119 , n23120 );
nand ( n23122 , n21768 , n21852 );
nand ( n23123 , n23121 , n23122 );
not ( n23124 , n23123 );
or ( n23125 , n23118 , n23124 );
not ( n23126 , n21853 );
not ( n23127 , n21831 );
or ( n23128 , n23126 , n23127 );
nand ( n23129 , n21830 , n21852 );
nand ( n23130 , n23128 , n23129 );
nand ( n23131 , n23130 , n21846 );
nand ( n23132 , n23125 , n23131 );
and ( n23133 , n23117 , n23132 );
and ( n23134 , n23091 , n23116 );
or ( n23135 , n23133 , n23134 );
and ( n23136 , n22991 , n23135 );
and ( n23137 , n22954 , n22990 );
or ( n23138 , n23136 , n23137 );
and ( n23139 , n22952 , n23138 );
and ( n23140 , n22949 , n22951 );
or ( n23141 , n23139 , n23140 );
xor ( n23142 , n22947 , n23141 );
not ( n23143 , n22134 );
not ( n23144 , n22662 );
or ( n23145 , n23143 , n23144 );
nand ( n23146 , n22803 , n22166 );
nand ( n23147 , n23145 , n23146 );
not ( n23148 , n22811 );
not ( n23149 , n22645 );
or ( n23150 , n23148 , n23149 );
not ( n23151 , n22650 );
or ( n23152 , n23151 , n22643 );
nand ( n23153 , n23150 , n23152 );
xor ( n23154 , n23147 , n23153 );
not ( n23155 , n22051 );
or ( n23156 , n22833 , n23155 );
or ( n23157 , n22673 , n21845 );
nand ( n23158 , n23156 , n23157 );
xor ( n23159 , n23154 , n23158 );
xor ( n23160 , n22594 , n22604 );
xor ( n23161 , n23160 , n22623 );
not ( n23162 , n22121 );
not ( n23163 , n22845 );
not ( n23164 , n23163 );
or ( n23165 , n23162 , n23164 );
nand ( n23166 , n22689 , n22062 );
nand ( n23167 , n23165 , n23166 );
xor ( n23168 , n23161 , n23167 );
nor ( n23169 , n22936 , n22931 );
not ( n23170 , n21646 );
or ( n23171 , n22922 , n23170 );
not ( n23172 , n21577 );
or ( n23173 , n22760 , n23172 );
nand ( n23174 , n23171 , n23173 );
xor ( n23175 , n23169 , n23174 );
xor ( n23176 , n22739 , n22750 );
and ( n23177 , n23175 , n23176 );
and ( n23178 , n23169 , n23174 );
or ( n23179 , n23177 , n23178 );
not ( n23180 , n22702 );
or ( n23181 , n23180 , n22864 );
not ( n23182 , n22863 );
nand ( n23183 , n23182 , n19316 );
nand ( n23184 , n23181 , n23183 );
xor ( n23185 , n23179 , n23184 );
not ( n23186 , n21698 );
not ( n23187 , n22876 );
not ( n23188 , n23187 );
or ( n23189 , n23186 , n23188 );
nand ( n23190 , n22711 , n21837 );
nand ( n23191 , n23189 , n23190 );
and ( n23192 , n23185 , n23191 );
and ( n23193 , n23179 , n23184 );
or ( n23194 , n23192 , n23193 );
xor ( n23195 , n23168 , n23194 );
xor ( n23196 , n23159 , n23195 );
xor ( n23197 , n23179 , n23184 );
xor ( n23198 , n23197 , n23191 );
not ( n23199 , n23198 );
not ( n23200 , n21846 );
not ( n23201 , n22826 );
or ( n23202 , n23200 , n23201 );
nand ( n23203 , n23130 , n22051 );
nand ( n23204 , n23202 , n23203 );
not ( n23205 , n22645 );
and ( n23206 , n22178 , n22111 );
not ( n23207 , n22178 );
and ( n23208 , n23207 , n22114 );
nor ( n23209 , n23206 , n23208 );
not ( n23210 , n23209 );
or ( n23211 , n23205 , n23210 );
nand ( n23212 , n22818 , n22642 );
nand ( n23213 , n23211 , n23212 );
xor ( n23214 , n23204 , n23213 );
xor ( n23215 , n23102 , n23108 );
and ( n23216 , n23215 , n23115 );
and ( n23217 , n23102 , n23108 );
or ( n23218 , n23216 , n23217 );
and ( n23219 , n23214 , n23218 );
and ( n23220 , n23204 , n23213 );
or ( n23221 , n23219 , n23220 );
not ( n23222 , n23221 );
or ( n23223 , n23199 , n23222 );
or ( n23224 , n23221 , n23198 );
xor ( n23225 , n23169 , n23174 );
xor ( n23226 , n23225 , n23176 );
not ( n23227 , n22166 );
not ( n23228 , n22978 );
or ( n23229 , n23227 , n23228 );
nand ( n23230 , n22796 , n22134 );
nand ( n23231 , n23229 , n23230 );
xor ( n23232 , n23226 , n23231 );
not ( n23233 , n22062 );
not ( n23234 , n22851 );
or ( n23235 , n23233 , n23234 );
nand ( n23236 , n22969 , n22121 );
nand ( n23237 , n23235 , n23236 );
and ( n23238 , n23232 , n23237 );
and ( n23239 , n23226 , n23231 );
or ( n23240 , n23238 , n23239 );
nand ( n23241 , n23224 , n23240 );
nand ( n23242 , n23223 , n23241 );
xor ( n23243 , n23196 , n23242 );
xnor ( n23244 , n23142 , n23243 );
xor ( n23245 , n22949 , n22951 );
xor ( n23246 , n23245 , n23138 );
xor ( n23247 , n23198 , n23240 );
xnor ( n23248 , n23247 , n23221 );
not ( n23249 , n23248 );
or ( n23250 , n23246 , n23249 );
xor ( n23251 , n23226 , n23231 );
xor ( n23252 , n23251 , n23237 );
xor ( n23253 , n23204 , n23213 );
xor ( n23254 , n23253 , n23218 );
xor ( n23255 , n23252 , n23254 );
not ( n23256 , n22645 );
and ( n23257 , n22178 , n22150 );
not ( n23258 , n22178 );
and ( n23259 , n23258 , n22153 );
nor ( n23260 , n23257 , n23259 );
not ( n23261 , n23260 );
or ( n23262 , n23256 , n23261 );
nand ( n23263 , n23209 , n22642 );
nand ( n23264 , n23262 , n23263 );
xor ( n23265 , n23096 , n23097 );
xor ( n23266 , n23265 , n23099 );
not ( n23267 , n22166 );
and ( n23268 , n22137 , n22314 );
not ( n23269 , n22137 );
and ( n23270 , n23269 , n22317 );
nor ( n23271 , n23268 , n23270 );
not ( n23272 , n23271 );
or ( n23273 , n23267 , n23272 );
nand ( n23274 , n22985 , n22134 );
nand ( n23275 , n23273 , n23274 );
xor ( n23276 , n23266 , n23275 );
xor ( n23277 , n23005 , n23018 );
xor ( n23278 , n23277 , n23088 );
and ( n23279 , n23276 , n23278 );
and ( n23280 , n23266 , n23275 );
or ( n23281 , n23279 , n23280 );
xor ( n23282 , n23264 , n23281 );
not ( n23283 , n23059 );
not ( n23284 , n23034 );
or ( n23285 , n23283 , n23284 );
or ( n23286 , n23034 , n23059 );
nand ( n23287 , n23285 , n23286 );
not ( n23288 , n21577 );
not ( n23289 , n23071 );
or ( n23290 , n23288 , n23289 );
and ( n23291 , n21595 , n22737 );
not ( n23292 , n21595 );
and ( n23293 , n23292 , n22736 );
nor ( n23294 , n23291 , n23293 );
not ( n23295 , n23294 );
or ( n23296 , n23295 , n23170 );
nand ( n23297 , n23290 , n23296 );
and ( n23298 , n23287 , n23297 );
not ( n23299 , n21549 );
not ( n23300 , n23003 );
or ( n23301 , n23299 , n23300 );
and ( n23302 , n19319 , n22417 );
not ( n23303 , n19319 );
and ( n23304 , n23303 , n22418 );
nor ( n23305 , n23302 , n23304 );
nand ( n23306 , n23305 , n19316 );
nand ( n23307 , n23301 , n23306 );
xor ( n23308 , n23298 , n23307 );
xor ( n23309 , n23060 , n23073 );
xor ( n23310 , n23309 , n23085 );
and ( n23311 , n23308 , n23310 );
and ( n23312 , n23298 , n23307 );
or ( n23313 , n23311 , n23312 );
not ( n23314 , n22062 );
not ( n23315 , n22962 );
or ( n23316 , n23314 , n23315 );
not ( n23317 , n22071 );
not ( n23318 , n21620 );
or ( n23319 , n23317 , n23318 );
nand ( n23320 , n22974 , n22070 );
nand ( n23321 , n23319 , n23320 );
nand ( n23322 , n23321 , n22121 );
nand ( n23323 , n23316 , n23322 );
xor ( n23324 , n23313 , n23323 );
not ( n23325 , n21846 );
not ( n23326 , n23123 );
or ( n23327 , n23325 , n23326 );
not ( n23328 , n21851 );
not ( n23329 , n21546 );
or ( n23330 , n23328 , n23329 );
nand ( n23331 , n21543 , n21852 );
nand ( n23332 , n23330 , n23331 );
nand ( n23333 , n23332 , n22051 );
nand ( n23334 , n23327 , n23333 );
and ( n23335 , n23324 , n23334 );
and ( n23336 , n23313 , n23323 );
or ( n23337 , n23335 , n23336 );
and ( n23338 , n23282 , n23337 );
and ( n23339 , n23264 , n23281 );
or ( n23340 , n23338 , n23339 );
and ( n23341 , n23255 , n23340 );
and ( n23342 , n23252 , n23254 );
or ( n23343 , n23341 , n23342 );
nand ( n23344 , n23250 , n23343 );
nand ( n23345 , n23246 , n23249 );
and ( n23346 , n23344 , n23345 );
nand ( n23347 , n23244 , n23346 );
xor ( n23348 , n23343 , n23248 );
xor ( n23349 , n23348 , n23246 );
xor ( n23350 , n23252 , n23254 );
xor ( n23351 , n23350 , n23340 );
xor ( n23352 , n22954 , n22990 );
xor ( n23353 , n23352 , n23135 );
or ( n23354 , n23351 , n23353 );
xor ( n23355 , n22956 , n22971 );
xor ( n23356 , n23355 , n22987 );
xor ( n23357 , n23091 , n23116 );
xor ( n23358 , n23357 , n23132 );
xor ( n23359 , n23356 , n23358 );
not ( n23360 , n21837 );
not ( n23361 , n23010 );
or ( n23362 , n23360 , n23361 );
not ( n23363 , n21651 );
not ( n23364 , n22426 );
or ( n23365 , n23363 , n23364 );
nand ( n23366 , n22231 , n21834 );
nand ( n23367 , n23365 , n23366 );
nand ( n23368 , n23367 , n21698 );
nand ( n23369 , n23362 , n23368 );
not ( n23370 , n23369 );
not ( n23371 , n22134 );
not ( n23372 , n23271 );
or ( n23373 , n23371 , n23372 );
and ( n23374 , n22137 , n22273 );
not ( n23375 , n22137 );
and ( n23376 , n23375 , n22274 );
nor ( n23377 , n23374 , n23376 );
nand ( n23378 , n23377 , n22166 );
nand ( n23379 , n23373 , n23378 );
not ( n23380 , n23379 );
or ( n23381 , n23370 , n23380 );
or ( n23382 , n23369 , n23379 );
not ( n23383 , n19316 );
and ( n23384 , n19319 , n22535 );
not ( n23385 , n19319 );
and ( n23386 , n23385 , n22742 );
nor ( n23387 , n23384 , n23386 );
not ( n23388 , n23387 );
or ( n23389 , n23383 , n23388 );
nand ( n23390 , n23305 , n21549 );
nand ( n23391 , n23389 , n23390 );
and ( n23392 , n20871 , n20974 );
buf ( n23393 , n20971 );
xor ( n23394 , n23392 , n23393 );
not ( n23395 , n23394 );
or ( n23396 , n23395 , n22242 );
or ( n23397 , n23045 , n22224 );
nand ( n23398 , n23396 , n23397 );
and ( n23399 , n22277 , n23057 );
not ( n23400 , n22277 );
and ( n23401 , n23400 , n23056 );
nor ( n23402 , n23399 , n23401 );
or ( n23403 , n23402 , n22934 );
or ( n23404 , n23031 , n22265 );
nand ( n23405 , n23403 , n23404 );
xor ( n23406 , n23398 , n23405 );
not ( n23407 , n21646 );
not ( n23408 , n21595 );
not ( n23409 , n22926 );
or ( n23410 , n23408 , n23409 );
nand ( n23411 , n22884 , n21623 );
nand ( n23412 , n23410 , n23411 );
not ( n23413 , n23412 );
or ( n23414 , n23407 , n23413 );
nand ( n23415 , n23294 , n21577 );
nand ( n23416 , n23414 , n23415 );
and ( n23417 , n23406 , n23416 );
and ( n23418 , n23398 , n23405 );
or ( n23419 , n23417 , n23418 );
xor ( n23420 , n23391 , n23419 );
not ( n23421 , n21698 );
and ( n23422 , n21651 , n22241 );
not ( n23423 , n21651 );
and ( n23424 , n23423 , n22544 );
nor ( n23425 , n23422 , n23424 );
not ( n23426 , n23425 );
or ( n23427 , n23421 , n23426 );
nand ( n23428 , n23367 , n21837 );
nand ( n23429 , n23427 , n23428 );
and ( n23430 , n23420 , n23429 );
and ( n23431 , n23391 , n23419 );
or ( n23432 , n23430 , n23431 );
nand ( n23433 , n23382 , n23432 );
nand ( n23434 , n23381 , n23433 );
not ( n23435 , n23434 );
not ( n23436 , n22642 );
not ( n23437 , n23260 );
or ( n23438 , n23436 , n23437 );
and ( n23439 , n22178 , n21830 );
not ( n23440 , n22178 );
and ( n23441 , n23440 , n21831 );
nor ( n23442 , n23439 , n23441 );
nand ( n23443 , n23442 , n22645 );
nand ( n23444 , n23438 , n23443 );
not ( n23445 , n23444 );
or ( n23446 , n23435 , n23445 );
not ( n23447 , n23434 );
not ( n23448 , n23447 );
not ( n23449 , n23444 );
not ( n23450 , n23449 );
or ( n23451 , n23448 , n23450 );
not ( n23452 , n22051 );
not ( n23453 , n21853 );
not ( n23454 , n21459 );
or ( n23455 , n23453 , n23454 );
nand ( n23456 , n21456 , n21852 );
nand ( n23457 , n23455 , n23456 );
not ( n23458 , n23457 );
or ( n23459 , n23452 , n23458 );
nand ( n23460 , n23332 , n21846 );
nand ( n23461 , n23459 , n23460 );
xor ( n23462 , n23298 , n23307 );
xor ( n23463 , n23462 , n23310 );
xor ( n23464 , n23461 , n23463 );
not ( n23465 , n22062 );
not ( n23466 , n23321 );
or ( n23467 , n23465 , n23466 );
and ( n23468 , n22071 , n21636 );
not ( n23469 , n22071 );
and ( n23470 , n23469 , n21637 );
nor ( n23471 , n23468 , n23470 );
nand ( n23472 , n23471 , n22121 );
nand ( n23473 , n23467 , n23472 );
and ( n23474 , n23464 , n23473 );
and ( n23475 , n23461 , n23463 );
or ( n23476 , n23474 , n23475 );
nand ( n23477 , n23451 , n23476 );
nand ( n23478 , n23446 , n23477 );
and ( n23479 , n23359 , n23478 );
and ( n23480 , n23356 , n23358 );
or ( n23481 , n23479 , n23480 );
and ( n23482 , n23354 , n23481 );
and ( n23483 , n23353 , n23351 );
nor ( n23484 , n23482 , n23483 );
nand ( n23485 , n23349 , n23484 );
and ( n23486 , n23347 , n23485 );
not ( n23487 , n23486 );
xor ( n23488 , n23353 , n23351 );
xor ( n23489 , n23488 , n23481 );
xor ( n23490 , n23356 , n23358 );
xor ( n23491 , n23490 , n23478 );
xor ( n23492 , n23264 , n23281 );
xor ( n23493 , n23492 , n23337 );
or ( n23494 , n23491 , n23493 );
xor ( n23495 , n23266 , n23275 );
xor ( n23496 , n23495 , n23278 );
xor ( n23497 , n23313 , n23323 );
xor ( n23498 , n23497 , n23334 );
xor ( n23499 , n23496 , n23498 );
xor ( n23500 , n23369 , n23432 );
xnor ( n23501 , n23500 , n23379 );
not ( n23502 , n23501 );
not ( n23503 , n22642 );
not ( n23504 , n23442 );
or ( n23505 , n23503 , n23504 );
not ( n23506 , n22178 );
not ( n23507 , n21769 );
or ( n23508 , n23506 , n23507 );
nand ( n23509 , n21768 , n22179 );
nand ( n23510 , n23508 , n23509 );
nand ( n23511 , n23510 , n22645 );
nand ( n23512 , n23505 , n23511 );
not ( n23513 , n23512 );
not ( n23514 , n23513 );
or ( n23515 , n23502 , n23514 );
xor ( n23516 , n23297 , n23287 );
not ( n23517 , n22166 );
not ( n23518 , n22137 );
not ( n23519 , n22289 );
or ( n23520 , n23518 , n23519 );
nand ( n23521 , n22288 , n22136 );
nand ( n23522 , n23520 , n23521 );
not ( n23523 , n23522 );
or ( n23524 , n23517 , n23523 );
nand ( n23525 , n23377 , n22134 );
nand ( n23526 , n23524 , n23525 );
xor ( n23527 , n23516 , n23526 );
not ( n23528 , n22225 );
not ( n23529 , n23394 );
or ( n23530 , n23528 , n23529 );
nand ( n23531 , n20966 , n20970 );
not ( n23532 , n20956 );
and ( n23533 , n23531 , n23532 );
not ( n23534 , n23531 );
and ( n23535 , n23534 , n20956 );
nor ( n23536 , n23533 , n23535 );
not ( n23537 , n23536 );
or ( n23538 , n23537 , n22242 );
nand ( n23539 , n23530 , n23538 );
not ( n23540 , n22264 );
not ( n23541 , n23402 );
not ( n23542 , n23541 );
or ( n23543 , n23540 , n23542 );
and ( n23544 , n23046 , n22277 );
and ( n23545 , n23045 , n22268 );
nor ( n23546 , n23544 , n23545 );
or ( n23547 , n23546 , n22934 );
nand ( n23548 , n23543 , n23547 );
xor ( n23549 , n23539 , n23548 );
not ( n23550 , n21577 );
not ( n23551 , n23412 );
or ( n23552 , n23550 , n23551 );
not ( n23553 , n21595 );
not ( n23554 , n22892 );
or ( n23555 , n23553 , n23554 );
nand ( n23556 , n23027 , n21623 );
nand ( n23557 , n23555 , n23556 );
nand ( n23558 , n23557 , n21646 );
nand ( n23559 , n23552 , n23558 );
and ( n23560 , n23549 , n23559 );
and ( n23561 , n23539 , n23548 );
or ( n23562 , n23560 , n23561 );
not ( n23563 , n21549 );
not ( n23564 , n23387 );
or ( n23565 , n23563 , n23564 );
and ( n23566 , n19319 , n22611 );
not ( n23567 , n19319 );
and ( n23568 , n23567 , n22612 );
nor ( n23569 , n23566 , n23568 );
nand ( n23570 , n23569 , n19316 );
nand ( n23571 , n23565 , n23570 );
xor ( n23572 , n23562 , n23571 );
xor ( n23573 , n23398 , n23405 );
xor ( n23574 , n23573 , n23416 );
and ( n23575 , n23572 , n23574 );
and ( n23576 , n23562 , n23571 );
or ( n23577 , n23575 , n23576 );
and ( n23578 , n23527 , n23577 );
and ( n23579 , n23516 , n23526 );
or ( n23580 , n23578 , n23579 );
nand ( n23581 , n23515 , n23580 );
not ( n23582 , n23501 );
nand ( n23583 , n23582 , n23512 );
nand ( n23584 , n23581 , n23583 );
and ( n23585 , n23499 , n23584 );
and ( n23586 , n23496 , n23498 );
or ( n23587 , n23585 , n23586 );
nand ( n23588 , n23494 , n23587 );
nand ( n23589 , n23491 , n23493 );
nand ( n23590 , n23588 , n23589 );
or ( n23591 , n23489 , n23590 );
xor ( n23592 , n23493 , n23587 );
xnor ( n23593 , n23592 , n23491 );
not ( n23594 , n23434 );
not ( n23595 , n23449 );
or ( n23596 , n23594 , n23595 );
nand ( n23597 , n23447 , n23444 );
nand ( n23598 , n23596 , n23597 );
xnor ( n23599 , n23598 , n23476 );
not ( n23600 , n23599 );
xor ( n23601 , n23496 , n23498 );
xor ( n23602 , n23601 , n23584 );
not ( n23603 , n23602 );
not ( n23604 , n23603 );
or ( n23605 , n23600 , n23604 );
not ( n23606 , n22121 );
and ( n23607 , n22071 , n22314 );
not ( n23608 , n22071 );
and ( n23609 , n23608 , n22317 );
nor ( n23610 , n23607 , n23609 );
not ( n23611 , n23610 );
or ( n23612 , n23606 , n23611 );
nand ( n23613 , n23471 , n22062 );
nand ( n23614 , n23612 , n23613 );
xor ( n23615 , n23391 , n23419 );
xor ( n23616 , n23615 , n23429 );
xor ( n23617 , n23614 , n23616 );
not ( n23618 , n22051 );
and ( n23619 , n21851 , n22974 );
not ( n23620 , n21851 );
and ( n23621 , n23620 , n21620 );
nor ( n23622 , n23619 , n23621 );
not ( n23623 , n23622 );
or ( n23624 , n23618 , n23623 );
nand ( n23625 , n23457 , n21846 );
nand ( n23626 , n23624 , n23625 );
and ( n23627 , n23617 , n23626 );
and ( n23628 , n23614 , n23616 );
or ( n23629 , n23627 , n23628 );
xor ( n23630 , n23461 , n23463 );
xor ( n23631 , n23630 , n23473 );
xor ( n23632 , n23629 , n23631 );
and ( n23633 , n21651 , n22417 );
not ( n23634 , n21651 );
and ( n23635 , n23634 , n22418 );
nor ( n23636 , n23633 , n23635 );
not ( n23637 , n23636 );
not ( n23638 , n21698 );
or ( n23639 , n23637 , n23638 );
not ( n23640 , n23425 );
or ( n23641 , n23640 , n22877 );
nand ( n23642 , n23639 , n23641 );
xor ( n23643 , n20882 , n20914 );
xor ( n23644 , n23643 , n20953 );
buf ( n23645 , n23644 );
not ( n23646 , n23645 );
or ( n23647 , n23646 , n22242 );
or ( n23648 , n23537 , n22224 );
nand ( n23649 , n23647 , n23648 );
buf ( n23650 , n23394 );
and ( n23651 , n22277 , n23650 );
not ( n23652 , n22277 );
not ( n23653 , n23650 );
and ( n131208 , n23652 , n23653 );
nor ( n23654 , n23651 , n131208 );
or ( n23655 , n23654 , n22934 );
or ( n23656 , n23546 , n22265 );
nand ( n23657 , n23655 , n23656 );
xor ( n23658 , n23649 , n23657 );
not ( n23659 , n21577 );
not ( n23660 , n23557 );
or ( n23661 , n23659 , n23660 );
not ( n23662 , n21595 );
not ( n23663 , n23056 );
or ( n23664 , n23662 , n23663 );
not ( n23665 , n21595 );
nand ( n23666 , n23665 , n23057 );
nand ( n23667 , n23664 , n23666 );
nand ( n23668 , n23667 , n21646 );
nand ( n23669 , n23661 , n23668 );
and ( n23670 , n23658 , n23669 );
and ( n23671 , n23649 , n23657 );
or ( n23672 , n23670 , n23671 );
xor ( n23673 , n23539 , n23548 );
xor ( n23674 , n23673 , n23559 );
xor ( n23675 , n23672 , n23674 );
not ( n23676 , n19316 );
and ( n23677 , n19319 , n22737 );
not ( n23678 , n19319 );
and ( n23679 , n23678 , n22736 );
nor ( n23680 , n23677 , n23679 );
not ( n23681 , n23680 );
or ( n23682 , n23676 , n23681 );
nand ( n23683 , n23569 , n21549 );
nand ( n23684 , n23682 , n23683 );
and ( n23685 , n23675 , n23684 );
and ( n23686 , n23672 , n23674 );
or ( n23687 , n23685 , n23686 );
xor ( n23688 , n23642 , n23687 );
not ( n23689 , n22134 );
not ( n23690 , n23522 );
or ( n23691 , n23689 , n23690 );
and ( n23692 , n22137 , n22231 );
not ( n23693 , n22137 );
and ( n23694 , n23693 , n22426 );
nor ( n23695 , n23692 , n23694 );
nand ( n23696 , n23695 , n22166 );
nand ( n23697 , n23691 , n23696 );
and ( n23698 , n23688 , n23697 );
and ( n23699 , n23642 , n23687 );
or ( n23700 , n23698 , n23699 );
not ( n23701 , n23700 );
not ( n23702 , n22642 );
not ( n23703 , n23510 );
or ( n23704 , n23702 , n23703 );
and ( n23705 , n22178 , n21543 );
not ( n23706 , n22178 );
and ( n23707 , n23706 , n21546 );
nor ( n23708 , n23705 , n23707 );
nand ( n23709 , n23708 , n22645 );
nand ( n23710 , n23704 , n23709 );
not ( n23711 , n23710 );
or ( n23712 , n23701 , n23711 );
xor ( n23713 , n23562 , n23571 );
xor ( n23714 , n23713 , n23574 );
not ( n23715 , n22121 );
and ( n23716 , n22071 , n22273 );
not ( n23717 , n22071 );
and ( n23718 , n23717 , n22274 );
nor ( n23719 , n23716 , n23718 );
not ( n23720 , n23719 );
or ( n23721 , n23715 , n23720 );
not ( n23722 , n22061 );
buf ( n23723 , n23610 );
nand ( n23724 , n23722 , n23723 );
nand ( n23725 , n23721 , n23724 );
xor ( n23726 , n23714 , n23725 );
not ( n23727 , n21837 );
not ( n23728 , n23636 );
or ( n23729 , n23727 , n23728 );
and ( n23730 , n21651 , n22535 );
not ( n23731 , n21651 );
and ( n23732 , n23731 , n22742 );
or ( n23733 , n23730 , n23732 );
not ( n23734 , n23733 );
nand ( n23735 , n23734 , n21698 );
nand ( n23736 , n23729 , n23735 );
not ( n23737 , n22225 );
not ( n23738 , n23645 );
or ( n23739 , n23737 , n23738 );
not ( n23740 , n20943 );
not ( n23741 , n23740 );
not ( n23742 , n20950 );
nand ( n23743 , n20952 , n23742 );
not ( n23744 , n23743 );
or ( n23745 , n23741 , n23744 );
not ( n23746 , n23743 );
nand ( n23747 , n23746 , n20943 );
nand ( n23748 , n23745 , n23747 );
buf ( n23749 , n23748 );
not ( n23750 , n23749 );
or ( n23751 , n23750 , n22242 );
nand ( n23752 , n23739 , n23751 );
not ( n23753 , n22264 );
not ( n23754 , n23654 );
not ( n23755 , n23754 );
or ( n23756 , n23753 , n23755 );
buf ( n23757 , n23536 );
and ( n23758 , n22268 , n23757 );
not ( n23759 , n22268 );
and ( n23760 , n23759 , n23537 );
nor ( n23761 , n23758 , n23760 );
nand ( n23762 , n23761 , n22299 );
nand ( n23763 , n23756 , n23762 );
xor ( n23764 , n23752 , n23763 );
not ( n23765 , n21577 );
not ( n23766 , n23667 );
or ( n23767 , n23765 , n23766 );
not ( n23768 , n21595 );
not ( n23769 , n23045 );
or ( n23770 , n23768 , n23769 );
nand ( n23771 , n23046 , n21623 );
nand ( n23772 , n23770 , n23771 );
nand ( n23773 , n23772 , n21646 );
nand ( n23774 , n23767 , n23773 );
and ( n23775 , n23764 , n23774 );
and ( n23776 , n23752 , n23763 );
or ( n23777 , n23775 , n23776 );
xor ( n23778 , n23649 , n23657 );
xor ( n23779 , n23778 , n23669 );
xor ( n23780 , n23777 , n23779 );
not ( n23781 , n19316 );
not ( n23782 , n19319 );
not ( n23783 , n22926 );
or ( n23784 , n23782 , n23783 );
nand ( n23785 , n22884 , n19318 );
nand ( n23786 , n23784 , n23785 );
not ( n23787 , n23786 );
or ( n23788 , n23781 , n23787 );
nand ( n23789 , n23680 , n21549 );
nand ( n23790 , n23788 , n23789 );
and ( n23791 , n23780 , n23790 );
and ( n23792 , n23777 , n23779 );
or ( n23793 , n23791 , n23792 );
xor ( n23794 , n23736 , n23793 );
not ( n23795 , n22166 );
not ( n23796 , n22137 );
not ( n23797 , n22544 );
or ( n23798 , n23796 , n23797 );
nand ( n23799 , n22241 , n22136 );
nand ( n23800 , n23798 , n23799 );
not ( n23801 , n23800 );
or ( n23802 , n23795 , n23801 );
nand ( n23803 , n23695 , n22134 );
nand ( n23804 , n23802 , n23803 );
and ( n23805 , n23794 , n23804 );
and ( n23806 , n23736 , n23793 );
or ( n23807 , n23805 , n23806 );
and ( n23808 , n23726 , n23807 );
and ( n23809 , n23714 , n23725 );
or ( n23810 , n23808 , n23809 );
not ( n23811 , n23700 );
not ( n23812 , n23710 );
nand ( n23813 , n23811 , n23812 );
nand ( n23814 , n23810 , n23813 );
nand ( n23815 , n23712 , n23814 );
and ( n23816 , n23632 , n23815 );
and ( n23817 , n23629 , n23631 );
or ( n23818 , n23816 , n23817 );
nand ( n23819 , n23605 , n23818 );
not ( n23820 , n23599 );
nand ( n23821 , n23820 , n23602 );
and ( n23822 , n23819 , n23821 );
nand ( n23823 , n23593 , n23822 );
and ( n23824 , n23591 , n23823 );
not ( n23825 , n23824 );
xnor ( n23826 , n23599 , n23818 );
and ( n23827 , n23826 , n23603 );
not ( n23828 , n23826 );
and ( n23829 , n23828 , n23602 );
nor ( n23830 , n23827 , n23829 );
xor ( n23831 , n23629 , n23631 );
xor ( n23832 , n23831 , n23815 );
xor ( n23833 , n23516 , n23526 );
xor ( n23834 , n23833 , n23577 );
xor ( n23835 , n23614 , n23616 );
xor ( n23836 , n23835 , n23626 );
xor ( n23837 , n23834 , n23836 );
not ( n23838 , n22051 );
and ( n23839 , n21853 , n21636 );
not ( n23840 , n21853 );
and ( n23841 , n23840 , n21637 );
nor ( n23842 , n23839 , n23841 );
not ( n23843 , n23842 );
or ( n23844 , n23838 , n23843 );
nand ( n23845 , n23622 , n21846 );
nand ( n23846 , n23844 , n23845 );
xor ( n23847 , n23642 , n23687 );
xor ( n23848 , n23847 , n23697 );
xor ( n23849 , n23846 , n23848 );
not ( n23850 , n22642 );
not ( n23851 , n23708 );
or ( n23852 , n23850 , n23851 );
and ( n23853 , n22178 , n21456 );
not ( n23854 , n22178 );
and ( n23855 , n23854 , n21459 );
nor ( n23856 , n23853 , n23855 );
nand ( n23857 , n23856 , n22645 );
nand ( n23858 , n23852 , n23857 );
and ( n23859 , n23849 , n23858 );
and ( n23860 , n23846 , n23848 );
or ( n23861 , n23859 , n23860 );
and ( n23862 , n23837 , n23861 );
and ( n23863 , n23834 , n23836 );
or ( n23864 , n23862 , n23863 );
not ( n23865 , n23864 );
xor ( n23866 , n23513 , n23580 );
and ( n23867 , n23866 , n23582 );
not ( n23868 , n23866 );
and ( n23869 , n23868 , n23501 );
nor ( n23870 , n23867 , n23869 );
nand ( n23871 , n23865 , n23870 );
nand ( n23872 , n23832 , n23871 );
not ( n23873 , n23870 );
nand ( n23874 , n23873 , n23864 );
and ( n23875 , n23872 , n23874 );
nand ( n23876 , n23830 , n23875 );
and ( n23877 , n23870 , n23864 );
not ( n23878 , n23870 );
and ( n23879 , n23878 , n23865 );
or ( n23880 , n23877 , n23879 );
xnor ( n23881 , n23880 , n23832 );
xor ( n23882 , n23834 , n23836 );
xor ( n23883 , n23882 , n23861 );
not ( n23884 , n23883 );
not ( n23885 , n23884 );
xor ( n23886 , n23812 , n23700 );
xor ( n23887 , n23886 , n23810 );
not ( n23888 , n23887 );
and ( n23889 , n23885 , n23888 );
nand ( n23890 , n23884 , n23887 );
xor ( n23891 , n23672 , n23674 );
xor ( n23892 , n23891 , n23684 );
not ( n23893 , n22062 );
not ( n23894 , n23719 );
or ( n23895 , n23893 , n23894 );
and ( n23896 , n22071 , n22288 );
not ( n23897 , n22071 );
and ( n23898 , n23897 , n22289 );
nor ( n23899 , n23896 , n23898 );
nand ( n23900 , n23899 , n22121 );
nand ( n23901 , n23895 , n23900 );
xor ( n23902 , n23892 , n23901 );
not ( n23903 , n21846 );
not ( n23904 , n23842 );
or ( n23905 , n23903 , n23904 );
not ( n23906 , n21853 );
not ( n23907 , n22317 );
or ( n23908 , n23906 , n23907 );
nand ( n23909 , n22314 , n21852 );
nand ( n23910 , n23908 , n23909 );
nand ( n23911 , n23910 , n22051 );
nand ( n23912 , n23905 , n23911 );
and ( n23913 , n23902 , n23912 );
and ( n23914 , n23892 , n23901 );
or ( n23915 , n23913 , n23914 );
or ( n23916 , n23733 , n22877 );
not ( n23917 , n21651 );
not ( n23918 , n22612 );
or ( n23919 , n23917 , n23918 );
nand ( n23920 , n22611 , n21834 );
nand ( n23921 , n23919 , n23920 );
nand ( n23922 , n23921 , n21698 );
nand ( n23923 , n23916 , n23922 );
not ( n23924 , n22134 );
not ( n23925 , n23800 );
or ( n23926 , n23924 , n23925 );
not ( n23927 , n22137 );
not ( n23928 , n22418 );
or ( n23929 , n23927 , n23928 );
nand ( n23930 , n22417 , n22136 );
nand ( n23931 , n23929 , n23930 );
nand ( n23932 , n23931 , n22166 );
nand ( n23933 , n23926 , n23932 );
or ( n23934 , n23923 , n23933 );
not ( n23935 , n20928 );
not ( n23936 , n20941 );
or ( n23937 , n23935 , n23936 );
nand ( n23938 , n23937 , n20937 );
not ( n23939 , n20937 );
nand ( n23940 , n20941 , n20928 , n23939 );
nand ( n23941 , n23938 , n23940 );
not ( n23942 , n23941 );
or ( n23943 , n23942 , n22242 );
or ( n23944 , n23750 , n22224 );
nand ( n23945 , n23943 , n23944 );
not ( n23946 , n22264 );
not ( n23947 , n23761 );
or ( n23948 , n23946 , n23947 );
and ( n23949 , n22268 , n23645 );
not ( n23950 , n22268 );
not ( n23951 , n23644 );
and ( n23952 , n23950 , n23951 );
nor ( n23953 , n23949 , n23952 );
not ( n23954 , n23953 );
or ( n23955 , n23954 , n22934 );
nand ( n23956 , n23948 , n23955 );
xor ( n23957 , n23945 , n23956 );
not ( n23958 , n21577 );
not ( n23959 , n23772 );
or ( n23960 , n23958 , n23959 );
and ( n23961 , n21594 , n23395 );
not ( n23962 , n21594 );
and ( n23963 , n23962 , n23394 );
nor ( n23964 , n23961 , n23963 );
nand ( n23965 , n23964 , n21646 );
nand ( n23966 , n23960 , n23965 );
and ( n23967 , n23957 , n23966 );
and ( n23968 , n23945 , n23956 );
or ( n23969 , n23967 , n23968 );
xor ( n23970 , n23752 , n23763 );
xor ( n23971 , n23970 , n23774 );
xor ( n23972 , n23969 , n23971 );
not ( n23973 , n21549 );
not ( n23974 , n23786 );
or ( n23975 , n23973 , n23974 );
not ( n23976 , n19318 );
and ( n23977 , n23976 , n23027 );
not ( n23978 , n23976 );
and ( n23979 , n23978 , n22892 );
nor ( n23980 , n23977 , n23979 );
nand ( n23981 , n23980 , n19316 );
nand ( n23982 , n23975 , n23981 );
and ( n23983 , n23972 , n23982 );
and ( n23984 , n23969 , n23971 );
or ( n23985 , n23983 , n23984 );
nand ( n23986 , n23934 , n23985 );
nand ( n23987 , n23933 , n23923 );
nand ( n23988 , n23986 , n23987 );
xor ( n23989 , n23736 , n23793 );
xor ( n23990 , n23989 , n23804 );
xor ( n23991 , n23988 , n23990 );
xor ( n23992 , n23777 , n23779 );
xor ( n23993 , n23992 , n23790 );
not ( n23994 , n22225 );
not ( n23995 , n23941 );
or ( n23996 , n23994 , n23995 );
not ( n23997 , n20934 );
not ( n23998 , n20936 );
or ( n23999 , n23997 , n23998 );
nand ( n24000 , n23999 , n23939 );
not ( n24001 , n24000 );
not ( n24002 , n24001 );
or ( n24003 , n22242 , n24002 );
nand ( n24004 , n23996 , n24003 );
not ( n24005 , n22264 );
not ( n24006 , n23953 );
or ( n24007 , n24005 , n24006 );
and ( n24008 , n22268 , n23749 );
not ( n24009 , n22268 );
and ( n24010 , n24009 , n23750 );
nor ( n24011 , n24008 , n24010 );
nand ( n24012 , n24011 , n22299 );
nand ( n24013 , n24007 , n24012 );
xor ( n24014 , n24004 , n24013 );
not ( n24015 , n20935 );
not ( n24016 , n24015 );
or ( n24017 , n22242 , n24016 );
or ( n24018 , n24002 , n22224 );
nand ( n24019 , n24017 , n24018 );
not ( n24020 , n24011 );
not ( n24021 , n22264 );
or ( n24022 , n24020 , n24021 );
and ( n24023 , n22268 , n23941 );
not ( n24024 , n22268 );
buf ( n24025 , n23941 );
not ( n24026 , n24025 );
and ( n24027 , n24024 , n24026 );
nor ( n24028 , n24023 , n24027 );
nand ( n24029 , n24028 , n22299 );
nand ( n24030 , n24022 , n24029 );
xor ( n24031 , n24019 , n24030 );
and ( n24032 , n22225 , n24015 );
not ( n24033 , n22299 );
and ( n24034 , n22294 , n24002 );
not ( n24035 , n22294 );
and ( n24036 , n24035 , n24001 );
nor ( n24037 , n24034 , n24036 );
not ( n24038 , n24037 );
or ( n24039 , n24033 , n24038 );
nand ( n24040 , n24028 , n22264 );
nand ( n24041 , n24039 , n24040 );
xor ( n24042 , n24032 , n24041 );
and ( n24043 , n22259 , n24015 );
and ( n24044 , n22295 , n24016 );
nor ( n24045 , n24044 , n21594 );
nor ( n24046 , n24043 , n24045 , n22277 );
not ( n24047 , n22264 );
not ( n24048 , n24037 );
or ( n24049 , n24047 , n24048 );
or ( n24050 , n22268 , n24016 );
or ( n24051 , n22277 , n24015 );
nand ( n24052 , n24050 , n24051 );
nand ( n24053 , n22299 , n24052 );
nand ( n24054 , n24049 , n24053 );
and ( n24055 , n24046 , n24054 );
and ( n24056 , n24042 , n24055 );
and ( n24057 , n24032 , n24041 );
or ( n24058 , n24056 , n24057 );
and ( n24059 , n24031 , n24058 );
and ( n24060 , n24019 , n24030 );
or ( n24061 , n24059 , n24060 );
and ( n24062 , n24014 , n24061 );
and ( n24063 , n24004 , n24013 );
or ( n24064 , n24062 , n24063 );
xor ( n24065 , n23945 , n23956 );
xor ( n24066 , n24065 , n23966 );
xor ( n24067 , n24064 , n24066 );
not ( n24068 , n21549 );
not ( n24069 , n23980 );
or ( n24070 , n24068 , n24069 );
not ( n24071 , n23976 );
not ( n24072 , n23056 );
or ( n24073 , n24071 , n24072 );
nand ( n24074 , n23057 , n19318 );
nand ( n24075 , n24073 , n24074 );
nand ( n24076 , n24075 , n19316 );
nand ( n24077 , n24070 , n24076 );
and ( n24078 , n24067 , n24077 );
and ( n24079 , n24064 , n24066 );
or ( n24080 , n24078 , n24079 );
not ( n24081 , n21837 );
not ( n24082 , n23921 );
or ( n24083 , n24081 , n24082 );
not ( n24084 , n21651 );
not ( n24085 , n22736 );
or ( n24086 , n24084 , n24085 );
nand ( n24087 , n22737 , n21834 );
nand ( n24088 , n24086 , n24087 );
nand ( n24089 , n24088 , n21698 );
nand ( n24090 , n24083 , n24089 );
xor ( n24091 , n24080 , n24090 );
not ( n24092 , n22166 );
and ( n24093 , n22137 , n22535 );
not ( n24094 , n22137 );
and ( n24095 , n24094 , n22742 );
nor ( n24096 , n24093 , n24095 );
not ( n24097 , n24096 );
or ( n24098 , n24092 , n24097 );
nand ( n24099 , n23931 , n22134 );
nand ( n24100 , n24098 , n24099 );
and ( n24101 , n24091 , n24100 );
and ( n24102 , n24080 , n24090 );
or ( n24103 , n24101 , n24102 );
xor ( n24104 , n23993 , n24103 );
not ( n24105 , n22062 );
not ( n24106 , n23899 );
or ( n24107 , n24105 , n24106 );
and ( n24108 , n22071 , n22231 );
not ( n24109 , n22071 );
and ( n24110 , n24109 , n22426 );
nor ( n24111 , n24108 , n24110 );
nand ( n24112 , n24111 , n22121 );
nand ( n24113 , n24107 , n24112 );
and ( n24114 , n24104 , n24113 );
and ( n24115 , n23993 , n24103 );
or ( n24116 , n24114 , n24115 );
and ( n24117 , n23991 , n24116 );
and ( n24118 , n23988 , n23990 );
or ( n24119 , n24117 , n24118 );
xor ( n24120 , n23915 , n24119 );
xor ( n24121 , n23714 , n23725 );
xor ( n24122 , n24121 , n23807 );
and ( n24123 , n24120 , n24122 );
and ( n24124 , n23915 , n24119 );
or ( n24125 , n24123 , n24124 );
and ( n24126 , n23890 , n24125 );
nor ( n24127 , n23889 , n24126 );
nand ( n24128 , n23881 , n24127 );
and ( n24129 , n23876 , n24128 );
not ( n24130 , n24129 );
xnor ( n24131 , n23887 , n24125 );
and ( n24132 , n24131 , n23883 );
not ( n24133 , n24131 );
and ( n24134 , n24133 , n23884 );
nor ( n24135 , n24132 , n24134 );
xor ( n24136 , n23846 , n23848 );
xor ( n24137 , n24136 , n23858 );
not ( n24138 , n22642 );
not ( n24139 , n23856 );
or ( n24140 , n24138 , n24139 );
not ( n24141 , n22178 );
not ( n24142 , n21620 );
or ( n24143 , n24141 , n24142 );
nand ( n24144 , n21619 , n22179 );
nand ( n24145 , n24143 , n24144 );
nand ( n24146 , n24145 , n22645 );
nand ( n24147 , n24140 , n24146 );
xor ( n24148 , n23892 , n23901 );
xor ( n24149 , n24148 , n23912 );
xor ( n24150 , n24147 , n24149 );
xor ( n24151 , n23923 , n23985 );
xnor ( n24152 , n24151 , n23933 );
not ( n24153 , n24152 );
not ( n24154 , n24153 );
not ( n24155 , n21846 );
not ( n24156 , n23910 );
or ( n24157 , n24155 , n24156 );
not ( n24158 , n21853 );
not ( n24159 , n22274 );
or ( n24160 , n24158 , n24159 );
nand ( n24161 , n22273 , n21852 );
nand ( n24162 , n24160 , n24161 );
nand ( n24163 , n24162 , n22051 );
nand ( n24164 , n24157 , n24163 );
not ( n24165 , n24164 );
or ( n24166 , n24154 , n24165 );
or ( n24167 , n24164 , n24153 );
xor ( n24168 , n23969 , n23971 );
xor ( n24169 , n24168 , n23982 );
not ( n24170 , n22062 );
not ( n24171 , n24111 );
or ( n24172 , n24170 , n24171 );
and ( n24173 , n22071 , n22241 );
not ( n24174 , n22071 );
and ( n24175 , n24174 , n22544 );
nor ( n24176 , n24173 , n24175 );
nand ( n24177 , n24176 , n22121 );
nand ( n24178 , n24172 , n24177 );
xor ( n24179 , n24169 , n24178 );
xor ( n24180 , n24080 , n24090 );
xor ( n24181 , n24180 , n24100 );
and ( n24182 , n24179 , n24181 );
and ( n24183 , n24169 , n24178 );
or ( n24184 , n24182 , n24183 );
nand ( n24185 , n24167 , n24184 );
nand ( n24186 , n24166 , n24185 );
and ( n24187 , n24150 , n24186 );
and ( n24188 , n24147 , n24149 );
or ( n24189 , n24187 , n24188 );
xor ( n24190 , n24137 , n24189 );
xor ( n24191 , n23915 , n24119 );
xor ( n24192 , n24191 , n24122 );
and ( n24193 , n24190 , n24192 );
and ( n24194 , n24137 , n24189 );
or ( n24195 , n24193 , n24194 );
nor ( n24196 , n24135 , n24195 );
xor ( n24197 , n24137 , n24189 );
xor ( n24198 , n24197 , n24192 );
not ( n24199 , n22642 );
not ( n24200 , n24145 );
or ( n24201 , n24199 , n24200 );
and ( n24202 , n22178 , n21636 );
not ( n24203 , n22178 );
and ( n24204 , n24203 , n21637 );
nor ( n24205 , n24202 , n24204 );
nand ( n24206 , n24205 , n22645 );
nand ( n24207 , n24201 , n24206 );
xor ( n24208 , n23993 , n24103 );
xor ( n24209 , n24208 , n24113 );
xor ( n24210 , n24207 , n24209 );
not ( n24211 , n21837 );
not ( n24212 , n24088 );
or ( n24213 , n24211 , n24212 );
and ( n24214 , n21651 , n22884 );
not ( n24215 , n21651 );
and ( n24216 , n24215 , n22926 );
nor ( n24217 , n24214 , n24216 );
nand ( n24218 , n24217 , n21698 );
nand ( n24219 , n24213 , n24218 );
not ( n24220 , n24219 );
not ( n24221 , n22134 );
not ( n24222 , n24096 );
or ( n24223 , n24221 , n24222 );
and ( n24224 , n22137 , n22611 );
not ( n24225 , n22137 );
and ( n24226 , n24225 , n22612 );
nor ( n24227 , n24224 , n24226 );
nand ( n24228 , n24227 , n22166 );
nand ( n24229 , n24223 , n24228 );
not ( n24230 , n24229 );
or ( n24231 , n24220 , n24230 );
or ( n24232 , n24229 , n24219 );
not ( n24233 , n21549 );
not ( n24234 , n24075 );
or ( n24235 , n24233 , n24234 );
and ( n24236 , n23976 , n23046 );
not ( n24237 , n23976 );
and ( n24238 , n24237 , n23045 );
nor ( n24239 , n24236 , n24238 );
nand ( n24240 , n24239 , n19316 );
nand ( n24241 , n24235 , n24240 );
not ( n24242 , n24241 );
not ( n24243 , n21577 );
not ( n24244 , n23964 );
or ( n24245 , n24243 , n24244 );
xor ( n24246 , n21595 , n23757 );
nand ( n24247 , n24246 , n21646 );
nand ( n24248 , n24245 , n24247 );
not ( n24249 , n24248 );
nand ( n24250 , n24242 , n24249 );
xor ( n24251 , n24004 , n24013 );
xor ( n24252 , n24251 , n24061 );
and ( n24253 , n24250 , n24252 );
and ( n24254 , n24241 , n24248 );
nor ( n24255 , n24253 , n24254 );
not ( n24256 , n24255 );
nand ( n24257 , n24232 , n24256 );
nand ( n24258 , n24231 , n24257 );
not ( n24259 , n24258 );
not ( n24260 , n21846 );
not ( n24261 , n24162 );
or ( n24262 , n24260 , n24261 );
not ( n24263 , n21851 );
not ( n24264 , n22289 );
or ( n24265 , n24263 , n24264 );
nand ( n24266 , n22288 , n21852 );
nand ( n24267 , n24265 , n24266 );
nand ( n24268 , n24267 , n22051 );
nand ( n24269 , n24262 , n24268 );
not ( n24270 , n24269 );
or ( n24271 , n24259 , n24270 );
or ( n24272 , n24269 , n24258 );
xor ( n24273 , n24064 , n24066 );
xor ( n24274 , n24273 , n24077 );
xor ( n24275 , n24019 , n24030 );
xor ( n24276 , n24275 , n24058 );
not ( n24277 , n21577 );
not ( n24278 , n24246 );
or ( n24279 , n24277 , n24278 );
and ( n24280 , n21595 , n23644 );
not ( n24281 , n21595 );
and ( n24282 , n24281 , n23646 );
nor ( n24283 , n24280 , n24282 );
nand ( n24284 , n24283 , n21646 );
nand ( n24285 , n24279 , n24284 );
xor ( n24286 , n24276 , n24285 );
xor ( n24287 , n24032 , n24041 );
xor ( n24288 , n24287 , n24055 );
not ( n24289 , n21577 );
not ( n24290 , n24283 );
or ( n24291 , n24289 , n24290 );
and ( n24292 , n21595 , n23749 );
not ( n24293 , n21595 );
and ( n24294 , n24293 , n23750 );
nor ( n24295 , n24292 , n24294 );
nand ( n24296 , n24295 , n21646 );
nand ( n24297 , n24291 , n24296 );
xor ( n24298 , n24288 , n24297 );
xor ( n24299 , n24046 , n24054 );
not ( n24300 , n21577 );
not ( n24301 , n24295 );
or ( n24302 , n24300 , n24301 );
and ( n24303 , n21595 , n23941 );
not ( n24304 , n21595 );
and ( n24305 , n24304 , n23942 );
nor ( n24306 , n24303 , n24305 );
not ( n24307 , n24306 );
or ( n24308 , n24307 , n23170 );
nand ( n24309 , n24302 , n24308 );
xor ( n24310 , n24299 , n24309 );
nor ( n24311 , n22265 , n24016 );
not ( n24312 , n21577 );
not ( n24313 , n24306 );
or ( n24314 , n24312 , n24313 );
xnor ( n24315 , n21595 , n24002 );
nand ( n24316 , n24315 , n21646 );
nand ( n24317 , n24314 , n24316 );
xor ( n24318 , n24311 , n24317 );
and ( n24319 , n21572 , n24015 );
and ( n24320 , n21642 , n24016 );
nor ( n24321 , n24320 , n19318 );
nor ( n24322 , n24319 , n24321 , n21594 );
not ( n24323 , n21577 );
not ( n24324 , n24315 );
or ( n24325 , n24323 , n24324 );
or ( n24326 , n21595 , n24016 );
or ( n24327 , n21594 , n24015 );
nand ( n24328 , n24326 , n24327 );
nand ( n24329 , n21646 , n24328 );
nand ( n24330 , n24325 , n24329 );
and ( n24331 , n24322 , n24330 );
and ( n24332 , n24318 , n24331 );
and ( n24333 , n24311 , n24317 );
or ( n24334 , n24332 , n24333 );
and ( n24335 , n24310 , n24334 );
and ( n24336 , n24299 , n24309 );
or ( n24337 , n24335 , n24336 );
and ( n24338 , n24298 , n24337 );
and ( n24339 , n24288 , n24297 );
or ( n24340 , n24338 , n24339 );
and ( n24341 , n24286 , n24340 );
and ( n24342 , n24276 , n24285 );
or ( n24343 , n24341 , n24342 );
not ( n24344 , n21837 );
not ( n24345 , n24217 );
or ( n24346 , n24344 , n24345 );
and ( n24347 , n21651 , n23027 );
not ( n24348 , n21651 );
and ( n24349 , n24348 , n22892 );
nor ( n24350 , n24347 , n24349 );
nand ( n24351 , n24350 , n21698 );
nand ( n24352 , n24346 , n24351 );
xor ( n24353 , n24343 , n24352 );
and ( n24354 , n24252 , n24249 );
not ( n24355 , n24252 );
and ( n24356 , n24355 , n24248 );
nor ( n24357 , n24354 , n24356 );
not ( n24358 , n24357 );
not ( n24359 , n24241 );
or ( n24360 , n24358 , n24359 );
or ( n24361 , n24241 , n24357 );
nand ( n24362 , n24360 , n24361 );
and ( n24363 , n24353 , n24362 );
and ( n24364 , n24343 , n24352 );
or ( n24365 , n24363 , n24364 );
xor ( n24366 , n24274 , n24365 );
not ( n24367 , n22062 );
not ( n24368 , n24176 );
or ( n24369 , n24367 , n24368 );
and ( n24370 , n22071 , n22417 );
not ( n24371 , n22071 );
and ( n24372 , n24371 , n22418 );
nor ( n24373 , n24370 , n24372 );
nand ( n24374 , n24373 , n22121 );
nand ( n24375 , n24369 , n24374 );
and ( n24376 , n24366 , n24375 );
and ( n24377 , n24274 , n24365 );
or ( n24378 , n24376 , n24377 );
nand ( n24379 , n24272 , n24378 );
nand ( n24380 , n24271 , n24379 );
and ( n24381 , n24210 , n24380 );
and ( n24382 , n24207 , n24209 );
or ( n24383 , n24381 , n24382 );
xor ( n24384 , n23988 , n23990 );
xor ( n24385 , n24384 , n24116 );
xor ( n24386 , n24383 , n24385 );
xor ( n24387 , n24147 , n24149 );
xor ( n24388 , n24387 , n24186 );
and ( n24389 , n24386 , n24388 );
and ( n24390 , n24383 , n24385 );
or ( n24391 , n24389 , n24390 );
nor ( n24392 , n24198 , n24391 );
nor ( n24393 , n24196 , n24392 );
not ( n24394 , n24393 );
xor ( n24395 , n24383 , n24385 );
xor ( n24396 , n24395 , n24388 );
xor ( n24397 , n24207 , n24209 );
xor ( n24398 , n24397 , n24380 );
and ( n24399 , n24164 , n24152 );
not ( n24400 , n24164 );
and ( n24401 , n24400 , n24153 );
or ( n24402 , n24399 , n24401 );
not ( n24403 , n24184 );
and ( n24404 , n24402 , n24403 );
not ( n24405 , n24402 );
and ( n24406 , n24405 , n24184 );
nor ( n24407 , n24404 , n24406 );
not ( n24408 , n24407 );
or ( n24409 , n24398 , n24408 );
not ( n24410 , n22645 );
not ( n24411 , n22178 );
not ( n24412 , n22317 );
or ( n24413 , n24411 , n24412 );
nand ( n24414 , n22314 , n22179 );
nand ( n24415 , n24413 , n24414 );
not ( n24416 , n24415 );
or ( n24417 , n24410 , n24416 );
nand ( n24418 , n24205 , n22642 );
nand ( n24419 , n24417 , n24418 );
not ( n24420 , n24419 );
xor ( n24421 , n24169 , n24178 );
xor ( n24422 , n24421 , n24181 );
not ( n24423 , n24422 );
or ( n24424 , n24420 , n24423 );
or ( n24425 , n24419 , n24422 );
xor ( n24426 , n24219 , n24255 );
xor ( n24427 , n24426 , n24229 );
not ( n24428 , n24427 );
not ( n24429 , n24428 );
not ( n24430 , n21846 );
not ( n24431 , n24267 );
or ( n24432 , n24430 , n24431 );
and ( n24433 , n22231 , n21853 );
not ( n24434 , n22231 );
and ( n24435 , n24434 , n21852 );
nor ( n24436 , n24433 , n24435 );
nand ( n24437 , n24436 , n22051 );
nand ( n24438 , n24432 , n24437 );
not ( n24439 , n24438 );
or ( n24440 , n24429 , n24439 );
or ( n24441 , n24438 , n24428 );
not ( n24442 , n21549 );
not ( n24443 , n24239 );
or ( n24444 , n24442 , n24443 );
and ( n24445 , n19318 , n23650 );
not ( n24446 , n19318 );
and ( n24447 , n24446 , n23653 );
nor ( n24448 , n24445 , n24447 );
or ( n24449 , n24448 , n22573 );
nand ( n24450 , n24444 , n24449 );
xor ( n24451 , n24276 , n24285 );
xor ( n24452 , n24451 , n24340 );
xor ( n24453 , n24450 , n24452 );
not ( n24454 , n21698 );
xor ( n24455 , n21651 , n23055 );
not ( n24456 , n24455 );
or ( n24457 , n24454 , n24456 );
nand ( n24458 , n24350 , n21837 );
nand ( n24459 , n24457 , n24458 );
and ( n24460 , n24453 , n24459 );
and ( n24461 , n24450 , n24452 );
or ( n24462 , n24460 , n24461 );
not ( n24463 , n22134 );
not ( n24464 , n24227 );
or ( n24465 , n24463 , n24464 );
and ( n24466 , n22137 , n22737 );
not ( n24467 , n22137 );
and ( n24468 , n24467 , n22736 );
nor ( n24469 , n24466 , n24468 );
nand ( n24470 , n24469 , n22166 );
nand ( n24471 , n24465 , n24470 );
xor ( n24472 , n24462 , n24471 );
not ( n24473 , n22062 );
not ( n24474 , n24373 );
or ( n24475 , n24473 , n24474 );
and ( n24476 , n22071 , n22535 );
not ( n24477 , n22071 );
and ( n24478 , n24477 , n22742 );
nor ( n24479 , n24476 , n24478 );
nand ( n24480 , n24479 , n22121 );
nand ( n24481 , n24475 , n24480 );
and ( n24482 , n24472 , n24481 );
and ( n24483 , n24462 , n24471 );
or ( n24484 , n24482 , n24483 );
nand ( n24485 , n24441 , n24484 );
nand ( n24486 , n24440 , n24485 );
nand ( n24487 , n24425 , n24486 );
nand ( n24488 , n24424 , n24487 );
nand ( n24489 , n24409 , n24488 );
nand ( n24490 , n24398 , n24408 );
nand ( n24491 , n24489 , n24490 );
xor ( n24492 , n24396 , n24491 );
xor ( n24493 , n24488 , n24407 );
xor ( n24494 , n24493 , n24398 );
xor ( n24495 , n24269 , n24258 );
xnor ( n24496 , n24495 , n24378 );
xor ( n24497 , n24343 , n24352 );
xor ( n24498 , n24497 , n24362 );
not ( n24499 , n21846 );
not ( n24500 , n24436 );
or ( n24501 , n24499 , n24500 );
and ( n24502 , n21853 , n22241 );
not ( n24503 , n21853 );
and ( n24504 , n24503 , n22544 );
nor ( n24505 , n24502 , n24504 );
nand ( n24506 , n24505 , n22051 );
nand ( n24507 , n24501 , n24506 );
xor ( n24508 , n24498 , n24507 );
not ( n24509 , n21549 );
not ( n24510 , n24448 );
not ( n24511 , n24510 );
or ( n24512 , n24509 , n24511 );
and ( n24513 , n23976 , n23536 );
not ( n24514 , n23976 );
and ( n24515 , n24514 , n23537 );
nor ( n24516 , n24513 , n24515 );
nand ( n24517 , n24516 , n19316 );
nand ( n24518 , n24512 , n24517 );
xor ( n24519 , n24288 , n24297 );
xor ( n24520 , n24519 , n24337 );
xor ( n24521 , n24518 , n24520 );
not ( n24522 , n21837 );
not ( n24523 , n24455 );
or ( n24524 , n24522 , n24523 );
and ( n24525 , n21834 , n23046 );
not ( n24526 , n21834 );
and ( n24527 , n24526 , n23045 );
nor ( n24528 , n24525 , n24527 );
not ( n24529 , n24528 );
nand ( n24530 , n24529 , n21698 );
nand ( n24531 , n24524 , n24530 );
and ( n24532 , n24521 , n24531 );
and ( n24533 , n24518 , n24520 );
or ( n24534 , n24532 , n24533 );
not ( n24535 , n22134 );
not ( n24536 , n24469 );
or ( n24537 , n24535 , n24536 );
buf ( n24538 , n21692 );
and ( n24539 , n24538 , n22884 );
not ( n24540 , n24538 );
and ( n24541 , n24540 , n22926 );
nor ( n24542 , n24539 , n24541 );
nand ( n24543 , n24542 , n22166 );
nand ( n24544 , n24537 , n24543 );
xor ( n24545 , n24534 , n24544 );
xor ( n24546 , n24450 , n24452 );
xor ( n24547 , n24546 , n24459 );
and ( n24548 , n24545 , n24547 );
and ( n24549 , n24534 , n24544 );
or ( n24550 , n24548 , n24549 );
and ( n24551 , n24508 , n24550 );
and ( n24552 , n24498 , n24507 );
or ( n24553 , n24551 , n24552 );
xor ( n24554 , n24274 , n24365 );
xor ( n24555 , n24554 , n24375 );
xor ( n24556 , n24553 , n24555 );
not ( n24557 , n22645 );
and ( n24558 , n22273 , n22178 );
not ( n24559 , n22273 );
and ( n24560 , n24559 , n22179 );
nor ( n24561 , n24558 , n24560 );
not ( n24562 , n24561 );
or ( n24563 , n24557 , n24562 );
nand ( n24564 , n24415 , n22642 );
nand ( n24565 , n24563 , n24564 );
and ( n24566 , n24556 , n24565 );
and ( n24567 , n24553 , n24555 );
or ( n24568 , n24566 , n24567 );
not ( n24569 , n24568 );
xor ( n24570 , n24496 , n24569 );
xor ( n24571 , n24419 , n24422 );
xnor ( n24572 , n24571 , n24486 );
and ( n24573 , n24570 , n24572 );
and ( n24574 , n24496 , n24569 );
or ( n24575 , n24573 , n24574 );
nand ( n24576 , n24494 , n24575 );
xor ( n24577 , n24496 , n24569 );
xor ( n24578 , n24577 , n24572 );
xor ( n24579 , n24553 , n24555 );
xor ( n24580 , n24579 , n24565 );
not ( n24581 , n22642 );
not ( n24582 , n24561 );
or ( n24583 , n24581 , n24582 );
not ( n24584 , n22178 );
not ( n24585 , n22289 );
or ( n24586 , n24584 , n24585 );
nand ( n24587 , n22288 , n22179 );
nand ( n24588 , n24586 , n24587 );
nand ( n24589 , n24588 , n22645 );
nand ( n24590 , n24583 , n24589 );
xor ( n24591 , n24462 , n24471 );
xor ( n24592 , n24591 , n24481 );
xor ( n24593 , n24590 , n24592 );
xor ( n24594 , n24299 , n24309 );
xor ( n24595 , n24594 , n24334 );
not ( n24596 , n24595 );
not ( n24597 , n21549 );
not ( n24598 , n24516 );
or ( n24599 , n24597 , n24598 );
and ( n24600 , n23976 , n23644 );
not ( n24601 , n23976 );
and ( n24602 , n24601 , n23646 );
nor ( n24603 , n24600 , n24602 );
nand ( n24604 , n24603 , n19316 );
nand ( n24605 , n24599 , n24604 );
not ( n24606 , n24605 );
or ( n24607 , n24596 , n24606 );
or ( n24608 , n24605 , n24595 );
xor ( n24609 , n24311 , n24317 );
xor ( n24610 , n24609 , n24331 );
not ( n24611 , n21549 );
not ( n24612 , n24603 );
or ( n24613 , n24611 , n24612 );
and ( n24614 , n23976 , n23749 );
not ( n24615 , n23976 );
and ( n24616 , n24615 , n23750 );
or ( n24617 , n24614 , n24616 );
not ( n24618 , n24617 );
nand ( n24619 , n24618 , n19316 );
nand ( n24620 , n24613 , n24619 );
xor ( n24621 , n24610 , n24620 );
xor ( n24622 , n24322 , n24330 );
and ( n24623 , n23976 , n23941 );
not ( n24624 , n23976 );
and ( n24625 , n24624 , n23942 );
nor ( n24626 , n24623 , n24625 );
not ( n24627 , n24626 );
or ( n24628 , n24627 , n22573 );
or ( n24629 , n24617 , n22864 );
nand ( n24630 , n24628 , n24629 );
xor ( n24631 , n24622 , n24630 );
and ( n24632 , n21577 , n24015 );
and ( n24633 , n19283 , n24015 );
nor ( n24634 , n24633 , n19318 );
or ( n24635 , n19283 , n24015 );
nand ( n24636 , n24635 , n21651 );
and ( n24637 , n24634 , n24636 );
not ( n24638 , n21549 );
and ( n24639 , n19311 , n24001 );
not ( n24640 , n19311 );
and ( n24641 , n24640 , n24002 );
nor ( n24642 , n24639 , n24641 );
not ( n24643 , n24642 );
or ( n24644 , n24638 , n24643 );
and ( n24645 , n19318 , n24015 );
and ( n24646 , n19311 , n24016 );
nor ( n24647 , n24645 , n24646 );
not ( n24648 , n24647 );
nand ( n24649 , n24648 , n19316 );
nand ( n24650 , n24644 , n24649 );
and ( n24651 , n24637 , n24650 );
xor ( n24652 , n24632 , n24651 );
not ( n24653 , n21549 );
not ( n24654 , n24626 );
or ( n24655 , n24653 , n24654 );
nand ( n24656 , n24642 , n19316 );
nand ( n24657 , n24655 , n24656 );
and ( n24658 , n24652 , n24657 );
or ( n24660 , n24658 , C0 );
and ( n24661 , n24631 , n24660 );
and ( n24662 , n24622 , n24630 );
or ( n24663 , n24661 , n24662 );
and ( n24664 , n24621 , n24663 );
and ( n24665 , n24610 , n24620 );
or ( n24666 , n24664 , n24665 );
nand ( n24667 , n24608 , n24666 );
nand ( n24668 , n24607 , n24667 );
xor ( n24669 , n24518 , n24520 );
xor ( n24670 , n24669 , n24531 );
xor ( n24671 , n24668 , n24670 );
not ( n24672 , n22166 );
not ( n24673 , n22137 );
not ( n24674 , n22892 );
or ( n24675 , n24673 , n24674 );
nand ( n24676 , n23027 , n22136 );
nand ( n24677 , n24675 , n24676 );
not ( n24678 , n24677 );
or ( n24679 , n24672 , n24678 );
nand ( n24680 , n24542 , n22134 );
nand ( n24681 , n24679 , n24680 );
and ( n24682 , n24671 , n24681 );
and ( n24683 , n24668 , n24670 );
or ( n24684 , n24682 , n24683 );
not ( n24685 , n22062 );
not ( n24686 , n24479 );
or ( n24687 , n24685 , n24686 );
not ( n24688 , n22071 );
not ( n24689 , n22612 );
or ( n24690 , n24688 , n24689 );
nand ( n24691 , n22611 , n22070 );
nand ( n24692 , n24690 , n24691 );
nand ( n24693 , n24692 , n22121 );
nand ( n24694 , n24687 , n24693 );
xor ( n24695 , n24684 , n24694 );
not ( n24696 , n22051 );
and ( n24697 , n21853 , n22417 );
not ( n24698 , n21853 );
and ( n24699 , n24698 , n22418 );
nor ( n24700 , n24697 , n24699 );
not ( n24701 , n24700 );
or ( n24702 , n24696 , n24701 );
nand ( n24703 , n24505 , n21846 );
nand ( n24704 , n24702 , n24703 );
and ( n24705 , n24695 , n24704 );
and ( n24706 , n24684 , n24694 );
or ( n24707 , n24705 , n24706 );
and ( n24708 , n24593 , n24707 );
and ( n24709 , n24590 , n24592 );
or ( n24710 , n24708 , n24709 );
not ( n24711 , n24710 );
and ( n24712 , n24484 , n24427 );
not ( n24713 , n24484 );
and ( n24714 , n24713 , n24428 );
or ( n24715 , n24712 , n24714 );
not ( n24716 , n24438 );
and ( n24717 , n24715 , n24716 );
not ( n24718 , n24715 );
and ( n24719 , n24718 , n24438 );
nor ( n24720 , n24717 , n24719 );
nand ( n24721 , n24711 , n24720 );
and ( n24722 , n24580 , n24721 );
not ( n24723 , n24710 );
nor ( n24724 , n24723 , n24720 );
nor ( n24725 , n24722 , n24724 );
nand ( n24726 , n24578 , n24725 );
and ( n24727 , n24576 , n24726 );
not ( n24728 , n24727 );
xor ( n24729 , n24498 , n24507 );
xor ( n24730 , n24729 , n24550 );
not ( n24731 , n24730 );
not ( n24732 , n24731 );
xor ( n24733 , n24534 , n24544 );
xor ( n24734 , n24733 , n24547 );
not ( n24735 , n22062 );
not ( n24736 , n24692 );
or ( n24737 , n24735 , n24736 );
not ( n24738 , n22071 );
not ( n24739 , n22736 );
or ( n24740 , n24738 , n24739 );
nand ( n24741 , n22737 , n22070 );
nand ( n24742 , n24740 , n24741 );
nand ( n24743 , n24742 , n22121 );
nand ( n24744 , n24737 , n24743 );
not ( n24745 , n24744 );
not ( n24746 , n24528 );
not ( n24747 , n22877 );
and ( n24748 , n24746 , n24747 );
and ( n24749 , n21651 , n23650 );
not ( n24750 , n21651 );
and ( n24751 , n24750 , n23395 );
nor ( n24752 , n24749 , n24751 );
and ( n24753 , n24752 , n21698 );
nor ( n24754 , n24748 , n24753 );
xor ( n24755 , n24605 , n24595 );
xnor ( n24756 , n24755 , n24666 );
xor ( n24757 , n24754 , n24756 );
and ( n24758 , n24677 , n22134 );
and ( n24759 , n24538 , n23056 );
not ( n24760 , n24538 );
and ( n24761 , n24760 , n23055 );
or ( n24762 , n24759 , n24761 );
and ( n24763 , n24762 , n22166 );
nor ( n24764 , n24758 , n24763 );
and ( n24765 , n24757 , n24764 );
and ( n24766 , n24754 , n24756 );
or ( n24767 , n24765 , n24766 );
nand ( n24768 , n24745 , n24767 );
not ( n24769 , n24768 );
xor ( n24770 , n24668 , n24670 );
xor ( n24771 , n24770 , n24681 );
not ( n24772 , n24771 );
or ( n24773 , n24769 , n24772 );
not ( n24774 , n24767 );
nand ( n24775 , n24744 , n24774 );
nand ( n24776 , n24773 , n24775 );
xor ( n24777 , n24734 , n24776 );
and ( n24778 , n22178 , n22231 );
not ( n24779 , n22178 );
and ( n24780 , n24779 , n22426 );
nor ( n24781 , n24778 , n24780 );
not ( n24782 , n24781 );
not ( n24783 , n22645 );
or ( n24784 , n24782 , n24783 );
not ( n24785 , n24588 );
or ( n24786 , n24785 , n22643 );
nand ( n24787 , n24784 , n24786 );
and ( n24788 , n24777 , n24787 );
and ( n24789 , n24734 , n24776 );
or ( n24790 , n24788 , n24789 );
not ( n24791 , n24790 );
not ( n24792 , n24791 );
or ( n24793 , n24732 , n24792 );
xor ( n24794 , n24590 , n24592 );
xor ( n24795 , n24794 , n24707 );
nand ( n24796 , n24793 , n24795 );
nand ( n24797 , n24790 , n24730 );
nand ( n24798 , n24796 , n24797 );
not ( n24799 , n24720 );
not ( n24800 , n24710 );
and ( n24801 , n24799 , n24800 );
and ( n24802 , n24720 , n24710 );
nor ( n24803 , n24801 , n24802 );
xnor ( n24804 , n24580 , n24803 );
xor ( n24805 , n24798 , n24804 );
not ( n24806 , n21698 );
and ( n24807 , n21651 , n23536 );
not ( n24808 , n21651 );
and ( n24809 , n24808 , n23537 );
nor ( n24810 , n24807 , n24809 );
not ( n24811 , n24810 );
or ( n24812 , n24806 , n24811 );
nand ( n24813 , n24752 , n21837 );
nand ( n24814 , n24812 , n24813 );
xor ( n24815 , n24610 , n24620 );
xor ( n24816 , n24815 , n24663 );
xor ( n24817 , n24814 , n24816 );
not ( n24818 , n22134 );
not ( n24819 , n24762 );
or ( n24820 , n24818 , n24819 );
and ( n24821 , n24538 , n23046 );
not ( n24822 , n24538 );
and ( n24823 , n24822 , n23045 );
nor ( n24824 , n24821 , n24823 );
nand ( n24825 , n24824 , n22166 );
nand ( n24826 , n24820 , n24825 );
and ( n24827 , n24817 , n24826 );
and ( n24828 , n24814 , n24816 );
or ( n24829 , n24827 , n24828 );
not ( n24830 , n22062 );
not ( n24831 , n24742 );
or ( n24832 , n24830 , n24831 );
and ( n24833 , n22071 , n22884 );
not ( n24834 , n22071 );
and ( n24835 , n24834 , n22926 );
or ( n24836 , n24833 , n24835 );
not ( n24837 , n24836 );
nand ( n24838 , n24837 , n22121 );
nand ( n24839 , n24832 , n24838 );
xor ( n24840 , n24829 , n24839 );
not ( n24841 , n21846 );
not ( n24842 , n21853 );
not ( n24843 , n22742 );
or ( n24844 , n24842 , n24843 );
nand ( n24845 , n22535 , n21852 );
nand ( n24846 , n24844 , n24845 );
not ( n24847 , n24846 );
or ( n24848 , n24841 , n24847 );
and ( n24849 , n21853 , n22612 );
not ( n24850 , n21853 );
and ( n24851 , n24850 , n22611 );
or ( n24852 , n24849 , n24851 );
nand ( n24853 , n24852 , n22050 );
nand ( n24854 , n24848 , n24853 );
xor ( n24855 , n24840 , n24854 );
not ( n24856 , n21846 );
not ( n24857 , n24852 );
or ( n24858 , n24856 , n24857 );
not ( n24859 , n21853 );
not ( n24860 , n22736 );
or ( n24861 , n24859 , n24860 );
nand ( n24862 , n22735 , n21852 );
nand ( n24863 , n24861 , n24862 );
nand ( n24864 , n24863 , n22050 );
nand ( n24865 , n24858 , n24864 );
not ( n24866 , n22166 );
and ( n24867 , n24538 , n23650 );
not ( n24868 , n24538 );
and ( n24869 , n24868 , n23653 );
nor ( n24870 , n24867 , n24869 );
not ( n24871 , n24870 );
or ( n24872 , n24866 , n24871 );
nand ( n24873 , n24824 , n22134 );
nand ( n24874 , n24872 , n24873 );
xor ( n24875 , n24622 , n24630 );
xor ( n24876 , n24875 , n24660 );
not ( n24877 , n21837 );
not ( n24878 , n24810 );
or ( n24879 , n24877 , n24878 );
and ( n24880 , n21651 , n23644 );
not ( n24881 , n21651 );
and ( n24882 , n24881 , n23646 );
nor ( n24883 , n24880 , n24882 );
not ( n24884 , n24883 );
or ( n24885 , n24884 , n22871 );
nand ( n24886 , n24879 , n24885 );
xor ( n24887 , n24876 , n24886 );
xor ( n24888 , n24632 , n24651 );
xor ( n24889 , n24888 , n24657 );
not ( n24890 , n21837 );
not ( n24891 , n24883 );
or ( n24892 , n24890 , n24891 );
and ( n24893 , n21651 , n23749 );
not ( n24894 , n21651 );
and ( n24895 , n24894 , n23750 );
nor ( n24896 , n24893 , n24895 );
nand ( n24897 , n24896 , n21698 );
nand ( n24898 , n24892 , n24897 );
xor ( n24899 , n24889 , n24898 );
xor ( n24900 , n24637 , n24650 );
not ( n24901 , n21837 );
not ( n24902 , n24896 );
or ( n24903 , n24901 , n24902 );
and ( n24904 , n21651 , n24025 );
not ( n24905 , n21651 );
and ( n24906 , n24905 , n23942 );
nor ( n24907 , n24904 , n24906 );
nand ( n24908 , n24907 , n21698 );
nand ( n24909 , n24903 , n24908 );
xor ( n24910 , n24900 , n24909 );
and ( n24911 , n21549 , n24015 );
not ( n24912 , n21837 );
not ( n24913 , n24907 );
or ( n24914 , n24912 , n24913 );
and ( n24915 , n21651 , n24001 );
not ( n24916 , n21651 );
and ( n24917 , n24916 , n24002 );
nor ( n24918 , n24915 , n24917 );
nand ( n24919 , n24918 , n21698 );
nand ( n24920 , n24914 , n24919 );
xor ( n24921 , n24911 , n24920 );
or ( n24922 , n24015 , n21658 );
nand ( n24923 , n24922 , n24538 );
nand ( n24924 , n24015 , n21658 );
and ( n24925 , n24923 , n21651 , n24924 );
not ( n24926 , n21837 );
not ( n24927 , n24918 );
or ( n24928 , n24926 , n24927 );
or ( n24929 , n21651 , n24016 );
or ( n24930 , n21650 , n24015 );
nand ( n24931 , n24929 , n24930 );
nand ( n24932 , n21697 , n24931 );
nand ( n24933 , n24928 , n24932 );
and ( n24934 , n24925 , n24933 );
and ( n24935 , n24921 , n24934 );
and ( n24936 , n24911 , n24920 );
or ( n24937 , n24935 , n24936 );
and ( n24938 , n24910 , n24937 );
and ( n24939 , n24900 , n24909 );
or ( n24940 , n24938 , n24939 );
and ( n24941 , n24899 , n24940 );
and ( n24942 , n24889 , n24898 );
or ( n24943 , n24941 , n24942 );
xor ( n24944 , n24887 , n24943 );
xor ( n24945 , n24874 , n24944 );
not ( n24946 , n22121 );
and ( n24947 , n22071 , n23055 );
not ( n24948 , n22071 );
and ( n24949 , n24948 , n23056 );
nor ( n24950 , n24947 , n24949 );
not ( n24951 , n24950 );
or ( n24952 , n24946 , n24951 );
not ( n24953 , n22071 );
not ( n24954 , n22892 );
or ( n24955 , n24953 , n24954 );
nand ( n24956 , n23027 , n22070 );
nand ( n24957 , n24955 , n24956 );
nand ( n24958 , n24957 , n22062 );
nand ( n24959 , n24952 , n24958 );
and ( n24960 , n24945 , n24959 );
and ( n24961 , n24874 , n24944 );
or ( n24962 , n24960 , n24961 );
xor ( n24963 , n24865 , n24962 );
and ( n24964 , n22179 , n22418 );
not ( n24965 , n22179 );
and ( n24966 , n24965 , n22417 );
nor ( n24967 , n24964 , n24966 );
not ( n24968 , n24967 );
not ( n24969 , n22642 );
or ( n24970 , n24968 , n24969 );
and ( n24971 , n22178 , n22535 );
not ( n24972 , n22178 );
and ( n24973 , n24972 , n22742 );
nor ( n24974 , n24971 , n24973 );
nand ( n24975 , n24974 , n22645 );
nand ( n24976 , n24970 , n24975 );
and ( n24977 , n24963 , n24976 );
and ( n24978 , n24865 , n24962 );
or ( n24979 , n24977 , n24978 );
xor ( n24980 , n24855 , n24979 );
xor ( n24981 , n24876 , n24886 );
and ( n24982 , n24981 , n24943 );
and ( n24983 , n24876 , n24886 );
or ( n24984 , n24982 , n24983 );
not ( n24985 , n24957 );
not ( n24986 , n22121 );
or ( n24987 , n24985 , n24986 );
or ( n24988 , n24836 , n22061 );
nand ( n24989 , n24987 , n24988 );
xor ( n24990 , n24984 , n24989 );
xor ( n24991 , n24814 , n24816 );
xor ( n24992 , n24991 , n24826 );
and ( n24993 , n24990 , n24992 );
and ( n24994 , n24984 , n24989 );
or ( n24995 , n24993 , n24994 );
not ( n24996 , n24995 );
xor ( n24997 , n24754 , n24756 );
xor ( n24998 , n24997 , n24764 );
not ( n24999 , n24998 );
and ( n25000 , n24996 , n24999 );
and ( n25001 , n24995 , n24998 );
nor ( n25002 , n25000 , n25001 );
and ( n25003 , n22178 , n22241 );
not ( n25004 , n22178 );
and ( n25005 , n25004 , n22544 );
nor ( n25006 , n25003 , n25005 );
not ( n25007 , n25006 );
not ( n25008 , n22642 );
or ( n25009 , n25007 , n25008 );
nand ( n25010 , n24967 , n22645 );
nand ( n25011 , n25009 , n25010 );
not ( n25012 , n25011 );
and ( n25013 , n25002 , n25012 );
not ( n25014 , n25002 );
and ( n25015 , n25014 , n25011 );
nor ( n25016 , n25013 , n25015 );
and ( n25017 , n24980 , n25016 );
and ( n25018 , n24855 , n24979 );
or ( n25019 , n25017 , n25018 );
not ( n25020 , n25019 );
and ( n25021 , n24744 , n24774 );
not ( n25022 , n24744 );
and ( n25023 , n25022 , n24767 );
nor ( n25024 , n25021 , n25023 );
xnor ( n25025 , n25024 , n24771 );
not ( n25026 , n24998 );
not ( n25027 , n25012 );
or ( n25028 , n25026 , n25027 );
nand ( n25029 , n25028 , n24995 );
not ( n25030 , n24998 );
nand ( n25031 , n25030 , n25011 );
and ( n25032 , n25029 , n25031 );
xor ( n25033 , n25025 , n25032 );
not ( n25034 , n21846 );
not ( n25035 , n24700 );
or ( n25036 , n25034 , n25035 );
nand ( n25037 , n24846 , n22051 );
nand ( n25038 , n25036 , n25037 );
not ( n25039 , n22642 );
not ( n25040 , n24781 );
or ( n25041 , n25039 , n25040 );
nand ( n25042 , n25006 , n22645 );
nand ( n25043 , n25041 , n25042 );
xor ( n25044 , n25038 , n25043 );
xor ( n25045 , n24829 , n24839 );
and ( n25046 , n25045 , n24854 );
and ( n25047 , n24829 , n24839 );
or ( n25048 , n25046 , n25047 );
xnor ( n25049 , n25044 , n25048 );
xor ( n25050 , n25033 , n25049 );
nand ( n25051 , n25020 , n25050 );
not ( n25052 , n25051 );
xor ( n25053 , n24984 , n24989 );
xor ( n25054 , n25053 , n24992 );
not ( n25055 , n21846 );
not ( n25056 , n24863 );
or ( n25057 , n25055 , n25056 );
and ( n25058 , n22883 , n21852 );
not ( n25059 , n22883 );
and ( n25060 , n25059 , n21851 );
or ( n25061 , n25058 , n25060 );
nand ( n25062 , n25061 , n22050 );
nand ( n25063 , n25057 , n25062 );
not ( n25064 , n22134 );
not ( n25065 , n24870 );
or ( n25066 , n25064 , n25065 );
and ( n25067 , n24538 , n23536 );
not ( n25068 , n24538 );
and ( n25069 , n25068 , n23537 );
nor ( n25070 , n25067 , n25069 );
nand ( n25071 , n25070 , n22165 );
nand ( n25072 , n25066 , n25071 );
xor ( n25073 , n24889 , n24898 );
xor ( n25074 , n25073 , n24940 );
xor ( n25075 , n25072 , n25074 );
not ( n25076 , n22062 );
not ( n25077 , n24950 );
or ( n25078 , n25076 , n25077 );
not ( n25079 , n22071 );
not ( n25080 , n23045 );
or ( n25081 , n25079 , n25080 );
nand ( n25082 , n23046 , n22070 );
nand ( n25083 , n25081 , n25082 );
nand ( n25084 , n25083 , n22121 );
nand ( n25085 , n25078 , n25084 );
and ( n25086 , n25075 , n25085 );
and ( n25087 , n25072 , n25074 );
or ( n25088 , n25086 , n25087 );
xor ( n25089 , n25063 , n25088 );
not ( n25090 , n21846 );
not ( n25091 , n25061 );
or ( n25092 , n25090 , n25091 );
and ( n25093 , n22891 , n21852 );
not ( n25094 , n22891 );
and ( n25095 , n25094 , n21851 );
or ( n25096 , n25093 , n25095 );
nand ( n25097 , n25096 , n22050 );
nand ( n25098 , n25092 , n25097 );
not ( n25099 , n25098 );
xor ( n25100 , n24900 , n24909 );
xor ( n25101 , n25100 , n24937 );
not ( n25102 , n22134 );
not ( n25103 , n25070 );
or ( n25104 , n25102 , n25103 );
not ( n25105 , n24538 );
not ( n25106 , n23951 );
or ( n25107 , n25105 , n25106 );
nand ( n25108 , n23645 , n22136 );
nand ( n25109 , n25107 , n25108 );
nand ( n25110 , n25109 , n22165 );
nand ( n25111 , n25104 , n25110 );
xor ( n25112 , n25101 , n25111 );
xor ( n25113 , n24911 , n24920 );
xor ( n25114 , n25113 , n24934 );
not ( n25115 , n22134 );
not ( n25116 , n25109 );
or ( n25117 , n25115 , n25116 );
xor ( n25118 , n21692 , n23740 );
xor ( n25119 , n25118 , n23746 );
nand ( n25120 , n25119 , n22165 );
nand ( n25121 , n25117 , n25120 );
xor ( n25122 , n25114 , n25121 );
xor ( n25123 , n24925 , n24933 );
not ( n25124 , n22134 );
not ( n25125 , n25119 );
or ( n25126 , n25124 , n25125 );
and ( n25127 , n24538 , n23941 );
not ( n25128 , n24538 );
and ( n25129 , n25128 , n23942 );
nor ( n25130 , n25127 , n25129 );
nand ( n25131 , n25130 , n22165 );
nand ( n25132 , n25126 , n25131 );
xor ( n25133 , n25123 , n25132 );
and ( n25134 , n21837 , n24015 );
not ( n25135 , n22134 );
not ( n25136 , n25130 );
or ( n25137 , n25135 , n25136 );
and ( n25138 , n22162 , n24000 );
not ( n25139 , n22162 );
and ( n25140 , n25139 , n24001 );
or ( n25141 , n25138 , n25140 );
nand ( n25142 , n25141 , n22165 );
nand ( n25143 , n25137 , n25142 );
xor ( n25144 , n25134 , n25143 );
not ( n25145 , n22133 );
not ( n25146 , n25141 );
or ( n25147 , n25145 , n25146 );
not ( n25148 , n22162 );
not ( n25149 , n20935 );
or ( n25150 , n25148 , n25149 );
or ( n25151 , n24016 , n24538 );
nand ( n25152 , n25150 , n25151 );
nand ( n25153 , n22165 , n25152 );
nand ( n25154 , n25147 , n25153 );
or ( n25155 , n22132 , n24015 );
nand ( n25156 , n25155 , n22069 );
nand ( n25157 , n22132 , n24015 );
and ( n25158 , n25156 , n22162 , n25157 );
and ( n25159 , n25154 , n25158 );
and ( n25160 , n25144 , n25159 );
and ( n25161 , n25134 , n25143 );
or ( n25162 , n25160 , n25161 );
and ( n25163 , n25133 , n25162 );
and ( n25164 , n25123 , n25132 );
or ( n25165 , n25163 , n25164 );
and ( n25166 , n25122 , n25165 );
and ( n25167 , n25114 , n25121 );
or ( n25168 , n25166 , n25167 );
and ( n25169 , n25112 , n25168 );
and ( n25170 , n25101 , n25111 );
or ( n25171 , n25169 , n25170 );
not ( n25172 , n25171 );
nand ( n25173 , n25099 , n25172 );
not ( n25174 , n25173 );
xor ( n25175 , n25072 , n25074 );
xor ( n25176 , n25175 , n25085 );
not ( n25177 , n25176 );
or ( n25178 , n25174 , n25177 );
nand ( n25179 , n25098 , n25171 );
nand ( n25180 , n25178 , n25179 );
and ( n25181 , n25089 , n25180 );
and ( n25182 , n25063 , n25088 );
or ( n25183 , n25181 , n25182 );
xor ( n25184 , n25054 , n25183 );
xor ( n25185 , n24865 , n24962 );
xor ( n25186 , n25185 , n24976 );
and ( n25187 , n25184 , n25186 );
and ( n25188 , n25054 , n25183 );
or ( n25189 , n25187 , n25188 );
xor ( n25190 , n24855 , n24979 );
xor ( n25191 , n25190 , n25016 );
xor ( n25192 , n25189 , n25191 );
xor ( n25193 , n24874 , n24944 );
xor ( n25194 , n25193 , n24959 );
not ( n25195 , n22642 );
not ( n25196 , n24974 );
or ( n25197 , n25195 , n25196 );
and ( n25198 , n22610 , n22179 );
not ( n25199 , n22610 );
and ( n25200 , n25199 , n22178 );
or ( n25201 , n25198 , n25200 );
nand ( n25202 , n25201 , n22645 );
nand ( n25203 , n25197 , n25202 );
xor ( n25204 , n25194 , n25203 );
xor ( n25205 , n25063 , n25088 );
xor ( n25206 , n25205 , n25180 );
and ( n25207 , n25204 , n25206 );
and ( n25208 , n25194 , n25203 );
or ( n25209 , n25207 , n25208 );
xor ( n25210 , n25054 , n25183 );
xor ( n25211 , n25210 , n25186 );
xor ( n25212 , n25209 , n25211 );
xor ( n25213 , n25098 , n25172 );
xor ( n25214 , n25213 , n25176 );
and ( n25215 , n23394 , n22070 );
not ( n25216 , n23394 );
not ( n25217 , n22070 );
and ( n25218 , n25216 , n25217 );
or ( n25219 , n25215 , n25218 );
not ( n25220 , n25219 );
not ( n25221 , n22121 );
or ( n25222 , n25220 , n25221 );
not ( n25223 , n25083 );
or ( n25224 , n25223 , n22061 );
nand ( n25225 , n25222 , n25224 );
not ( n25226 , n25225 );
and ( n25227 , n25096 , n21846 );
and ( n25228 , n23055 , n21852 );
not ( n25229 , n23055 );
and ( n25230 , n25229 , n21851 );
or ( n25231 , n25228 , n25230 );
not ( n25232 , n25231 );
nor ( n25233 , n25232 , n22049 );
nor ( n25234 , n25227 , n25233 );
nand ( n25235 , n25226 , n25234 );
xor ( n25236 , n25101 , n25111 );
xor ( n25237 , n25236 , n25168 );
and ( n25238 , n25235 , n25237 );
not ( n25239 , n25225 );
nor ( n25240 , n25239 , n25234 );
nor ( n25241 , n25238 , n25240 );
and ( n25242 , n25201 , n22642 );
and ( n25243 , n22735 , n22179 );
not ( n25244 , n22735 );
and ( n25245 , n25244 , n22178 );
or ( n25246 , n25243 , n25245 );
not ( n25247 , n25246 );
nor ( n25248 , n25247 , n22644 );
nor ( n25249 , n25242 , n25248 );
and ( n25250 , n25241 , n25249 );
or ( n25251 , n25214 , n25250 );
or ( n25252 , n25249 , n25241 );
nand ( n25253 , n25251 , n25252 );
xor ( n25254 , n25194 , n25203 );
xor ( n25255 , n25254 , n25206 );
xor ( n25256 , n25253 , n25255 );
xor ( n25257 , n25234 , n25237 );
xnor ( n25258 , n25257 , n25225 );
not ( n25259 , n25258 );
not ( n25260 , n22642 );
not ( n25261 , n25246 );
or ( n25262 , n25260 , n25261 );
and ( n25263 , n22883 , n22179 );
not ( n25264 , n22883 );
and ( n25265 , n25264 , n22178 );
or ( n25266 , n25263 , n25265 );
nand ( n25267 , n25266 , n22645 );
nand ( n25268 , n25262 , n25267 );
not ( n25269 , n22062 );
not ( n25270 , n25219 );
or ( n25271 , n25269 , n25270 );
xor ( n25272 , n25217 , n23536 );
nand ( n25273 , n25272 , n22121 );
nand ( n25274 , n25271 , n25273 );
xor ( n25275 , n25114 , n25121 );
xor ( n25276 , n25275 , n25165 );
xor ( n25277 , n25274 , n25276 );
not ( n25278 , n22050 );
not ( n25279 , n21851 );
not ( n25280 , n23045 );
or ( n25281 , n25279 , n25280 );
nand ( n25282 , n23044 , n21852 );
nand ( n25283 , n25281 , n25282 );
not ( n25284 , n25283 );
or ( n25285 , n25278 , n25284 );
nand ( n25286 , n25231 , n21846 );
nand ( n25287 , n25285 , n25286 );
and ( n25288 , n25277 , n25287 );
and ( n25289 , n25274 , n25276 );
or ( n25290 , n25288 , n25289 );
not ( n25291 , n25290 );
and ( n25292 , n25268 , n25291 );
not ( n25293 , n25268 );
and ( n25294 , n25293 , n25290 );
nor ( n25295 , n25292 , n25294 );
not ( n25296 , n25295 );
xor ( n25297 , n25123 , n25132 );
xor ( n25298 , n25297 , n25162 );
not ( n25299 , n22062 );
not ( n25300 , n25272 );
or ( n25301 , n25299 , n25300 );
and ( n25302 , n23644 , n22070 );
not ( n25303 , n23644 );
and ( n25304 , n25303 , n25217 );
or ( n25305 , n25302 , n25304 );
nand ( n25306 , n25305 , n22121 );
nand ( n25307 , n25301 , n25306 );
xor ( n25308 , n25298 , n25307 );
xor ( n25309 , n25134 , n25143 );
xor ( n25310 , n25309 , n25159 );
not ( n25311 , n22062 );
not ( n25312 , n25305 );
or ( n25313 , n25311 , n25312 );
not ( n25314 , n25217 );
not ( n25315 , n23748 );
not ( n25316 , n25315 );
or ( n25317 , n25314 , n25316 );
nand ( n25318 , n23749 , n22070 );
nand ( n25319 , n25317 , n25318 );
nand ( n25320 , n25319 , n22121 );
nand ( n25321 , n25313 , n25320 );
xor ( n25322 , n25310 , n25321 );
not ( n25323 , n25158 );
not ( n25324 , n25154 );
or ( n25325 , n25323 , n25324 );
or ( n25326 , n25154 , n25158 );
nand ( n25327 , n25325 , n25326 );
not ( n25328 , n25327 );
not ( n25329 , n25328 );
not ( n25330 , n22062 );
not ( n25331 , n25319 );
or ( n25332 , n25330 , n25331 );
not ( n25333 , n25217 );
not ( n25334 , n23942 );
or ( n25335 , n25333 , n25334 );
nand ( n25336 , n23941 , n22070 );
nand ( n25337 , n25335 , n25336 );
nand ( n25338 , n25337 , n22120 );
nand ( n25339 , n25332 , n25338 );
not ( n25340 , n25339 );
or ( n25341 , n25329 , n25340 );
not ( n25342 , n25339 );
nand ( n25343 , n25342 , n25327 );
nand ( n25344 , n22133 , n24015 );
not ( n25345 , n25344 );
not ( n25346 , n25345 );
not ( n25347 , n22062 );
not ( n25348 , n25337 );
or ( n25349 , n25347 , n25348 );
not ( n25350 , n25217 );
not ( n25351 , n24000 );
or ( n25352 , n25350 , n25351 );
nand ( n25353 , n24001 , n22070 );
nand ( n25354 , n25352 , n25353 );
nand ( n25355 , n25354 , n22120 );
nand ( n25356 , n25349 , n25355 );
not ( n25357 , n25356 );
or ( n25358 , n25346 , n25357 );
not ( n25359 , n25344 );
not ( n25360 , n25356 );
not ( n25361 , n25360 );
or ( n25362 , n25359 , n25361 );
not ( n25363 , n22062 );
not ( n25364 , n25354 );
or ( n25365 , n25363 , n25364 );
or ( n25366 , n25217 , n24016 );
or ( n25367 , n22070 , n24015 );
nand ( n25368 , n25366 , n25367 );
nand ( n25369 , n22120 , n25368 );
nand ( n25370 , n25365 , n25369 );
or ( n25371 , n22056 , n24015 );
nand ( n25372 , n25371 , n21851 );
nand ( n25373 , n22056 , n24015 );
and ( n25374 , n25217 , n25372 , n25373 );
and ( n25375 , n25370 , n25374 );
nand ( n25376 , n25362 , n25375 );
nand ( n25377 , n25358 , n25376 );
nand ( n25378 , n25343 , n25377 );
nand ( n25379 , n25341 , n25378 );
and ( n25380 , n25322 , n25379 );
and ( n25381 , n25310 , n25321 );
or ( n25382 , n25380 , n25381 );
and ( n25383 , n25308 , n25382 );
and ( n25384 , n25298 , n25307 );
or ( n25385 , n25383 , n25384 );
not ( n25386 , n22642 );
not ( n25387 , n25266 );
or ( n25388 , n25386 , n25387 );
and ( n25389 , n22891 , n22179 );
not ( n25390 , n22891 );
and ( n25391 , n25390 , n22178 );
or ( n25392 , n25389 , n25391 );
nand ( n25393 , n25392 , n22645 );
nand ( n25394 , n25388 , n25393 );
xor ( n25395 , n25385 , n25394 );
xor ( n25396 , n25274 , n25276 );
xor ( n25397 , n25396 , n25287 );
and ( n25398 , n25395 , n25397 );
and ( n25399 , n25385 , n25394 );
or ( n25400 , n25398 , n25399 );
not ( n25401 , n25400 );
and ( n25402 , n25296 , n25401 );
and ( n25403 , n25400 , n25295 );
nor ( n25404 , n25402 , n25403 );
nand ( n25405 , n25259 , n25404 );
and ( n25406 , n25283 , n21846 );
xor ( n25407 , n21851 , n23394 );
not ( n25408 , n25407 );
nor ( n25409 , n25408 , n22049 );
nor ( n25410 , n25406 , n25409 );
not ( n25411 , n25410 );
not ( n25412 , n22642 );
not ( n25413 , n25392 );
or ( n25414 , n25412 , n25413 );
xor ( n25415 , n22178 , n23055 );
nand ( n25416 , n25415 , n22645 );
nand ( n25417 , n25414 , n25416 );
not ( n25418 , n25417 );
not ( n25419 , n25418 );
or ( n25420 , n25411 , n25419 );
xor ( n25421 , n25298 , n25307 );
xor ( n25422 , n25421 , n25382 );
nand ( n25423 , n25420 , n25422 );
not ( n25424 , n25410 );
nand ( n25425 , n25424 , n25417 );
nand ( n25426 , n25423 , n25425 );
xor ( n25427 , n25385 , n25394 );
xor ( n25428 , n25427 , n25397 );
xor ( n25429 , n25426 , n25428 );
not ( n25430 , n21846 );
not ( n25431 , n25407 );
or ( n25432 , n25430 , n25431 );
and ( n25433 , n23536 , n21852 );
not ( n25434 , n23536 );
and ( n25435 , n25434 , n21851 );
or ( n25436 , n25433 , n25435 );
nand ( n25437 , n25436 , n22050 );
nand ( n25438 , n25432 , n25437 );
xor ( n25439 , n25310 , n25321 );
xor ( n25440 , n25439 , n25379 );
xor ( n25441 , n25438 , n25440 );
not ( n25442 , n22645 );
and ( n25443 , n23044 , n22179 );
not ( n25444 , n23044 );
and ( n25445 , n25444 , n22178 );
or ( n25446 , n25443 , n25445 );
not ( n25447 , n25446 );
or ( n25448 , n25442 , n25447 );
nand ( n25449 , n25415 , n22642 );
nand ( n25450 , n25448 , n25449 );
and ( n25451 , n25441 , n25450 );
and ( n25452 , n25438 , n25440 );
or ( n25453 , n25451 , n25452 );
not ( n25454 , n25453 );
not ( n25455 , n25410 );
not ( n25456 , n25422 );
or ( n25457 , n25455 , n25456 );
or ( n25458 , n25422 , n25410 );
nand ( n25459 , n25457 , n25458 );
not ( n25460 , n25459 );
not ( n25461 , n25418 );
and ( n25462 , n25460 , n25461 );
and ( n25463 , n25459 , n25418 );
nor ( n25464 , n25462 , n25463 );
nand ( n25465 , n25454 , n25464 );
not ( n25466 , n25465 );
not ( n25467 , n25328 );
not ( n25468 , n25342 );
or ( n25469 , n25467 , n25468 );
nand ( n25470 , n25339 , n25327 );
nand ( n25471 , n25469 , n25470 );
xnor ( n25472 , n25471 , n25377 );
not ( n25473 , n25472 );
not ( n25474 , n25473 );
not ( n25475 , n21846 );
not ( n25476 , n25436 );
or ( n25477 , n25475 , n25476 );
and ( n25478 , n23644 , n22046 );
not ( n25479 , n23644 );
and ( n25480 , n25479 , n21851 );
or ( n25481 , n25478 , n25480 );
nand ( n25482 , n25481 , n22050 );
nand ( n25483 , n25477 , n25482 );
not ( n25484 , n25483 );
or ( n25485 , n25474 , n25484 );
not ( n25486 , n25345 );
not ( n25487 , n25360 );
or ( n25488 , n25486 , n25487 );
nand ( n25489 , n25356 , n25344 );
nand ( n25490 , n25488 , n25489 );
xnor ( n25491 , n25490 , n25375 );
not ( n25492 , n25491 );
not ( n25493 , n21846 );
not ( n25494 , n25481 );
or ( n25495 , n25493 , n25494 );
not ( n25496 , n21851 );
not ( n25497 , n25315 );
or ( n25498 , n25496 , n25497 );
nand ( n25499 , n23749 , n22046 );
nand ( n25500 , n25498 , n25499 );
nand ( n25501 , n25500 , n22050 );
nand ( n25502 , n25495 , n25501 );
not ( n25503 , n25502 );
not ( n25504 , n25503 );
or ( n25505 , n25492 , n25504 );
xor ( n25506 , n25374 , n25370 );
not ( n25507 , n21846 );
not ( n25508 , n25500 );
or ( n25509 , n25507 , n25508 );
not ( n25510 , n21851 );
not ( n25511 , n23942 );
or ( n25512 , n25510 , n25511 );
nand ( n25513 , n24025 , n22046 );
nand ( n25514 , n25512 , n25513 );
nand ( n25515 , n25514 , n22050 );
nand ( n25516 , n25509 , n25515 );
xor ( n25517 , n25506 , n25516 );
nor ( n25518 , n22061 , n24016 );
or ( n25519 , n24015 , n21842 );
nand ( n25520 , n25519 , n22178 );
nand ( n25521 , n24015 , n21842 );
and ( n25522 , n25520 , n21851 , n25521 );
or ( n25523 , n21851 , n24016 );
or ( n25524 , n22046 , n24015 );
nand ( n25525 , n25523 , n25524 );
nand ( n25526 , n22050 , n25525 );
not ( n25527 , n21851 );
not ( n25528 , n24000 );
or ( n25529 , n25527 , n25528 );
nand ( n25530 , n24001 , n22046 );
nand ( n25531 , n25529 , n25530 );
nand ( n25532 , n21846 , n25531 );
nand ( n25533 , n25526 , n25532 );
and ( n25534 , n25522 , n25533 );
xor ( n25535 , n25518 , n25534 );
not ( n25536 , n22050 );
not ( n25537 , n25531 );
or ( n25538 , n25536 , n25537 );
nand ( n25539 , n25514 , n21846 );
nand ( n25540 , n25538 , n25539 );
and ( n25541 , n25535 , n25540 );
or ( n25543 , n25541 , C0 );
and ( n25544 , n25517 , n25543 );
and ( n25545 , n25506 , n25516 );
or ( n25546 , n25544 , n25545 );
nand ( n25547 , n25505 , n25546 );
not ( n25548 , n25491 );
nand ( n25549 , n25548 , n25502 );
nand ( n25550 , n25547 , n25549 );
not ( n25551 , n25483 );
nand ( n25552 , n25551 , n25472 );
nand ( n25553 , n25550 , n25552 );
nand ( n25554 , n25485 , n25553 );
xor ( n25555 , n25438 , n25440 );
xor ( n25556 , n25555 , n25450 );
xor ( n25557 , n25554 , n25556 );
not ( n25558 , n25446 );
or ( n25559 , n25558 , n22643 );
and ( n25560 , n22179 , n23650 );
not ( n25561 , n22179 );
and ( n25562 , n25561 , n23653 );
nor ( n25563 , n25560 , n25562 );
or ( n25564 , n25563 , n22644 );
nand ( n25565 , n25559 , n25564 );
not ( n25566 , n25565 );
not ( n25567 , n25550 );
not ( n25568 , n25483 );
not ( n25569 , n25472 );
and ( n25570 , n25568 , n25569 );
and ( n25571 , n25483 , n25472 );
nor ( n25572 , n25570 , n25571 );
not ( n25573 , n25572 );
and ( n25574 , n25567 , n25573 );
and ( n25575 , n25550 , n25572 );
nor ( n25576 , n25574 , n25575 );
nand ( n25577 , n25566 , n25576 );
not ( n25578 , n25577 );
xnor ( n25579 , n25491 , n25502 );
not ( n25580 , n25546 );
and ( n25581 , n25579 , n25580 );
not ( n25582 , n25579 );
and ( n25583 , n25582 , n25546 );
nor ( n25584 , n25581 , n25583 );
not ( n25585 , n25563 );
not ( n25586 , n22643 );
and ( n25587 , n25585 , n25586 );
and ( n25588 , n22178 , n23537 );
not ( n25589 , n22178 );
and ( n25590 , n25589 , n23757 );
nor ( n25591 , n25588 , n25590 );
not ( n25592 , n25591 );
and ( n25593 , n25592 , n22645 );
nor ( n25594 , n25587 , n25593 );
and ( n25595 , n25584 , n25594 );
or ( n25596 , n25591 , n22643 );
and ( n25597 , n22178 , n23646 );
not ( n25598 , n22178 );
and ( n25599 , n25598 , n23645 );
nor ( n25600 , n25597 , n25599 );
or ( n25601 , n25600 , n22644 );
nand ( n25602 , n25596 , n25601 );
xor ( n25603 , n25506 , n25516 );
xor ( n25604 , n25603 , n25543 );
nor ( n25605 , n25602 , n25604 );
xor ( n25606 , n25522 , n25533 );
and ( n25607 , n22178 , n25315 );
not ( n25608 , n22178 );
and ( n25609 , n25608 , n23749 );
nor ( n25610 , n25607 , n25609 );
or ( n25611 , n25610 , n22643 );
and ( n25612 , n23942 , n22178 );
not ( n25613 , n23942 );
and ( n25614 , n25613 , n22179 );
nor ( n25615 , n25612 , n25614 );
or ( n25616 , n25615 , n22644 );
nand ( n25617 , n25611 , n25616 );
xor ( n25618 , n25606 , n25617 );
nor ( n25619 , n21845 , n24016 );
not ( n25620 , n24015 );
not ( n25621 , n22644 );
and ( n25622 , n25620 , n25621 );
and ( n25623 , n24001 , n22179 );
not ( n25624 , n24001 );
and ( n25625 , n25624 , n22178 );
or ( n25626 , n25623 , n25625 );
and ( n25627 , n25626 , n22642 );
nor ( n25628 , n25622 , n25627 );
nand ( n25629 , n24015 , n22642 );
nand ( n25630 , n25629 , n22178 );
nor ( n25631 , n25628 , n25630 );
xor ( n25632 , n25619 , n25631 );
not ( n25633 , n22645 );
not ( n25634 , n25626 );
or ( n25635 , n25633 , n25634 );
or ( n25636 , n25615 , n22643 );
nand ( n25637 , n25635 , n25636 );
and ( n25638 , n25632 , n25637 );
or ( n25640 , n25638 , C0 );
and ( n25641 , n25618 , n25640 );
and ( n25642 , n25606 , n25617 );
or ( n25643 , n25641 , n25642 );
or ( n25644 , n25600 , n22643 );
or ( n25645 , n25610 , n22644 );
nand ( n25646 , n25644 , n25645 );
or ( n25647 , n25643 , n25646 );
xor ( n25648 , n25518 , n25534 );
xor ( n25649 , n25648 , n25540 );
nand ( n25650 , n25647 , n25649 );
nand ( n25651 , n25643 , n25646 );
and ( n25652 , n25650 , n25651 );
or ( n25653 , n25605 , n25652 );
nand ( n25654 , n25602 , n25604 );
nand ( n25655 , n25653 , n25654 );
not ( n25656 , n25655 );
or ( n25657 , n25595 , n25656 );
or ( n25658 , n25584 , n25594 );
nand ( n25659 , n25657 , n25658 );
not ( n25660 , n25659 );
or ( n25661 , n25578 , n25660 );
not ( n25662 , n25576 );
nand ( n25663 , n25662 , n25565 );
nand ( n25664 , n25661 , n25663 );
and ( n25665 , n25557 , n25664 );
and ( n25666 , n25554 , n25556 );
or ( n25667 , n25665 , n25666 );
not ( n25668 , n25667 );
or ( n25669 , n25466 , n25668 );
not ( n25670 , n25464 );
nand ( n25671 , n25670 , n25453 );
nand ( n25672 , n25669 , n25671 );
and ( n25673 , n25429 , n25672 );
and ( n25674 , n25426 , n25428 );
or ( n25675 , n25673 , n25674 );
nand ( n25676 , n25405 , n25675 );
not ( n25677 , n25214 );
xor ( n25678 , n25241 , n25249 );
not ( n25679 , n25678 );
and ( n25680 , n25677 , n25679 );
and ( n25681 , n25214 , n25678 );
nor ( n25682 , n25680 , n25681 );
not ( n25683 , n25268 );
nand ( n25684 , n25683 , n25291 );
and ( n25685 , n25400 , n25684 );
nor ( n25686 , n25683 , n25291 );
nor ( n25687 , n25685 , n25686 );
and ( n25688 , n25682 , n25687 );
or ( n25689 , n25676 , n25688 );
not ( n25690 , n25404 );
nand ( n25691 , n25690 , n25258 );
or ( n25692 , n25688 , n25691 );
or ( n25693 , n25682 , n25687 );
nand ( n25694 , n25689 , n25692 , n25693 );
and ( n25695 , n25256 , n25694 );
and ( n25696 , n25253 , n25255 );
or ( n25697 , n25695 , n25696 );
and ( n25698 , n25212 , n25697 );
and ( n25699 , n25209 , n25211 );
or ( n25700 , n25698 , n25699 );
and ( n25701 , n25192 , n25700 );
and ( n25702 , n25189 , n25191 );
or ( n25703 , n25701 , n25702 );
not ( n25704 , n25703 );
or ( n25705 , n25052 , n25704 );
not ( n25706 , n25050 );
nand ( n25707 , n25706 , n25019 );
nand ( n25708 , n25705 , n25707 );
not ( n25709 , n25708 );
not ( n25710 , n24730 );
not ( n25711 , n24791 );
or ( n25712 , n25710 , n25711 );
nand ( n25713 , n24790 , n24731 );
nand ( n25714 , n25712 , n25713 );
not ( n25715 , n24795 );
and ( n25716 , n25714 , n25715 );
not ( n25717 , n25714 );
and ( n25718 , n25717 , n24795 );
nor ( n25719 , n25716 , n25718 );
xor ( n25720 , n24684 , n24694 );
xor ( n25721 , n25720 , n24704 );
not ( n25722 , n25721 );
not ( n25723 , n25038 );
not ( n25724 , n25043 );
or ( n25725 , n25723 , n25724 );
or ( n25726 , n25043 , n25038 );
nand ( n25727 , n25726 , n25048 );
nand ( n25728 , n25725 , n25727 );
not ( n25729 , n25728 );
or ( n25730 , n25722 , n25729 );
or ( n25731 , n25728 , n25721 );
xor ( n25732 , n24734 , n24776 );
xor ( n25733 , n25732 , n24787 );
nand ( n25734 , n25731 , n25733 );
nand ( n25735 , n25730 , n25734 );
not ( n25736 , n25735 );
nand ( n25737 , n25719 , n25736 );
xor ( n25738 , n25721 , n25728 );
xnor ( n25739 , n25738 , n25733 );
xor ( n25740 , n25025 , n25032 );
and ( n25741 , n25740 , n25049 );
and ( n25742 , n25025 , n25032 );
or ( n25743 , n25741 , n25742 );
nand ( n25744 , n25739 , n25743 );
and ( n25745 , n25737 , n25744 );
not ( n25746 , n25745 );
or ( n25747 , n25709 , n25746 );
nor ( n25748 , n25739 , n25743 );
and ( n25749 , n25737 , n25748 );
nor ( n25750 , n25719 , n25736 );
nor ( n25751 , n25749 , n25750 );
nand ( n25752 , n25747 , n25751 );
and ( n25753 , n24805 , n25752 );
and ( n25754 , n24798 , n24804 );
or ( n25755 , n25753 , n25754 );
not ( n25756 , n25755 );
or ( n25757 , n24728 , n25756 );
nor ( n25758 , n24578 , n24725 );
and ( n25759 , n24576 , n25758 );
nor ( n25760 , n24494 , n24575 );
nor ( n25761 , n25759 , n25760 );
nand ( n25762 , n25757 , n25761 );
and ( n25763 , n24492 , n25762 );
and ( n25764 , n24396 , n24491 );
or ( n25765 , n25763 , n25764 );
not ( n25766 , n25765 );
or ( n25767 , n24394 , n25766 );
not ( n25768 , n24196 );
and ( n25769 , n24198 , n24391 );
and ( n25770 , n25768 , n25769 );
and ( n25771 , n24195 , n24135 );
nor ( n25772 , n25770 , n25771 );
nand ( n25773 , n25767 , n25772 );
not ( n25774 , n25773 );
or ( n25775 , n24130 , n25774 );
nor ( n25776 , n23881 , n24127 );
and ( n25777 , n23876 , n25776 );
nor ( n25778 , n23830 , n23875 );
nor ( n25779 , n25777 , n25778 );
nand ( n25780 , n25775 , n25779 );
not ( n25781 , n25780 );
or ( n25782 , n23825 , n25781 );
nor ( n25783 , n23593 , n23822 );
and ( n25784 , n23591 , n25783 );
and ( n25785 , n23489 , n23590 );
nor ( n25786 , n25784 , n25785 );
nand ( n25787 , n25782 , n25786 );
not ( n25788 , n25787 );
or ( n25789 , n23487 , n25788 );
nor ( n25790 , n23349 , n23484 );
and ( n25791 , n23347 , n25790 );
nor ( n25792 , n23244 , n23346 );
nor ( n25793 , n25791 , n25792 );
nand ( n25794 , n25789 , n25793 );
buf ( n25795 , n25794 );
xor ( n25796 , n22664 , n22654 );
xor ( n25797 , n25796 , n22676 );
xor ( n25798 , n22577 , n22591 );
xor ( n25799 , n25798 , n22626 );
xor ( n25800 , n23147 , n23153 );
and ( n25801 , n25800 , n23158 );
and ( n25802 , n23147 , n23153 );
or ( n25803 , n25801 , n25802 );
xor ( n25804 , n25799 , n25803 );
xor ( n25805 , n25797 , n25804 );
xor ( n25806 , n23161 , n23167 );
and ( n25807 , n25806 , n23194 );
and ( n25808 , n23161 , n23167 );
or ( n25809 , n25807 , n25808 );
xor ( n25810 , n22693 , n22695 );
xor ( n25811 , n25810 , n22769 );
xor ( n25812 , n25809 , n25811 );
xor ( n25813 , n22790 , n22838 );
and ( n25814 , n25813 , n22946 );
and ( n25815 , n22790 , n22838 );
or ( n25816 , n25814 , n25815 );
xor ( n25817 , n25812 , n25816 );
xor ( n25818 , n25805 , n25817 );
xor ( n25819 , n23159 , n23195 );
and ( n25820 , n25819 , n23242 );
and ( n25821 , n23159 , n23195 );
or ( n25822 , n25820 , n25821 );
xor ( n25823 , n25818 , n25822 );
buf ( n25824 , n22947 );
or ( n25825 , n23243 , n25824 );
nand ( n25826 , n25825 , n23141 );
nand ( n25827 , n23243 , n25824 );
nand ( n25828 , n25826 , n25827 );
nor ( n25829 , n25823 , n25828 );
xor ( n25830 , n22772 , n22774 );
xor ( n25831 , n25830 , n22777 );
not ( n25832 , n25831 );
xor ( n25833 , n25809 , n25811 );
and ( n25834 , n25833 , n25816 );
and ( n25835 , n25809 , n25811 );
or ( n25836 , n25834 , n25835 );
not ( n25837 , n25836 );
not ( n25838 , n25797 );
not ( n25839 , n25803 );
not ( n25840 , n25839 );
and ( n25841 , n25838 , n25840 );
nand ( n25842 , n25797 , n25839 );
not ( n25843 , n25799 );
and ( n25844 , n25842 , n25843 );
nor ( n25845 , n25841 , n25844 );
not ( n25846 , n25845 );
and ( n25847 , n25837 , n25846 );
and ( n25848 , n25836 , n25845 );
nor ( n25849 , n25847 , n25848 );
not ( n25850 , n25849 );
or ( n25851 , n25832 , n25850 );
or ( n25852 , n25831 , n25849 );
nand ( n25853 , n25851 , n25852 );
xor ( n25854 , n25805 , n25817 );
and ( n25855 , n25854 , n25822 );
and ( n25856 , n25805 , n25817 );
or ( n25857 , n25855 , n25856 );
nor ( n25858 , n25853 , n25857 );
nor ( n25859 , n25829 , n25858 );
and ( n25860 , n25795 , n25859 );
nand ( n25861 , n25823 , n25828 );
or ( n25862 , n25861 , n25858 );
nand ( n25863 , n25853 , n25857 );
nand ( n25864 , n25862 , n25863 );
nor ( n25865 , n25860 , n25864 );
not ( n25866 , n22683 );
not ( n25867 , n22782 );
or ( n25868 , n25866 , n25867 );
nand ( n25869 , n22636 , n22682 );
nand ( n25870 , n25868 , n25869 );
not ( n25871 , n22780 );
and ( n25872 , n25870 , n25871 );
not ( n25873 , n25870 );
and ( n25874 , n25873 , n22780 );
nor ( n25875 , n25872 , n25874 );
not ( n25876 , n25836 );
not ( n25877 , n25876 );
not ( n25878 , n25845 );
and ( n25879 , n25877 , n25878 );
nand ( n25880 , n25876 , n25845 );
and ( n25881 , n25831 , n25880 );
nor ( n25882 , n25879 , n25881 );
nand ( n25883 , n25875 , n25882 );
not ( n25884 , n25883 );
or ( n25885 , n25865 , n25884 );
or ( n25886 , n25875 , n25882 );
nand ( n25887 , n25885 , n25886 );
xor ( n25888 , n22788 , n25887 );
or ( n25889 , n25888 , n19220 );
nand ( n25890 , n19222 , n25889 );
not ( n25891 , n19220 );
not ( n25892 , n18434 );
buf ( n25893 , n18971 );
not ( n25894 , n25893 );
or ( n25895 , n25892 , n25894 );
not ( n25896 , n18367 );
not ( n25897 , n18361 );
nor ( n25898 , n25896 , n25897 );
nand ( n25899 , n25895 , n25898 );
not ( n25900 , n18977 );
nand ( n25901 , n25900 , n18404 );
not ( n25902 , n25901 );
and ( n25903 , n25899 , n25902 );
not ( n25904 , n25899 );
and ( n25905 , n25904 , n25901 );
nor ( n25906 , n25903 , n25905 );
not ( n25907 , n25906 );
or ( n25908 , n25891 , n25907 );
not ( n25909 , n25778 );
nand ( n25910 , n25909 , n23876 );
not ( n25911 , n25910 );
not ( n25912 , n25773 );
not ( n25913 , n24128 );
or ( n25914 , n25912 , n25913 );
not ( n25915 , n25776 );
nand ( n25916 , n25914 , n25915 );
not ( n25917 , n25916 );
or ( n25918 , n25911 , n25917 );
or ( n25919 , n25916 , n25910 );
nand ( n25920 , n25918 , n25919 );
nand ( n25921 , n25920 , n19221 );
nand ( n25922 , n25908 , n25921 );
not ( n25923 , n18432 );
not ( n25924 , n25893 );
or ( n25925 , n25923 , n25924 );
not ( n25926 , n18340 );
nand ( n25927 , n25925 , n25926 );
buf ( n25928 , n18364 );
nand ( n25929 , n18273 , n25928 );
xor ( n25930 , n25927 , n25929 );
or ( n25931 , n25930 , n19221 );
not ( n25932 , n25768 );
nor ( n25933 , n25932 , n25771 );
not ( n25934 , n24392 );
and ( n25935 , n25765 , n25934 );
nor ( n25936 , n25935 , n25769 );
xor ( n25937 , n25933 , n25936 );
or ( n25938 , n25937 , n19220 );
nand ( n25939 , n25931 , n25938 );
not ( n25940 , n18431 );
not ( n25941 , n25940 );
not ( n25942 , n25893 );
or ( n25943 , n25941 , n25942 );
nand ( n25944 , n25943 , n18337 );
not ( n25945 , n18290 );
nand ( n25946 , n25945 , n18339 );
xor ( n25947 , n25944 , n25946 );
or ( n25948 , n25947 , n19221 );
not ( n25949 , n25769 );
nand ( n25950 , n25949 , n25934 );
xor ( n25951 , n25950 , n25765 );
or ( n25952 , n25951 , n19220 );
nand ( n25953 , n25948 , n25952 );
nand ( n25954 , n25940 , n18337 );
xor ( n25955 , n25954 , n18971 );
or ( n25956 , n25955 , n19221 );
xor ( n25957 , n24396 , n24491 );
xor ( n25958 , n25957 , n25762 );
not ( n25959 , n25958 );
or ( n25960 , n25959 , n19220 );
nand ( n25961 , n25956 , n25960 );
buf ( n25962 , n18496 );
not ( n25963 , n25962 );
buf ( n25964 , n18962 );
not ( n25965 , n25964 );
or ( n25966 , n25963 , n25965 );
nand ( n25967 , n25966 , n18966 );
nor ( n25968 , n18504 , n18969 );
and ( n25969 , n25967 , n25968 );
not ( n25970 , n25967 );
not ( n25971 , n25968 );
and ( n25972 , n25970 , n25971 );
or ( n25973 , n25969 , n25972 );
or ( n25974 , n25973 , n19221 );
not ( n25975 , n24576 );
nor ( n25976 , n25975 , n25760 );
and ( n25977 , n25755 , n24726 );
nor ( n25978 , n25977 , n25758 );
xor ( n25979 , n25976 , n25978 );
or ( n25980 , n25979 , n19220 );
nand ( n25981 , n25974 , n25980 );
not ( n25982 , n19220 );
not ( n25983 , n19191 );
not ( n25984 , n25983 );
not ( n25985 , n19179 );
or ( n25986 , n25984 , n25985 );
nand ( n25987 , n25986 , n19207 );
not ( n25988 , n25987 );
buf ( n25989 , n25988 );
not ( n25990 , n25989 );
not ( n25991 , n18990 );
or ( n25992 , n25990 , n25991 );
nor ( n25993 , n19178 , n19191 );
or ( n25994 , n25993 , n19203 );
nand ( n25995 , n25994 , n19194 );
not ( n25996 , n25995 );
nand ( n25997 , n25992 , n25996 );
not ( n25998 , n25997 );
xor ( n25999 , n19130 , n19170 );
and ( n26000 , n25999 , n19177 );
and ( n26001 , n19130 , n19170 );
or ( n26002 , n26000 , n26001 );
buf ( n26003 , n19129 );
and ( n26004 , n26003 , n471 );
xor ( n26005 , n19172 , n19173 );
and ( n26006 , n26005 , n19176 );
and ( n26007 , n19172 , n19173 );
or ( n26008 , n26006 , n26007 );
xor ( n26009 , n26004 , n26008 );
not ( n26010 , n9907 );
nand ( n26011 , n16722 , n17577 );
not ( n26012 , n16205 );
and ( n26013 , n26012 , n17582 );
and ( n26014 , n26011 , n26013 );
not ( n26015 , n26011 );
not ( n26016 , n26013 );
and ( n26017 , n26015 , n26016 );
nor ( n26018 , n26014 , n26017 );
not ( n26019 , n26018 );
or ( n26020 , n26010 , n26019 );
nor ( n26021 , n19119 , n19080 );
nor ( n26022 , n19062 , n26021 );
not ( n26023 , n26022 );
not ( n26024 , n15409 );
or ( n26025 , n26023 , n26024 );
and ( n26026 , n19073 , n19120 );
not ( n26027 , n19121 );
nor ( n26028 , n26026 , n26027 );
nand ( n26029 , n26025 , n26028 );
xor ( n26030 , n19098 , n19113 );
and ( n26031 , n26030 , n19118 );
and ( n26032 , n19098 , n19113 );
or ( n26033 , n26031 , n26032 );
or ( n26034 , n3288 , n3955 );
nand ( n26035 , n26034 , n541 );
not ( n26036 , n3103 );
not ( n26037 , n19086 );
or ( n26038 , n26036 , n26037 );
not ( n26039 , n539 );
not ( n26040 , n17972 );
or ( n26041 , n26039 , n26040 );
nand ( n26042 , n17971 , n3069 );
nand ( n26043 , n26041 , n26042 );
nand ( n26044 , n26043 , n14397 );
nand ( n26045 , n26038 , n26044 );
xor ( n26046 , n26035 , n26045 );
and ( n26047 , n537 , n17985 );
xor ( n26048 , n26046 , n26047 );
not ( n26049 , n11729 );
not ( n26050 , n19095 );
or ( n26051 , n26049 , n26050 );
xor ( n26052 , n537 , n14354 );
nand ( n26053 , n26052 , n3134 );
nand ( n26054 , n26051 , n26053 );
not ( n26055 , n19103 );
xor ( n26056 , n26054 , n26055 );
xor ( n26057 , n19081 , n19090 );
and ( n26058 , n26057 , n19097 );
and ( n26059 , n19081 , n19090 );
or ( n26060 , n26058 , n26059 );
xor ( n26061 , n26056 , n26060 );
xor ( n26062 , n26048 , n26061 );
xor ( n26063 , n19103 , n19107 );
and ( n26064 , n26063 , n19112 );
and ( n26065 , n19103 , n19107 );
or ( n26066 , n26064 , n26065 );
xor ( n26067 , n26062 , n26066 );
nor ( n26068 , n26033 , n26067 );
not ( n26069 , n26068 );
nand ( n26070 , n26033 , n26067 );
nand ( n26071 , n26069 , n26070 );
and ( n26072 , n454 , n26071 );
and ( n26073 , n26029 , n26072 );
not ( n26074 , n26029 );
not ( n26075 , n454 );
nor ( n26076 , n26075 , n26071 );
and ( n26077 , n26074 , n26076 );
nor ( n26078 , n26073 , n26077 );
nand ( n26079 , n26020 , n26078 );
and ( n26080 , n26079 , n472 );
and ( n26081 , n19175 , n469 );
xor ( n26082 , n26080 , n26081 );
and ( n26083 , n19166 , n470 );
xor ( n26084 , n26082 , n26083 );
xor ( n26085 , n26009 , n26084 );
nand ( n26086 , n26002 , n26085 );
buf ( n26087 , n26086 );
not ( n26088 , n26087 );
nor ( n26089 , n26021 , n26068 );
not ( n26090 , n26089 );
not ( n26091 , n19075 );
or ( n26092 , n26090 , n26091 );
and ( n26093 , n26027 , n26069 );
not ( n26094 , n26070 );
nor ( n26095 , n26093 , n26094 );
nand ( n26096 , n26092 , n26095 );
xor ( n26097 , n26048 , n26061 );
and ( n26098 , n26097 , n26066 );
and ( n26099 , n26048 , n26061 );
or ( n26100 , n26098 , n26099 );
xor ( n26101 , n26035 , n26045 );
and ( n26102 , n26101 , n26047 );
and ( n26103 , n26035 , n26045 );
or ( n26104 , n26102 , n26103 );
not ( n26105 , n3134 );
not ( n26106 , n537 );
not ( n26107 , n14323 );
or ( n26108 , n26106 , n26107 );
nand ( n26109 , n14326 , n3177 );
nand ( n26110 , n26108 , n26109 );
not ( n26111 , n26110 );
or ( n26112 , n26105 , n26111 );
nand ( n26113 , n26052 , n11729 );
nand ( n26114 , n26112 , n26113 );
and ( n26115 , n14419 , n537 );
xor ( n26116 , n26114 , n26115 );
and ( n26117 , n26043 , n3103 );
nor ( n26118 , n26117 , n11416 );
xor ( n26119 , n26116 , n26118 );
xor ( n26120 , n26104 , n26119 );
xor ( n26121 , n26054 , n26055 );
and ( n26122 , n26121 , n26060 );
and ( n26123 , n26054 , n26055 );
or ( n26124 , n26122 , n26123 );
xor ( n26125 , n26120 , n26124 );
nor ( n26126 , n26100 , n26125 );
not ( n26127 , n26126 );
nand ( n26128 , n26100 , n26125 );
nand ( n26129 , n26127 , n26128 );
not ( n26130 , n26129 );
and ( n26131 , n26096 , n26130 );
not ( n26132 , n454 );
nor ( n26133 , n26131 , n26132 );
not ( n26134 , n26133 );
not ( n26135 , n26096 );
nand ( n26136 , n26135 , n26129 );
not ( n26137 , n26136 );
or ( n26138 , n26134 , n26137 );
not ( n26139 , n454 );
not ( n26140 , n26012 );
not ( n26141 , n17578 );
or ( n26142 , n26140 , n26141 );
nand ( n26143 , n26142 , n17582 );
not ( n26144 , n17581 );
nand ( n26145 , n26144 , n17584 );
not ( n26146 , n26145 );
and ( n26147 , n26143 , n26146 );
not ( n26148 , n26143 );
and ( n26149 , n26148 , n26145 );
nor ( n26150 , n26147 , n26149 );
nand ( n26151 , n26139 , n26150 );
nand ( n26152 , n26138 , n26151 );
buf ( n26153 , n26152 );
and ( n26154 , n26153 , n472 );
xor ( n26155 , n26080 , n26081 );
and ( n26156 , n26155 , n26083 );
and ( n26157 , n26080 , n26081 );
or ( n26158 , n26156 , n26157 );
xor ( n26159 , n26154 , n26158 );
and ( n26160 , n26079 , n471 );
not ( n26161 , n19166 );
nor ( n26162 , n26161 , n17873 );
xor ( n26163 , n26160 , n26162 );
and ( n26164 , n19129 , n470 );
xor ( n26165 , n26163 , n26164 );
xor ( n26166 , n26159 , n26165 );
xor ( n26167 , n26004 , n26008 );
and ( n26168 , n26167 , n26084 );
and ( n26169 , n26004 , n26008 );
or ( n26170 , n26168 , n26169 );
nor ( n26171 , n26166 , n26170 );
not ( n26172 , n26171 );
buf ( n26173 , n26166 );
nand ( n26174 , n26173 , n26170 );
nand ( n26175 , n26172 , n26174 );
nor ( n26176 , n26088 , n26175 );
nand ( n26177 , n25998 , n26176 );
or ( n26178 , n26002 , n26085 );
nand ( n26179 , n25997 , n26178 , n26175 );
and ( n26180 , n26175 , n26087 );
not ( n26181 , n26175 );
not ( n26182 , n26178 );
nand ( n26183 , n26182 , n26087 );
and ( n26184 , n26181 , n26183 );
or ( n26185 , n26180 , n26184 );
nand ( n26186 , n26177 , n26179 , n26185 );
not ( n26187 , n26186 );
or ( n26188 , n25982 , n26187 );
or ( n26189 , n22317 , n22242 );
or ( n26190 , n21637 , n22224 );
nand ( n26191 , n26189 , n26190 );
or ( n26192 , n22121 , n22062 );
nand ( n26193 , n26192 , n22071 );
xor ( n26194 , n26191 , n26193 );
not ( n26195 , n21577 );
not ( n26196 , n21595 );
not ( n26197 , n21769 );
or ( n26198 , n26196 , n26197 );
nand ( n26199 , n21768 , n21623 );
nand ( n26200 , n26198 , n26199 );
not ( n26201 , n26200 );
or ( n26202 , n26195 , n26201 );
and ( n26203 , n21595 , n21543 );
not ( n26204 , n21595 );
and ( n26205 , n26204 , n21546 );
nor ( n26206 , n26203 , n26205 );
nand ( n26207 , n26206 , n21646 );
nand ( n26208 , n26202 , n26207 );
xor ( n26209 , n26194 , n26208 );
not ( n26210 , n22225 );
not ( n26211 , n22314 );
or ( n26212 , n26210 , n26211 );
nand ( n26213 , n22273 , n22243 );
nand ( n26214 , n26212 , n26213 );
not ( n26215 , n22299 );
not ( n26216 , n22268 );
not ( n26217 , n21620 );
or ( n26218 , n26216 , n26217 );
nand ( n26219 , n22974 , n22277 );
nand ( n26220 , n26218 , n26219 );
not ( n26221 , n26220 );
or ( n26222 , n26215 , n26221 );
not ( n26223 , n22268 );
not ( n26224 , n21459 );
or ( n26225 , n26223 , n26224 );
nand ( n26226 , n21456 , n22277 );
nand ( n26227 , n26225 , n26226 );
nand ( n26228 , n26227 , n22266 );
nand ( n26229 , n26222 , n26228 );
xor ( n26230 , n26214 , n26229 );
not ( n26231 , n21549 );
not ( n26232 , n19319 );
not ( n26233 , n22153 );
or ( n26234 , n26232 , n26233 );
nand ( n26235 , n22150 , n19318 );
nand ( n26236 , n26234 , n26235 );
not ( n26237 , n26236 );
or ( n26238 , n26231 , n26237 );
and ( n26239 , n19319 , n21830 );
not ( n26240 , n19319 );
and ( n26241 , n26240 , n21831 );
nor ( n26242 , n26239 , n26241 );
nand ( n26243 , n26242 , n19316 );
nand ( n26244 , n26238 , n26243 );
xor ( n26245 , n26230 , n26244 );
xor ( n26246 , n26209 , n26245 );
not ( n26247 , n22071 );
not ( n26248 , n22062 );
or ( n26249 , n26247 , n26248 );
nand ( n26250 , n22479 , n22121 );
nand ( n26251 , n26249 , n26250 );
xor ( n26252 , n22341 , n22346 );
and ( n26253 , n26252 , n22362 );
and ( n26254 , n22341 , n22346 );
or ( n26255 , n26253 , n26254 );
xor ( n26256 , n26251 , n26255 );
not ( n26257 , n19316 );
not ( n26258 , n22381 );
or ( n26259 , n26257 , n26258 );
nand ( n26260 , n26242 , n21549 );
nand ( n26261 , n26259 , n26260 );
and ( n26262 , n26256 , n26261 );
and ( n26263 , n26251 , n26255 );
or ( n26264 , n26262 , n26263 );
xor ( n26265 , n26246 , n26264 );
not ( n26266 , n21837 );
not ( n26267 , n21651 );
not ( n26268 , n22114 );
or ( n26269 , n26267 , n26268 );
nand ( n26270 , n22111 , n21834 );
nand ( n26271 , n26269 , n26270 );
not ( n26272 , n26271 );
or ( n26273 , n26266 , n26272 );
nand ( n26274 , n22489 , n21698 );
nand ( n26275 , n26273 , n26274 );
not ( n26276 , n22134 );
and ( n26277 , n22137 , n22038 );
not ( n26278 , n22137 );
and ( n26279 , n26278 , n22041 );
nor ( n26280 , n26277 , n26279 );
not ( n26281 , n26280 );
or ( n26282 , n26276 , n26281 );
nand ( n26283 , n22498 , n22166 );
nand ( n26284 , n26282 , n26283 );
xor ( n26285 , n26275 , n26284 );
xor ( n26286 , n22376 , n22385 );
and ( n26287 , n26286 , n22395 );
and ( n26288 , n22376 , n22385 );
or ( n26289 , n26287 , n26288 );
and ( n26290 , n26285 , n26289 );
and ( n26291 , n26275 , n26284 );
or ( n26292 , n26290 , n26291 );
not ( n26293 , n21698 );
not ( n26294 , n26271 );
or ( n26295 , n26293 , n26294 );
not ( n26296 , n21651 );
not ( n26297 , n22086 );
or ( n26298 , n26296 , n26297 );
nand ( n26299 , n22083 , n21834 );
nand ( n26300 , n26298 , n26299 );
nand ( n26301 , n26300 , n21837 );
nand ( n26302 , n26295 , n26301 );
not ( n26303 , n22166 );
not ( n26304 , n26280 );
or ( n26305 , n26303 , n26304 );
not ( n26306 , n22137 );
not ( n26307 , n22021 );
or ( n26308 , n26306 , n26307 );
nand ( n26309 , n22018 , n22136 );
nand ( n26310 , n26308 , n26309 );
nand ( n26311 , n26310 , n22134 );
nand ( n26312 , n26305 , n26311 );
xor ( n26313 , n26302 , n26312 );
not ( n26314 , n26214 );
not ( n26315 , n21646 );
not ( n26316 , n22391 );
or ( n26317 , n26315 , n26316 );
nand ( n26318 , n26206 , n21577 );
nand ( n26319 , n26317 , n26318 );
xor ( n26320 , n26314 , n26319 );
not ( n26321 , n22266 );
not ( n26322 , n26220 );
or ( n26323 , n26321 , n26322 );
nand ( n26324 , n22353 , n22299 );
nand ( n26325 , n26323 , n26324 );
and ( n26326 , n26320 , n26325 );
and ( n26327 , n26314 , n26319 );
or ( n26328 , n26326 , n26327 );
xor ( n26329 , n26313 , n26328 );
xor ( n26330 , n26292 , n26329 );
xor ( n26331 , n26314 , n26319 );
xor ( n26332 , n26331 , n26325 );
xor ( n26333 , n22481 , n22491 );
and ( n26334 , n26333 , n22502 );
and ( n26335 , n22481 , n22491 );
or ( n26336 , n26334 , n26335 );
xor ( n26337 , n26332 , n26336 );
xor ( n26338 , n26251 , n26255 );
xor ( n26339 , n26338 , n26261 );
and ( n26340 , n26337 , n26339 );
and ( n26341 , n26332 , n26336 );
or ( n26342 , n26340 , n26341 );
xor ( n26343 , n26330 , n26342 );
xor ( n26344 , n26265 , n26343 );
xor ( n26345 , n26275 , n26284 );
xor ( n26346 , n26345 , n26289 );
xor ( n26347 , n22341 , n22346 );
xor ( n26348 , n26347 , n22362 );
and ( n26349 , n22375 , n26348 );
xor ( n26350 , n22341 , n22346 );
xor ( n26351 , n26350 , n22362 );
and ( n26352 , n22396 , n26351 );
and ( n26353 , n22375 , n22396 );
or ( n26354 , n26349 , n26352 , n26353 );
xor ( n26355 , n26346 , n26354 );
xor ( n26356 , n22467 , n22471 );
and ( n26357 , n26356 , n22503 );
and ( n26358 , n22467 , n22471 );
or ( n26359 , n26357 , n26358 );
and ( n26360 , n26355 , n26359 );
and ( n26361 , n26346 , n26354 );
or ( n26362 , n26360 , n26361 );
xor ( n26363 , n26344 , n26362 );
xor ( n26364 , n26332 , n26336 );
xor ( n26365 , n26364 , n26339 );
xor ( n26366 , n26346 , n26354 );
xor ( n26367 , n26366 , n26359 );
xor ( n26368 , n26365 , n26367 );
xor ( n26369 , n22398 , n22462 );
and ( n26370 , n26369 , n22504 );
and ( n26371 , n22398 , n22462 );
or ( n26372 , n26370 , n26371 );
and ( n26373 , n26368 , n26372 );
and ( n26374 , n26365 , n26367 );
or ( n26375 , n26373 , n26374 );
nand ( n26376 , n26363 , n26375 );
nor ( n26377 , n26363 , n26375 );
not ( n26378 , n26377 );
nand ( n26379 , n26376 , n26378 );
not ( n26380 , n26379 );
and ( n26381 , n22787 , n25859 , n25883 );
not ( n26382 , n26381 );
not ( n26383 , n25794 );
or ( n26384 , n26382 , n26383 );
not ( n26385 , n25883 );
not ( n26386 , n25864 );
or ( n26387 , n26385 , n26386 );
nand ( n26388 , n26387 , n25886 );
and ( n26389 , n26388 , n22787 );
nor ( n26390 , n26389 , n22785 );
nand ( n26391 , n26384 , n26390 );
xor ( n26392 , n26365 , n26367 );
xor ( n26393 , n26392 , n26372 );
or ( n26394 , n22633 , n22339 );
nand ( n26395 , n26394 , n22505 );
nand ( n26396 , n22633 , n22339 );
nand ( n26397 , n26395 , n26396 );
or ( n26398 , n26393 , n26397 );
nand ( n26399 , n26391 , n26398 );
nand ( n26400 , n26393 , n26397 );
nand ( n26401 , n26399 , n26400 );
not ( n26402 , n26401 );
or ( n26403 , n26380 , n26402 );
or ( n26404 , n26401 , n26379 );
nand ( n26405 , n26403 , n26404 );
nand ( n26406 , n26405 , n19221 );
nand ( n26407 , n26188 , n26406 );
nand ( n26408 , n25962 , n18966 );
not ( n26409 , n26408 );
and ( n26410 , n25964 , n26409 );
not ( n26411 , n25964 );
and ( n26412 , n26411 , n26408 );
or ( n26413 , n26410 , n26412 );
or ( n26414 , n26413 , n19221 );
not ( n26415 , n25758 );
nand ( n26416 , n26415 , n24726 );
xor ( n26417 , n26416 , n25755 );
or ( n26418 , n26417 , n19220 );
nand ( n26419 , n26414 , n26418 );
not ( n26420 , n18546 );
not ( n26421 , n26420 );
not ( n26422 , n18953 );
or ( n26423 , n26421 , n26422 );
nand ( n26424 , n26423 , n18957 );
or ( n26425 , n18960 , n18529 );
xor ( n26426 , n26424 , n26425 );
or ( n26427 , n26426 , n19221 );
xor ( n26428 , n24798 , n24804 );
xor ( n26429 , n26428 , n25752 );
not ( n26430 , n26429 );
or ( n26431 , n26430 , n19220 );
nand ( n26432 , n26427 , n26431 );
nand ( n26433 , n26420 , n18957 );
xor ( n26434 , n18953 , n26433 );
or ( n26435 , n26434 , n19221 );
not ( n26436 , n25750 );
nand ( n26437 , n26436 , n25737 );
and ( n26438 , n25703 , n25051 );
not ( n26439 , n25707 );
nor ( n26440 , n26438 , n26439 );
not ( n26441 , n25744 );
or ( n26442 , n26440 , n26441 );
not ( n26443 , n25748 );
nand ( n26444 , n26442 , n26443 );
xor ( n26445 , n26437 , n26444 );
or ( n26446 , n26445 , n19220 );
nand ( n26447 , n26435 , n26446 );
nand ( n26448 , n26178 , n26086 );
xor ( n26449 , n25997 , n26448 );
or ( n26450 , n26449 , n19221 );
nand ( n26451 , n26400 , n26398 );
buf ( n26452 , n26391 );
xor ( n26453 , n26451 , n26452 );
or ( n26454 , n26453 , n19220 );
nand ( n26455 , n26450 , n26454 );
not ( n26456 , n18943 );
not ( n26457 , n26456 );
buf ( n26458 , n18921 );
not ( n26459 , n26458 );
or ( n26460 , n26457 , n26459 );
nand ( n26461 , n26460 , n18948 );
not ( n26462 , n18951 );
nand ( n26463 , n26462 , n18947 );
xor ( n26464 , n26461 , n26463 );
or ( n26465 , n26464 , n19221 );
nor ( n26466 , n26441 , n25748 );
xor ( n26467 , n26466 , n26440 );
or ( n26468 , n26467 , n19220 );
nand ( n26469 , n26465 , n26468 );
nand ( n26470 , n18948 , n26456 );
not ( n26471 , n26470 );
and ( n26472 , n26458 , n26471 );
not ( n26473 , n26458 );
and ( n26474 , n26473 , n26470 );
or ( n26475 , n26472 , n26474 );
or ( n26476 , n26475 , n19221 );
nand ( n26477 , n25707 , n25051 );
xor ( n26478 , n26477 , n25703 );
or ( n26479 , n26478 , n19220 );
nand ( n26480 , n26476 , n26479 );
not ( n26481 , n18648 );
not ( n26482 , n26481 );
not ( n26483 , n18912 );
or ( n26484 , n26482 , n26483 );
nand ( n26485 , n26484 , n18916 );
nor ( n26486 , n18919 , n18601 );
not ( n26487 , n26486 );
and ( n26488 , n26485 , n26487 );
not ( n26489 , n26485 );
and ( n26490 , n26489 , n26486 );
nor ( n26491 , n26488 , n26490 );
or ( n26492 , n26491 , n19221 );
xor ( n26493 , n25189 , n25191 );
xor ( n26494 , n26493 , n25700 );
not ( n26495 , n26494 );
or ( n26496 , n26495 , n19220 );
nand ( n26497 , n26492 , n26496 );
nand ( n26498 , n26481 , n18916 );
xor ( n26499 , n26498 , n18912 );
or ( n26500 , n26499 , n19221 );
xor ( n26501 , n25209 , n25211 );
xor ( n26502 , n26501 , n25697 );
not ( n26503 , n26502 );
or ( n26504 , n26503 , n19220 );
nand ( n26505 , n26500 , n26504 );
not ( n26506 , n18712 );
not ( n26507 , n18697 );
not ( n26508 , n18901 );
or ( n26509 , n26507 , n26508 );
nand ( n26510 , n26509 , n18905 );
not ( n26511 , n26510 );
or ( n26512 , n26506 , n26511 );
nand ( n26513 , n26512 , n18907 );
not ( n26514 , n18904 );
nor ( n26515 , n26514 , n18910 );
not ( n26516 , n26515 );
and ( n26517 , n26513 , n26516 );
not ( n26518 , n26513 );
and ( n26519 , n26518 , n26515 );
nor ( n26520 , n26517 , n26519 );
or ( n26521 , n26520 , n19221 );
xor ( n26522 , n25253 , n25255 );
xor ( n26523 , n26522 , n25694 );
not ( n26524 , n26523 );
or ( n26525 , n26524 , n19220 );
nand ( n26526 , n26521 , n26525 );
buf ( n26527 , n18420 );
not ( n26528 , n26527 );
not ( n26529 , n18972 );
not ( n26530 , n26529 );
not ( n26531 , n18435 );
not ( n26532 , n26531 );
or ( n26533 , n26530 , n26532 );
nor ( n26534 , n18417 , n18988 );
nand ( n26535 , n26533 , n26534 );
not ( n26536 , n26535 );
or ( n26537 , n26528 , n26536 );
not ( n26538 , n17928 );
nand ( n26539 , n26537 , n26538 );
not ( n26540 , n18179 );
not ( n26541 , n26540 );
or ( n26542 , n18050 , n18055 );
nand ( n26543 , n26541 , n26542 );
and ( n26544 , n26539 , n26543 );
not ( n26545 , n26539 );
not ( n26546 , n26543 );
and ( n26547 , n26545 , n26546 );
nor ( n26548 , n26544 , n26547 );
or ( n26549 , n26548 , n19221 );
not ( n26550 , n25861 );
nor ( n26551 , n26550 , n25829 );
and ( n26552 , n26551 , n25795 );
not ( n26553 , n26551 );
not ( n26554 , n25795 );
and ( n26555 , n26553 , n26554 );
or ( n26556 , n26552 , n26555 );
or ( n26557 , n26556 , n19220 );
nand ( n26558 , n26549 , n26557 );
nand ( n26559 , n18773 , n18894 );
xor ( n26560 , n18891 , n26559 );
not ( n26561 , n19220 );
or ( n26562 , n26560 , n26561 );
xor ( n26563 , n25554 , n25556 );
xor ( n26564 , n26563 , n25664 );
not ( n26565 , n26564 );
or ( n26566 , n26565 , n19220 );
nand ( n26567 , n26562 , n26566 );
not ( n26568 , n19220 );
or ( n26569 , n17887 , n17821 );
nand ( n26570 , n26569 , n17927 );
not ( n26571 , n26570 );
not ( n26572 , n18419 );
not ( n26573 , n26572 );
not ( n26574 , n26535 );
or ( n26575 , n26573 , n26574 );
buf ( n26576 , n17925 );
nand ( n26577 , n26575 , n26576 );
not ( n26578 , n26577 );
or ( n26579 , n26571 , n26578 );
or ( n26580 , n26577 , n26570 );
nand ( n26581 , n26579 , n26580 );
not ( n26582 , n26581 );
or ( n26583 , n26568 , n26582 );
not ( n26584 , n25792 );
nand ( n26585 , n26584 , n23347 );
not ( n26586 , n26585 );
not ( n26587 , n23485 );
not ( n26588 , n25787 );
or ( n26589 , n26587 , n26588 );
not ( n26590 , n25790 );
nand ( n26591 , n26589 , n26590 );
not ( n26592 , n26591 );
or ( n26593 , n26586 , n26592 );
or ( n26594 , n26591 , n26585 );
nand ( n26595 , n26593 , n26594 );
nand ( n26596 , n26595 , n19221 );
nand ( n26597 , n26583 , n26596 );
not ( n26598 , n19220 );
nand ( n26599 , n26576 , n26572 );
not ( n26600 , n26599 );
and ( n26601 , n26535 , n26600 );
not ( n26602 , n26535 );
and ( n26603 , n26602 , n26599 );
nor ( n26604 , n26601 , n26603 );
not ( n26605 , n26604 );
or ( n26606 , n26598 , n26605 );
nand ( n26607 , n23485 , n26590 );
not ( n26608 , n26607 );
not ( n26609 , n25787 );
or ( n26610 , n26608 , n26609 );
or ( n26611 , n25787 , n26607 );
nand ( n26612 , n26610 , n26611 );
nand ( n26613 , n26612 , n19221 );
nand ( n26614 , n26606 , n26613 );
not ( n26615 , n25595 );
nand ( n26616 , n26615 , n25658 );
xor ( n26617 , n25655 , n26616 );
or ( n26618 , n26617 , n19220 );
nand ( n26619 , n18846 , n18886 );
xnor ( n26620 , n26619 , n18883 );
nand ( n26621 , n19220 , n26620 );
nand ( n26622 , n26618 , n26621 );
not ( n26623 , n6587 );
nand ( n26624 , n26623 , n454 );
not ( n26625 , n6595 );
nand ( n26626 , n26625 , n6597 );
or ( n26627 , n26624 , n26626 );
not ( n26628 , n9757 );
nand ( n26629 , n26628 , n9797 );
xor ( n26630 , n26629 , n9795 );
or ( n26631 , n454 , n26630 );
nand ( n26632 , n26626 , n6587 , n454 );
nand ( n26633 , n26627 , n26631 , n26632 );
not ( n26634 , n26633 );
not ( n26635 , n19220 );
and ( n26636 , n22573 , n22864 );
nor ( n26637 , n26636 , n19318 );
not ( n26638 , n21831 );
not ( n26639 , n22242 );
and ( n26640 , n26638 , n26639 );
and ( n26641 , n22150 , n22225 );
nor ( n26642 , n26640 , n26641 );
xor ( n26643 , n26637 , n26642 );
not ( n26644 , n21595 );
not ( n26645 , n22041 );
or ( n26646 , n26644 , n26645 );
nand ( n26647 , n22038 , n21623 );
nand ( n26648 , n26646 , n26647 );
not ( n26649 , n26648 );
not ( n26650 , n26649 );
not ( n26651 , n23170 );
and ( n26652 , n26650 , n26651 );
and ( n26653 , n21595 , n22018 );
not ( n26654 , n21595 );
and ( n26655 , n26654 , n22021 );
nor ( n26656 , n26653 , n26655 );
and ( n26657 , n26656 , n21577 );
nor ( n26658 , n26652 , n26657 );
xor ( n26659 , n26643 , n26658 );
not ( n26660 , n19316 );
not ( n26661 , n19319 );
not ( n26662 , n22021 );
or ( n26663 , n26661 , n26662 );
nand ( n26664 , n19318 , n22018 );
nand ( n26665 , n26663 , n26664 );
not ( n26666 , n26665 );
or ( n26667 , n26660 , n26666 );
nand ( n26668 , n21549 , n19319 );
nand ( n26669 , n26667 , n26668 );
not ( n26670 , n22225 );
not ( n26671 , n21768 );
or ( n26672 , n26670 , n26671 );
nand ( n26673 , n21543 , n22243 );
nand ( n26674 , n26672 , n26673 );
not ( n26675 , n26674 );
and ( n26676 , n22871 , n22877 );
nor ( n26677 , n26676 , n21834 );
nand ( n26678 , n26675 , n26677 );
not ( n26679 , n26678 );
not ( n26680 , n22299 );
and ( n26681 , n22268 , n21830 );
not ( n26682 , n22268 );
and ( n26683 , n26682 , n21831 );
nor ( n26684 , n26681 , n26683 );
not ( n26685 , n26684 );
or ( n26686 , n26680 , n26685 );
not ( n26687 , n22268 );
not ( n26688 , n22153 );
or ( n26689 , n26687 , n26688 );
nand ( n26690 , n22150 , n22277 );
nand ( n26691 , n26689 , n26690 );
nand ( n26692 , n26691 , n22266 );
nand ( n26693 , n26686 , n26692 );
not ( n26694 , n26693 );
or ( n26695 , n26679 , n26694 );
not ( n26696 , n26677 );
nand ( n26697 , n26696 , n26674 );
nand ( n26698 , n26695 , n26697 );
not ( n26699 , n26698 );
xor ( n26700 , n26669 , n26699 );
not ( n26701 , n22243 );
not ( n26702 , n21456 );
or ( n26703 , n26701 , n26702 );
nand ( n26704 , n21543 , n22225 );
nand ( n26705 , n26703 , n26704 );
not ( n26706 , n19316 );
not ( n26707 , n19319 );
not ( n26708 , n22041 );
or ( n26709 , n26707 , n26708 );
nand ( n26710 , n22038 , n19318 );
nand ( n26711 , n26709 , n26710 );
not ( n26712 , n26711 );
or ( n26713 , n26706 , n26712 );
nand ( n26714 , n26665 , n21549 );
nand ( n26715 , n26713 , n26714 );
xor ( n26716 , n26705 , n26715 );
not ( n26717 , n21646 );
not ( n26718 , n21595 );
not ( n26719 , n22114 );
or ( n26720 , n26718 , n26719 );
nand ( n26721 , n22111 , n21623 );
nand ( n26722 , n26720 , n26721 );
not ( n26723 , n26722 );
or ( n26724 , n26717 , n26723 );
not ( n26725 , n21595 );
not ( n26726 , n22086 );
or ( n26727 , n26725 , n26726 );
nand ( n26728 , n22083 , n21623 );
nand ( n26729 , n26727 , n26728 );
nand ( n26730 , n26729 , n21577 );
nand ( n26731 , n26724 , n26730 );
and ( n26732 , n26716 , n26731 );
and ( n26733 , n26705 , n26715 );
or ( n26734 , n26732 , n26733 );
not ( n26735 , n26734 );
and ( n26736 , n26700 , n26735 );
and ( n26737 , n26669 , n26699 );
or ( n26738 , n26736 , n26737 );
xor ( n26739 , n26659 , n26738 );
and ( n26740 , n22277 , n22086 );
not ( n26741 , n22277 );
and ( n26742 , n26741 , n22083 );
nor ( n26743 , n26740 , n26742 );
not ( n26744 , n26743 );
not ( n26745 , n22266 );
or ( n26746 , n26744 , n26745 );
and ( n26747 , n22277 , n22111 );
not ( n26748 , n22277 );
and ( n26749 , n26748 , n22114 );
nor ( n26750 , n26747 , n26749 );
not ( n26751 , n26750 );
nand ( n26752 , n26751 , n22299 );
nand ( n26753 , n26746 , n26752 );
xor ( n26754 , n26753 , n26669 );
not ( n26755 , n22225 );
not ( n26756 , n21830 );
or ( n26757 , n26755 , n26756 );
or ( n26758 , n21769 , n22242 );
nand ( n26759 , n26757 , n26758 );
not ( n26760 , n21646 );
not ( n26761 , n26729 );
or ( n26762 , n26760 , n26761 );
nand ( n26763 , n26648 , n21577 );
nand ( n26764 , n26762 , n26763 );
xor ( n26765 , n26759 , n26764 );
not ( n26766 , n26691 );
or ( n26767 , n26766 , n22934 );
or ( n26768 , n26750 , n22265 );
nand ( n26769 , n26767 , n26768 );
and ( n26770 , n26765 , n26769 );
and ( n26771 , n26759 , n26764 );
or ( n26772 , n26770 , n26771 );
xor ( n26773 , n26754 , n26772 );
not ( n26774 , n26773 );
and ( n26775 , n26739 , n26774 );
and ( n26776 , n26659 , n26738 );
or ( n26777 , n26775 , n26776 );
xor ( n26778 , n26637 , n26642 );
and ( n26779 , n26778 , n26658 );
and ( n26780 , n26637 , n26642 );
or ( n26781 , n26779 , n26780 );
and ( n26782 , n22150 , n22243 );
and ( n26783 , n22111 , n22225 );
nor ( n26784 , n26782 , n26783 );
not ( n26785 , n26656 );
not ( n26786 , n21646 );
or ( n26787 , n26785 , n26786 );
nand ( n26788 , n21577 , n21595 );
nand ( n26789 , n26787 , n26788 );
xor ( n26790 , n26784 , n26789 );
and ( n26791 , n26743 , n22299 );
and ( n26792 , n22268 , n22041 );
not ( n26793 , n22268 );
and ( n26794 , n26793 , n22038 );
nor ( n26795 , n26792 , n26794 );
not ( n26796 , n26795 );
and ( n26797 , n26796 , n22266 );
nor ( n26798 , n26791 , n26797 );
xor ( n26799 , n26790 , n26798 );
xor ( n26800 , n26781 , n26799 );
xor ( n26801 , n26753 , n26669 );
and ( n26802 , n26801 , n26772 );
and ( n26803 , n26753 , n26669 );
nor ( n26804 , n26802 , n26803 );
xor ( n26805 , n26800 , n26804 );
nand ( n26806 , n26777 , n26805 );
not ( n26807 , n26806 );
not ( n26808 , n22299 );
not ( n26809 , n26227 );
or ( n26810 , n26808 , n26809 );
and ( n26811 , n22268 , n21543 );
not ( n26812 , n22268 );
and ( n26813 , n26812 , n21546 );
nor ( n26814 , n26811 , n26813 );
nand ( n26815 , n26814 , n22266 );
nand ( n26816 , n26810 , n26815 );
or ( n26817 , n22166 , n22134 );
nand ( n26818 , n26817 , n22137 );
not ( n26819 , n22225 );
not ( n26820 , n21456 );
or ( n26821 , n26819 , n26820 );
nand ( n26822 , n22974 , n22243 );
nand ( n26823 , n26821 , n26822 );
xor ( n26824 , n26818 , n26823 );
not ( n26825 , n22266 );
and ( n26826 , n22268 , n21768 );
not ( n26827 , n22268 );
and ( n26828 , n26827 , n21769 );
nor ( n26829 , n26826 , n26828 );
not ( n26830 , n26829 );
or ( n26831 , n26825 , n26830 );
nand ( n26832 , n26814 , n22299 );
nand ( n26833 , n26831 , n26832 );
xor ( n26834 , n26824 , n26833 );
xor ( n26835 , n26816 , n26834 );
not ( n26836 , n22225 );
not ( n26837 , n22974 );
or ( n26838 , n26836 , n26837 );
or ( n26839 , n21637 , n22242 );
nand ( n26840 , n26838 , n26839 );
not ( n26841 , n22166 );
not ( n26842 , n26310 );
or ( n26843 , n26841 , n26842 );
nand ( n26844 , n22134 , n22137 );
nand ( n26845 , n26843 , n26844 );
xor ( n26846 , n26840 , n26845 );
not ( n26847 , n21577 );
not ( n26848 , n21595 );
not ( n26849 , n21831 );
or ( n26850 , n26848 , n26849 );
nand ( n26851 , n21830 , n21623 );
nand ( n26852 , n26850 , n26851 );
not ( n26853 , n26852 );
or ( n26854 , n26847 , n26853 );
nand ( n26855 , n26200 , n21646 );
nand ( n26856 , n26854 , n26855 );
and ( n26857 , n26846 , n26856 );
and ( n26858 , n26840 , n26845 );
or ( n26859 , n26857 , n26858 );
and ( n26860 , n26835 , n26859 );
and ( n26861 , n26816 , n26834 );
or ( n26862 , n26860 , n26861 );
not ( n26863 , n21837 );
not ( n26864 , n21651 );
not ( n26865 , n22021 );
or ( n26866 , n26864 , n26865 );
nand ( n26867 , n22018 , n21834 );
nand ( n26868 , n26866 , n26867 );
not ( n26869 , n26868 );
or ( n26870 , n26863 , n26869 );
not ( n26871 , n21651 );
not ( n26872 , n22041 );
or ( n26873 , n26871 , n26872 );
nand ( n26874 , n22038 , n21834 );
nand ( n26875 , n26873 , n26874 );
nand ( n26876 , n26875 , n21698 );
nand ( n26877 , n26870 , n26876 );
not ( n26878 , n19316 );
and ( n26879 , n19319 , n22111 );
not ( n26880 , n19319 );
and ( n26881 , n26880 , n22114 );
nor ( n26882 , n26879 , n26881 );
not ( n26883 , n26882 );
or ( n26884 , n26878 , n26883 );
not ( n26885 , n19319 );
not ( n26886 , n22086 );
or ( n26887 , n26885 , n26886 );
nand ( n26888 , n22083 , n19318 );
nand ( n26889 , n26887 , n26888 );
nand ( n26890 , n26889 , n21549 );
nand ( n26891 , n26884 , n26890 );
xor ( n26892 , n26877 , n26891 );
not ( n26893 , n21646 );
not ( n26894 , n26852 );
or ( n26895 , n26893 , n26894 );
not ( n26896 , n21595 );
not ( n26897 , n22153 );
or ( n26898 , n26896 , n26897 );
nand ( n26899 , n21623 , n22150 );
nand ( n26900 , n26898 , n26899 );
nand ( n26901 , n26900 , n21577 );
nand ( n26902 , n26895 , n26901 );
and ( n26903 , n26892 , n26902 );
and ( n26904 , n26877 , n26891 );
or ( n26905 , n26903 , n26904 );
not ( n26906 , n21698 );
not ( n26907 , n26868 );
or ( n26908 , n26906 , n26907 );
nand ( n26909 , n21837 , n21651 );
nand ( n26910 , n26908 , n26909 );
not ( n26911 , n21549 );
not ( n26912 , n26711 );
or ( n26913 , n26911 , n26912 );
nand ( n26914 , n26889 , n19316 );
nand ( n26915 , n26913 , n26914 );
xor ( n26916 , n26910 , n26915 );
not ( n26917 , n22266 );
not ( n26918 , n26684 );
or ( n26919 , n26917 , n26918 );
nand ( n26920 , n26829 , n22299 );
nand ( n26921 , n26919 , n26920 );
xor ( n26922 , n26916 , n26921 );
xor ( n26923 , n26905 , n26922 );
not ( n26924 , n26705 );
not ( n26925 , n21577 );
not ( n26926 , n26722 );
or ( n26927 , n26925 , n26926 );
nand ( n26928 , n26900 , n21646 );
nand ( n26929 , n26927 , n26928 );
xor ( n26930 , n26924 , n26929 );
xor ( n26931 , n26818 , n26823 );
and ( n26932 , n26931 , n26833 );
and ( n26933 , n26818 , n26823 );
or ( n26934 , n26932 , n26933 );
xor ( n26935 , n26930 , n26934 );
xor ( n26936 , n26923 , n26935 );
xor ( n26937 , n26862 , n26936 );
xor ( n26938 , n26877 , n26891 );
xor ( n26939 , n26938 , n26902 );
not ( n26940 , n26939 );
not ( n26941 , n19316 );
not ( n26942 , n26236 );
or ( n26943 , n26941 , n26942 );
nand ( n26944 , n26882 , n21549 );
nand ( n26945 , n26943 , n26944 );
not ( n26946 , n21837 );
not ( n26947 , n26875 );
or ( n26948 , n26946 , n26947 );
nand ( n26949 , n26300 , n21698 );
nand ( n26950 , n26948 , n26949 );
or ( n26951 , n26945 , n26950 );
not ( n26952 , n26816 );
nand ( n26953 , n26951 , n26952 );
nand ( n26954 , n26945 , n26950 );
nand ( n26955 , n26953 , n26954 );
not ( n26956 , n26955 );
nand ( n26957 , n26940 , n26956 );
not ( n26958 , n26957 );
xor ( n26959 , n26816 , n26834 );
xor ( n26960 , n26959 , n26859 );
not ( n26961 , n26960 );
or ( n26962 , n26958 , n26961 );
nand ( n26963 , n26939 , n26955 );
nand ( n26964 , n26962 , n26963 );
xor ( n26965 , n26937 , n26964 );
xor ( n26966 , n26214 , n26229 );
and ( n26967 , n26966 , n26244 );
and ( n26968 , n26214 , n26229 );
or ( n26969 , n26967 , n26968 );
not ( n26970 , n26969 );
not ( n26971 , n26970 );
xor ( n26972 , n26945 , n26950 );
and ( n26973 , n26972 , n26816 );
not ( n26974 , n26972 );
and ( n26975 , n26974 , n26952 );
nor ( n26976 , n26973 , n26975 );
not ( n26977 , n26976 );
or ( n26978 , n26971 , n26977 );
xor ( n26979 , n26191 , n26193 );
and ( n26980 , n26979 , n26208 );
and ( n26981 , n26191 , n26193 );
or ( n26982 , n26980 , n26981 );
nand ( n26983 , n26978 , n26982 );
not ( n26984 , n26976 );
nand ( n26985 , n26984 , n26969 );
nand ( n26986 , n26983 , n26985 );
not ( n26987 , n26986 );
not ( n26988 , n26987 );
xor ( n26989 , n26956 , n26939 );
xor ( n26990 , n26989 , n26960 );
not ( n26991 , n26990 );
or ( n26992 , n26988 , n26991 );
xor ( n26993 , n26840 , n26845 );
xor ( n26994 , n26993 , n26856 );
xor ( n26995 , n26302 , n26312 );
and ( n26996 , n26995 , n26328 );
and ( n26997 , n26302 , n26312 );
or ( n26998 , n26996 , n26997 );
xor ( n26999 , n26994 , n26998 );
xor ( n27000 , n26209 , n26245 );
and ( n27001 , n27000 , n26264 );
and ( n27002 , n26209 , n26245 );
or ( n27003 , n27001 , n27002 );
and ( n27004 , n26999 , n27003 );
and ( n27005 , n26994 , n26998 );
or ( n27006 , n27004 , n27005 );
nand ( n27007 , n26992 , n27006 );
not ( n27008 , n26990 );
nand ( n27009 , n27008 , n26986 );
nand ( n27010 , n27007 , n27009 );
or ( n27011 , n26965 , n27010 );
xor ( n27012 , n26862 , n26936 );
and ( n27013 , n27012 , n26964 );
and ( n27014 , n26862 , n26936 );
or ( n27015 , n27013 , n27014 );
xor ( n27016 , n26924 , n26929 );
and ( n27017 , n27016 , n26934 );
and ( n27018 , n26924 , n26929 );
or ( n27019 , n27017 , n27018 );
xor ( n27020 , n26905 , n26922 );
and ( n27021 , n27020 , n26935 );
and ( n27022 , n26905 , n26922 );
or ( n27023 , n27021 , n27022 );
xor ( n27024 , n27019 , n27023 );
not ( n27025 , n26674 );
not ( n27026 , n26677 );
and ( n27027 , n27025 , n27026 );
and ( n27028 , n26674 , n26677 );
nor ( n27029 , n27027 , n27028 );
not ( n27030 , n27029 );
not ( n27031 , n26693 );
or ( n27032 , n27030 , n27031 );
or ( n27033 , n26693 , n27029 );
nand ( n27034 , n27032 , n27033 );
xor ( n27035 , n26705 , n26715 );
xor ( n27036 , n27035 , n26731 );
xor ( n27037 , n27034 , n27036 );
xor ( n27038 , n26910 , n26915 );
and ( n27039 , n27038 , n26921 );
and ( n27040 , n26910 , n26915 );
or ( n27041 , n27039 , n27040 );
xor ( n27042 , n27037 , n27041 );
xor ( n27043 , n27024 , n27042 );
nor ( n27044 , n27015 , n27043 );
not ( n27045 , n27044 );
and ( n27046 , n27011 , n27045 );
xor ( n27047 , n27019 , n27023 );
and ( n27048 , n27047 , n27042 );
and ( n27049 , n27019 , n27023 );
or ( n27050 , n27048 , n27049 );
not ( n27051 , n27050 );
xor ( n27052 , n26759 , n26764 );
xor ( n27053 , n27052 , n26769 );
not ( n27054 , n27053 );
not ( n27055 , n27054 );
xor ( n27056 , n26669 , n26699 );
xor ( n27057 , n27056 , n26735 );
not ( n27058 , n27057 );
not ( n27059 , n27058 );
or ( n27060 , n27055 , n27059 );
nand ( n27061 , n27057 , n27053 );
nand ( n27062 , n27060 , n27061 );
xor ( n27063 , n27034 , n27036 );
and ( n27064 , n27063 , n27041 );
and ( n27065 , n27034 , n27036 );
or ( n27066 , n27064 , n27065 );
not ( n27067 , n27066 );
xor ( n27068 , n27062 , n27067 );
nand ( n27069 , n27051 , n27068 );
not ( n27070 , n27054 );
not ( n27071 , n27057 );
or ( n27072 , n27070 , n27071 );
nand ( n27073 , n27072 , n27066 );
nand ( n27074 , n27058 , n27053 );
nand ( n27075 , n27073 , n27074 );
not ( n27076 , n27075 );
xor ( n27077 , n26659 , n26738 );
xor ( n27078 , n27077 , n26774 );
nand ( n27079 , n27076 , n27078 );
nand ( n27080 , n27069 , n27079 );
not ( n27081 , n27080 );
and ( n27082 , n27046 , n27081 );
not ( n27083 , n27082 );
not ( n27084 , n26970 );
not ( n27085 , n26982 );
and ( n27086 , n27084 , n27085 );
and ( n27087 , n26970 , n26982 );
nor ( n27088 , n27086 , n27087 );
and ( n27089 , n27088 , n26984 );
not ( n27090 , n27088 );
and ( n27091 , n27090 , n26976 );
nor ( n27092 , n27089 , n27091 );
xor ( n27093 , n26994 , n26998 );
xor ( n27094 , n27093 , n27003 );
xor ( n27095 , n27092 , n27094 );
xor ( n27096 , n26292 , n26329 );
and ( n27097 , n27096 , n26342 );
and ( n27098 , n26292 , n26329 );
or ( n27099 , n27097 , n27098 );
xor ( n27100 , n27095 , n27099 );
or ( n27101 , n26265 , n26343 );
and ( n27102 , n27101 , n26362 );
and ( n27103 , n26265 , n26343 );
nor ( n27104 , n27102 , n27103 );
nand ( n27105 , n27100 , n27104 );
not ( n27106 , n27092 );
not ( n27107 , n27094 );
not ( n27108 , n27107 );
or ( n27109 , n27106 , n27108 );
nand ( n27110 , n27109 , n27099 );
not ( n27111 , n27092 );
nand ( n27112 , n27111 , n27094 );
nand ( n27113 , n27110 , n27112 );
not ( n27114 , n27113 );
xor ( n27115 , n26987 , n27006 );
xor ( n27116 , n27115 , n27008 );
nand ( n27117 , n27114 , n27116 );
nand ( n27118 , n26378 , n26398 , n27105 , n27117 );
not ( n27119 , n27118 );
not ( n27120 , n27119 );
not ( n27121 , n26391 );
or ( n27122 , n27120 , n27121 );
not ( n27123 , n27117 );
not ( n27124 , n27105 );
or ( n27125 , n26377 , n26400 );
nand ( n27126 , n27125 , n26376 );
not ( n27127 , n27126 );
or ( n27128 , n27124 , n27127 );
or ( n27129 , n27100 , n27104 );
nand ( n27130 , n27128 , n27129 );
not ( n27131 , n27130 );
or ( n27132 , n27123 , n27131 );
not ( n27133 , n27116 );
nand ( n27134 , n27133 , n27113 );
nand ( n27135 , n27132 , n27134 );
not ( n27136 , n27135 );
nand ( n27137 , n27122 , n27136 );
not ( n27138 , n27137 );
or ( n27139 , n27083 , n27138 );
nand ( n27140 , n26965 , n27010 );
or ( n27141 , n27140 , n27044 );
nand ( n27142 , n27015 , n27043 );
nand ( n27143 , n27141 , n27142 );
and ( n27144 , n27143 , n27081 );
not ( n27145 , n27068 );
nand ( n27146 , n27145 , n27050 );
not ( n27147 , n27079 );
or ( n27148 , n27146 , n27147 );
not ( n27149 , n27078 );
nand ( n27150 , n27149 , n27075 );
nand ( n27151 , n27148 , n27150 );
nor ( n27152 , n27144 , n27151 );
nand ( n27153 , n27139 , n27152 );
not ( n27154 , n27153 );
or ( n27155 , n26807 , n27154 );
nor ( n27156 , n26777 , n26805 );
not ( n27157 , n27156 );
nand ( n27158 , n27155 , n27157 );
xor ( n27159 , n26781 , n26799 );
and ( n27160 , n27159 , n26804 );
and ( n27161 , n26781 , n26799 );
or ( n27162 , n27160 , n27161 );
not ( n27163 , n26789 );
and ( n27164 , n23170 , n21576 );
nor ( n27165 , n27164 , n21623 );
not ( n27166 , n22114 );
not ( n27167 , n22242 );
and ( n27168 , n27166 , n27167 );
and ( n27169 , n22083 , n22225 );
nor ( n27170 , n27168 , n27169 );
xor ( n27171 , n27165 , n27170 );
or ( n27172 , n26795 , n22934 );
and ( n27173 , n22268 , n22021 );
not ( n27174 , n22268 );
and ( n27175 , n27174 , n22018 );
nor ( n27176 , n27173 , n27175 );
or ( n27177 , n27176 , n22265 );
nand ( n27178 , n27172 , n27177 );
not ( n27179 , n27178 );
xor ( n27180 , n27171 , n27179 );
xor ( n27181 , n27163 , n27180 );
xor ( n27182 , n26784 , n26789 );
and ( n27183 , n27182 , n26798 );
and ( n27184 , n26784 , n26789 );
or ( n27185 , n27183 , n27184 );
xor ( n27186 , n27181 , n27185 );
nor ( n27187 , n27162 , n27186 );
not ( n27188 , n27187 );
nand ( n27189 , n27162 , n27186 );
nand ( n27190 , n27188 , n27189 );
xnor ( n27191 , n27158 , n27190 );
nand ( n27192 , n26635 , n27191 );
not ( n27193 , n19220 );
and ( n27194 , n26153 , n471 );
xor ( n27195 , n26160 , n26162 );
and ( n27196 , n27195 , n26164 );
and ( n27197 , n26160 , n26162 );
or ( n27198 , n27196 , n27197 );
xor ( n27199 , n27194 , n27198 );
and ( n27200 , n26079 , n470 );
not ( n27201 , n19129 );
nor ( n27202 , n27201 , n17873 );
xor ( n27203 , n27200 , n27202 );
not ( n27204 , n454 );
nor ( n27205 , n26068 , n26126 );
not ( n27206 , n27205 );
nor ( n27207 , n27206 , n19121 );
or ( n27208 , n26070 , n26126 );
nand ( n27209 , n27208 , n26128 );
nor ( n27210 , n27207 , n27209 );
xor ( n27211 , n26104 , n26119 );
and ( n27212 , n27211 , n26124 );
and ( n27213 , n26104 , n26119 );
or ( n27214 , n27212 , n27213 );
not ( n27215 , n26118 );
or ( n27216 , n3103 , n3026 );
nand ( n27217 , n27216 , n539 );
not ( n27218 , n11729 );
not ( n27219 , n26110 );
or ( n27220 , n27218 , n27219 );
xor ( n27221 , n537 , n17971 );
nand ( n27222 , n3186 , n27221 );
nand ( n27223 , n27220 , n27222 );
xor ( n27224 , n27217 , n27223 );
and ( n27225 , n537 , n14354 );
xor ( n27226 , n27224 , n27225 );
xor ( n27227 , n27215 , n27226 );
xor ( n27228 , n26114 , n26115 );
and ( n27229 , n27228 , n26118 );
and ( n27230 , n26114 , n26115 );
or ( n27231 , n27229 , n27230 );
xor ( n27232 , n27227 , n27231 );
nor ( n27233 , n27214 , n27232 );
not ( n27234 , n27233 );
nand ( n27235 , n27214 , n27232 );
and ( n27236 , n27234 , n27235 );
and ( n27237 , n27210 , n27236 );
not ( n27238 , n27237 );
nor ( n27239 , n27206 , n26021 );
nand ( n27240 , n19075 , n27239 );
not ( n27241 , n27240 );
or ( n27242 , n27238 , n27241 );
not ( n27243 , n27210 );
not ( n27244 , n27240 );
or ( n27245 , n27243 , n27244 );
not ( n27246 , n27236 );
nand ( n27247 , n27245 , n27246 );
nand ( n27248 , n27242 , n27247 );
not ( n27249 , n27248 );
or ( n27250 , n27204 , n27249 );
nand ( n27251 , n27250 , n17645 );
and ( n27252 , n27251 , n472 );
xor ( n27253 , n27203 , n27252 );
xor ( n27254 , n27199 , n27253 );
xor ( n27255 , n26154 , n26158 );
and ( n27256 , n27255 , n26165 );
and ( n27257 , n26154 , n26158 );
or ( n27258 , n27256 , n27257 );
or ( n27259 , n27254 , n27258 );
nand ( n27260 , n27254 , n27258 );
buf ( n27261 , n27260 );
nand ( n27262 , n27259 , n27261 );
not ( n27263 , n27262 );
or ( n27264 , n26085 , n26002 );
or ( n27265 , n26166 , n26170 );
nand ( n27266 , n27264 , n27265 );
nor ( n27267 , n27266 , n25987 );
not ( n27268 , n27267 );
nand ( n27269 , n18188 , n18423 , n18974 , n18989 );
not ( n27270 , n27269 );
or ( n27271 , n27268 , n27270 );
not ( n27272 , n26085 );
not ( n27273 , n26002 );
and ( n27274 , n27272 , n27273 );
not ( n27275 , n26166 );
not ( n27276 , n26170 );
and ( n27277 , n27275 , n27276 );
nor ( n27278 , n27274 , n27277 );
nand ( n27279 , n25995 , n27278 );
nor ( n27280 , n26171 , n26086 );
not ( n27281 , n27280 );
nand ( n27282 , n27279 , n27281 , n26174 );
not ( n27283 , n27282 );
nand ( n27284 , n27271 , n27283 );
not ( n27285 , n27284 );
or ( n27286 , n27263 , n27285 );
or ( n27287 , n27262 , n27284 );
nand ( n27288 , n27286 , n27287 );
not ( n27289 , n27288 );
or ( n27290 , n27193 , n27289 );
not ( n27291 , n19220 );
and ( n27292 , n27129 , n27105 );
not ( n27293 , n27292 );
nor ( n27294 , n26399 , n26377 );
or ( n27295 , n27294 , n27126 );
not ( n27296 , n27295 );
not ( n27297 , n27296 );
or ( n27298 , n27293 , n27297 );
or ( n27299 , n27296 , n27292 );
nand ( n27300 , n27298 , n27299 );
nand ( n27301 , n27291 , n27300 );
nand ( n27302 , n27290 , n27301 );
not ( n27303 , n25605 );
nand ( n27304 , n27303 , n25654 );
xor ( n27305 , n25652 , n27304 );
and ( n27306 , n26561 , n27305 );
not ( n27307 , n26561 );
not ( n27308 , n18880 );
not ( n27309 , n27308 );
not ( n27310 , n18852 );
nand ( n27311 , n27310 , n18882 );
not ( n27312 , n27311 );
or ( n27313 , n27309 , n27312 );
or ( n27314 , n27308 , n27311 );
nand ( n27315 , n27313 , n27314 );
and ( n27316 , n27307 , n27315 );
or ( n27317 , n27306 , n27316 );
nor ( n27318 , n22021 , n22242 );
not ( n27319 , n27318 );
and ( n27320 , n22038 , n22243 );
and ( n27321 , n22018 , n22225 );
nor ( n27322 , n27320 , n27321 );
and ( n27323 , n22934 , n22265 );
nor ( n27324 , n27323 , n22277 );
xor ( n27325 , n27322 , n27324 );
not ( n27326 , n22041 );
not ( n27327 , n22224 );
and ( n27328 , n27326 , n27327 );
and ( n27329 , n22083 , n22243 );
nor ( n27330 , n27328 , n27329 );
and ( n27331 , n27325 , n27330 );
and ( n27332 , n27322 , n27324 );
or ( n27333 , n27331 , n27332 );
not ( n27334 , n27333 );
or ( n27335 , n27319 , n27334 );
or ( n27336 , n27333 , n27318 );
nand ( n27337 , n27335 , n27336 );
not ( n27338 , n27337 );
or ( n27339 , n27176 , n22934 );
or ( n27340 , n22265 , n22277 );
nand ( n27341 , n27339 , n27340 );
xor ( n27342 , n27341 , n27330 );
xor ( n27343 , n27165 , n27170 );
and ( n27344 , n27343 , n27179 );
and ( n27345 , n27165 , n27170 );
or ( n27346 , n27344 , n27345 );
not ( n27347 , n27346 );
and ( n27348 , n27342 , n27347 );
and ( n27349 , n27341 , n27330 );
or ( n27350 , n27348 , n27349 );
not ( n27351 , n27350 );
xor ( n27352 , n27322 , n27324 );
xor ( n27353 , n27352 , n27330 );
nand ( n27354 , n27351 , n27353 );
xor ( n27355 , n27341 , n27330 );
not ( n27356 , n27346 );
xor ( n27357 , n27355 , n27356 );
not ( n27358 , n27357 );
xor ( n27359 , n27163 , n27180 );
and ( n27360 , n27359 , n27185 );
and ( n27361 , n27163 , n27180 );
or ( n27362 , n27360 , n27361 );
nand ( n27363 , n27358 , n27362 );
nand ( n27364 , n26806 , n27189 , n27363 );
nor ( n27365 , n27080 , n27364 );
nand ( n27366 , n27046 , n27354 , n27365 );
nor ( n27367 , n27366 , n27118 );
not ( n27368 , n27367 );
not ( n27369 , n26391 );
or ( n27370 , n27368 , n27369 );
not ( n27371 , n27366 );
and ( n27372 , n27135 , n27371 );
not ( n27373 , n27354 );
not ( n27374 , n27365 );
not ( n27375 , n27143 );
or ( n27376 , n27374 , n27375 );
not ( n27377 , n27364 );
and ( n27378 , n27151 , n27377 );
and ( n27379 , n27189 , n27156 );
nor ( n27380 , n27379 , n27187 );
not ( n27381 , n27363 );
or ( n27382 , n27380 , n27381 );
not ( n27383 , n27362 );
nand ( n27384 , n27383 , n27357 );
nand ( n27385 , n27382 , n27384 );
nor ( n27386 , n27378 , n27385 );
nand ( n27387 , n27376 , n27386 );
not ( n27388 , n27387 );
or ( n27389 , n27373 , n27388 );
or ( n27390 , n27351 , n27353 );
nand ( n27391 , n27389 , n27390 );
nor ( n27392 , n27372 , n27391 );
nand ( n27393 , n27370 , n27392 );
not ( n27394 , n27393 );
or ( n27395 , n27338 , n27394 );
or ( n27396 , n27337 , n27393 );
nand ( n27397 , n27395 , n27396 );
not ( n27398 , n27397 );
nor ( n27399 , n27398 , n19220 );
xor ( n27400 , n27217 , n27223 );
and ( n27401 , n27400 , n27225 );
and ( n27402 , n27217 , n27223 );
or ( n27403 , n27401 , n27402 );
xor ( n27404 , n27215 , n27226 );
and ( n27405 , n27404 , n27231 );
and ( n27406 , n27215 , n27226 );
or ( n27407 , n27405 , n27406 );
not ( n27408 , n27221 );
or ( n27409 , n27408 , n14865 );
or ( n27410 , n10598 , n3177 );
nand ( n27411 , n27409 , n27410 );
nand ( n27412 , n14326 , n537 );
xor ( n27413 , n27411 , n27412 );
xor ( n27414 , n27413 , n27403 );
xor ( n27415 , n27411 , n27412 );
and ( n27416 , n27415 , n27403 );
and ( n27417 , n27411 , n27412 );
or ( n27418 , n27416 , n27417 );
not ( n27419 , n27209 );
not ( n27420 , n27234 );
or ( n27421 , n27419 , n27420 );
nand ( n27422 , n27421 , n27235 );
nor ( n27423 , n27207 , n27422 );
not ( n27424 , n27214 );
not ( n27425 , n27232 );
and ( n27426 , n27424 , n27425 );
nor ( n27427 , n27407 , n27414 );
nor ( n27428 , n27426 , n27427 );
nand ( n27429 , n27205 , n27428 );
or ( n27430 , n27429 , n19121 );
nand ( n27431 , n27407 , n27414 );
nand ( n27432 , n27430 , n27431 );
not ( n27433 , n6583 );
not ( n27434 , n6586 );
nand ( n27435 , n27434 , n6562 );
not ( n27436 , n27435 );
or ( n27437 , n27433 , n27436 );
or ( n27438 , n6583 , n27435 );
nand ( n27439 , n27437 , n27438 );
xor ( n27440 , n6564 , n6575 );
xor ( n27441 , n27440 , n6580 );
and ( n27442 , n6572 , n6574 );
nor ( n27443 , n27442 , n6575 );
or ( n27444 , n11729 , n3186 );
nand ( n27445 , n27444 , n537 );
not ( n27446 , n27412 );
and ( n27447 , n537 , n17971 );
not ( n27448 , n6573 );
not ( n27449 , n27422 );
nand ( n27450 , n27449 , n27233 );
xor ( n27451 , n27445 , n27447 );
xor ( n27452 , n27451 , n27446 );
and ( n27454 , n27158 , n27189 );
nor ( n27455 , n27454 , n27187 );
nand ( n27456 , n27354 , n27390 );
not ( n27457 , n27456 );
not ( n27458 , n27365 );
not ( n27459 , n27046 );
not ( n27460 , n27137 );
or ( n27461 , n27459 , n27460 );
not ( n27462 , n27143 );
nand ( n27463 , n27461 , n27462 );
not ( n27464 , n27463 );
or ( n27465 , n27458 , n27464 );
nand ( n27466 , n27465 , n27386 );
not ( n27467 , n27466 );
or ( n27468 , n27457 , n27467 );
or ( n27469 , n27456 , n27466 );
nand ( n27470 , n27468 , n27469 );
not ( n27471 , n27153 );
not ( n27472 , n27069 );
not ( n27473 , n27463 );
or ( n27474 , n27472 , n27473 );
nand ( n27475 , n27474 , n27146 );
nand ( n27476 , n27295 , n27105 );
nand ( n27477 , n27476 , n27129 );
not ( n27478 , n27137 );
not ( n27479 , n27011 );
or ( n27480 , n27478 , n27479 );
nand ( n27481 , n27480 , n27140 );
or ( n27482 , n26554 , n25829 );
nand ( n27483 , n27482 , n25861 );
not ( n27484 , n23823 );
not ( n27485 , n25780 );
or ( n27486 , n27484 , n27485 );
not ( n27487 , n25783 );
nand ( n27488 , n27486 , n27487 );
nor ( n27489 , n25776 , n25913 );
and ( n27490 , n27489 , n25773 );
not ( n27491 , n27489 );
and ( n27492 , n27491 , n25912 );
nor ( n27493 , n27490 , n27492 );
not ( n27494 , n25688 );
nand ( n27495 , n27494 , n25693 );
not ( n27496 , n27495 );
nand ( n27497 , n25676 , n25691 );
not ( n27498 , n27497 );
or ( n27499 , n27496 , n27498 );
or ( n27500 , n27497 , n27495 );
nand ( n27501 , n27499 , n27500 );
not ( n27502 , n25858 );
nand ( n27503 , n27502 , n25863 );
not ( n27504 , n25785 );
nand ( n27505 , n27504 , n23591 );
and ( n27506 , n25886 , n25883 );
not ( n27507 , n25675 );
nand ( n27508 , n25691 , n25405 );
not ( n27509 , n27508 );
or ( n27510 , n27507 , n27509 );
or ( n27511 , n27508 , n25675 );
nand ( n27512 , n27510 , n27511 );
nand ( n27513 , n27487 , n23823 );
xor ( n27514 , n25426 , n25428 );
xor ( n27515 , n27514 , n25672 );
not ( n27516 , n25667 );
nand ( n27517 , n25671 , n25465 );
not ( n27518 , n27517 );
or ( n27519 , n27516 , n27518 );
or ( n27520 , n27517 , n25667 );
nand ( n27521 , n27519 , n27520 );
nand ( n27522 , n27134 , n27117 );
not ( n27523 , n27140 );
nor ( n27524 , n27523 , n27479 );
not ( n27525 , n25659 );
nand ( n27526 , n25663 , n25577 );
not ( n27527 , n27526 );
or ( n27528 , n27525 , n27527 );
or ( n27529 , n27526 , n25659 );
nand ( n27530 , n27528 , n27529 );
nand ( n27531 , n27146 , n27069 );
not ( n27532 , n27147 );
nand ( n27533 , n27532 , n27150 );
nand ( n27534 , n27045 , n27142 );
and ( n27535 , n26806 , n27157 );
nand ( n27536 , n27363 , n27384 );
not ( n27537 , n25643 );
not ( n27538 , n25649 );
not ( n27539 , n25646 );
or ( n27540 , n27538 , n27539 );
or ( n27541 , n25646 , n25649 );
nand ( n27542 , n27540 , n27541 );
not ( n27543 , n27542 );
or ( n27544 , n27537 , n27543 );
or ( n27545 , n27542 , n25643 );
nand ( n27546 , n27544 , n27545 );
xor ( n27547 , n25606 , n25617 );
xor ( n27548 , n27547 , n25640 );
xor ( n27549 , n25619 , n25631 );
xor ( n27550 , n27549 , n25637 );
xnor ( n27551 , n27477 , n27522 );
xor ( n27552 , n27455 , n27536 );
xor ( n27554 , n17589 , n17599 );
and ( n27555 , n27554 , n17604 );
and ( n27556 , n17589 , n17599 );
or ( n27557 , n27555 , n27556 );
xor ( n27558 , n17616 , n17620 );
and ( n27559 , n27558 , n17625 );
and ( n27560 , n17616 , n17620 );
or ( n27561 , n27559 , n27560 );
xor ( n27562 , n17605 , n17626 );
and ( n27563 , n27562 , n17631 );
and ( n27564 , n17605 , n17626 );
or ( n27565 , n27563 , n27564 );
or ( n27566 , n7405 , n7371 );
nand ( n27567 , n27566 , n493 );
and ( n27568 , n489 , n15788 );
xor ( n27569 , n27567 , n27568 );
not ( n27570 , n6867 );
not ( n27571 , n17610 );
or ( n27572 , n27570 , n27571 );
xor ( n27573 , n489 , n15904 );
nand ( n27574 , n27573 , n6848 );
nand ( n27575 , n27572 , n27574 );
xor ( n27576 , n27569 , n27575 );
xor ( n27577 , n27567 , n27568 );
and ( n27578 , n27577 , n27575 );
and ( n27579 , n27567 , n27568 );
or ( n27580 , n27578 , n27579 );
not ( n27581 , n6842 );
and ( n27582 , n491 , n15760 );
not ( n27583 , n491 );
and ( n27584 , n27583 , n15761 );
or ( n27585 , n27582 , n27584 );
not ( n27586 , n27585 );
or ( n27587 , n27581 , n27586 );
nand ( n27588 , n17595 , n6719 );
nand ( n27589 , n27587 , n27588 );
not ( n27590 , n17616 );
xor ( n27591 , n27589 , n27590 );
xor ( n27592 , n27591 , n27576 );
xor ( n27593 , n27589 , n27590 );
and ( n27594 , n27593 , n27576 );
and ( n27595 , n27589 , n27590 );
or ( n27596 , n27594 , n27595 );
xor ( n27597 , n27557 , n27592 );
xor ( n27598 , n27597 , n27561 );
xor ( n27599 , n27557 , n27592 );
and ( n27600 , n27599 , n27561 );
and ( n27601 , n27557 , n27592 );
or ( n27602 , n27600 , n27601 );
not ( n27603 , n6848 );
not ( n27604 , n489 );
not ( n27605 , n15886 );
or ( n27606 , n27604 , n27605 );
nand ( n27607 , n15887 , n4046 );
nand ( n27608 , n27606 , n27607 );
not ( n27609 , n27608 );
or ( n27610 , n27603 , n27609 );
nand ( n27611 , n27573 , n6867 );
nand ( n27612 , n27610 , n27611 );
not ( n27613 , n6719 );
not ( n27614 , n27585 );
or ( n27615 , n27613 , n27614 );
nand ( n27616 , n27615 , n12976 );
xor ( n27617 , n27612 , n27616 );
nand ( n27618 , n15844 , n489 );
xor ( n27619 , n27617 , n27618 );
xor ( n27620 , n27612 , n27616 );
and ( n27621 , n27620 , n27618 );
and ( n27622 , n27612 , n27616 );
or ( n27623 , n27621 , n27622 );
xor ( n27624 , n27580 , n27619 );
xor ( n27625 , n27624 , n27596 );
xor ( n27626 , n27580 , n27619 );
and ( n27627 , n27626 , n27596 );
and ( n27628 , n27580 , n27619 );
or ( n27629 , n27627 , n27628 );
or ( n27630 , n6719 , n6842 );
nand ( n27631 , n27630 , n491 );
and ( n27632 , n489 , n15904 );
xor ( n27633 , n27631 , n27632 );
not ( n27634 , n6867 );
not ( n27635 , n27608 );
or ( n27636 , n27634 , n27635 );
xor ( n27637 , n489 , n15761 );
nand ( n27638 , n27637 , n6848 );
nand ( n27639 , n27636 , n27638 );
xor ( n27640 , n27633 , n27639 );
xor ( n27641 , n27631 , n27632 );
and ( n27642 , n27641 , n27639 );
and ( n27643 , n27631 , n27632 );
or ( n27644 , n27642 , n27643 );
not ( n27645 , n27618 );
xor ( n27646 , n27645 , n27640 );
xor ( n27647 , n27646 , n27623 );
xor ( n27648 , n27645 , n27640 );
and ( n27649 , n27648 , n27623 );
and ( n27650 , n27645 , n27640 );
or ( n27651 , n27649 , n27650 );
not ( n27652 , n27637 );
or ( n27653 , n27652 , n7355 );
or ( n27654 , n6898 , n4046 );
nand ( n27655 , n27653 , n27654 );
not ( n27656 , n15886 );
nand ( n27657 , n27656 , n489 );
xor ( n27658 , n27655 , n27657 );
xor ( n27659 , n27658 , n27644 );
xor ( n27660 , n27655 , n27657 );
and ( n27661 , n27660 , n27644 );
and ( n27662 , n27655 , n27657 );
or ( n27663 , n27661 , n27662 );
not ( n27664 , n17576 );
nor ( n27665 , n27565 , n27598 );
not ( n27666 , n27665 );
nand ( n27667 , n27666 , n16206 , n17637 );
nor ( n27668 , n27664 , n27667 );
not ( n27669 , n27668 );
not ( n27670 , n17944 );
or ( n27671 , n27669 , n27670 );
or ( n27672 , n16722 , n27667 );
nand ( n27673 , n27671 , n27672 );
not ( n27674 , n17637 );
not ( n27675 , n17585 );
or ( n27676 , n27674 , n27675 );
nand ( n27677 , n27676 , n17638 );
not ( n27678 , n27677 );
or ( n27679 , n27678 , n27665 );
nand ( n27680 , n27598 , n27565 );
nand ( n27681 , n27679 , n27680 );
nor ( n27682 , n27602 , n27625 );
nor ( n27683 , n27665 , n27682 );
or ( n27684 , n27629 , n27647 );
nand ( n27685 , n27683 , n27684 );
not ( n27686 , n27685 );
not ( n27687 , n27686 );
not ( n27688 , n27677 );
or ( n27689 , n27687 , n27688 );
or ( n27690 , n27680 , n27682 );
nand ( n27691 , n27602 , n27625 );
nand ( n27692 , n27690 , n27691 );
and ( n27693 , n27692 , n27684 );
and ( n27694 , n27629 , n27647 );
nor ( n27695 , n27693 , n27694 );
nand ( n27696 , n27689 , n27695 );
not ( n27697 , n27696 );
and ( n27698 , n17637 , n27683 );
and ( n27699 , n17586 , n27698 );
not ( n27700 , n17638 );
not ( n27701 , n27700 );
not ( n27702 , n27683 );
or ( n27703 , n27701 , n27702 );
not ( n27704 , n27692 );
nand ( n27705 , n27703 , n27704 );
nor ( n27706 , n27699 , n27705 );
nand ( n27707 , n27666 , n27680 );
not ( n27708 , n27682 );
nand ( n27709 , n27708 , n27691 );
not ( n27710 , n9792 );
not ( n27711 , n9794 );
nand ( n27712 , n27711 , n9768 );
not ( n27713 , n27712 );
or ( n27714 , n27710 , n27713 );
or ( n27715 , n27712 , n9792 );
nand ( n27716 , n27714 , n27715 );
xor ( n27717 , n9770 , n9783 );
xor ( n27718 , n27717 , n9789 );
and ( n27719 , n9780 , n9782 );
nor ( n27720 , n27719 , n9783 );
or ( n27721 , n6867 , n6848 );
nand ( n27722 , n27721 , n489 );
not ( n27723 , n27657 );
and ( n27724 , n489 , n15761 );
xor ( n27725 , n27722 , n27724 );
xor ( n27726 , n27725 , n27723 );
xor ( n27727 , n27200 , n27202 );
and ( n27728 , n27727 , n27252 );
and ( n27729 , n27200 , n27202 );
or ( n27730 , n27728 , n27729 );
xor ( n27731 , n27194 , n27198 );
and ( n27732 , n27731 , n27253 );
and ( n27733 , n27194 , n27198 );
or ( n27734 , n27732 , n27733 );
and ( n27735 , n26079 , n469 );
nand ( n27736 , n27251 , n471 );
not ( n27737 , n27736 );
xor ( n27738 , n27735 , n27737 );
and ( n27739 , n26152 , n470 );
xor ( n27740 , n27738 , n27739 );
xor ( n27741 , n27735 , n27737 );
and ( n27742 , n27741 , n27739 );
and ( n27743 , n27735 , n27737 );
or ( n27744 , n27742 , n27743 );
not ( n27745 , n27423 );
not ( n27746 , n27240 );
or ( n27747 , n27745 , n27746 );
nand ( n27748 , n27747 , n27450 );
or ( n27749 , n27407 , n27414 );
nand ( n27750 , n27749 , n27431 );
and ( n27751 , n27748 , n27750 );
not ( n27752 , n27748 );
not ( n27753 , n27750 );
and ( n27754 , n27752 , n27753 );
nor ( n27755 , n27751 , n27754 );
nand ( n27756 , n27755 , n454 );
and ( n27757 , n16206 , n17637 );
not ( n27758 , n27757 );
not ( n27759 , n17578 );
or ( n27760 , n27758 , n27759 );
nand ( n27761 , n27760 , n27678 );
xnor ( n27762 , n27761 , n27707 );
nand ( n27763 , n27762 , n9907 );
nand ( n27764 , n27756 , n27763 );
and ( n27765 , n27764 , n472 );
xor ( n27766 , n27765 , n27730 );
xor ( n27767 , n27766 , n27740 );
xor ( n27768 , n27765 , n27730 );
and ( n27769 , n27768 , n27740 );
and ( n27770 , n27765 , n27730 );
or ( n27771 , n27769 , n27770 );
not ( n27772 , n472 );
nor ( n27773 , n27709 , n27681 );
not ( n27774 , n27773 );
not ( n27775 , n27673 );
not ( n27776 , n27775 );
or ( n27777 , n27774 , n27776 );
buf ( n27778 , n27681 );
or ( n27779 , n27778 , n27673 );
nand ( n27780 , n27779 , n27709 );
nand ( n27781 , n27777 , n27780 );
nand ( n27782 , n27781 , n9907 );
not ( n27783 , n27782 );
not ( n27784 , n27783 );
or ( n27785 , n27772 , n27784 );
nor ( n27786 , n27429 , n26021 );
not ( n27787 , n27786 );
not ( n27788 , n19075 );
or ( n27789 , n27787 , n27788 );
and ( n27790 , n27422 , n27749 );
nor ( n27791 , n27790 , n27432 );
nand ( n27792 , n27789 , n27791 );
or ( n27793 , n27452 , n27418 );
nand ( n27794 , n27418 , n27452 );
nand ( n27795 , n27793 , n27794 );
not ( n27796 , n27795 );
and ( n27797 , n27792 , n27796 );
not ( n27798 , n27792 );
and ( n27799 , n27798 , n27795 );
nor ( n27800 , n27797 , n27799 );
not ( n27801 , n454 );
nor ( n27802 , n27801 , n6725 );
nand ( n27803 , n27800 , n27802 );
nand ( n27804 , n27785 , n27803 );
nand ( n27805 , n26136 , n26133 );
and ( n27806 , n27805 , n26151 );
nor ( n27807 , n27806 , n17873 );
xor ( n27808 , n27804 , n27807 );
and ( n27809 , n27251 , n470 );
xor ( n27810 , n27808 , n27809 );
xor ( n27811 , n27804 , n27807 );
and ( n27812 , n27811 , n27809 );
and ( n27813 , n27804 , n27807 );
or ( n27814 , n27812 , n27813 );
and ( n27815 , n27764 , n471 );
xor ( n27816 , n27815 , n27744 );
xor ( n27817 , n27816 , n27810 );
xor ( n27818 , n27815 , n27744 );
and ( n27819 , n27818 , n27810 );
and ( n27820 , n27815 , n27744 );
or ( n27821 , n27819 , n27820 );
and ( n27822 , n16206 , n17637 , n27683 );
not ( n27823 , n27822 );
not ( n27824 , n17578 );
or ( n27825 , n27823 , n27824 );
nand ( n27826 , n27825 , n27706 );
not ( n27827 , n27694 );
nand ( n27828 , n27827 , n27684 );
not ( n27829 , n27828 );
and ( n27830 , n27826 , n27829 );
not ( n27831 , n27826 );
and ( n27832 , n27831 , n27828 );
nor ( n27833 , n27830 , n27832 );
not ( n27834 , n454 );
nand ( n27835 , n27833 , n27834 );
not ( n27836 , n27835 );
and ( n27837 , n27836 , n472 );
and ( n27838 , n27251 , n469 );
xor ( n27839 , n27837 , n27838 );
and ( n27840 , n27756 , n27763 );
not ( n27841 , n470 );
nor ( n27842 , n27840 , n27841 );
xor ( n27843 , n27839 , n27842 );
xor ( n27844 , n27837 , n27838 );
and ( n27845 , n27844 , n27842 );
and ( n27846 , n27837 , n27838 );
or ( n27847 , n27845 , n27846 );
not ( n27848 , n454 );
not ( n27849 , n27848 );
nand ( n27850 , n27849 , n27795 );
nand ( n27851 , n27792 , n27850 );
not ( n27852 , n27851 );
not ( n27853 , n27792 );
or ( n27854 , n27795 , n27848 );
nand ( n27855 , n27853 , n27854 );
not ( n27856 , n27855 );
or ( n27857 , n27852 , n27856 );
nand ( n27858 , n27857 , n27782 );
and ( n27859 , n27858 , n471 );
xor ( n27860 , n27859 , n27814 );
xor ( n27861 , n27860 , n27843 );
xor ( n27862 , n27859 , n27814 );
and ( n27863 , n27862 , n27843 );
and ( n27864 , n27859 , n27814 );
or ( n27865 , n27863 , n27864 );
and ( n27866 , n27836 , n471 );
not ( n27867 , n27757 );
nor ( n27868 , n27867 , n27685 );
not ( n27869 , n27868 );
not ( n27870 , n17578 );
or ( n27871 , n27869 , n27870 );
nand ( n27872 , n27871 , n27697 );
and ( n27873 , n27651 , n27659 );
not ( n27874 , n27873 );
or ( n27875 , n27651 , n27659 );
nand ( n27876 , n27874 , n27875 );
not ( n27877 , n27876 );
and ( n27878 , n27872 , n27877 );
not ( n27879 , n27872 );
and ( n27880 , n27879 , n27876 );
nor ( n27881 , n27878 , n27880 );
and ( n27882 , n27834 , n472 , n27881 );
xor ( n27883 , n27866 , n27882 );
and ( n27884 , n27858 , n470 );
xor ( n27885 , n27883 , n27884 );
xor ( n27886 , n27866 , n27882 );
and ( n27887 , n27886 , n27884 );
and ( n27888 , n27866 , n27882 );
or ( n27889 , n27887 , n27888 );
and ( n27890 , n27764 , n469 );
xor ( n27891 , n27890 , n27885 );
xor ( n27892 , n27891 , n27847 );
xor ( n27893 , n27890 , n27885 );
and ( n27894 , n27893 , n27847 );
and ( n27895 , n27890 , n27885 );
or ( n27896 , n27894 , n27895 );
xor ( n27897 , n27663 , n27726 );
and ( n27898 , n27897 , n27834 );
not ( n27899 , n27898 );
not ( n27900 , n27875 );
nor ( n27901 , n27867 , n27685 , n27900 );
not ( n27902 , n27901 );
not ( n27903 , n17578 );
or ( n27904 , n27902 , n27903 );
and ( n27905 , n27875 , n27696 );
nor ( n27906 , n27905 , n27873 );
nand ( n27907 , n27904 , n27906 );
not ( n27908 , n27907 );
not ( n27909 , n27908 );
or ( n27910 , n27899 , n27909 );
not ( n27911 , n27834 );
nor ( n27912 , n27911 , n27897 );
nand ( n27913 , n27907 , n27912 );
nand ( n27914 , n27910 , n27913 );
and ( n27915 , n27914 , n472 );
and ( n27916 , n27836 , n470 );
xor ( n27917 , n27915 , n27916 );
nand ( n27918 , n27881 , n27834 );
not ( n27919 , n27918 );
and ( n27920 , n27919 , n471 );
xor ( n27921 , n27917 , n27920 );
xor ( n27922 , n27915 , n27916 );
and ( n27923 , n27922 , n27920 );
and ( n27924 , n27915 , n27916 );
or ( n27925 , n27923 , n27924 );
and ( n27926 , n27858 , n469 );
xor ( n27927 , n27926 , n27921 );
xor ( n27928 , n27927 , n27889 );
xor ( n27929 , n27926 , n27921 );
and ( n27930 , n27929 , n27889 );
and ( n27931 , n27926 , n27921 );
or ( n27932 , n27930 , n27931 );
and ( n27933 , n27919 , n470 );
nand ( n27934 , n27914 , n471 );
not ( n27935 , n27934 );
and ( n27936 , n27834 , n469 );
nand ( n27937 , n27833 , n27936 );
not ( n27938 , n27937 );
not ( n27939 , n27938 );
or ( n27940 , n27935 , n27939 );
or ( n27941 , n27934 , n27938 );
nand ( n27942 , n27940 , n27941 );
xor ( n27943 , n27933 , n27942 );
xor ( n27944 , n27943 , n27925 );
xor ( n27945 , n27933 , n27942 );
and ( n27946 , n27945 , n27925 );
and ( n27947 , n27933 , n27942 );
or ( n27948 , n27946 , n27947 );
and ( n27949 , n27914 , n470 );
and ( n27950 , n27919 , n469 );
xor ( n27951 , n27949 , n27950 );
nor ( n27952 , n27934 , n27937 );
xor ( n27953 , n27951 , n27952 );
xor ( n27954 , n27949 , n27950 );
and ( n27955 , n27954 , n27952 );
and ( n27956 , n27949 , n27950 );
or ( n27957 , n27955 , n27956 );
and ( n27958 , n26527 , n26542 );
not ( n27959 , n27958 );
not ( n27960 , n26535 );
or ( n27961 , n27959 , n27960 );
not ( n27962 , n26542 );
not ( n27963 , n17928 );
or ( n27964 , n27962 , n27963 );
nand ( n27965 , n27964 , n26541 );
not ( n27966 , n27965 );
nand ( n27967 , n27961 , n27966 );
xor ( n27968 , n18736 , n18738 );
xor ( n27969 , n27968 , n18898 );
xor ( n27970 , n18753 , n18755 );
xor ( n27971 , n27970 , n18895 );
nand ( n27972 , n27861 , n27821 );
not ( n27973 , n27972 );
not ( n27974 , n27928 );
not ( n27975 , n27974 );
not ( n27976 , n27896 );
not ( n27977 , n27976 );
or ( n27978 , n27975 , n27977 );
not ( n27979 , n27892 );
not ( n27980 , n27979 );
or ( n27981 , n27980 , n27865 );
nand ( n27982 , n27978 , n27981 );
nor ( n27983 , n27932 , n27944 );
nor ( n27984 , n27982 , n27983 );
not ( n27985 , n27948 );
not ( n27986 , n27953 );
nand ( n27987 , n27985 , n27986 );
nand ( n27988 , n27984 , n27987 );
not ( n27989 , n27988 );
nand ( n27990 , n27973 , n27989 );
not ( n27991 , n27865 );
nor ( n27992 , n27979 , n27991 );
not ( n27993 , n27992 );
nand ( n27994 , n27976 , n27974 );
not ( n27995 , n27994 );
or ( n27996 , n27993 , n27995 );
nand ( n27997 , n27928 , n27896 );
nand ( n27998 , n27996 , n27997 );
not ( n27999 , n27998 );
buf ( n28000 , n27999 );
nand ( n28001 , n18697 , n18905 );
nand ( n28002 , n18712 , n18907 );
nand ( n28003 , n27979 , n27991 );
not ( n28004 , n27992 );
nand ( n28005 , n28003 , n28004 );
not ( n28006 , n27861 );
not ( n28007 , n27821 );
nand ( n28008 , n28006 , n28007 );
buf ( n28009 , n28008 );
nand ( n28010 , n28009 , n27972 );
not ( n28011 , n27817 );
not ( n28012 , n27771 );
nand ( n28013 , n28011 , n28012 );
nand ( n28014 , n27817 , n27771 );
nand ( n28015 , n28013 , n28014 );
not ( n28016 , n27982 );
not ( n28017 , n26174 );
xor ( n28018 , n18859 , n18861 );
xor ( n28019 , n28018 , n18874 );
nand ( n28020 , n27932 , n27944 );
and ( n28021 , n27914 , n469 );
nor ( n28022 , n27957 , n28021 );
not ( n28023 , n28022 );
nand ( n28024 , n27957 , n28021 );
nand ( n28025 , n28023 , n28024 );
and ( n28026 , n18806 , n472 );
and ( n28027 , n14012 , n471 );
nor ( n28028 , n28026 , n28027 );
not ( n28029 , n27254 );
not ( n28030 , n27258 );
and ( n28031 , n28029 , n28030 );
nor ( n28032 , n27767 , n27734 );
nor ( n28033 , n28031 , n28032 );
nand ( n28034 , n28033 , n27278 );
not ( n28035 , n27817 );
nand ( n28036 , n28035 , n28012 );
nand ( n28037 , n28006 , n28007 );
nand ( n28038 , n28036 , n25988 , n28037 );
nor ( n28039 , n28034 , n28038 );
nand ( n28040 , n27269 , n28039 );
not ( n28041 , n28040 );
nand ( n28042 , n28041 , n27989 );
and ( n28043 , n18802 , n18890 );
xor ( n28044 , n18887 , n28043 );
xnor ( n28045 , n18901 , n28001 );
xnor ( n28046 , n26510 , n28002 );
not ( n28047 , n27983 );
nand ( n28048 , n28047 , n28020 );
xor ( n28049 , n27534 , n27481 );
xor ( n28050 , n27503 , n27483 );
xor ( n28051 , n27524 , n27478 );
nand ( n28052 , n27948 , n27953 );
xnor ( n28053 , n27531 , n27463 );
not ( n28054 , n19221 );
nand ( n28055 , n28054 , n27994 , n27997 );
not ( n28056 , n28003 );
not ( n28057 , n28039 );
not ( n28058 , n27269 );
or ( n28059 , n28057 , n28058 );
nand ( n28060 , n28013 , n28033 );
not ( n28061 , n27861 );
nand ( n28062 , n28007 , n28061 );
not ( n28063 , n28062 );
nor ( n28064 , n28060 , n28063 );
nand ( n28065 , n27282 , n28064 );
nand ( n28066 , n28059 , n28065 );
not ( n28067 , n28066 );
not ( n28068 , n28013 );
nor ( n28069 , n27767 , n27734 );
or ( n28070 , n27260 , n28069 );
nand ( n28071 , n27767 , n27734 );
nand ( n28072 , n28070 , n28071 );
not ( n28073 , n28072 );
or ( n28074 , n28068 , n28073 );
nand ( n28075 , n28074 , n28014 );
nand ( n28076 , n28075 , n28009 );
nand ( n28077 , n27972 , n28076 );
not ( n28078 , n28077 );
nand ( n28079 , n28067 , n28078 );
not ( n28080 , n28079 );
or ( n28081 , n28056 , n28080 );
buf ( n28082 , n28004 );
nand ( n28083 , n28081 , n28082 );
or ( n28084 , n28055 , n28083 );
and ( n28085 , n27994 , n27997 );
nor ( n28086 , n28085 , n19221 );
nand ( n28087 , n28083 , n28086 );
xor ( n28088 , n27533 , n27475 );
or ( n28089 , n28088 , n19220 );
nand ( n28090 , n28084 , n28087 , n28089 );
or ( n28091 , n28015 , n19221 );
not ( n28092 , n27254 );
not ( n28093 , n27258 );
and ( n28094 , n28092 , n28093 );
buf ( n28095 , n28032 );
nor ( n28096 , n28094 , n28095 );
not ( n28097 , n28096 );
not ( n28098 , n27284 );
or ( n28099 , n28097 , n28098 );
buf ( n28100 , n28072 );
not ( n28101 , n28100 );
nand ( n28102 , n28099 , n28101 );
not ( n28103 , n28015 );
nor ( n28104 , n28103 , n19221 );
nand ( n28105 , n28102 , n28104 );
or ( n28106 , n28051 , n19220 );
not ( n28107 , n27259 );
not ( n28108 , n27284 );
or ( n28109 , n28107 , n28108 );
nand ( n28110 , n28109 , n27261 );
not ( n28111 , n28069 );
buf ( n28112 , n28071 );
nand ( n28113 , n28111 , n28112 );
or ( n28114 , n28113 , n19221 );
or ( n28115 , n28110 , n28114 );
not ( n28116 , n28113 );
nor ( n28117 , n28116 , n19221 );
nand ( n28118 , n28110 , n28117 );
not ( n28119 , n19220 );
nand ( n28120 , n28119 , n27551 );
nand ( n28121 , n28115 , n28118 , n28120 );
not ( n28122 , n28066 );
not ( n28123 , n28122 );
not ( n28124 , n28078 );
or ( n28125 , n28123 , n28124 );
not ( n28126 , n28005 );
nor ( n28127 , n28126 , n26561 );
nand ( n28128 , n28125 , n28127 );
nor ( n28129 , n28005 , n26561 );
nand ( n28130 , n28122 , n28078 , n28129 );
nand ( n28131 , n28053 , n26561 );
nand ( n28132 , n28128 , n28130 , n28131 );
or ( n28133 , n28048 , n19221 );
not ( n28134 , n28016 );
not ( n28135 , n28079 );
or ( n28136 , n28134 , n28135 );
nand ( n28137 , n28136 , n28000 );
or ( n28138 , n28133 , n28137 );
not ( n28139 , n28048 );
nor ( n28140 , n28139 , n19221 );
nand ( n28141 , n28137 , n28140 );
xor ( n28142 , n27535 , n27471 );
or ( n28143 , n28142 , n19220 );
nand ( n28144 , n28138 , n28141 , n28143 );
or ( n28145 , n28025 , n19221 );
or ( n28146 , n28010 , n19221 );
nand ( n28147 , n27267 , n27269 );
not ( n28148 , n28060 );
not ( n28149 , n28148 );
or ( n28150 , n28147 , n28149 );
not ( n28151 , n27279 );
nor ( n28152 , n28151 , n27280 );
or ( n28153 , n28149 , n28152 );
not ( n28154 , n28149 );
nand ( n28155 , n28154 , n28017 );
not ( n28156 , n28013 );
not ( n28157 , n28072 );
or ( n28158 , n28156 , n28157 );
nand ( n28159 , n28158 , n28014 );
not ( n28160 , n28159 );
nand ( n28161 , n28150 , n28153 , n28155 , n28160 );
or ( n28162 , n28146 , n28161 );
not ( n28163 , n28010 );
nor ( n28164 , n28163 , n19221 );
nand ( n28165 , n28161 , n28164 );
or ( n28166 , n28049 , n19220 );
nand ( n28167 , n28162 , n28165 , n28166 );
not ( n28168 , n27987 );
not ( n28169 , n28168 );
nand ( n28170 , n28169 , n28052 );
not ( n28171 , n28170 );
nand ( n28172 , n28171 , n19220 );
nor ( n28173 , n27944 , n27932 );
nand ( n28174 , n18181 , n18185 );
or ( n28175 , n28174 , n19221 );
or ( n28176 , n27967 , n28175 );
not ( n28177 , n28174 );
nor ( n28178 , n28177 , n19221 );
nand ( n28179 , n27967 , n28178 );
or ( n28180 , n28050 , n19220 );
nand ( n28181 , n28176 , n28179 , n28180 );
not ( n28182 , n27983 );
not ( n28183 , n27972 );
and ( n28184 , n27976 , n27974 );
nor ( n28185 , n28184 , n28173 );
nand ( n28186 , n28183 , n28185 , n28003 );
not ( n28187 , n27948 );
not ( n28188 , n25899 );
and ( n28189 , n19207 , n19203 );
not ( n28190 , n27984 );
not ( n28191 , n28066 );
or ( n28192 , n28190 , n28191 );
and ( n28193 , n28185 , n28003 , n28062 );
not ( n28194 , n28193 );
not ( n28195 , n28159 );
or ( n28196 , n28194 , n28195 );
nand ( n28197 , n28196 , n28186 );
not ( n28198 , n28182 );
not ( n28199 , n27998 );
or ( n28200 , n28198 , n28199 );
nand ( n28201 , n28200 , n28020 );
nor ( n28202 , n28197 , n28201 );
nand ( n28203 , n28192 , n28202 );
not ( n28204 , n19220 );
nor ( n28205 , n28168 , n28022 , n28204 );
not ( n28206 , n18404 );
not ( n28207 , n25899 );
or ( n28208 , n28206 , n28207 );
nand ( n28209 , n28208 , n25900 );
or ( n28210 , n28091 , n28102 );
nand ( n28211 , n28210 , n28105 , n28106 );
or ( n28212 , n18873 , n18871 );
not ( n28213 , n18871 );
and ( n28214 , n18867 , n28213 );
not ( n28215 , n18866 );
nor ( n28216 , n28213 , n28215 , n18864 );
nor ( n28217 , n28214 , n28216 );
nand ( n28218 , n28215 , n18871 , n18864 );
nand ( n28219 , n28212 , n28217 , n28218 );
not ( n28220 , n18864 );
nand ( n28221 , n18273 , n25927 );
and ( n28222 , n28221 , n25928 );
not ( n28223 , n18360 );
nor ( n28224 , n28223 , n18366 );
or ( n28225 , n28222 , n28224 , n26561 );
and ( n28226 , n28224 , n25928 , n19220 );
and ( n28227 , n28221 , n28226 );
and ( n28228 , n27493 , n19221 );
nor ( n28229 , n28227 , n28228 );
nand ( n28230 , n28225 , n28229 );
not ( n28231 , n28065 );
not ( n28232 , n28076 );
or ( n28233 , n28231 , n28232 );
nand ( n28234 , n28233 , n27989 );
not ( n28235 , n28187 );
not ( n28236 , n27986 );
and ( n28237 , n28235 , n28236 );
and ( n28238 , n28201 , n27987 );
nor ( n28239 , n28237 , n28238 );
nand ( n28240 , n28234 , n27990 , n28042 , n28239 );
not ( n28241 , n28025 );
nor ( n28242 , n28241 , n19221 );
nand ( n28243 , n28240 , n28242 );
or ( n28244 , n28172 , n28203 );
and ( n28245 , n19220 , n28170 );
nand ( n28246 , n28203 , n28245 );
nand ( n28247 , n28244 , n28246 , n27192 );
buf ( n28248 , n18413 );
nand ( n28249 , n28248 , n18982 );
or ( n28250 , n28249 , n19221 );
or ( n28251 , n28209 , n28250 );
not ( n28252 , n28209 );
nand ( n28253 , n28249 , n19220 );
or ( n28254 , n28252 , n28253 );
xor ( n28255 , n27513 , n25780 );
or ( n28256 , n28255 , n19220 );
nand ( n28257 , n28251 , n28254 , n28256 );
buf ( n28258 , n18414 );
nor ( n28259 , n28258 , n19221 );
nand ( n28260 , n18387 , n18987 );
nand ( n28261 , n28259 , n28260 );
or ( n28262 , n28188 , n28261 );
buf ( n28263 , n18983 );
buf ( n28264 , n28263 );
not ( n28265 , n28264 );
not ( n28266 , n28265 );
nor ( n28267 , n28266 , n28260 , n19221 );
nand ( n28268 , n28188 , n28267 );
nor ( n28269 , n28265 , n19221 );
and ( n28270 , n28269 , n28260 );
not ( n28271 , n19221 );
nand ( n28272 , n28265 , n28258 , n28271 );
or ( n28273 , n28272 , n28260 );
xor ( n28274 , n27505 , n27488 );
or ( n28275 , n28274 , n19220 );
nand ( n28276 , n28273 , n28275 );
nor ( n28277 , n28270 , n28276 );
nand ( n28278 , n28262 , n28268 , n28277 );
and ( n28279 , n25628 , n25630 );
nor ( n28280 , n28279 , n25631 );
not ( n28281 , n28280 );
not ( n28282 , n19220 );
and ( n28283 , n28281 , n28282 );
and ( n28284 , n28028 , n19220 );
nor ( n28285 , n28283 , n28284 );
not ( n28286 , n19220 );
nand ( n28287 , n27552 , n28286 );
nor ( n28288 , n28189 , n19221 );
and ( n28289 , n19220 , n18863 );
not ( n28290 , n19220 );
and ( n28291 , n28290 , n25629 );
nor ( n28292 , n28289 , n28291 );
and ( n28293 , n28220 , n19220 );
not ( n28294 , n28285 );
nor ( n28295 , n28293 , n28294 );
and ( n28296 , n27441 , n454 );
and ( n28297 , n27718 , n17777 );
nor ( n28298 , n28296 , n28297 );
and ( n28299 , n27448 , n454 );
and ( n28300 , n9781 , n17777 );
nor ( n28301 , n28299 , n28300 );
and ( n28302 , n27439 , n454 );
and ( n28303 , n27716 , n17777 );
nor ( n28304 , n28302 , n28303 );
and ( n28305 , n454 , n27443 );
and ( n28306 , n27720 , n17777 );
nor ( n28307 , n28305 , n28306 );
not ( n28308 , n28307 );
not ( n28309 , n28205 );
not ( n28310 , n28203 );
or ( n28311 , n28309 , n28310 );
and ( n28312 , n27470 , n19221 );
or ( n28313 , n28022 , n28052 );
nand ( n28314 , n28313 , n28024 );
and ( n28315 , n28314 , n19220 );
nor ( n28316 , n28312 , n28315 );
nand ( n28317 , n28311 , n28316 );
not ( n28318 , n19220 );
not ( n28319 , n27971 );
or ( n28320 , n28318 , n28319 );
nand ( n28321 , n27521 , n26561 );
nand ( n28322 , n28320 , n28321 );
not ( n28323 , n19220 );
not ( n28324 , n28046 );
or ( n28325 , n28323 , n28324 );
nand ( n28326 , n27501 , n26561 );
nand ( n28327 , n28325 , n28326 );
not ( n28328 , n19220 );
not ( n28329 , n28044 );
or ( n28330 , n28328 , n28329 );
nand ( n28331 , n27530 , n26561 );
nand ( n28332 , n28330 , n28331 );
not ( n28333 , n19220 );
not ( n28334 , n28045 );
or ( n28335 , n28333 , n28334 );
nand ( n28336 , n27512 , n26561 );
nand ( n28337 , n28335 , n28336 );
not ( n28338 , n19220 );
not ( n28339 , n27969 );
or ( n28340 , n28338 , n28339 );
nand ( n28341 , n27515 , n26561 );
nand ( n28342 , n28340 , n28341 );
not ( n28343 , n19220 );
not ( n28344 , n28219 );
or ( n28345 , n28343 , n28344 );
nand ( n28346 , n27550 , n26561 );
nand ( n28347 , n28345 , n28346 );
not ( n28348 , n19220 );
xor ( n28349 , n18854 , n18856 );
xor ( n28350 , n28349 , n18877 );
not ( n28351 , n28350 );
or ( n28352 , n28348 , n28351 );
nand ( n28353 , n27546 , n26561 );
nand ( n28354 , n28352 , n28353 );
not ( n28355 , n28301 );
not ( n28356 , n28298 );
not ( n28357 , n28304 );
not ( n28358 , n28288 );
not ( n28359 , n18991 );
or ( n28360 , n28358 , n28359 );
and ( n28361 , n18992 , n28189 , n19220 );
not ( n28362 , n25865 );
and ( n28363 , n28362 , n27506 );
not ( n28364 , n27506 );
and ( n28365 , n25865 , n28364 );
nor ( n28366 , n28363 , n28365 , n19220 );
nor ( n28367 , n28361 , n28366 );
nand ( n28368 , n28360 , n28367 );
not ( n28369 , n19220 );
not ( n28370 , n28019 );
or ( n28371 , n28369 , n28370 );
nand ( n28372 , n27548 , n26561 );
nand ( n28373 , n28371 , n28372 );
or ( n28375 , n28240 , n28145 );
nand ( n28376 , n28375 , n28243 , n28287 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
