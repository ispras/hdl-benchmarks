// IWLS benchmark module "x4" printed on Wed May 29 17:30:39 2002
module x4(a, b, g, h, i, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5);
input
  a,
  b,
  g,
  h,
  i,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  a1,
  a2,
  b0,
  b1,
  b2,
  c0,
  c1,
  c2,
  d0,
  d1,
  d2,
  e0,
  e1,
  e2,
  f0,
  f1,
  f2,
  g0,
  g1,
  g2,
  h0,
  h1,
  h2,
  i0,
  i1,
  i2,
  j1,
  j2,
  k0,
  k1,
  k2,
  l0,
  l1,
  l2,
  m0,
  m1,
  m2,
  n0,
  n1,
  n2,
  o0,
  o1,
  o2,
  p0,
  p1,
  p2,
  q0,
  q1,
  q2,
  r0,
  r1,
  r2,
  s0,
  s1,
  s2,
  t0,
  t1,
  t2,
  u0,
  u1,
  u2,
  v0,
  v1,
  v2,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1,
  z0,
  z1;
output
  a3,
  a4,
  a5,
  b3,
  b4,
  b5,
  c3,
  c4,
  c5,
  d3,
  d4,
  d5,
  e3,
  e4,
  e5,
  f3,
  f4,
  f5,
  g3,
  g4,
  g5,
  h3,
  h4,
  h5,
  i3,
  i4,
  i5,
  j3,
  j4,
  j5,
  k3,
  k4,
  k5,
  l3,
  l4,
  l5,
  m3,
  m4,
  m5,
  n3,
  n4,
  n5,
  o3,
  o4,
  o5,
  p3,
  p4,
  q3,
  q4,
  r3,
  r4,
  s3,
  s4,
  t3,
  t4,
  u3,
  u4,
  v3,
  v4,
  w2,
  w3,
  w4,
  x2,
  x3,
  x4,
  y2,
  y3,
  y4,
  z2,
  z3,
  z4;
wire
  \[59] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  l10,
  l11,
  \[60] ,
  \[61] ,
  \[62] ,
  \[0] ,
  \[63] ,
  \[1] ,
  \[64] ,
  \[20] ,
  \[2] ,
  \[65] ,
  \[21] ,
  \[3] ,
  \[66] ,
  \[22] ,
  \[4] ,
  \[67] ,
  \[23] ,
  \[5] ,
  \[68] ,
  \[24] ,
  \[6] ,
  \[69] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  \[28] ,
  \[29] ,
  \[70] ,
  \[72] ,
  \[73] ,
  z13,
  \[74] ,
  i11,
  \[30] ,
  \[75] ,
  \[31] ,
  \[76] ,
  \[32] ,
  \[77] ,
  \[33] ,
  v10,
  \[78] ,
  \[34] ,
  e11,
  \[79] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  n10,
  \[80] ,
  \[81] ,
  \[83] ,
  \[84] ,
  \[40] ,
  \[85] ,
  \[41] ,
  \[42] ,
  \[87] ,
  \[43] ,
  \[44] ,
  \[89] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  k11,
  \[50] ,
  \[51] ,
  \[52] ,
  \[97] ,
  \[53] ,
  \[98] ,
  \[54] ,
  \[10] ,
  \[55] ,
  \[11] ,
  \[56] ,
  \[12] ,
  \[57] ,
  \[13] ,
  \[58] ,
  \[14] ;
assign
  \[59]  = (\[89]  & (~k2 & ~c1)) | (\[98]  & ~\[89] ),
  \[15]  = \[81]  & s0,
  \[16]  = \[81]  & t0,
  \[17]  = b & ~i0,
  \[18]  = a & ~i0,
  \[19]  = ~i0 & v0,
  l10 = \[92]  & (~p2 & o2),
  l11 = ~\[72]  | k11,
  \[60]  = (z13 & (l2 & (~k2 & ~c1))) | ((\[98]  & (~\[59]  & ~l2)) | (z13 & (\[59]  & l2))),
  \[61]  = (\[98]  & (~\[59]  & (~m2 & l2))) | ((m2 & (~l2 & ~c1)) | (\[60]  & m2)),
  \[62]  = (~\[27]  & (n2 & ~c1)) | (\[27]  & ~n2),
  \[0]  = ~f1,
  \[63]  = (~\[27]  & (o2 & ~c1)) | ((\[27]  & (~o2 & n2)) | (\[93]  & ~n2)),
  \[1]  = ~g1,
  \[64]  = (\[93]  & ~\[78] ) | (\[87]  & p2),
  \[20]  = ~i0 & w0,
  \[2]  = ~h1,
  \[65]  = (\[93]  & (~\[63]  & (~q2 & p2))) | ((\[27]  & (q2 & ~p2)) | (\[87]  & q2)),
  \[21]  = ~i0 & x0,
  \[3]  = ~i1,
  \[66]  = (\[93]  & (~\[90]  & (~\[63]  & ~r2))) | ((\[90]  & (r2 & ~c1)) | (\[64]  & r2)),
  \[22]  = ~i0 & y0,
  \[4]  = ~j1,
  \[67]  = (\[72]  & (b1 & ~i0)) | (\[73]  & n1),
  \[23]  = ~i0 & z0,
  \[5]  = ~k1,
  \[68]  = (~\[91]  & (~t2 & ~c1)) | (\[91]  & (t2 & ~c1)),
  \[24]  = ~i0 & a1,
  \[6]  = (~\[83]  & (~t2 & (~i0 & ~h0))) | ((~\[83]  & (t2 & (~i0 & h0))) | (\[83]  & (s2 & ~i0))),
  \[69]  = (z13 & (u2 & ~i0)) | (\[17]  & ~u0),
  \[25]  = (v2 & f0) | (\[97]  | ~\[83] ),
  \[7]  = (~k11 & (v2 & (~c1 & g0))) | ((v2 & (~c1 & f0)) | (~c1 & k0)),
  \[26]  = ~e11 & (v10 & (v2 & (~m1 & ~g0))),
  \[8]  = (\[92]  & (~\[79]  & (~l10 & ~c1))) | (~c1 & l0),
  \[27]  = (~z13 & ~c1) | ((e1 & ~c1) | (d1 & ~c1)),
  \[9]  = (~v10 & m0) | \[97] ,
  \[28]  = (\[85]  & f1) | (\[84]  & o0),
  \[29]  = (\[85]  & g1) | (\[84]  & p0),
  \[70]  = (~v10 & (v2 & ~f0)) | (~\[83]  & ~v10),
  \[72]  = ~e1 | m0,
  \[73]  = ~\[72]  & ~i0,
  z13 = k2 | (~l2 | ~m2),
  \[74]  = ~e11 & g0,
  i11 = i0 | (~m1 | ~v2),
  \[30]  = (\[85]  & h1) | (\[84]  & q0),
  \[75]  = ~l11 & ~i0,
  \[31]  = (\[85]  & i1) | (\[84]  & r0),
  \[76]  = \[74]  & ~i11,
  \[32]  = (\[85]  & j1) | (\[84]  & s0),
  \[77]  = \[73]  & ~k11,
  \[33]  = (\[85]  & k1) | (\[84]  & t0),
  v10 = (g0 & v2) | i0,
  \[78]  = p2 | ~n2,
  \[34]  = (\[92]  & (~\[79]  & (~l10 & ~c1))) | (l1 & ~c1),
  e11 = ~g & (~h & (~i & h0)),
  a3 = \[4] ,
  a4 = \[30] ,
  a5 = \[56] ,
  \[79]  = \[78]  | ~e1,
  \[35]  = (~z13 & (~v10 & (~h & ~g))) | (~v10 & m1),
  b3 = \[5] ,
  b4 = \[31] ,
  b5 = \[57] ,
  \[36]  = (k11 & (~i11 & i)) | ((\[77]  & ~o1) | (\[75]  & n1)),
  c3 = \[6] ,
  c4 = \[32] ,
  c5 = \[58] ,
  \[37]  = (~i11 & (~e11 & v10)) | ((~l11 & o1) | ((l11 & ~p1) | i0)),
  d3 = \[7] ,
  d4 = \[33] ,
  d5 = \[59] ,
  \[38]  = (\[77]  & q1) | ((\[76]  & k) | (\[75]  & p1)),
  e3 = \[8] ,
  e4 = \[34] ,
  e5 = \[60] ,
  \[39]  = (\[77]  & r1) | ((\[76]  & l) | (\[75]  & q1)),
  f3 = \[9] ,
  f4 = \[35] ,
  f5 = \[61] ,
  g3 = \[10] ,
  g4 = \[36] ,
  g5 = \[62] ,
  h3 = \[11] ,
  h4 = \[37] ,
  h5 = \[63] ,
  n10 = ~l10 | (n2 | ~e1),
  \[80]  = \[79]  | o2,
  i3 = \[12] ,
  i4 = \[38] ,
  i5 = \[64] ,
  \[81]  = ~c1 & ~i0,
  j3 = \[13] ,
  j4 = \[39] ,
  j5 = \[65] ,
  k3 = \[14] ,
  k4 = \[40] ,
  k5 = \[66] ,
  \[83]  = (~q2 & ~i) | (\[80]  | ~r2),
  l3 = \[15] ,
  l4 = \[41] ,
  l5 = \[67] ,
  \[84]  = ~n10 & ~c1,
  \[40]  = (\[77]  & s1) | ((\[76]  & m) | (\[75]  & r1)),
  m3 = \[16] ,
  m4 = \[42] ,
  m5 = \[68] ,
  \[85]  = n10 & ~c1,
  \[41]  = (\[77]  & t1) | ((\[76]  & n) | (\[75]  & s1)),
  n3 = \[17] ,
  n4 = \[43] ,
  n5 = \[69] ,
  \[42]  = (\[77]  & u1) | ((\[76]  & o) | (\[75]  & t1)),
  o3 = \[18] ,
  o4 = \[44] ,
  o5 = \[70] ,
  \[87]  = (~o2 & ~c1) | \[63] ,
  \[43]  = (\[77]  & v1) | ((\[76]  & p) | (\[75]  & u1)),
  p3 = \[19] ,
  p4 = \[45] ,
  \[44]  = (\[77]  & w1) | ((\[76]  & q) | (\[75]  & v1)),
  q3 = \[20] ,
  q4 = \[46] ,
  \[89]  = (~u0 & b) | u2,
  \[45]  = (\[77]  & x1) | ((\[76]  & r) | (\[75]  & w1)),
  r3 = \[21] ,
  r4 = \[47] ,
  \[46]  = (\[77]  & y1) | ((\[76]  & s) | (\[75]  & x1)),
  s3 = \[22] ,
  s4 = \[48] ,
  \[47]  = (\[77]  & z1) | ((\[76]  & t) | (\[75]  & y1)),
  t3 = \[23] ,
  t4 = \[49] ,
  \[48]  = (\[77]  & a2) | ((\[76]  & u) | (\[75]  & z1)),
  u3 = \[24] ,
  u4 = \[50] ,
  \[49]  = (\[77]  & b2) | ((\[76]  & v) | (\[75]  & a2)),
  v3 = \[25] ,
  v4 = \[51] ,
  w2 = \[0] ,
  w3 = \[26] ,
  w4 = \[52] ,
  x2 = \[1] ,
  x3 = \[27] ,
  x4 = \[53] ,
  \[90]  = ~q2 | ~p2,
  y2 = \[2] ,
  y3 = \[28] ,
  y4 = \[54] ,
  \[91]  = ~s2 | ~l1,
  z2 = \[3] ,
  z3 = \[29] ,
  z4 = \[55] ,
  \[92]  = ~r2 & ~q2,
  \[93]  = \[27]  & o2,
  k11 = \[74]  & (v2 & m1),
  \[50]  = (\[77]  & c2) | ((\[76]  & w) | (\[75]  & b2)),
  \[51]  = (\[77]  & d2) | ((\[76]  & \x ) | (\[75]  & c2)),
  \[52]  = (\[77]  & e2) | ((\[76]  & y) | (\[75]  & d2)),
  \[97]  = (e11 & v10) | ((v10 & ~m1) | i0),
  \[53]  = (\[77]  & f2) | ((\[76]  & z) | (\[75]  & e2)),
  \[98]  = k2 & ~c1,
  \[54]  = (\[77]  & g2) | ((\[76]  & a0) | (\[75]  & f2)),
  \[10]  = (\[92]  & (\[81]  & ~\[80] )) | (\[81]  & n0),
  \[55]  = (\[77]  & h2) | ((\[76]  & b0) | (\[75]  & g2)),
  \[11]  = \[81]  & o0,
  \[56]  = (\[77]  & i2) | ((\[76]  & c0) | (\[75]  & h2)),
  \[12]  = \[81]  & p0,
  \[57]  = (\[77]  & j2) | ((\[76]  & d0) | (\[75]  & i2)),
  \[13]  = \[81]  & q0,
  \[58]  = (\[76]  & e0) | (\[75]  & j2),
  \[14]  = \[81]  & r0;
endmodule

