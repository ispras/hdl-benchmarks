//NOTE: no-implementation module stub

module daddr (
    input wire SYSCLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire CLMI_RHOLD,
    input wire REGA_E_R,
    input wire REGBI_E_R,
    input wire REGBR_E_R,
    input wire WIDTH_E_P,
    input wire DBYEN_E,
    output wire DADALERR_E,
    output wire DADDR_E,
    output wire DWORD_E,
    output wire ADATAREG_M_R
);

endmodule
