// IWLS benchmark module "cordic" printed on Wed May 29 16:31:29 2002
module cordic(a6, a4, a3, a2, a5, v, x0, x1, x2, x3, y0, y1, y2, y3, z0, z1, z2, ex0, ex1, ex2, ey0, ey1, ey2, d, dn);
input
  v,
  ex0,
  ex1,
  ex2,
  ey0,
  ey1,
  ey2,
  a2,
  a3,
  a4,
  a5,
  a6,
  x0,
  x1,
  x2,
  x3,
  y0,
  y1,
  y2,
  y3,
  z0,
  z1,
  z2;
output
  d,
  dn;
wire
  \[120] ,
  \[638] ,
  \[590] ,
  \[566] ,
  \[398] ,
  \[345] ,
  \[592] ,
  \[568] ,
  \[514] ,
  \[123] ,
  \[346] ,
  \[124] ,
  \[347] ,
  \[594] ,
  \[540] ,
  \[516] ,
  \[348] ,
  \[614] ,
  \[349] ,
  \[596] ,
  \[542] ,
  \[128] ,
  \[640] ,
  \[375] ,
  \[616] ,
  \[321] ,
  \[598] ,
  \[544] ,
  \[77] ,
  \[129] ,
  \[376] ,
  \[250] ,
  \[78] ,
  \[642] ,
  \[618] ,
  \[570] ,
  \[546] ,
  \[644] ,
  \[572] ,
  \[157] ,
  \[350] ,
  \[646] ,
  \[351] ,
  \[327] ,
  \[574] ,
  \[352] ,
  \[328] ,
  \[130] ,
  \[353] ,
  \[329] ,
  \[576] ,
  \[522] ,
  \[578] ,
  \[524] ,
  \[526] ,
  \[358] ,
  \[359] ,
  \[552] ,
  \[626] ,
  \[554] ,
  \[628] ,
  \[580] ,
  \[237] ,
  \[557] ,
  \[503] ,
  \[335] ,
  \[582] ,
  \[360] ,
  \[336] ,
  \[505] ,
  \[361] ,
  \[337] ,
  \[584] ,
  \[362] ,
  \[338] ,
  \[363] ,
  \[339] ,
  \[586] ,
  \[532] ,
  \[508] ,
  \[117] ,
  \[90] ,
  \[118] ,
  \[630] ,
  \[588] ,
  \[91] ,
  \[119] ,
  \[535] ,
  \[632] ,
  \[367] ,
  \[608] ,
  \[560] ,
  \[392] ,
  \[368] ,
  \[537] ,
  \[0] ,
  \[634] ,
  \[1] ,
  \[340] ,
  \[563] ,
  \[636] ,
  \[511] ;
assign
  \[120]  = ~\[339]  & (~\[338]  & ~\[340] ),
  \[638]  = ~x3 | ~\[361] ,
  \[590]  = ~\[566]  | ~\[368] ,
  \[566]  = ~\[367] ,
  \[398]  = ~v,
  \[345]  = ~y0,
  \[592]  = ~x2 | ~\[362] ,
  \[568]  = ~\[540]  | ~\[398] ,
  \[514]  = ~\[608]  | ~\[398] ,
  \[123]  = ~\[338]  & ~\[77] ,
  \[346]  = ~y1,
  \[124]  = ~\[78]  & ~ex1,
  \[347]  = ~\[646]  | ~\[644] ,
  \[594]  = ~x3 | ~\[361] ,
  \[540]  = ~\[570]  | (~\[508]  | ~\[505] ),
  \[516]  = ~\[618]  | (~\[616]  | (~\[237]  | ~\[614] )),
  \[348]  = ~y2,
  \[614]  = ~ey1 | ~\[522] ,
  d = \[0] ,
  \[349]  = ~y3,
  \[596]  = ~\[359]  | ~\[358] ,
  \[542]  = ~\[574]  | ~\[572] ,
  \[128]  = ~\[352]  & (~z1 & ~z2),
  \[640]  = ~x0 | ~\[359] ,
  \[375]  = ~\[586]  | ~\[584] ,
  \[616]  = ~\[524]  | ~\[335] ,
  \[321]  = ~a5 & ~a2,
  \[598]  = ~x1 | ~x0,
  \[544]  = ~\[578]  | ~\[576] ,
  \[77]  = ~\[340]  & ~\[339] ,
  \[129]  = ~\[353]  & (~z0 & ~\[351] ),
  \[376]  = ~\[582]  | ~\[580] ,
  \[250]  = ~\[129]  & (~\[128]  & ~\[130] ),
  \[78]  = ~ex2 & ~ex0,
  \[642]  = ~x1 | ~\[358] ,
  \[618]  = ~\[526]  | ~\[508] ,
  \[570]  = ~\[542]  | (~\[544]  | (~\[157]  | ~\[546] )),
  \[546]  = ~\[590]  | ~\[588] ,
  \[644]  = ~y0 | ~\[346] ,
  \[572]  = ~z0 | ~\[552] ,
  \[157]  = ~\[90]  & ~\[91] ,
  \[350]  = ~\[634]  | ~\[632] ,
  \[646]  = ~y1 | ~\[345] ,
  \[351]  = ~z2,
  \[327]  = ~a3,
  \[574]  = ~\[554]  | ~\[352] ,
  \[352]  = ~z0,
  \[328]  = ~a6,
  \[130]  = ~\[350]  & ~\[537] ,
  \[353]  = ~z1,
  \[329]  = ~a4,
  \[576]  = ~\[557]  | ~\[375] ,
  \[522]  = ~ey2 | ~ey0,
  \[578]  = ~\[560]  | ~\[376] ,
  \[524]  = ~\[337]  | ~\[336] ,
  \[526]  = ~\[628]  | (~\[626]  | (~\[630]  | ~\[250] )),
  \[358]  = ~x0,
  \[359]  = ~x1,
  \[552]  = ~\[351]  | ~\[353] ,
  dn = \[1] ,
  \[626]  = ~\[537]  | ~\[350] ,
  \[554]  = ~z1 | ~z2,
  \[628]  = ~\[532]  | ~\[360] ,
  \[580]  = ~y2 | ~\[349] ,
  \[237]  = ~\[124]  & ~\[123] ,
  \[557]  = ~\[376] ,
  \[503]  = ~\[514]  | ~\[511] ,
  \[335]  = ~ey1,
  \[582]  = ~y3 | ~\[348] ,
  \[360]  = ~\[642]  | ~\[640] ,
  \[336]  = ~ey0,
  \[505]  = ~\[392]  | (~\[327]  | (~a4 | ~a6)),
  \[361]  = ~x2,
  \[337]  = ~ey2,
  \[584]  = ~\[346]  | ~\[345] ,
  \[362]  = ~x3,
  \[338]  = ~ex1,
  \[363]  = ~\[638]  | ~\[636] ,
  \[339]  = ~ex0,
  \[586]  = ~y1 | ~y0,
  \[532]  = ~\[363] ,
  \[508]  = ~a3 | (~\[392]  | (~a6 | ~\[329] )),
  \[117]  = ~ey1 & (~ey0 & ~ey2),
  \[90]  = ~\[118]  & ~\[117] ,
  \[118]  = ~\[336]  & (~\[335]  & ~\[337] ),
  \[630]  = ~\[535]  | ~\[363] ,
  \[588]  = ~\[563]  | ~\[367] ,
  \[91]  = ~\[120]  & ~\[119] ,
  \[119]  = ~ex1 & (~ex0 & ~ex2),
  \[535]  = ~\[360] ,
  \[632]  = ~y2 | ~\[349] ,
  \[367]  = ~\[598]  | ~\[596] ,
  \[608]  = ~\[516]  | ~\[505] ,
  \[560]  = ~\[375] ,
  \[392]  = ~a2,
  \[368]  = ~\[594]  | ~\[592] ,
  \[537]  = ~\[347] ,
  \[0]  = ~\[503] ,
  \[634]  = ~y3 | ~\[348] ,
  \[1]  = ~\[568]  | ~\[511] ,
  \[340]  = ~ex2,
  \[563]  = ~\[368] ,
  \[636]  = ~x2 | ~\[362] ,
  \[511]  = ~\[329]  | (~\[328]  | (~\[327]  | ~\[321] ));
endmodule

