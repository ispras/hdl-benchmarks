// IWLS benchmark module "i7" printed on Wed May 29 17:26:51 2002
module i7(\V199(1) , \V32(27) , \V199(0) , \V32(26) , \V32(25) , \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V96(27) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V128(27) , \V199(4) , \V128(26) , \V128(25) , \V128(24) , \V128(23) , \V128(22) , \V128(21) , \V128(20) , \V128(19) , \V128(18) , \V128(17) , \V128(16) , \V128(15) , \V128(14) , \V128(13) , \V128(12) , \V128(11) , \V128(10) , \V128(9) , \V128(8) , \V128(7) , \V128(6) , \V128(5) , \V128(4) , \V128(3) , \V128(2) , \V128(1) , \V128(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V192(27) , \V192(26) , \V192(25) , \V192(24) , \V192(23) , \V192(22) , \V192(21) , \V192(20) , \V192(19) , \V192(18) , \V192(17) , \V192(16) , \V192(15) , \V192(14) , \V192(13) , \V192(12) , \V192(11) , \V192(10) , \V192(9) , \V192(8) , \V192(7) , \V192(6) , \V192(5) , \V192(4) , \V192(3) , \V192(2) , \V192(1) , \V192(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V160(27) , \V160(26) , \V160(25) , \V160(24) , \V160(23) , \V160(22) , \V160(21) , \V160(20) , \V160(19) , \V160(18) , \V160(17) , \V160(16) , \V160(15) , \V160(14) , \V160(13) , \V160(12) , \V160(11) , \V160(10) , \V160(9) , \V160(8) , \V160(7) , \V160(6) , \V160(5) , \V160(4) , \V160(3) , \V160(2) , \V160(1) , \V160(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V128(31) , \V199(3) , \V128(30) , \V128(29) , \V128(28) , \V195(0) , \V194(1) , \V194(0) , \V192(31) , \V192(30) , \V192(29) , \V192(28) , \V160(31) , \V160(30) , \V160(29) , \V160(28) , \V227(27) , \V227(26) , \V227(25) , \V227(24) , \V227(23) , \V227(22) , \V227(21) , \V227(20) , \V227(19) , \V227(18) , \V227(17) , \V227(16) , \V227(15) , \V227(14) , \V227(13) , \V227(12) , \V227(11) , \V227(10) , \V227(9) , \V227(8) , \V227(7) , \V227(6) , \V227(5) , \V227(4) , \V227(3) , \V227(2) , \V227(1) , \V227(0) , \V259(31) , \V259(30) , \V259(29) , \V259(28) , \V259(27) , \V259(26) , \V259(25) , \V259(24) , \V259(23) , \V259(22) , \V259(21) , \V259(20) , \V259(19) , \V259(18) , \V259(17) , \V259(16) , \V259(15) , \V259(14) , \V259(13) , \V259(12) , \V259(11) , \V259(10) , \V259(9) , \V259(8) , \V259(7) , \V259(6) , \V259(5) , \V259(4) , \V259(3) , \V259(2) , \V259(1) , \V259(0) , \V266(6) , \V266(5) , \V266(4) , \V266(3) , \V266(2) , \V266(1) , \V266(0) );
input
  \V32(30) ,
  \V199(1) ,
  \V199(0) ,
  \V128(21) ,
  \V128(20) ,
  \V192(31) ,
  \V128(23) ,
  \V192(30) ,
  \V128(22) ,
  \V160(3) ,
  \V128(25) ,
  \V160(2) ,
  \V128(24) ,
  \V160(5) ,
  \V128(17) ,
  \V160(4) ,
  \V128(16) ,
  \V128(19) ,
  \V128(18) ,
  \V160(1) ,
  \V160(0) ,
  \V160(7) ,
  \V128(11) ,
  \V160(6) ,
  \V128(10) ,
  \V160(9) ,
  \V128(13) ,
  \V160(8) ,
  \V160(31) ,
  \V128(12) ,
  \V160(30) ,
  \V128(15) ,
  \V128(3) ,
  \V128(14) ,
  \V128(2) ,
  \V128(5) ,
  \V128(4) ,
  \V128(1) ,
  \V128(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V128(7) ,
  \V32(4) ,
  \V128(6) ,
  \V32(5) ,
  \V128(9) ,
  \V32(6) ,
  \V128(8) ,
  \V32(7) ,
  \V32(8) ,
  \V32(9) ,
  \V96(0) ,
  \V96(1) ,
  \V96(2) ,
  \V96(3) ,
  \V96(4) ,
  \V96(13) ,
  \V96(5) ,
  \V128(31) ,
  \V96(12) ,
  \V96(6) ,
  \V128(30) ,
  \V96(15) ,
  \V96(7) ,
  \V96(14) ,
  \V96(8) ,
  \V96(9) ,
  \V96(11) ,
  \V96(10) ,
  \V96(17) ,
  \V96(16) ,
  \V96(19) ,
  \V96(18) ,
  \V96(23) ,
  \V96(22) ,
  \V64(13) ,
  \V96(25) ,
  \V64(12) ,
  \V96(24) ,
  \V64(15) ,
  \V64(14) ,
  \V192(27) ,
  \V96(21) ,
  \V192(26) ,
  \V96(20) ,
  \V192(29) ,
  \V64(11) ,
  \V192(28) ,
  \V64(10) ,
  \V192(3) ,
  \V192(2) ,
  \V192(5) ,
  \V96(27) ,
  \V192(4) ,
  \V96(26) ,
  \V64(17) ,
  \V96(29) ,
  \V64(16) ,
  \V96(28) ,
  \V192(21) ,
  \V64(19) ,
  \V192(1) ,
  \V192(20) ,
  \V64(18) ,
  \V192(0) ,
  \V192(23) ,
  \V64(23) ,
  \V192(22) ,
  \V64(22) ,
  \V32(13) ,
  \V192(25) ,
  \V64(25) ,
  \V32(12) ,
  \V192(24) ,
  \V64(24) ,
  \V32(15) ,
  \V192(17) ,
  \V192(7) ,
  \V32(14) ,
  \V96(31) ,
  \V192(16) ,
  \V160(27) ,
  \V192(6) ,
  \V96(30) ,
  \V192(19) ,
  \V64(21) ,
  \V160(26) ,
  \V192(9) ,
  \V192(18) ,
  \V64(20) ,
  \V160(29) ,
  \V192(8) ,
  \V32(11) ,
  \V160(28) ,
  \V32(10) ,
  \V194(1) ,
  \V194(0) ,
  \V64(27) ,
  \V64(26) ,
  \V32(17) ,
  \V192(11) ,
  \V64(29) ,
  \V32(16) ,
  \V192(10) ,
  \V64(28) ,
  \V160(21) ,
  \V32(19) ,
  \V192(13) ,
  \V160(20) ,
  \V32(18) ,
  \V192(12) ,
  \V160(23) ,
  \V32(23) ,
  \V64(0) ,
  \V192(15) ,
  \V160(22) ,
  \V195(0) ,
  \V32(22) ,
  \V64(1) ,
  \V192(14) ,
  \V160(25) ,
  \V32(25) ,
  \V64(2) ,
  \V160(24) ,
  \V32(24) ,
  \V64(3) ,
  \V160(17) ,
  \V64(4) ,
  \V64(31) ,
  \V160(16) ,
  \V64(5) ,
  \V64(30) ,
  \V160(19) ,
  \V32(21) ,
  \V64(6) ,
  \V160(18) ,
  \V32(20) ,
  \V64(7) ,
  \V64(8) ,
  \V64(9) ,
  \V32(27) ,
  \V32(26) ,
  \V160(11) ,
  \V32(29) ,
  \V160(10) ,
  \V32(28) ,
  \V160(13) ,
  \V160(12) ,
  \V128(27) ,
  \V160(15) ,
  \V128(26) ,
  \V160(14) ,
  \V128(29) ,
  \V199(3) ,
  \V128(28) ,
  \V32(31) ,
  \V199(4) ;
output
  \V259(27) ,
  \V259(26) ,
  \V259(29) ,
  \V227(3) ,
  \V259(28) ,
  \V227(2) ,
  \V227(5) ,
  \V227(4) ,
  \V227(1) ,
  \V227(0) ,
  \V259(21) ,
  \V259(20) ,
  \V259(23) ,
  \V259(22) ,
  \V259(25) ,
  \V227(7) ,
  \V259(24) ,
  \V227(6) ,
  \V259(17) ,
  \V227(9) ,
  \V259(16) ,
  \V227(8) ,
  \V227(27) ,
  \V259(19) ,
  \V227(26) ,
  \V259(18) ,
  \V259(11) ,
  \V259(10) ,
  \V227(21) ,
  \V259(13) ,
  \V227(20) ,
  \V259(12) ,
  \V227(23) ,
  \V266(3) ,
  \V259(15) ,
  \V227(22) ,
  \V266(2) ,
  \V259(14) ,
  \V227(25) ,
  \V266(5) ,
  \V227(24) ,
  \V266(4) ,
  \V227(17) ,
  \V227(16) ,
  \V227(19) ,
  \V266(1) ,
  \V227(18) ,
  \V266(0) ,
  \V266(6) ,
  \V227(11) ,
  \V227(10) ,
  \V227(13) ,
  \V227(12) ,
  \V227(15) ,
  \V227(14) ,
  \V259(31) ,
  \V259(30) ,
  \V259(3) ,
  \V259(2) ,
  \V259(5) ,
  \V259(4) ,
  \V259(1) ,
  \V259(0) ,
  \V259(7) ,
  \V259(6) ,
  \V259(9) ,
  \V259(8) ;
wire
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[70] ,
  \[5] ,
  \[71] ,
  \[6] ,
  \[72] ,
  \[7] ,
  \[73] ,
  \[8] ,
  \[74] ,
  \[9] ,
  \[75] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  V572,
  \[35] ,
  V586,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ;
assign
  \[60]  = \V195(0)  & (\V199(3)  & ~\V199(0) ),
  \[61]  = (\[74]  & \V194(1) ) | ((~\V194(1)  & \V199(1) ) | (\[73]  | V586)),
  \[62]  = (\[74]  & \V194(0) ) | ((~\V194(0)  & \V199(1) ) | (\[73]  | V586)),
  \[63]  = (\[75]  & \V128(31) ) | ((\[74]  & \V192(31) ) | ((\[68]  & ~\V192(31) ) | ((V586 & \V160(31) ) | \[73] ))),
  \[64]  = (\[75]  & \V128(30) ) | ((\[74]  & \V192(30) ) | ((\[68]  & ~\V192(30) ) | ((V586 & \V160(30) ) | \[73] ))),
  \[65]  = (\[75]  & \V128(29) ) | ((\[74]  & \V192(29) ) | ((\[68]  & ~\V192(29) ) | ((V586 & \V160(29) ) | \[73] ))),
  \[66]  = (\[75]  & \V128(28) ) | ((\[74]  & \V192(28) ) | ((\[68]  & ~\V192(28) ) | ((V586 & \V160(28) ) | \[73] ))),
  \[67]  = ~\V199(0)  & ~\V199(1) ,
  \[68]  = ~\V199(0)  & \V199(1) ,
  \[69]  = \V199(0)  & ~\V199(1) ,
  \[0]  = (\[70]  & \V64(27) ) | ((\[69]  & \V32(27) ) | ((\[68]  & ~\V96(27) ) | (\[67]  & \V96(27) ))),
  \[1]  = (\[70]  & \V64(26) ) | ((\[69]  & \V32(26) ) | ((\[68]  & ~\V96(26) ) | (\[67]  & \V96(26) ))),
  \[2]  = (\[70]  & \V64(25) ) | ((\[69]  & \V32(25) ) | ((\[68]  & ~\V96(25) ) | (\[67]  & \V96(25) ))),
  \[3]  = (\[70]  & \V64(24) ) | ((\[69]  & \V32(24) ) | ((\[68]  & ~\V96(24) ) | (\[67]  & \V96(24) ))),
  \[4]  = (\[70]  & \V64(23) ) | ((\[69]  & \V32(23) ) | ((\[68]  & ~\V96(23) ) | (\[67]  & \V96(23) ))),
  \[70]  = \V199(0)  & \V199(1) ,
  \[5]  = (\[70]  & \V64(22) ) | ((\[69]  & \V32(22) ) | ((\[68]  & ~\V96(22) ) | (\[67]  & \V96(22) ))),
  \[71]  = \[69]  & \V199(4) ,
  \[6]  = (\[70]  & \V64(21) ) | ((\[69]  & \V32(21) ) | ((\[68]  & ~\V96(21) ) | (\[67]  & \V96(21) ))),
  \[72]  = \[67]  & \V199(4) ,
  \[7]  = (\[70]  & \V64(20) ) | ((\[69]  & \V32(20) ) | ((\[68]  & ~\V96(20) ) | (\[67]  & \V96(20) ))),
  \[73]  = ~\V199(3)  & \V199(1) ,
  \[8]  = (\[70]  & \V64(19) ) | ((\[69]  & \V32(19) ) | ((\[68]  & ~\V96(19) ) | (\[67]  & \V96(19) ))),
  \[74]  = \[67]  & \V199(3) ,
  \[9]  = (\[70]  & \V64(18) ) | ((\[69]  & \V32(18) ) | ((\[68]  & ~\V96(18) ) | (\[67]  & \V96(18) ))),
  \[75]  = \[69]  & \V199(3) ,
  \V259(27)  = \[32] ,
  \V259(26)  = \[33] ,
  \V259(29)  = \[30] ,
  \V227(3)  = \[24] ,
  \V259(28)  = \[31] ,
  \V227(2)  = \[25] ,
  \V227(5)  = \[22] ,
  \V227(4)  = \[23] ,
  \V227(1)  = \[26] ,
  \V227(0)  = \[27] ,
  \V259(21)  = \[38] ,
  \V259(20)  = \[39] ,
  \V259(23)  = \[36] ,
  \V259(22)  = \[37] ,
  \V259(25)  = \[34] ,
  \V227(7)  = \[20] ,
  \V259(24)  = \[35] ,
  \V227(6)  = \[21] ,
  \V259(17)  = \[42] ,
  \V227(9)  = \[18] ,
  \V259(16)  = \[43] ,
  \V227(8)  = \[19] ,
  \V227(27)  = \[0] ,
  \V259(19)  = \[40] ,
  \V227(26)  = \[1] ,
  \[10]  = (\[70]  & \V64(17) ) | ((\[69]  & \V32(17) ) | ((\[68]  & ~\V96(17) ) | (\[67]  & \V96(17) ))),
  \V259(18)  = \[41] ,
  \[11]  = (\[70]  & \V64(16) ) | ((\[69]  & \V32(16) ) | ((\[68]  & ~\V96(16) ) | (\[67]  & \V96(16) ))),
  \[12]  = (\[70]  & \V64(15) ) | ((\[69]  & \V32(15) ) | ((\[68]  & ~\V96(15) ) | (\[67]  & \V96(15) ))),
  \[13]  = (\[70]  & \V64(14) ) | ((\[69]  & \V32(14) ) | ((\[68]  & ~\V96(14) ) | (\[67]  & \V96(14) ))),
  \[14]  = (\[70]  & \V64(13) ) | ((\[69]  & \V32(13) ) | ((\[68]  & ~\V96(13) ) | (\[67]  & \V96(13) ))),
  \[15]  = (\[70]  & \V64(12) ) | ((\[69]  & \V32(12) ) | ((\[68]  & ~\V96(12) ) | (\[67]  & \V96(12) ))),
  \[16]  = (\[70]  & \V64(11) ) | ((\[69]  & \V32(11) ) | ((\[68]  & ~\V96(11) ) | (\[67]  & \V96(11) ))),
  \[17]  = (\[70]  & \V64(10) ) | ((\[69]  & \V32(10) ) | ((\[68]  & ~\V96(10) ) | (\[67]  & \V96(10) ))),
  \V259(11)  = \[48] ,
  \[18]  = (\[70]  & \V64(9) ) | ((\[69]  & \V32(9) ) | ((\[68]  & ~\V96(9) ) | (\[67]  & \V96(9) ))),
  \V259(10)  = \[49] ,
  \V227(21)  = \[6] ,
  \[19]  = (\[70]  & \V64(8) ) | ((\[69]  & \V32(8) ) | ((\[68]  & ~\V96(8) ) | (\[67]  & \V96(8) ))),
  \V259(13)  = \[46] ,
  \V227(20)  = \[7] ,
  \V259(12)  = \[47] ,
  \V227(23)  = \[4] ,
  \V266(3)  = \[63] ,
  \V259(15)  = \[44] ,
  \V227(22)  = \[5] ,
  \V266(2)  = \[64] ,
  \V259(14)  = \[45] ,
  \V227(25)  = \[2] ,
  \V266(5)  = \[61] ,
  \V227(24)  = \[3] ,
  \V266(4)  = \[62] ,
  \V227(17)  = \[10] ,
  \V227(16)  = \[11] ,
  \[20]  = (\[70]  & \V64(7) ) | ((\[69]  & \V32(7) ) | ((\[68]  & ~\V96(7) ) | (\[67]  & \V96(7) ))),
  \V227(19)  = \[8] ,
  \V266(1)  = \[65] ,
  \[21]  = (\[70]  & \V64(6) ) | ((\[69]  & \V32(6) ) | ((\[68]  & ~\V96(6) ) | (\[67]  & \V96(6) ))),
  \V227(18)  = \[9] ,
  \V266(0)  = \[66] ,
  \[22]  = (\[70]  & \V64(5) ) | ((\[69]  & \V32(5) ) | ((\[68]  & ~\V96(5) ) | (\[67]  & \V96(5) ))),
  \[23]  = (\[70]  & \V64(4) ) | ((\[69]  & \V32(4) ) | ((\[68]  & ~\V96(4) ) | (\[67]  & \V96(4) ))),
  \[24]  = (\[70]  & \V64(3) ) | ((\[69]  & \V32(3) ) | ((\[68]  & ~\V96(3) ) | (\[67]  & \V96(3) ))),
  \[25]  = (\[70]  & \V64(2) ) | ((\[69]  & \V32(2) ) | ((\[68]  & ~\V96(2) ) | (\[67]  & \V96(2) ))),
  \[26]  = (\[70]  & \V64(1) ) | ((\[69]  & \V32(1) ) | ((\[68]  & ~\V96(1) ) | (\[67]  & \V96(1) ))),
  \[27]  = (\[70]  & \V64(0) ) | ((\[69]  & \V32(0) ) | ((\[68]  & ~\V96(0) ) | (\[67]  & \V96(0) ))),
  \V266(6)  = \[60] ,
  \[28]  = (\[72]  & \V192(27) ) | ((\[71]  & \V128(27) ) | ((\[70]  & \V160(27) ) | ((\[68]  & ~\V192(27) ) | V572))),
  \V227(11)  = \[16] ,
  \[29]  = (\[72]  & \V192(26) ) | ((\[71]  & \V128(26) ) | ((\[70]  & \V160(26) ) | ((\[68]  & ~\V192(26) ) | V572))),
  \V227(10)  = \[17] ,
  \V227(13)  = \[14] ,
  \V227(12)  = \[15] ,
  \V227(15)  = \[12] ,
  \V227(14)  = \[13] ,
  \[30]  = (\[72]  & \V192(25) ) | ((\[71]  & \V128(25) ) | ((\[70]  & \V160(25) ) | ((\[68]  & ~\V192(25) ) | V572))),
  \[31]  = (\[72]  & \V192(24) ) | ((\[71]  & \V128(24) ) | ((\[70]  & \V160(24) ) | ((\[68]  & ~\V192(24) ) | V572))),
  \[32]  = (\[72]  & \V192(23) ) | ((\[71]  & \V128(23) ) | ((\[70]  & \V160(23) ) | ((\[68]  & ~\V192(23) ) | V572))),
  \[33]  = (\[72]  & \V192(22) ) | ((\[71]  & \V128(22) ) | ((\[70]  & \V160(22) ) | ((\[68]  & ~\V192(22) ) | V572))),
  \[34]  = (\[72]  & \V192(21) ) | ((\[71]  & \V128(21) ) | ((\[70]  & \V160(21) ) | ((\[68]  & ~\V192(21) ) | V572))),
  V572 = ~\V199(4)  & \V199(1) ,
  \[35]  = (\[72]  & \V192(20) ) | ((\[71]  & \V128(20) ) | ((\[70]  & \V160(20) ) | ((\[68]  & ~\V192(20) ) | V572))),
  V586 = \[70] ,
  \[36]  = (\[72]  & \V192(19) ) | ((\[71]  & \V128(19) ) | ((\[70]  & \V160(19) ) | ((\[68]  & ~\V192(19) ) | V572))),
  \[37]  = (\[72]  & \V192(18) ) | ((\[71]  & \V128(18) ) | ((\[70]  & \V160(18) ) | ((\[68]  & ~\V192(18) ) | V572))),
  \V259(31)  = \[28] ,
  \[38]  = (\[72]  & \V192(17) ) | ((\[71]  & \V128(17) ) | ((\[70]  & \V160(17) ) | ((\[68]  & ~\V192(17) ) | V572))),
  \V259(30)  = \[29] ,
  \[39]  = (\[72]  & \V192(16) ) | ((\[71]  & \V128(16) ) | ((\[70]  & \V160(16) ) | ((\[68]  & ~\V192(16) ) | V572))),
  \[40]  = (\[72]  & \V192(15) ) | ((\[71]  & \V128(15) ) | ((\[70]  & \V160(15) ) | ((\[68]  & ~\V192(15) ) | V572))),
  \[41]  = (\[72]  & \V192(14) ) | ((\[71]  & \V128(14) ) | ((\[70]  & \V160(14) ) | ((\[68]  & ~\V192(14) ) | V572))),
  \[42]  = (\[72]  & \V192(13) ) | ((\[71]  & \V128(13) ) | ((\[70]  & \V160(13) ) | ((\[68]  & ~\V192(13) ) | V572))),
  \[43]  = (\[72]  & \V192(12) ) | ((\[71]  & \V128(12) ) | ((\[70]  & \V160(12) ) | ((\[68]  & ~\V192(12) ) | V572))),
  \[44]  = (\[72]  & \V192(11) ) | ((\[71]  & \V128(11) ) | ((\[70]  & \V160(11) ) | ((\[68]  & ~\V192(11) ) | V572))),
  \V259(3)  = \[56] ,
  \[45]  = (\[72]  & \V192(10) ) | ((\[71]  & \V128(10) ) | ((\[70]  & \V160(10) ) | ((\[68]  & ~\V192(10) ) | V572))),
  \V259(2)  = \[57] ,
  \[46]  = (\[72]  & \V192(9) ) | ((\[71]  & \V128(9) ) | ((\[70]  & \V160(9) ) | ((\[68]  & ~\V192(9) ) | V572))),
  \V259(5)  = \[54] ,
  \[47]  = (\[72]  & \V192(8) ) | ((\[71]  & \V128(8) ) | ((\[70]  & \V160(8) ) | ((\[68]  & ~\V192(8) ) | V572))),
  \V259(4)  = \[55] ,
  \[48]  = (\[72]  & \V192(7) ) | ((\[71]  & \V128(7) ) | ((\[70]  & \V160(7) ) | ((\[68]  & ~\V192(7) ) | V572))),
  \[49]  = (\[72]  & \V192(6) ) | ((\[71]  & \V128(6) ) | ((\[70]  & \V160(6) ) | ((\[68]  & ~\V192(6) ) | V572))),
  \V259(1)  = \[58] ,
  \V259(0)  = \[59] ,
  \[50]  = (\[72]  & \V192(5) ) | ((\[71]  & \V128(5) ) | ((\[70]  & \V160(5) ) | ((\[68]  & ~\V192(5) ) | V572))),
  \V259(7)  = \[52] ,
  \[51]  = (\[72]  & \V192(4) ) | ((\[71]  & \V128(4) ) | ((\[70]  & \V160(4) ) | ((\[68]  & ~\V192(4) ) | V572))),
  \V259(6)  = \[53] ,
  \[52]  = (\[72]  & \V192(3) ) | ((\[71]  & \V128(3) ) | ((\[70]  & \V160(3) ) | ((\[68]  & ~\V192(3) ) | V572))),
  \V259(9)  = \[50] ,
  \[53]  = (\[72]  & \V192(2) ) | ((\[71]  & \V128(2) ) | ((\[70]  & \V160(2) ) | ((\[68]  & ~\V192(2) ) | V572))),
  \V259(8)  = \[51] ,
  \[54]  = (\[72]  & \V192(1) ) | ((\[71]  & \V128(1) ) | ((\[70]  & \V160(1) ) | ((\[68]  & ~\V192(1) ) | V572))),
  \[55]  = (\[72]  & \V192(0) ) | ((\[71]  & \V128(0) ) | ((\[70]  & \V160(0) ) | ((\[68]  & ~\V192(0) ) | V572))),
  \[56]  = (\[72]  & \V96(31) ) | ((\[71]  & \V32(31) ) | ((\[70]  & \V64(31) ) | ((\[68]  & ~\V96(31) ) | V572))),
  \[57]  = (\[72]  & \V96(30) ) | ((\[71]  & \V32(30) ) | ((\[70]  & \V64(30) ) | ((\[68]  & ~\V96(30) ) | V572))),
  \[58]  = (\[72]  & \V96(29) ) | ((\[71]  & \V32(29) ) | ((\[70]  & \V64(29) ) | ((\[68]  & ~\V96(29) ) | V572))),
  \[59]  = (\[72]  & \V96(28) ) | ((\[71]  & \V32(28) ) | ((\[70]  & \V64(28) ) | ((\[68]  & ~\V96(28) ) | V572)));
endmodule

