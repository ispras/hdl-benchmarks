// IWLS benchmark module "pcle_cl" printed on Wed May 29 17:28:07 2002
module pcle_cl(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s;
output
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0;
wire
  \[7] ,
  \[8] ,
  \[9] ,
  \[10] ,
  \[0] ,
  \[11] ,
  \[1] ,
  u0,
  \[2] ,
  \[3] ,
  \[4] ,
  x0,
  \[5] ,
  \[6] ;
assign
  \[7]  = (~\[10]  & (u0 & ~r)) | ((\[10]  & (u0 & r)) | (i & g)),
  \[8]  = (~\[10]  & (u0 & (~\[0]  & r))) | ((u0 & (~\[0]  & s)) | (i & h)),
  \[9]  = ~m | ~l,
  \[10]  = ~x0 | ~q,
  \[0]  = ~\[10]  & (u0 & (s & r)),
  \[11]  = \[9]  | ~n,
  \[1]  = (u0 & ~l) | (i & a),
  u0 = ~k & (j & ~i),
  t = \[0] ,
  \[2]  = (~m & (l & u0)) | ((m & (~l & u0)) | (i & b)),
  u = \[1] ,
  v = \[2] ,
  w = \[3] ,
  \x  = \[4] ,
  y = \[5] ,
  z = \[6] ,
  \[3]  = (~\[9]  & (u0 & ~n)) | ((\[9]  & (u0 & n)) | (i & c)),
  \[4]  = (~\[11]  & (u0 & ~o)) | ((\[11]  & (u0 & o)) | (i & d)),
  a0 = \[7] ,
  x0 = ~\[11]  & (p & o),
  \[5]  = (~\[11]  & (~x0 & (u0 & o))) | ((~x0 & (u0 & p)) | (i & e)),
  b0 = \[8] ,
  \[6]  = (~x0 & (q & u0)) | ((x0 & (~q & u0)) | (i & f));
endmodule

