// IWLS benchmark module "term1" printed on Wed May 29 17:29:18 2002
module term1(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0;
output
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0;
wire
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  a2,
  a3,
  a4,
  a7,
  b3,
  b4,
  b5,
  b6,
  b7,
  c3,
  c4,
  c5,
  c6,
  d2,
  d3,
  d4,
  d6,
  e1,
  e2,
  e3,
  e4,
  e6,
  e7,
  f1,
  f2,
  f3,
  f4,
  f5,
  f6,
  f7,
  g2,
  g3,
  g4,
  g5,
  g6,
  g7,
  h1,
  h2,
  h3,
  h4,
  h5,
  h6,
  i2,
  i3,
  i4,
  i5,
  i6,
  i7,
  j1,
  j3,
  j4,
  j5,
  j6,
  j7,
  k2,
  k3,
  k4,
  k5,
  k6,
  k7,
  l2,
  l3,
  l4,
  l6,
  l7,
  m2,
  m3,
  m4,
  m5,
  m6,
  n2,
  n3,
  n4,
  n5,
  n6,
  o3,
  o4,
  o5,
  o6,
  o7,
  p3,
  p4,
  p5,
  p6,
  p7,
  q2,
  q3,
  q4,
  q5,
  q6,
  q7,
  r2,
  r3,
  r4,
  r5,
  s1,
  s2,
  s3,
  s4,
  s5,
  s6,
  t1,
  t2,
  t3,
  t4,
  t5,
  t6,
  u1,
  u2,
  u4,
  u5,
  u6,
  v2,
  v4,
  v5,
  v6,
  w1,
  w2,
  w3,
  w4,
  w5,
  w6,
  x1,
  x4,
  x5,
  y1,
  y2,
  y3,
  y4,
  y5,
  y6,
  z1,
  z2,
  z3,
  z4,
  z5,
  z6;
assign
  \[0]  = ~h0,
  \[1]  = (~t6 & ~c) | ((~t6 & d) | (~t6 & ~h0)),
  \[2]  = (y6 & (~v6 & b)) | (~w6 & (~v6 & ~b)),
  \[3]  = ~f1 & (~e1 & b),
  \[4]  = ~t1 & (~s1 & b),
  \[5]  = ~f2 & (~s1 & b),
  \[6]  = ~t2 & (~s1 & b),
  \[7]  = (~j3 & (q & u)) | ((~k3 & p) | ~l3),
  \[8]  = ~w3 & (a & ~a0),
  \[9]  = ~h5 & (a & ~a0),
  a2 = (~d2 & (p & t)) | ((~d2 & (p & y)) | ((~d2 & (u & t)) | (~d2 & (u & y)))),
  a3 = (~d3 & (~c3 & ~b3)) | ((~d3 & (~c3 & ~s)) | ((~d3 & (~c3 & ~w)) | ((~d3 & (~r & ~b3)) | ((~d3 & (~r & ~s)) | (~d3 & (~r & ~w)))))),
  a4 = (~m4 & ~r) | ((~l4 & ~q) | ~n4),
  a7 = (~b7 & ~d) | ((~b7 & ~e) | (~b7 & ~h)),
  b3 = t | y,
  b4 = ~k4 & (q & r),
  b5 = ~q | (~r | ~s),
  b6 = ~f0 | ~g0,
  b7 = (~e7 & d) | ((~e7 & e) | (~e7 & h)),
  c3 = (\x  & y) | ((\x  & t) | ((s & y) | (s & t))),
  c4 = (~f4 & (~e4 & ~d4)) | ((~f4 & (~e4 & ~e0)) | ((~f4 & (~e4 & ~f0)) | ((~f4 & (q & ~d4)) | ((~f4 & (q & ~e0)) | (~f4 & (q & ~f0)))))),
  c5 = (~f0 & (~d0 & ~c0)) | (~f0 & ~e0),
  c6 = (~l6 & q) | ((~s5 & ~q) | ~m6),
  d2 = (~w & ~r) | ((~v & ~q) | (~\x  & ~s)),
  d3 = (\x  & (t & w)) | ((\x  & (y & w)) | (e0 & (d0 & c0))),
  d4 = c0 | d0,
  d6 = f0 | g0,
  e1 = ~z | (a0 | c0),
  e2 = (~w & ~r) | ((~\x  & ~s) | (~u & ~p)),
  e3 = c0 & (d0 & e0),
  e4 = ~r | (~s | ~t),
  e6 = (d0 & e0) | ((~i6 & r) | ~j6),
  e7 = (e & h) | ((e & d) | (h & d)),
  f1 = (d & c) | ~h1,
  f2 = (~i2 & (~h2 & ~w1)) | ((~i2 & (~h2 & ~g2)) | ((~i2 & (~h2 & ~c0)) | ((~i2 & (c & ~w1)) | ((~i2 & (c & ~g2)) | ((~i2 & (c & ~c0)) | ((~i2 & (~e0 & ~w1)) | ((~i2 & (~e0 & ~g2)) | (~i2 & (~e0 & ~c0))))))))),
  f3 = (~g3 & (s & w)) | ((~h3 & r) | ~i3),
  f4 = (~f0 & (~d0 & ~c0)) | ((~f0 & ~e0) | ~g4),
  f5 = ~c0 & ~d0,
  f6 = ~g6 | (f0 | g0),
  f7 = (~g7 & ~d) | ((~g7 & e) | (~g7 & h)),
  g2 = d0 & ~e0,
  g3 = ~t & ~y,
  g4 = (~h4 & (t & r)) | (~h4 & s),
  g5 = (e0 & d0) | ((e0 & c0) | f0),
  g6 = (~h6 & (~d0 & ~c0)) | (~h6 & ~e0),
  g7 = (e & h) | ((e & ~d) | (h & ~d)),
  h1 = (~t & ~y) | ((~s & ~\x ) | ~j1),
  h2 = (~z1 & ~d0) | (~r2 & ~c0),
  h3 = (~\x  & ~s) | (~y & ~t),
  h4 = (~r & ~t) | (~i4 | ~g0),
  h5 = (~n5 & (~m5 & ~k5)) | ((~n5 & (~m5 & ~j5)) | ((~n5 & (~m5 & ~i5)) | ((~n5 & (~p & ~k5)) | ((~n5 & (~p & ~j5)) | ((~n5 & (~p & ~i5)) | ((~n5 & (i0 & ~k5)) | ((~n5 & (i0 & ~j5)) | (~n5 & (i0 & ~i5))))))))),
  h6 = ~s5 | (~l | q),
  i2 = ~k2 & (~d & e0),
  i3 = (~e0 & (~y & ~t)) | ((~d0 & (~y & ~t)) | ((~c0 & (~y & ~t)) | ((~e0 & ~\x ) | ((~e0 & ~w) | ((~d0 & ~\x ) | ((~d0 & ~w) | ((~c0 & ~\x ) | (~c0 & ~w)))))))),
  i4 = ~j4 | (~s | ~t),
  i5 = ~s6 & (k & ~p),
  i6 = (n & ~s) | ((o & ~t) | (~t & ~s)),
  i7 = (~q7 & (~p7 & ~o7)) | ((~q7 & (~p7 & d)) | ((~q7 & (~p7 & ~f)) | ((~q7 & (e & ~o7)) | ((~q7 & (e & d)) | ((~q7 & (e & ~f)) | ((~q7 & (~h & ~o7)) | ((~q7 & (~h & d)) | (~q7 & (~h & ~f))))))))),
  j0 = \[0] ,
  j1 = (w & (v & u)) | ((w & (v & p)) | ((w & (q & u)) | ((w & (q & p)) | ((r & (v & u)) | ((r & (v & p)) | ((r & (q & u)) | (r & (q & p)))))))),
  j3 = (~w & ~r) | ((~\x  & ~s) | (~y & ~t)),
  j4 = ~k & (q & r),
  j5 = q & (r & s),
  j6 = (~k6 & (s & ~c0)) | ((~k6 & (s & ~e0)) | ((~k6 & (t & ~c0)) | (~k6 & (t & ~e0)))),
  j7 = (~h & (~g & ~e)) | ((~h & (~e & c)) | ((h & (~g & e)) | (h & (e & c)))),
  k0 = \[1] ,
  k2 = (~m2 & ~l2) | ((~m2 & c0) | ((d0 & ~l2) | (d0 & c0))),
  k3 = (~s3 & (~m3 & ~c3)) | ((~s3 & (~m3 & ~r)) | ((~s3 & (~m3 & ~v)) | ((~s3 & (~q & ~c3)) | ((~s3 & (~q & ~r)) | (~s3 & (~q & ~v)))))),
  k4 = ~s | ~t,
  k5 = (~q6 & (~f0 & ~g0)) | (~f5 & (~b6 & e0)),
  k6 = (t & (s & ~m)) | ((~t & ~r) | ((~s & ~r) | (~r & ~m))),
  k7 = (~l7 & ~e) | (~l7 & ~h),
  l0 = \[2] ,
  l2 = (~t & ~y) | ((~r & ~w) | ~q2),
  l3 = (~o3 & (~n3 & ~m3)) | ((~o3 & (~n3 & ~u)) | ((~o3 & (~n3 & ~v)) | ((~o3 & (~g0 & ~m3)) | ((~o3 & (~g0 & ~u)) | (~o3 & (~g0 & ~v)))))),
  l4 = ~k4 & (~l & r),
  l6 = (~m4 & ~r) | ~n4,
  l7 = (g & ~c) | ((~h & ~e) | (f & ~d)),
  m0 = \[3] ,
  m2 = (~p & ~u) | ((~t & ~y) | ~n2),
  m3 = (w & (\x  & y)) | ((w & (\x  & t)) | ((w & (s & y)) | ((w & (s & t)) | ((r & (\x  & y)) | ((r & (\x  & t)) | ((r & (s & y)) | (r & (s & t)))))))),
  m4 = ~m & (s & t),
  m5 = (~e6 & (~d6 & q)) | ((~c6 & (~b6 & e0)) | ~f6),
  m6 = (~n6 & (s & c0)) | ((~n6 & (s & d0)) | ((~n6 & (t & c0)) | (~n6 & (t & d0)))),
  n0 = \[4] ,
  n2 = (v & (w & \x )) | ((v & (w & s)) | ((v & (r & \x )) | ((v & (r & s)) | ((q & (w & \x )) | ((q & (w & s)) | ((q & (r & \x )) | (q & (r & s)))))))),
  n3 = ~r3 | (~c0 | ~d0),
  n4 = (s & t) | ((s & ~o) | (t & ~n)),
  n5 = ~o5 & i0,
  n6 = (~t & ~r) | ((~s & ~r) | ~o6),
  o0 = \[5] ,
  o3 = ~p3 | (~z | ~b),
  o4 = ~k | (p | ~q),
  o5 = (~r5 & (~q5 & ~p5)) | ((~r5 & (~q5 & ~p)) | (~r5 & (~p5 & p))),
  o6 = ~p6 | ~t,
  o7 = (~h & ~e) | (h & e),
  p0 = \[6] ,
  p3 = (~q3 & (~a0 & ~c)) | (~q3 & (~a0 & ~d)),
  p4 = (~f5 & (e0 & f0)) | ~g5,
  p5 = (~z5 & (~y5 & ~x5)) | ((~z5 & (~y5 & q)) | ((~z5 & (r & ~x5)) | (~z5 & (r & q)))),
  p6 = ~l & (r & s),
  p7 = d | ~f,
  q0 = \[7] ,
  q2 = (\x  & (v & u)) | ((\x  & (v & p)) | ((\x  & (q & u)) | ((\x  & (q & p)) | ((s & (v & u)) | ((s & (v & p)) | ((s & (q & u)) | (s & (q & p)))))))),
  q3 = ~z2 & (f0 & ~g0),
  q4 = ~l | (~p | q),
  q5 = ~w5 | (~q | ~r),
  q6 = (e0 & d0) | (e0 & c0),
  q7 = (e & (~h & ~f)) | (e & (~h & d)),
  r0 = \[8] ,
  r2 = (~s2 & (t & r)) | ((~s2 & (t & w)) | ((~s2 & (y & r)) | (~s2 & (y & w)))),
  r3 = e0 & f0,
  r4 = (~x4 & (~w4 & ~t4)) | ((~x4 & (~w4 & ~s4)) | ((~x4 & (~v4 & ~t4)) | ((~x4 & (~v4 & ~s4)) | (~x4 & ~u4)))),
  r5 = (~f5 & (e0 & ~g0)) | ((~s5 & ~q) | ~t5),
  s0 = \[9] ,
  s1 = ~z | a0,
  s2 = (~\x  & ~s) | ((~v & ~q) | (~u & ~p)),
  s3 = (~t3 & t) | (~t3 & y),
  s4 = m & (p & q),
  s5 = r & (s & t),
  s6 = ~t | i0,
  t1 = (~w1 & ~u1) | ((~w1 & ~d0) | ((~w1 & c0) | ((~u1 & d0) | ((~u1 & ~c0) | ((~d0 & ~c0) | (d0 & c0)))))),
  t2 = (~w2 & (~v2 & ~w1)) | ((~w2 & (~v2 & ~u2)) | ((~w2 & (~v2 & ~c0)) | ((~w2 & (c & ~w1)) | ((~w2 & (c & ~u2)) | ((~w2 & (c & ~c0)) | ((~w2 & (~f0 & ~w1)) | ((~w2 & (~f0 & ~u2)) | (~w2 & (~f0 & ~c0))))))))),
  t3 = (~\x  & ~s) | (~v | ~w),
  t4 = ~r & (s & t),
  t5 = (~u5 & (s & r)) | (~u5 & t),
  t6 = (~u6 & c) | ((~u6 & ~d) | (~u6 & h0)),
  u1 = (~a2 & ~d) | (~z1 & ~c),
  u2 = d0 & (e0 & ~f0),
  u4 = (~c5 & ~d4) | ((~c5 & ~e0) | (~c5 & ~f0)),
  u5 = (~e4 & (~k & q)) | ((~r & ~s) | ~v5),
  u6 = (c & ~i0) | ((c & ~d) | (~i0 & ~d)),
  v2 = (~e3 & (~v & ~q)) | ((~e3 & (~u & ~p)) | ~f3),
  v4 = n & (p & q),
  v5 = (f0 & (e0 & d0)) | ((f0 & (e0 & c0)) | (~g0 & ~f0)),
  v6 = ~i | j,
  w1 = (~x1 & ~d) | (~x1 & ~c),
  w2 = ~y2 & (~d & f0),
  w3 = (~z3 & ~y3) | ((~z3 & h0) | ((~z3 & ~g0) | ((~y3 & ~h0) | (~h0 & ~g0)))),
  w4 = r & (~s & t),
  w5 = s & t,
  w6 = (~k7 & (~j7 & ~i7)) | ((~k7 & (~j7 & c)) | ((~k7 & (~j7 & ~g)) | ((~k7 & (d & ~i7)) | ((~k7 & (d & c)) | ((~k7 & (d & ~g)) | ((~k7 & (~f & ~i7)) | ((~k7 & (~f & c)) | (~k7 & (~f & ~g))))))))),
  x1 = (~y1 & (q & r)) | ((~y1 & (q & w)) | ((~y1 & (v & r)) | (~y1 & (v & w)))),
  x4 = (~y4 & (~d4 & f0)) | ((~y4 & (~d4 & e0)) | ((~y4 & (~f0 & e0)) | (~y4 & (f0 & ~e0)))),
  x5 = ~w5 | (l | ~r),
  y1 = (~\x  & ~s) | ((~y & ~t) | (~u & ~p)),
  y2 = (~a3 & (v & u)) | ((~a3 & (v & p)) | ((~a3 & (q & u)) | ((~a3 & (q & p)) | (~a3 & ~z2)))),
  y3 = (~q4 & (~p4 & ~e4)) | ((~p4 & (~o4 & ~e4)) | ~r4),
  y4 = (~c0 & (~d0 & ~f0)) | (~z4 | t),
  y5 = m | (~s | ~t),
  y6 = (~a7 & ~z6) | ((~a7 & c) | (~z6 & ~c)),
  z1 = (~e2 & (q & t)) | ((~e2 & (q & y)) | ((~e2 & (v & t)) | (~e2 & (v & y)))),
  z2 = ~c0 | (~d0 | ~e0),
  z3 = (~b4 & ~p) | ((~a4 & p) | ~c4),
  z4 = ~b5 & (o & p),
  z5 = (n & ~s) | ((o & ~t) | (~t & ~s)),
  z6 = (~f7 & d) | ((~f7 & ~e) | (~f7 & ~h));
endmodule

