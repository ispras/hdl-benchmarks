//NOTE: no-implementation module stub

module REG16L (
    input wire DSPCLK,
    input wire CLKAY1renb,
    input wire GO_C,
    input wire [15:0] AYin,
    output reg [15:0] AY1r,
    input wire SCAN_TEST
);

endmodule
