module reduce_xor_9s_1(a, b);
  input signed [8:0] a;
  output b;
  assign b = ^a;
endmodule
