//NOTE: no-implementation module stub

module GTECH_MUXI2 (
    input wire A,
    input wire B,
    input wire S,
    output wire Z
);

endmodule
