// IWLS benchmark module "k2" printed on Wed May 29 17:27:51 2002
module k2(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0,
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  m0,
  n0,
  o0,
  p0,
  q0,
  r0,
  s0;
output
  z0,
  z1,
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2,
  g1,
  g2,
  h1,
  h2,
  i1,
  i2,
  j1,
  j2,
  k1,
  k2,
  l1,
  l2,
  m1,
  n1,
  o1,
  p1,
  q1,
  r1,
  s1,
  t0,
  t1,
  u0,
  u1,
  v0,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1;
wire
  \[60] ,
  z5,
  \[61] ,
  \[146] ,
  \[62] ,
  \[147] ,
  \[63] ,
  r11,
  \[148] ,
  \[64] ,
  \[149] ,
  \[65] ,
  \[66] ,
  z10,
  z11,
  \[67] ,
  \[245] ,
  \[68] ,
  \[246] ,
  \[69] ,
  \[247] ,
  \[150] ,
  \[0] ,
  \[151] ,
  \[1] ,
  \[152] ,
  \[2] ,
  \[153] ,
  \[3] ,
  \[154] ,
  \[4] ,
  \[70] ,
  k12,
  \[155] ,
  \[5] ,
  \[156] ,
  \[6] ,
  \[157] ,
  \[7] ,
  \[158] ,
  \[8] ,
  \[252] ,
  \[159] ,
  \[9] ,
  \[75] ,
  \[255] ,
  \[78] ,
  \[256] ,
  \[79] ,
  \[257] ,
  \[259] ,
  \[160] ,
  \[161] ,
  d12,
  \[162] ,
  \[163] ,
  \[164] ,
  \[80] ,
  l11,
  \[165] ,
  \[81] ,
  \[260] ,
  \[167] ,
  \[261] ,
  t11,
  t12,
  \[168] ,
  \[84] ,
  \[262] ,
  \[169] ,
  \[85] ,
  \[263] ,
  \[86] ,
  \[264] ,
  \[87] ,
  \[265] ,
  \[88] ,
  \[266] ,
  \[89] ,
  \[267] ,
  \[268] ,
  \[269] ,
  \[170] ,
  \[10] ,
  e10,
  e11,
  e12,
  \[172] ,
  \[11] ,
  \[173] ,
  \[12] ,
  \[174] ,
  \[13] ,
  m12,
  \[175] ,
  \[14] ,
  \[91] ,
  \[176] ,
  \[15] ,
  \[92] ,
  \[270] ,
  \[177] ,
  \[16] ,
  \[271] ,
  \[178] ,
  \[17] ,
  \[94] ,
  \[272] ,
  \[179] ,
  \[18] ,
  \[95] ,
  \[273] ,
  \[19] ,
  \[96] ,
  \[274] ,
  \[97] ,
  \[275] ,
  \[98] ,
  \[276] ,
  \[100] ,
  \[277] ,
  \[101] ,
  \[278] ,
  \[102] ,
  \[279] ,
  \[103] ,
  \[180] ,
  \[104] ,
  \[181] ,
  \[20] ,
  f10,
  f12,
  \[105] ,
  \[182] ,
  \[21] ,
  \[183] ,
  \[22] ,
  \[200] ,
  \[107] ,
  \[23] ,
  \[201] ,
  n10,
  n11,
  \[108] ,
  \[202] ,
  \[109] ,
  \[25] ,
  \[280] ,
  \[187] ,
  \[26] ,
  \[281] ,
  v12,
  \[188] ,
  \[27] ,
  \[282] ,
  \[189] ,
  \[28] ,
  \[283] ,
  \[29] ,
  \[207] ,
  \[284] ,
  \[208] ,
  \[209] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[30] ,
  g12,
  \[31] ,
  \[116] ,
  \[32] ,
  \[33] ,
  \[211] ,
  \[118] ,
  \[195] ,
  \[34] ,
  \[212] ,
  \[196] ,
  \[35] ,
  \[213] ,
  \[197] ,
  \[36] ,
  \[214] ,
  w11,
  \[198] ,
  \[37] ,
  \[215] ,
  \[199] ,
  \[38] ,
  \[216] ,
  \[39] ,
  \[217] ,
  \[218] ,
  \[219] ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \[40] ,
  h12,
  \[125] ,
  \[41] ,
  \[126] ,
  \[42] ,
  \[220] ,
  \[127] ,
  \[43] ,
  \[221] ,
  p12,
  \[128] ,
  \[222] ,
  \[129] ,
  \[45] ,
  \[223] ,
  \[46] ,
  x11,
  \[47] ,
  \[225] ,
  a7,
  a8,
  \[48] ,
  \[226] ,
  b6,
  b7,
  b8,
  b9,
  \[49] ,
  \[227] ,
  c7,
  \[228] ,
  d5,
  d7,
  d8,
  \[229] ,
  e6,
  e8,
  e9,
  \[130] ,
  f7,
  f8,
  \[131] ,
  a10,
  a11,
  a12,
  g7,
  g8,
  g9,
  \[132] ,
  h8,
  i7,
  i8,
  \[50] ,
  i10,
  j8,
  i12,
  \[51] ,
  k6,
  k8,
  k9,
  \[136] ,
  \[52] ,
  \[230] ,
  l6,
  l8,
  \[137] ,
  \[53] ,
  \[231] ,
  m6,
  m8,
  m9,
  q11,
  q12,
  \[138] ,
  \[54] ,
  \[232] ,
  n7,
  n8,
  n9,
  \[139] ,
  \[55] ,
  o6,
  o7,
  o8,
  \[56] ,
  p6,
  p7,
  p9,
  y10,
  \[57] ,
  \[235] ,
  q7,
  q8,
  \[58] ,
  \[236] ,
  r8,
  \[59] ,
  s6,
  s7,
  s8,
  \[238] ,
  t8,
  t9,
  u7,
  u8,
  u9,
  \[140] ,
  w9,
  \[142] ,
  \[144] ;
assign
  z0 = \[6] ,
  \[60]  = ~e0 & ~d0,
  z1 = \[32] ,
  z5 = \[274]  & (\[221]  & \[69] ),
  \[61]  = \[54]  & \[51] ,
  \[146]  = (\[278]  & \[58] ) | ((\[220]  & \[58] ) | (\[116]  | y10)),
  \[62]  = \[53]  & \[50] ,
  \[147]  = (\[277]  & (\[127]  & ~u)) | ((\[277]  & (\[57]  & ~u)) | ((\[223]  & (\[58]  & z)) | (\[283]  | \[122] ))),
  \[63]  = \[55]  & \[52] ,
  r11 = \[131]  & \[87] ,
  \[148]  = \[53]  & t,
  \[64]  = \[50]  & \[48] ,
  \[149]  = \[89]  & a,
  \[65]  = \[48]  & t,
  \[66]  = \[53]  & ~t,
  z10 = \[223]  & (\[157]  & \[80] ),
  z11 = \[213]  & y,
  \[67]  = \[56]  & c0,
  \[245]  = \[123]  | f10,
  \[68]  = \[59]  & \[49] ,
  \[246]  = \[124]  | \[97] ,
  \[69]  = \[45]  & a,
  \[247]  = \[164]  | \[124] ,
  \[150]  = \[55]  & \[49] ,
  \[0]  = e10 | (m9 | (g9 | \[4] )),
  \[151]  = \[66]  & ~c0,
  \[1]  = l11 | g9,
  \[152]  = \[112]  & ~g0,
  \[2]  = 0,
  \[153]  = \[56]  & \[54] ,
  \[3]  = n9 | m9,
  \[154]  = a0 & l,
  \[4]  = l11 | (n9 | l6),
  \[70]  = c0 & w,
  k12 = \[269]  & a,
  \[155]  = \[61]  & ~l,
  \[5]  = (\[227]  & \[69] ) | ((\[149]  & y) | (f10 | m6)),
  \[156]  = \[59]  & u,
  \[6]  = \[230]  | (\[229]  | (\[195]  | (\[183]  | (q12 | \[8] )))),
  \[157]  = \[103]  & \[69] ,
  \[7]  = \[231]  | (e6 | (p6 | (z10 | b9))),
  \[158]  = \[86]  & e0,
  \[8]  = \[232]  | (\[231]  | (\[207]  | (z5 | (e6 | (k6 | s6))))),
  \[252]  = \[197]  | z11,
  \[159]  = u7 | d8,
  \[9]  = g8 | (d12 | x11),
  \[75]  = (\[181]  & (\[60]  & (a0 & r))) | (\[221]  & (\[60]  & a0)),
  \[255]  = (\[177]  & \[130] ) | (\[200]  | \[43] ),
  \[78]  = (\[156]  & (\[57]  & \[52] )) | ((\[155]  & (\[47]  & z)) | ((\[279]  & ~a0) | ((\[279]  & y) | ((\[278]  & \[47] ) | ((\[227]  & \[47] ) | ((\[220]  & \[47] ) | o6)))))),
  \[256]  = (\[158]  & (w & u)) | ((\[270]  & w) | (\[213]  & a0)),
  \[79]  = ~c0 & ~b0,
  \[257]  = (\[281]  & \[80] ) | ((\[281]  & ~z) | (\[273]  & f)),
  \[259]  = \[207]  | (\[183]  | \[5] ),
  \[160]  = s7 | o7,
  \[161]  = (\[112]  & (g0 & ~f0)) | i7,
  d12 = \[222]  & (\[127]  & \[56] ),
  \[162]  = (\[176]  & i0) | g7,
  \[163]  = (\[179]  & (\[55]  & \[45] )) | (\[265]  & k0),
  \[164]  = \[94]  | i8,
  \[80]  = z & k,
  l11 = \[228]  & (\[227]  & y),
  \[165]  = \[120]  | \[97] ,
  \[81]  = (\[178]  & (~u & b)) | p9,
  \[260]  = \[188]  | (\[187]  | \[160] ),
  \[167]  = \[136]  | t9,
  \[261]  = \[208]  | (\[199]  | (\[198]  | \[189] )),
  t11 = \[272]  & (\[222]  & ~f),
  t12 = \[217]  & (\[52]  & f),
  \[168]  = \[140]  | \[126] ,
  \[84]  = (~q & h) | (q & i),
  \[262]  = (\[226]  & \[111] ) | ((\[131]  & \[111] ) | ((\[111]  & \[67] ) | (\[196]  | l6))),
  \[169]  = \[147]  | \[146] ,
  \[85]  = (\[284]  & \[271] ) | ((\[217]  & \[87] ) | ((\[151]  & \[87] ) | g12)),
  \[263]  = \[110]  & c,
  \[86]  = \[50]  & v,
  \[264]  = \[153]  & ~r,
  \[87]  = \[58]  & ~s,
  \[265]  = \[212]  & ~j0,
  \[88]  = \[57]  & ~j,
  \[266]  = \[218]  & ~o0,
  \[89]  = \[51]  & \[49] ,
  \[267]  = \[49]  & d,
  \[268]  = \[209]  & a,
  \[269]  = \[174]  & \[67] ,
  \[170]  = (\[102]  & m0) | (\[144]  | \[132] ),
  \[10]  = \[202]  | (\[165]  | (\[124]  | (\[123]  | (\[104]  | (i8 | (m8 | e11)))))),
  e10 = \[228]  & \[220] ,
  e11 = \[155]  & (\[58]  & a0),
  e12 = \[180]  & \[45] ,
  \[172]  = \[128]  & ~q0,
  \[11]  = \[201]  | (\[165]  | (\[123]  | o7)),
  \[173]  = \[64]  & b0,
  \[12]  = \[246]  | (\[201]  | (\[167]  | (\[123]  | (p7 | (q7 | (d8 | (f8 | i8))))))),
  \[174]  = \[110]  & ~c,
  \[13]  = \[247]  | (\[200]  | (\[167]  | (\[132]  | (\[125]  | (\[96]  | (\[81]  | (u8 | (r8 | u7)))))))),
  m12 = \[148]  & (\[49]  & w),
  \[175]  = \[64]  & (c0 & ~b0),
  \[14]  = \[247]  | (\[144]  | (\[137]  | (\[122]  | (\[116]  | (\[96]  | (t9 | p9)))))),
  \[91]  = r11 | a11,
  \[176]  = \[152]  & \[129] ,
  \[15]  = \[252]  | (\[246]  | (\[245]  | (\[198]  | (\[162]  | (\[160]  | (\[107]  | (\[81]  | (n7 | (i10 | (m8 | (\[33]  | \[27] ))))))))))),
  \[92]  = (\[276]  & (w & b)) | i12,
  \[270]  = \[182]  & \[66] ,
  \[177]  = \[62]  & \[45] ,
  \[16]  = \[247]  | (\[202]  | (\[197]  | (\[142]  | (\[121]  | (\[109]  | (\[95]  | (q8 | (a12 | (d5 | (e12 | (\[27]  | \[23] ))))))))))),
  \[271]  = \[62]  & \[58] ,
  \[178]  = \[68]  & \[57] ,
  \[17]  = \[260]  | (\[252]  | (\[169]  | (\[167]  | (\[164]  | (\[163]  | (\[140]  | (\[137]  | (\[123]  | (\[120]  | (\[118]  | (\[108]  | (\[78]  | (\[75]  | (g7 | e9)))))))))))))),
  \[94]  = (\[267]  & \[131] ) | (\[174]  & \[131] ),
  \[272]  = \[151]  & ~d,
  \[179]  = c0 & s,
  \[18]  = \[252]  | (\[245]  | (\[199]  | (\[142]  | (\[126]  | (\[120]  | (\[92]  | (\[78]  | (b7 | (i7 | (m12 | h8)))))))))),
  \[95]  = (\[153]  & (\[45]  & (a0 & r))) | (\[284]  & \[177] ),
  \[273]  = \[178]  & u,
  \[19]  = \[245]  | (\[189]  | (\[168]  | (\[165]  | (\[161]  | (\[160]  | (\[121]  | (\[94]  | (d5 | (e8 | (p12 | i12)))))))))),
  \[96]  = \[75]  | h8,
  \[274]  = a0 & ~l,
  \[97]  = \[78]  | \[23] ,
  \[275]  = \[180]  & \[58] ,
  \[98]  = \[85]  | d7,
  \[276]  = \[148]  & \[52] ,
  \[100]  = (\[271]  & z) | ((\[271]  & w) | ((\[221]  & \[101] ) | (\[21]  | \[20] ))),
  \[277]  = \[59]  & \[52] ,
  \[101]  = \[47]  & a0,
  \[278]  = \[61]  & w,
  \[102]  = \[88]  & \[63] ,
  \[279]  = \[52]  & \[51] ,
  \[103]  = ~p & ~f,
  \[180]  = \[79]  & \[64] ,
  \[104]  = (\[154]  & (\[61]  & \[58] )) | (\[283]  & a0),
  \[181]  = \[67]  & s,
  \[20]  = \[264]  & (\[58]  & a0),
  f10 = \[220]  & \[69] ,
  f12 = \[269]  & g,
  \[105]  = (\[226]  & \[52] ) | (\[67]  & \[52] ),
  \[182]  = e0 & s,
  \[21]  = \[181]  & \[101] ,
  \[183]  = (\[157]  & (\[154]  & \[61] )) | (\[154]  & \[149] ),
  \[22]  = \[261]  | (\[260]  | (\[255]  | (\[246]  | (\[202]  | (\[201]  | (\[196]  | (\[167]  | (\[138]  | (\[98]  | (\[94]  | (\[81]  | (f10 | (\[33]  | \[27] ))))))))))))),
  \[200]  = \[168]  | \[142] ,
  \[107]  = \[95]  | m12,
  \[23]  = (\[223]  & \[101] ) | ((\[155]  & \[101] ) | e9),
  \[201]  = \[169]  | \[121] ,
  n10 = \[215]  & (p & ~f),
  n11 = \[269]  & ~g,
  \[108]  = \[100]  | \[91] ,
  \[202]  = \[170]  | \[159] ,
  \[109]  = (\[264]  & (\[45]  & a0)) | ((\[177]  & \[80] ) | (\[177]  & w)),
  \[25]  = \[256]  | (\[255]  | (\[208]  | (n7 | u8))),
  \[280]  = \[216]  & \[60] ,
  \[187]  = (\[214]  & w) | p7,
  \[26]  = (\[217]  & \[49] ) | ((\[213]  & \[127] ) | ((\[151]  & \[49] ) | e12)),
  \[281]  = \[215]  & f,
  v12 = \[222]  & (\[217]  & ~f),
  \[188]  = q8 | n7,
  \[27]  = \[236]  | (\[235]  | (u9 | (t12 | (f12 | (q11 | (g8 | (k12 | x11))))))),
  \[282]  = \[179]  & \[51] ,
  \[189]  = (\[152]  & (h0 & ~f0)) | a12,
  \[28]  = (\[282]  & \[84] ) | (\[261]  | (\[257]  | (\[256]  | (\[187]  | (\[167]  | (\[147]  | (f7 | (k9 | (a7 | (d5 | s7)))))))))),
  \[283]  = \[87]  & \[51] ,
  \[29]  = \[259]  | (\[231]  | (\[230]  | (\[195]  | (z10 | b9)))),
  \[207]  = (\[157]  & (\[155]  & a0)) | ((\[278]  & \[157] ) | ((\[274]  & \[149] ) | ((\[149]  & w) | (k12 | (t11 | \[41] ))))),
  \[284]  = ~c0 & a0,
  \[208]  = (\[157]  & (\[130]  & \[61] )) | ((\[130]  & (\[51]  & ~s)) | ((\[281]  & \[130] ) | ((\[270]  & \[130] ) | ((\[219]  & \[130] ) | ((\[214]  & \[130] ) | b7))))),
  \[209]  = \[62]  & \[47] ,
  \[110]  = \[49]  & ~d,
  \[111]  = \[60]  & ~s,
  \[112]  = \[63]  & \x ,
  \[113]  = \[102]  & ~m0,
  \[30]  = \[238]  | (\[232]  | (e6 | p6)),
  g12 = \[153]  & (\[101]  & r),
  \[31]  = (\[274]  & (\[181]  & \[69] )) | ((\[221]  & (\[154]  & \[69] )) | (\[232]  | (z5 | s6))),
  \[116]  = (\[156]  & (\[87]  & \[57] )) | e11,
  \[32]  = \[280]  & (v & (~n & ~m)),
  \[33]  = \[236]  | (f8 | (i8 | g8)),
  \[211]  = \[150]  & (\[57]  & j),
  \[118]  = (\[182]  & (\[56]  & w)) | p12,
  \[195]  = (g12 & a) | (b6 | v12),
  \[34]  = \[262]  | (\[170]  | (\[146]  | (\[98]  | (\[94]  | (\[75]  | (a8 | (b8 | (l8 | (o7 | (m8 | (o6 | (n8 | (k12 | (x11 | (m6 | (\[31]  | \[3] )))))))))))))))),
  \[212]  = \[176]  & ~i0,
  \[196]  = \[137]  | i10,
  \[35]  = \[259]  | (\[238]  | (\[236]  | (\[229]  | (\[195]  | (\[188]  | (\[165]  | (\[159]  | (\[126]  | (\[107]  | (\[94]  | (\[91]  | (n11 | (h12 | (w11 | (l8 | (z11 | (h8 | (d12 | x11)))))))))))))))))),
  \[213]  = \[56]  & \[49] ,
  \[197]  = \[138]  | u8,
  \[36]  = (\[282]  & ~\[84] ) | (\[262]  | (\[195]  | (\[139]  | (\[121]  | (\[97]  | (n10 | (c7 | (a10 | (w9 | (t8 | (s8 | (q8 | (y10 | (u7 | (a11 | (g8 | (d12 | (t11 | (\[32]  | \[30] ))))))))))))))))))),
  \[214]  = \[158]  & ~u,
  w11 = \[226]  & \[174] ,
  \[198]  = (\[112]  & f0) | \[161] ,
  \[37]  = (\[158]  & a0) | (\[282]  | (\[262]  | (\[261]  | (\[260]  | (\[259]  | (\[257]  | (\[256]  | (\[255]  | (\[238]  | (\[235]  | (\[230]  | (\[229]  | (\[202]  | (\[201]  | (\[164]  | (\[139]  | (\[138]  | (\[136]  | (\[85]  | (n10 | (c7 | (a10 | (w9 | (t8 | (s8 | (n11 | (h12 | (w11 | (a8 | (b8 | (l8 | (f7 | (k9 | (a7 | (o8 | (f12 | (q11 | (r11 | (b6 | (v12 | (\[39]  | \[32] ))))))))))))))))))))))))))))))))))))))))),
  \[215]  = \[61]  & \[45] ,
  \[199]  = \[163]  | \[162] ,
  \[38]  = (\[103]  & (\[49]  & (w & (v & (u & ~a))))) | ((\[65]  & (\[52]  & (w & (~f & ~a)))) | ((\[272]  & (\[52]  & (~f & ~a))) | ((\[228]  & (\[103]  & (\[54]  & \[46] ))) | ((\[177]  & (c0 & (a0 & ~a))) | ((\[173]  & (~d0 & (d & ~a))) | ((\[127]  & (\[68]  & (~u & ~b))) | ((\[127]  & (\[56]  & (\[52]  & ~a))) | ((\[101]  & (\[62]  & (~c0 & ~a))) | ((\[276]  & (\x  & ~b)) | ((\[276]  & (w & ~b)) | ((\[275]  & (~f & ~a)) | ((\[263]  & (\[67]  & ~a)) | ((\[228]  & (\[181]  & \[154] )) | ((\[209]  & (z & ~a)) | ((\[209]  & (w & ~a)) | ((\[178]  & (~u & ~b)) | ((\[153]  & (\[101]  & ~a)) | ((\[131]  & (\[52]  & ~a)) | ((\[89]  & (a0 & ~a)) | ((\[89]  & (z & ~a)) | ((\[89]  & (w & ~a)) | ((\[68]  & (c0 & ~a)) | ((w11 & ~a) | (j8 | (e10 | \[1] ))))))))))))))))))))))))),
  \[216]  = \[79]  & ~o,
  \[39]  = \[165]  | (\[105]  | (\[100]  | (\[92]  | (k8 | (u9 | (t12 | (d7 | a11))))))),
  \[217]  = \[65]  & \[57] ,
  \[218]  = \[172]  & ~n0,
  \[219]  = \[68]  & ~c0,
  \[120]  = \[81]  | f8,
  \[121]  = \[96]  | m8,
  \[122]  = (\[87]  & (\[59]  & c0)) | \[104] ,
  \[123]  = \[105]  | \[98] ,
  \[124]  = \[108]  | \[92] ,
  \[40]  = \[257]  | (\[235]  | (o8 | t12)),
  h12 = \[267]  & (\[67]  & ~g),
  \[125]  = (\[211]  & (\[129]  & n0)) | ((\[87]  & (\[57]  & \[55] )) | (\[172]  & n0)),
  \[41]  = \[273]  & (\[103]  & a),
  \[126]  = (\[148]  & (\[49]  & \x )) | (\[109]  | \[26] ),
  \[42]  = 0,
  \[220]  = \[55]  & \[54] ,
  \[127]  = ~c0 & \x ,
  \[43]  = z11 | d5,
  \[221]  = \[62]  & c0,
  p12 = \[127]  & (\[65]  & \[49] ),
  \[128]  = \[113]  & ~p0,
  \[222]  = \[52]  & a,
  \[129]  = ~h0 & ~f0,
  \[45]  = e0 & ~d0,
  \[223]  = \[61]  & l,
  \[46]  = v & ~t,
  x11 = \[263]  & (\[226]  & a),
  \[47]  = ~e0 & d0,
  a1 = \[7] ,
  a2 = \[33] ,
  \[225]  = \[156]  & (\[111]  & \[70] ),
  a7 = \[225]  & (q & i),
  a8 = \[211]  & (\[129]  & ~n0),
  \[48]  = ~v & u,
  b1 = \[8] ,
  b2 = \[34] ,
  \[226]  = \[66]  & c0,
  b6 = \[101]  & (\[62]  & (~c0 & a)),
  b7 = \[270]  & \[80] ,
  b8 = \[211]  & f0,
  b9 = \[149]  & (\[80]  & l),
  \[49]  = \[45]  & ~s,
  c1 = \[9] ,
  c2 = \[35] ,
  \[227]  = \[86]  & u,
  c7 = \[225]  & (~q & ~h),
  d1 = \[10] ,
  d2 = \[36] ,
  \[228]  = \[45]  & ~a,
  d5 = \[213]  & w,
  d7 = \[87]  & (\[56]  & ~c0),
  d8 = \[150]  & \[88] ,
  e1 = \[11] ,
  e2 = \[37] ,
  \[229]  = \[31]  | \[7] ,
  e6 = p6 & ~l,
  e8 = \[173]  & (\[47]  & ~c0),
  e9 = \[279]  & a0,
  \[130]  = z & ~k,
  f1 = \[12] ,
  f2 = \[38] ,
  f7 = \[265]  & (~l0 & ~k0),
  f8 = \[173]  & \[45] ,
  \[131]  = \[70]  & \[65] ,
  g1 = \[13] ,
  g2 = \[39] ,
  a10 = \[225]  & (q & ~i),
  a11 = \[223]  & (\[47]  & z),
  a12 = \[56]  & (\[52]  & y),
  g7 = \[265]  & (l0 & ~k0),
  g8 = \[173]  & (\[60]  & (d & a)),
  g9 = \[89]  & (y & ~a),
  \[132]  = (\[128]  & (q0 & ~n0)) | q7,
  h1 = \[14] ,
  h2 = \[40] ,
  h8 = \[173]  & (\[60]  & ~d),
  i1 = \[15] ,
  i2 = \[41] ,
  i7 = \[212]  & j0,
  i8 = \[175]  & \[58] ,
  \[50]  = t & s,
  j1 = \[16] ,
  j2 = \[42] ,
  i10 = \[179]  & (\[60]  & \[55] ),
  j8 = \[175]  & (\[47]  & (~e & ~a)),
  i12 = \[276]  & (\x  & b),
  \[51]  = \[46]  & u,
  k1 = \[17] ,
  k2 = \[43] ,
  k6 = \[268]  & w,
  k8 = \[175]  & (\[47]  & e),
  k9 = \[225]  & (~q & h),
  \[136]  = (\[227]  & \[58] ) | (\[214]  & \[80] ),
  \[52]  = \[47]  & ~s,
  l1 = \[18] ,
  l2 = d5,
  \[230]  = n8 | \[9] ,
  l6 = \[219]  & y,
  l8 = \[175]  & \[45] ,
  \[137]  = (\[218]  & o0) | (\[211]  & h0),
  \[53]  = ~v & ~u,
  m1 = \[19] ,
  \[231]  = (\[157]  & (\[155]  & \[80] )) | (\[149]  & (\[80]  & ~l)),
  m6 = \[68]  & (c0 & a),
  m8 = \[175]  & \[60] ,
  m9 = \[219]  & \[80] ,
  q11 = \[267]  & (\[67]  & g),
  q12 = \[264]  & (\[101]  & a),
  \[138]  = e8 | r8,
  \[54]  = ~c0 & s,
  n1 = \[20] ,
  \[232]  = (\[222]  & \[131] ) | j8,
  n7 = \[150]  & \x ,
  n8 = \[275]  & (~f & a),
  n9 = \[219]  & a0,
  \[139]  = (\[280]  & (~v & n)) | \[3] ,
  \[55]  = \[46]  & ~u,
  o1 = \[21] ,
  o6 = \[277]  & c0,
  o7 = \[266]  & (~s0 & r0),
  o8 = \[275]  & f,
  \[56]  = \[48]  & ~t,
  p1 = \[22] ,
  p6 = \[268]  & \[80] ,
  p7 = \[266]  & (~s0 & ~r0),
  p9 = \[127]  & (\[68]  & (~u & b)),
  y10 = \[155]  & (\[58]  & z),
  \[57]  = ~c0 & w,
  q1 = \[23] ,
  \[235]  = (\[272]  & (\[52]  & f)) | (\[151]  & (\[52]  & d)),
  q7 = \[266]  & (s0 & ~r0),
  q8 = \[180]  & \[47] ,
  \[58]  = e0 & d0,
  r1 = d5,
  \[236]  = k8 | o8,
  r8 = \[79]  & (\[60]  & o),
  \[59]  = v & t,
  s1 = \[25] ,
  s6 = \[181]  & (\[154]  & \[69] ),
  s7 = \[70]  & (\[55]  & (e0 & ~s)),
  s8 = \[216]  & (\[111]  & (\[56]  & ~\x )),
  t0 = \[0] ,
  t1 = \[26] ,
  \[238]  = k6 | q12,
  t8 = \[66]  & (\[60]  & (\[54]  & (~b0 & ~o))),
  t9 = \[214]  & a0,
  u0 = \[1] ,
  u1 = \[27] ,
  u7 = \[128]  & (q0 & n0),
  u8 = \[280]  & (v & n),
  u9 = \[263]  & \[131] ,
  \[140]  = (\[182]  & (\[56]  & \x )) | \[107] ,
  v0 = \[2] ,
  v1 = \[28] ,
  w0 = \[3] ,
  w1 = \[29] ,
  w9 = \[273]  & (p & ~f),
  \[142]  = (\[284]  & (\[65]  & \[49] )) | \[118] ,
  x0 = \[4] ,
  x1 = \[30] ,
  y0 = \[5] ,
  y1 = \[31] ,
  \[144]  = (\[113]  & p0) | \[125] ;
endmodule

