module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 ;
output g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( n246 , g245 );
buf ( n247 , g246 );
buf ( n248 , g247 );
buf ( n249 , g248 );
buf ( n250 , g249 );
buf ( n251 , g250 );
buf ( n252 , g251 );
buf ( n253 , g252 );
buf ( n254 , g253 );
buf ( n255 , g254 );
buf ( n256 , g255 );
buf ( n257 , g256 );
buf ( n258 , g257 );
buf ( n259 , g258 );
buf ( n260 , g259 );
buf ( n261 , g260 );
buf ( n262 , g261 );
buf ( n263 , g262 );
buf ( n264 , g263 );
buf ( n265 , g264 );
buf ( n266 , g265 );
buf ( n267 , g266 );
buf ( n268 , g267 );
buf ( n269 , g268 );
buf ( n270 , g269 );
buf ( n271 , g270 );
buf ( n272 , g271 );
buf ( n273 , g272 );
buf ( n274 , g273 );
buf ( n275 , g274 );
buf ( n276 , g275 );
buf ( n277 , g276 );
buf ( n278 , g277 );
buf ( n279 , g278 );
buf ( n280 , g279 );
buf ( n281 , g280 );
buf ( n282 , g281 );
buf ( n283 , g282 );
buf ( n284 , g283 );
buf ( n285 , g284 );
buf ( n286 , g285 );
buf ( n287 , g286 );
buf ( n288 , g287 );
buf ( n289 , g288 );
buf ( n290 , g289 );
buf ( n291 , g290 );
buf ( n292 , g291 );
buf ( n293 , g292 );
buf ( n294 , g293 );
buf ( n295 , g294 );
buf ( n296 , g295 );
buf ( n297 , g296 );
buf ( n298 , g297 );
buf ( n299 , g298 );
buf ( n300 , g299 );
buf ( n301 , g300 );
buf ( n302 , g301 );
buf ( n303 , g302 );
buf ( n304 , g303 );
buf ( n305 , g304 );
buf ( n306 , g305 );
buf ( n307 , g306 );
buf ( n308 , g307 );
buf ( n309 , g308 );
buf ( n310 , g309 );
buf ( n311 , g310 );
buf ( n312 , g311 );
buf ( n313 , g312 );
buf ( n314 , g313 );
buf ( n315 , g314 );
buf ( n316 , g315 );
buf ( n317 , g316 );
buf ( n318 , g317 );
buf ( n319 , g318 );
buf ( n320 , g319 );
buf ( n321 , g320 );
buf ( n322 , g321 );
buf ( n323 , g322 );
buf ( n324 , g323 );
buf ( n325 , g324 );
buf ( n326 , g325 );
buf ( n327 , g326 );
buf ( n328 , g327 );
buf ( n329 , g328 );
buf ( n330 , g329 );
buf ( n331 , g330 );
buf ( n332 , g331 );
buf ( n333 , g332 );
buf ( n334 , g333 );
buf ( n335 , g334 );
buf ( n336 , g335 );
buf ( n337 , g336 );
buf ( n338 , g337 );
buf ( n339 , g338 );
buf ( n340 , g339 );
buf ( n341 , g340 );
buf ( n342 , g341 );
buf ( n343 , g342 );
buf ( n344 , g343 );
buf ( n345 , g344 );
buf ( n346 , g345 );
buf ( n347 , g346 );
buf ( n348 , g347 );
buf ( n349 , g348 );
buf ( n350 , g349 );
buf ( n351 , g350 );
buf ( n352 , g351 );
buf ( n353 , g352 );
buf ( n354 , g353 );
buf ( n355 , g354 );
buf ( n356 , g355 );
buf ( n357 , g356 );
buf ( n358 , g357 );
buf ( n359 , g358 );
buf ( n360 , g359 );
buf ( n361 , g360 );
buf ( n362 , g361 );
buf ( n363 , g362 );
buf ( n364 , g363 );
buf ( n365 , g364 );
buf ( n366 , g365 );
buf ( n367 , g366 );
buf ( n368 , g367 );
buf ( n369 , g368 );
buf ( n370 , g369 );
buf ( n371 , g370 );
buf ( n372 , g371 );
buf ( n373 , g372 );
buf ( n374 , g373 );
buf ( n375 , g374 );
buf ( n376 , g375 );
buf ( n377 , g376 );
buf ( n378 , g377 );
buf ( n379 , g378 );
buf ( n380 , g379 );
buf ( n381 , g380 );
buf ( n382 , g381 );
buf ( n383 , g382 );
buf ( n384 , g383 );
buf ( n385 , g384 );
buf ( n386 , g385 );
buf ( n387 , g386 );
buf ( n388 , g387 );
buf ( n389 , g388 );
buf ( n390 , g389 );
buf ( n391 , g390 );
buf ( n392 , g391 );
buf ( n393 , g392 );
buf ( n394 , g393 );
buf ( n395 , g394 );
buf ( n396 , g395 );
buf ( n397 , g396 );
buf ( n398 , g397 );
buf ( n399 , g398 );
buf ( n400 , g399 );
buf ( n401 , g400 );
buf ( n402 , g401 );
buf ( n403 , g402 );
buf ( n404 , g403 );
buf ( n405 , g404 );
buf ( n406 , g405 );
buf ( n407 , g406 );
buf ( n408 , g407 );
buf ( n409 , g408 );
buf ( n410 , g409 );
buf ( n411 , g410 );
buf ( g411 , n412 );
buf ( g412 , n413 );
buf ( g413 , n414 );
buf ( g414 , n415 );
buf ( g415 , n416 );
buf ( g416 , n417 );
buf ( g417 , n418 );
buf ( g418 , n419 );
buf ( g419 , n420 );
buf ( g420 , n421 );
buf ( g421 , n422 );
buf ( g422 , n423 );
buf ( g423 , n424 );
buf ( g424 , n425 );
buf ( g425 , n426 );
buf ( g426 , n427 );
buf ( g427 , n428 );
buf ( g428 , n429 );
buf ( g429 , n430 );
buf ( g430 , n431 );
buf ( g431 , n432 );
buf ( g432 , n433 );
buf ( g433 , n434 );
buf ( g434 , n435 );
buf ( g435 , n436 );
buf ( g436 , n437 );
buf ( g437 , n438 );
buf ( g438 , n439 );
buf ( g439 , n440 );
buf ( g440 , n441 );
buf ( g441 , n442 );
buf ( g442 , n443 );
buf ( g443 , n444 );
buf ( g444 , n445 );
buf ( g445 , n446 );
buf ( g446 , n447 );
buf ( g447 , n448 );
buf ( g448 , n449 );
buf ( g449 , n450 );
buf ( g450 , n451 );
buf ( g451 , n452 );
buf ( g452 , n453 );
buf ( g453 , n454 );
buf ( g454 , n455 );
buf ( g455 , n456 );
buf ( g456 , n457 );
buf ( g457 , n458 );
buf ( g458 , n459 );
buf ( g459 , n460 );
buf ( g460 , n461 );
buf ( g461 , n462 );
buf ( g462 , n463 );
buf ( g463 , n464 );
buf ( g464 , n465 );
buf ( g465 , n466 );
buf ( g466 , n467 );
buf ( g467 , n468 );
buf ( g468 , n469 );
buf ( g469 , n470 );
buf ( g470 , n471 );
buf ( g471 , n472 );
buf ( g472 , n473 );
buf ( g473 , n474 );
buf ( g474 , n475 );
buf ( g475 , n476 );
buf ( g476 , n477 );
buf ( g477 , n478 );
buf ( g478 , n479 );
buf ( g479 , n480 );
buf ( g480 , n481 );
buf ( g481 , n482 );
buf ( g482 , n483 );
buf ( g483 , n484 );
buf ( g484 , n485 );
buf ( g485 , n486 );
buf ( g486 , n487 );
buf ( g487 , n488 );
buf ( g488 , n489 );
buf ( g489 , n490 );
buf ( g490 , n491 );
buf ( g491 , n492 );
buf ( g492 , n493 );
buf ( g493 , n494 );
buf ( g494 , n495 );
buf ( g495 , n496 );
buf ( g496 , n497 );
buf ( g497 , n498 );
buf ( g498 , n499 );
buf ( g499 , n500 );
buf ( g500 , n501 );
buf ( g501 , n502 );
buf ( g502 , n503 );
buf ( g503 , n504 );
buf ( g504 , n505 );
buf ( g505 , n506 );
buf ( g506 , n507 );
buf ( g507 , n508 );
buf ( g508 , n509 );
buf ( g509 , n510 );
buf ( g510 , n511 );
buf ( g511 , n512 );
buf ( g512 , n513 );
buf ( g513 , n514 );
buf ( g514 , n515 );
buf ( g515 , n516 );
buf ( g516 , n517 );
buf ( g517 , n518 );
buf ( g518 , n519 );
buf ( g519 , n520 );
buf ( g520 , n521 );
buf ( g521 , n522 );
buf ( g522 , n523 );
buf ( g523 , n524 );
buf ( g524 , n525 );
buf ( g525 , n526 );
buf ( g526 , n527 );
buf ( g527 , n528 );
buf ( g528 , n529 );
buf ( g529 , n530 );
buf ( g530 , n531 );
buf ( g531 , n532 );
buf ( g532 , n533 );
buf ( g533 , n534 );
buf ( g534 , n535 );
buf ( g535 , n536 );
buf ( g536 , n537 );
buf ( g537 , n538 );
buf ( g538 , n539 );
buf ( n412 , n1405 );
buf ( n413 , n1457 );
buf ( n414 , n818 );
buf ( n415 , n788 );
buf ( n416 , n756 );
buf ( n417 , n1005 );
buf ( n418 , n848 );
buf ( n419 , n1487 );
buf ( n420 , n662 );
buf ( n421 , n706 );
buf ( n422 , n939 );
buf ( n423 , n1677 );
buf ( n424 , n1680 );
buf ( n425 , n1049 );
buf ( n426 , n1075 );
buf ( n427 , n913 );
buf ( n428 , n1108 );
buf ( n429 , n1137 );
buf ( n430 , n1214 );
buf ( n431 , n1162 );
buf ( n432 , n1378 );
buf ( n433 , n886 );
buf ( n434 , n965 );
buf ( n435 , n1250 );
buf ( n436 , n1431 );
buf ( n437 , n1279 );
buf ( n438 , n1345 );
buf ( n439 , n1312 );
buf ( n440 , n1683 );
buf ( n441 , n1686 );
buf ( n442 , n1691 );
buf ( n443 , n1650 );
buf ( n444 , n1657 );
buf ( n445 , n1707 );
buf ( n446 , n1664 );
buf ( n447 , n1549 );
buf ( n448 , n1697 );
buf ( n449 , n1701 );
buf ( n450 , n1185 );
buf ( n451 , n1627 );
buf ( n452 , n1803 );
buf ( n453 , n1554 );
buf ( n454 , n1634 );
buf ( n455 , n1621 );
buf ( n456 , n1801 );
buf ( n457 , n1706 );
buf ( n458 , n1787 );
buf ( n459 , n16 );
buf ( n460 , n16 );
buf ( n461 , n16 );
buf ( n462 , n16 );
buf ( n463 , n16 );
buf ( n464 , n16 );
buf ( n465 , n16 );
buf ( n466 , n16 );
buf ( n467 , n16 );
buf ( n468 , n16 );
buf ( n469 , n16 );
buf ( n470 , n16 );
buf ( n471 , n16 );
buf ( n472 , n16 );
buf ( n473 , n16 );
buf ( n474 , n16 );
buf ( n475 , n16 );
buf ( n476 , n16 );
buf ( n477 , n16 );
buf ( n478 , n16 );
buf ( n479 , n16 );
buf ( n480 , n16 );
buf ( n481 , n16 );
buf ( n482 , n16 );
buf ( n483 , n16 );
buf ( n484 , n16 );
buf ( n485 , n16 );
buf ( n486 , n16 );
buf ( n487 , n16 );
buf ( n488 , n16 );
buf ( n489 , n1734 );
buf ( n490 , n16 );
buf ( n491 , n16 );
buf ( n492 , n1732 );
buf ( n493 , n16 );
buf ( n494 , n16 );
buf ( n495 , n16 );
buf ( n496 , n16 );
buf ( n497 , n16 );
buf ( n498 , n16 );
buf ( n499 , n16 );
buf ( n500 , n16 );
buf ( n501 , n1792 );
buf ( n502 , n1793 );
buf ( n503 , n1790 );
buf ( n504 , n16 );
buf ( n505 , n1789 );
buf ( n506 , n16 );
buf ( n507 , n1785 );
buf ( n508 , n16 );
buf ( n509 , n1784 );
buf ( n510 , n16 );
buf ( n511 , n16 );
buf ( n512 , n16 );
buf ( n513 , n16 );
buf ( n514 , n1791 );
buf ( n515 , n16 );
buf ( n516 , n16 );
buf ( n517 , n16 );
buf ( n518 , n16 );
buf ( n519 , n16 );
buf ( n520 , n1743 );
buf ( n521 , n16 );
buf ( n522 , n16 );
buf ( n523 , n1755 );
buf ( n524 , n1759 );
buf ( n525 , n1716 );
buf ( n526 , n1720 );
buf ( n527 , n1712 );
buf ( n528 , n1747 );
buf ( n529 , n1728 );
buf ( n530 , n1763 );
buf ( n531 , n1751 );
buf ( n532 , n1767 );
buf ( n533 , n1738 );
buf ( n534 , n1724 );
buf ( n535 , n1771 );
buf ( n536 , n1775 );
buf ( n537 , n1779 );
buf ( n538 , n1742 );
buf ( n539 , n1783 );
not ( n542 , n119 );
not ( n543 , n2 );
not ( n544 , n3 );
and ( n545 , n543 , n544 );
and ( n546 , n2 , n3 );
nor ( n547 , n545 , n546 );
nor ( n548 , n4 , n5 );
not ( n549 , n6 );
nand ( n550 , n548 , n549 );
nor ( n551 , n547 , n550 );
not ( n552 , n16 );
and ( n553 , n551 , n552 );
not ( n554 , n553 );
or ( n555 , n542 , n554 );
xor ( n556 , n2 , n3 );
not ( n557 , n556 );
not ( n558 , n5 );
nor ( n559 , n558 , n6 , n4 );
and ( n560 , n557 , n559 );
nand ( n561 , n560 , n120 );
nand ( n562 , n555 , n561 );
not ( n563 , n117 );
not ( n564 , n3 );
nand ( n565 , n564 , n2 );
not ( n566 , n5 );
nor ( n567 , n566 , n4 );
not ( n568 , n2 );
nand ( n569 , n568 , n3 );
nand ( n570 , n565 , n567 , n569 , n6 );
not ( n571 , n570 );
not ( n572 , n571 );
or ( n573 , n563 , n572 );
not ( n574 , n6 );
nand ( n575 , n574 , n4 , n5 );
nor ( n576 , n575 , n556 );
buf ( n577 , n576 );
nand ( n578 , n577 , n115 );
nand ( n579 , n573 , n578 );
nor ( n580 , n562 , n579 );
not ( n581 , n580 );
not ( n582 , n118 );
nand ( n583 , n548 , n6 );
not ( n584 , n583 );
not ( n585 , n547 );
nand ( n586 , n584 , n585 );
buf ( n587 , n586 );
not ( n588 , n587 );
not ( n589 , n588 );
or ( n590 , n582 , n589 );
not ( n591 , n13 );
not ( n592 , n11 );
not ( n593 , n12 );
nand ( n594 , n591 , n592 , n593 );
buf ( n595 , n594 );
not ( n596 , n595 );
not ( n597 , n596 );
nand ( n598 , n590 , n597 );
nor ( n599 , n581 , n598 );
not ( n600 , n125 );
not ( n601 , n25 );
nor ( n602 , n601 , n26 );
nor ( n603 , n23 , n24 );
and ( n604 , n602 , n603 , n552 );
buf ( n605 , n604 );
not ( n606 , n605 );
or ( n607 , n600 , n606 );
nor ( n608 , n25 , n26 );
nor ( n609 , n24 , n16 );
and ( n610 , n608 , n609 , n23 );
buf ( n611 , n610 );
nand ( n612 , n611 , n127 );
nand ( n613 , n607 , n612 );
not ( n614 , n124 );
not ( n615 , n608 );
not ( n616 , n24 );
nor ( n617 , n616 , n23 );
not ( n618 , n617 );
or ( n619 , n615 , n618 );
not ( n620 , n16 );
nand ( n621 , n619 , n620 );
buf ( n622 , n621 );
not ( n623 , n622 );
or ( n624 , n614 , n623 );
not ( n625 , n16 );
not ( n626 , n20 );
not ( n627 , n21 );
nand ( n628 , n626 , n627 );
nand ( n629 , n625 , n628 );
buf ( n630 , n629 );
nand ( n631 , n624 , n630 );
not ( n632 , n26 );
nor ( n633 , n632 , n25 );
nand ( n634 , n633 , n603 , n620 );
not ( n635 , n634 );
and ( n636 , n635 , n126 );
or ( n637 , n613 , n631 , n636 );
nor ( n638 , n15 , n17 );
and ( n639 , n638 , n123 );
not ( n640 , n15 );
nor ( n641 , n640 , n17 );
and ( n642 , n641 , n121 );
and ( n643 , n17 , n122 );
nor ( n644 , n639 , n642 , n643 );
not ( n645 , n628 );
nor ( n646 , n645 , n16 );
nand ( n647 , n644 , n646 );
nand ( n648 , n637 , n647 );
or ( n649 , n599 , n648 );
nand ( n650 , n6 , n4 , n5 );
nor ( n651 , n547 , n650 );
not ( n652 , n651 );
nand ( n653 , n652 , n595 );
nand ( n654 , n653 , n116 );
not ( n655 , n654 );
not ( n656 , n580 );
or ( n657 , n655 , n656 );
nand ( n658 , n657 , n597 );
not ( n659 , n595 );
nor ( n660 , n587 , n659 );
nand ( n661 , n118 , n660 );
nand ( n662 , n649 , n658 , n661 );
not ( n663 , n130 );
not ( n664 , n553 );
or ( n665 , n663 , n664 );
nand ( n666 , n560 , n129 );
nand ( n667 , n665 , n666 );
not ( n668 , n131 );
not ( n669 , n571 );
or ( n670 , n668 , n669 );
not ( n671 , n576 );
not ( n672 , n671 );
nand ( n673 , n672 , n132 );
nand ( n674 , n670 , n673 );
nor ( n675 , n667 , n674 );
not ( n676 , n675 );
not ( n677 , n128 );
nor ( n678 , n677 , n587 );
not ( n679 , n678 );
buf ( n680 , n595 );
buf ( n681 , n680 );
nand ( n682 , n679 , n681 );
nor ( n683 , n676 , n682 );
nand ( n684 , n605 , n139 );
nand ( n685 , n622 , n136 );
nand ( n686 , n684 , n685 , n630 );
not ( n687 , n137 );
not ( n688 , n635 );
or ( n689 , n687 , n688 );
nand ( n690 , n611 , n138 );
nand ( n691 , n689 , n690 );
or ( n692 , n686 , n691 );
and ( n693 , n638 , n60 );
and ( n694 , n641 , n135 );
and ( n695 , n17 , n134 );
nor ( n696 , n693 , n694 , n695 );
nand ( n697 , n696 , n646 );
nand ( n698 , n692 , n697 );
or ( n699 , n683 , n698 );
not ( n700 , n675 );
and ( n701 , n653 , n133 );
nor ( n702 , n701 , n678 );
not ( n703 , n702 );
or ( n704 , n700 , n703 );
nand ( n705 , n704 , n680 );
nand ( n706 , n699 , n705 );
not ( n707 , n13 );
nor ( n708 , n11 , n12 );
nand ( n709 , n707 , n708 );
not ( n710 , n709 );
and ( n711 , n710 , n641 );
and ( n712 , n711 , n72 );
nand ( n713 , n710 , n17 );
not ( n714 , n713 );
and ( n715 , n714 , n73 );
nor ( n716 , n712 , n715 );
not ( n717 , n716 );
not ( n718 , n74 );
not ( n719 , n595 );
nand ( n720 , n719 , n638 );
nor ( n721 , n718 , n720 );
nand ( n722 , n629 , n710 );
not ( n723 , n722 );
nor ( n724 , n721 , n723 );
not ( n725 , n724 );
or ( n726 , n717 , n725 );
not ( n727 , n75 );
nand ( n728 , n727 , n630 );
not ( n729 , n728 );
not ( n730 , n622 );
nand ( n731 , n730 , n630 );
not ( n732 , n731 );
or ( n733 , n729 , n732 );
and ( n734 , n605 , n78 );
and ( n735 , n635 , n77 );
not ( n736 , n76 );
not ( n737 , n611 );
nor ( n738 , n736 , n737 );
nor ( n739 , n734 , n735 , n738 );
nand ( n740 , n733 , n739 );
nand ( n741 , n726 , n740 );
not ( n742 , n587 );
nand ( n743 , n742 , n70 );
buf ( n744 , n571 );
nand ( n745 , n744 , n69 );
buf ( n746 , n672 );
nand ( n747 , n746 , n67 );
nand ( n748 , n743 , n745 , n747 );
nand ( n749 , n748 , n597 );
and ( n750 , n560 , n595 );
and ( n751 , n750 , n71 );
and ( n752 , n651 , n709 );
buf ( n753 , n752 );
and ( n754 , n753 , n68 );
nor ( n755 , n751 , n754 );
nand ( n756 , n741 , n749 , n755 );
and ( n757 , n711 , n60 );
and ( n758 , n714 , n61 );
nor ( n759 , n757 , n758 );
not ( n760 , n759 );
not ( n761 , n62 );
nor ( n762 , n761 , n720 );
nor ( n763 , n762 , n723 );
not ( n764 , n763 );
or ( n765 , n760 , n764 );
not ( n766 , n63 );
nand ( n767 , n766 , n630 );
not ( n768 , n767 );
not ( n769 , n731 );
or ( n770 , n768 , n769 );
and ( n771 , n605 , n66 );
and ( n772 , n635 , n64 );
not ( n773 , n65 );
not ( n774 , n611 );
nor ( n775 , n773 , n774 );
nor ( n776 , n771 , n772 , n775 );
nand ( n777 , n770 , n776 );
nand ( n778 , n765 , n777 );
not ( n779 , n587 );
nand ( n780 , n779 , n58 );
nand ( n781 , n744 , n57 );
nand ( n782 , n746 , n55 );
nand ( n783 , n780 , n781 , n782 );
nand ( n784 , n783 , n597 );
and ( n785 , n750 , n59 );
and ( n786 , n753 , n56 );
nor ( n787 , n785 , n786 );
nand ( n788 , n778 , n784 , n787 );
and ( n789 , n711 , n48 );
and ( n790 , n714 , n49 );
nor ( n791 , n789 , n790 );
not ( n792 , n791 );
not ( n793 , n50 );
nor ( n794 , n793 , n720 );
nor ( n795 , n794 , n723 );
not ( n796 , n795 );
or ( n797 , n792 , n796 );
not ( n798 , n51 );
nand ( n799 , n798 , n630 );
not ( n800 , n799 );
not ( n801 , n731 );
or ( n802 , n800 , n801 );
and ( n803 , n605 , n52 );
and ( n804 , n635 , n53 );
not ( n805 , n54 );
nor ( n806 , n774 , n805 );
nor ( n807 , n803 , n804 , n806 );
nand ( n808 , n802 , n807 );
nand ( n809 , n797 , n808 );
nand ( n810 , n779 , n46 );
nand ( n811 , n744 , n45 );
nand ( n812 , n746 , n43 );
nand ( n813 , n810 , n811 , n812 );
nand ( n814 , n813 , n597 );
and ( n815 , n750 , n47 );
and ( n816 , n753 , n44 );
nor ( n817 , n815 , n816 );
nand ( n818 , n809 , n814 , n817 );
and ( n819 , n711 , n96 );
and ( n820 , n714 , n97 );
nor ( n821 , n819 , n820 );
not ( n822 , n821 );
not ( n823 , n98 );
nor ( n824 , n823 , n720 );
nor ( n825 , n824 , n723 );
not ( n826 , n825 );
or ( n827 , n822 , n826 );
not ( n828 , n99 );
nand ( n829 , n828 , n630 );
not ( n830 , n829 );
not ( n831 , n731 );
or ( n832 , n830 , n831 );
and ( n833 , n605 , n102 );
and ( n834 , n635 , n100 );
not ( n835 , n101 );
nor ( n836 , n774 , n835 );
nor ( n837 , n833 , n834 , n836 );
nand ( n838 , n832 , n837 );
nand ( n839 , n827 , n838 );
nand ( n840 , n588 , n94 );
nand ( n841 , n744 , n93 );
nand ( n842 , n746 , n91 );
nand ( n843 , n840 , n841 , n842 );
nand ( n844 , n843 , n597 );
and ( n845 , n750 , n95 );
and ( n846 , n753 , n92 );
nor ( n847 , n845 , n846 );
nand ( n848 , n839 , n844 , n847 );
nand ( n849 , n742 , n259 );
buf ( n850 , n560 );
nand ( n851 , n850 , n260 );
buf ( n852 , n651 );
nand ( n853 , n852 , n257 );
nand ( n854 , n849 , n851 , n853 );
nand ( n855 , n744 , n258 );
nand ( n856 , n746 , n256 );
not ( n857 , n659 );
nand ( n858 , n855 , n856 , n857 );
or ( n859 , n854 , n858 );
not ( n860 , n16 );
nand ( n861 , n860 , n628 );
not ( n862 , n861 );
nand ( n863 , n862 , n719 , n17 );
or ( n864 , n863 , n261 );
nand ( n865 , n859 , n864 );
not ( n866 , n262 );
not ( n867 , n866 );
not ( n868 , n861 );
not ( n869 , n17 );
nand ( n870 , n868 , n710 , n869 );
not ( n871 , n870 );
not ( n872 , n871 );
or ( n873 , n867 , n872 );
not ( n874 , n730 );
not ( n875 , n263 );
not ( n876 , n875 );
and ( n877 , n874 , n876 );
not ( n878 , n611 );
not ( n879 , n265 );
nor ( n880 , n878 , n879 );
nor ( n881 , n877 , n880 );
nand ( n882 , n605 , n266 );
nand ( n883 , n635 , n264 );
nand ( n884 , n881 , n723 , n882 , n883 );
nand ( n885 , n873 , n884 );
nor ( n886 , n865 , n885 );
nand ( n887 , n742 , n186 );
nand ( n888 , n850 , n187 );
nand ( n889 , n852 , n184 );
nand ( n890 , n887 , n888 , n889 );
nand ( n891 , n744 , n185 );
nand ( n892 , n746 , n183 );
buf ( n893 , n595 );
nand ( n894 , n891 , n892 , n893 );
or ( n895 , n890 , n894 );
or ( n896 , n863 , n188 );
nand ( n897 , n895 , n896 );
not ( n898 , n189 );
not ( n899 , n898 );
not ( n900 , n871 );
or ( n901 , n899 , n900 );
not ( n902 , n730 );
not ( n903 , n190 );
not ( n904 , n903 );
and ( n905 , n902 , n904 );
not ( n906 , n192 );
nor ( n907 , n906 , n878 );
nor ( n908 , n905 , n907 );
nand ( n909 , n605 , n193 );
nand ( n910 , n635 , n191 );
nand ( n911 , n908 , n723 , n909 , n910 );
nand ( n912 , n901 , n911 );
nor ( n913 , n897 , n912 );
nand ( n914 , n742 , n143 );
nand ( n915 , n850 , n144 );
nand ( n916 , n141 , n852 );
nand ( n917 , n914 , n915 , n916 );
nand ( n918 , n744 , n142 );
nand ( n919 , n746 , n140 );
nand ( n920 , n918 , n919 , n857 );
or ( n921 , n917 , n920 );
or ( n922 , n863 , n38 );
nand ( n923 , n921 , n922 );
not ( n924 , n145 );
not ( n925 , n924 );
not ( n926 , n871 );
or ( n927 , n925 , n926 );
not ( n928 , n730 );
not ( n929 , n146 );
not ( n930 , n929 );
and ( n931 , n928 , n930 );
not ( n932 , n148 );
nor ( n933 , n932 , n878 );
nor ( n934 , n931 , n933 );
nand ( n935 , n605 , n149 );
nand ( n936 , n147 , n635 );
nand ( n937 , n934 , n723 , n935 , n936 );
nand ( n938 , n927 , n937 );
nor ( n939 , n923 , n938 );
nand ( n940 , n742 , n270 );
nand ( n941 , n850 , n271 );
nand ( n942 , n852 , n268 );
nand ( n943 , n940 , n941 , n942 );
nand ( n944 , n744 , n269 );
nand ( n945 , n746 , n267 );
nand ( n946 , n944 , n945 , n857 );
or ( n947 , n943 , n946 );
or ( n948 , n863 , n272 );
nand ( n949 , n947 , n948 );
not ( n950 , n273 );
not ( n951 , n950 );
not ( n952 , n871 );
or ( n953 , n951 , n952 );
not ( n954 , n730 );
not ( n955 , n274 );
not ( n956 , n955 );
and ( n957 , n954 , n956 );
not ( n958 , n276 );
nor ( n959 , n958 , n737 );
nor ( n960 , n957 , n959 );
nand ( n961 , n605 , n277 );
nand ( n962 , n635 , n275 );
nand ( n963 , n960 , n723 , n961 , n962 );
nand ( n964 , n953 , n963 );
nor ( n965 , n949 , n964 );
not ( n966 , n720 );
and ( n967 , n966 , n86 );
and ( n968 , n711 , n84 );
nor ( n969 , n967 , n968 );
not ( n970 , n969 );
not ( n971 , n85 );
nor ( n972 , n971 , n713 );
nor ( n973 , n972 , n723 );
not ( n974 , n973 );
or ( n975 , n970 , n974 );
not ( n976 , n87 );
nand ( n977 , n976 , n630 );
not ( n978 , n977 );
not ( n979 , n731 );
or ( n980 , n978 , n979 );
and ( n981 , n605 , n90 );
and ( n982 , n635 , n88 );
not ( n983 , n89 );
nor ( n984 , n983 , n774 );
nor ( n985 , n981 , n982 , n984 );
nand ( n986 , n980 , n985 );
nand ( n987 , n975 , n986 );
and ( n988 , n753 , n80 );
not ( n989 , n3 );
not ( n990 , n2 );
or ( n991 , n989 , n990 );
or ( n992 , n2 , n3 );
nand ( n993 , n991 , n992 );
nand ( n994 , n993 , n82 );
not ( n995 , n994 );
not ( n996 , n583 );
and ( n997 , n995 , n996 );
and ( n998 , n571 , n81 );
nor ( n999 , n997 , n998 );
nand ( n1000 , n577 , n79 );
and ( n1001 , n999 , n1000 );
nor ( n1002 , n1001 , n596 );
nor ( n1003 , n988 , n1002 );
nand ( n1004 , n83 , n750 );
nand ( n1005 , n987 , n1003 , n1004 );
and ( n1006 , n753 , n164 );
not ( n1007 , n166 );
not ( n1008 , n553 );
nor ( n1009 , n1008 , n596 );
not ( n1010 , n1009 );
or ( n1011 , n1007 , n1010 );
nand ( n1012 , n571 , n595 );
not ( n1013 , n1012 );
nand ( n1014 , n1013 , n162 );
nand ( n1015 , n1011 , n1014 );
nor ( n1016 , n1006 , n1015 );
not ( n1017 , n5 );
nand ( n1018 , n549 , n1017 , n4 );
nor ( n1019 , n1018 , n547 );
and ( n1020 , n1019 , n709 );
nand ( n1021 , n1020 , n16 );
nand ( n1022 , n871 , n168 );
and ( n1023 , n1021 , n1022 );
not ( n1024 , n165 );
not ( n1025 , n660 );
or ( n1026 , n1024 , n1025 );
nand ( n1027 , n622 , n861 );
not ( n1028 , n1027 );
not ( n1029 , n893 );
nand ( n1030 , n1028 , n1029 , n169 );
nand ( n1031 , n1026 , n1030 );
and ( n1032 , n850 , n161 );
and ( n1033 , n1019 , n167 );
nor ( n1034 , n1032 , n1033 );
nand ( n1035 , n577 , n163 );
and ( n1036 , n1034 , n1035 );
nor ( n1037 , n1036 , n596 );
nor ( n1038 , n1031 , n1037 );
nand ( n1039 , n635 , n170 );
nand ( n1040 , n605 , n172 );
nand ( n1041 , n611 , n171 );
nand ( n1042 , n1039 , n1040 , n1041 );
and ( n1043 , n1042 , n723 );
not ( n1044 , n861 );
nand ( n1045 , n659 , n1044 , n17 );
not ( n1046 , n1045 );
and ( n1047 , n1046 , n121 );
nor ( n1048 , n1043 , n1047 );
nand ( n1049 , n1016 , n1023 , n1038 , n1048 );
nand ( n1050 , n742 , n176 );
nand ( n1051 , n850 , n177 );
nand ( n1052 , n852 , n174 );
nand ( n1053 , n1050 , n1051 , n1052 );
nand ( n1054 , n744 , n175 );
nand ( n1055 , n577 , n173 );
nand ( n1056 , n1054 , n1055 , n857 );
or ( n1057 , n1053 , n1056 );
or ( n1058 , n863 , n135 );
nand ( n1059 , n1057 , n1058 );
not ( n1060 , n178 );
not ( n1061 , n1060 );
not ( n1062 , n871 );
or ( n1063 , n1061 , n1062 );
not ( n1064 , n730 );
not ( n1065 , n179 );
not ( n1066 , n1065 );
and ( n1067 , n1064 , n1066 );
not ( n1068 , n181 );
nor ( n1069 , n1068 , n878 );
nor ( n1070 , n1067 , n1069 );
nand ( n1071 , n605 , n182 );
nand ( n1072 , n635 , n180 );
nand ( n1073 , n1070 , n723 , n1071 , n1072 );
nand ( n1074 , n1063 , n1073 );
nor ( n1075 , n1059 , n1074 );
and ( n1076 , n753 , n200 );
nor ( n1077 , n16 , n195 );
not ( n1078 , n1077 );
not ( n1079 , n1078 );
not ( n1080 , n1020 );
or ( n1081 , n1079 , n1080 );
buf ( n1082 , n551 );
nand ( n1083 , n1082 , n595 );
not ( n1084 , n1083 );
nand ( n1085 , n1084 , n196 );
nand ( n1086 , n1081 , n1085 );
nor ( n1087 , n1076 , n1086 );
and ( n1088 , n871 , n201 );
not ( n1089 , n198 );
nor ( n1090 , n1089 , n1012 );
nor ( n1091 , n1088 , n1090 );
nand ( n1092 , n605 , n205 );
nand ( n1093 , n622 , n202 );
nand ( n1094 , n635 , n203 );
nand ( n1095 , n611 , n204 );
nand ( n1096 , n1092 , n1093 , n1094 , n1095 );
and ( n1097 , n1096 , n723 );
and ( n1098 , n1046 , n72 );
nor ( n1099 , n1097 , n1098 );
and ( n1100 , n588 , n194 );
not ( n1101 , n197 );
not ( n1102 , n850 );
or ( n1103 , n1101 , n1102 );
nand ( n1104 , n577 , n199 );
nand ( n1105 , n1103 , n1104 );
or ( n1106 , n1100 , n1105 );
nand ( n1107 , n1106 , n597 );
nand ( n1108 , n1087 , n1091 , n1099 , n1107 );
not ( n1109 , n1020 );
not ( n1110 , n1109 );
not ( n1111 , n16 );
not ( n1112 , n207 );
nand ( n1113 , n1111 , n1112 );
not ( n1114 , n1113 );
not ( n1115 , n1114 );
and ( n1116 , n1110 , n1115 );
and ( n1117 , n1046 , n213 );
nor ( n1118 , n1116 , n1117 );
and ( n1119 , n753 , n212 );
not ( n1120 , n208 );
nor ( n1121 , n1120 , n1083 );
nor ( n1122 , n1119 , n1121 );
nand ( n1123 , n779 , n206 );
nand ( n1124 , n571 , n210 );
nand ( n1125 , n850 , n209 );
nand ( n1126 , n577 , n211 );
nand ( n1127 , n1123 , n1124 , n1125 , n1126 );
nand ( n1128 , n1127 , n893 );
nand ( n1129 , n605 , n216 );
nand ( n1130 , n622 , n217 );
nand ( n1131 , n635 , n215 );
nand ( n1132 , n611 , n218 );
nand ( n1133 , n1129 , n1130 , n1131 , n1132 );
and ( n1134 , n1133 , n723 );
and ( n1135 , n871 , n214 );
nor ( n1136 , n1134 , n1135 );
nand ( n1137 , n1118 , n1122 , n1128 , n1136 );
not ( n1138 , n1109 );
nor ( n1139 , n16 , n233 );
not ( n1140 , n1139 );
and ( n1141 , n1138 , n1140 );
and ( n1142 , n1046 , n14 );
nor ( n1143 , n1141 , n1142 );
nand ( n1144 , n779 , n232 );
nand ( n1145 , n850 , n237 );
nand ( n1146 , n577 , n235 );
nand ( n1147 , n236 , n852 );
nand ( n1148 , n1144 , n1145 , n1146 , n1147 );
nand ( n1149 , n1148 , n893 );
nand ( n1150 , n605 , n241 );
nand ( n1151 , n622 , n242 );
nand ( n1152 , n635 , n243 );
nand ( n1153 , n611 , n240 );
nand ( n1154 , n1150 , n1151 , n1152 , n1153 );
and ( n1155 , n1154 , n723 );
and ( n1156 , n871 , n239 );
nor ( n1157 , n1155 , n1156 );
and ( n1158 , n1013 , n238 );
not ( n1159 , n234 );
nor ( n1160 , n1159 , n1083 );
nor ( n1161 , n1158 , n1160 );
nand ( n1162 , n1143 , n1149 , n1157 , n1161 );
not ( n1163 , n344 );
nor ( n1164 , n1163 , n16 );
and ( n1165 , n1164 , n345 );
and ( n1166 , n360 , n361 );
nand ( n1167 , n1165 , n1166 );
and ( n1168 , n1167 , n345 );
nand ( n1169 , n620 , n363 );
nor ( n1170 , n1168 , n1169 );
and ( n1171 , n345 , n364 );
nand ( n1172 , n1170 , n1171 );
not ( n1173 , n1172 );
and ( n1174 , n365 , n366 );
nand ( n1175 , n1173 , n1174 );
not ( n1176 , n16 );
nand ( n1177 , n1176 , n346 );
not ( n1178 , n1177 );
or ( n1179 , n1175 , n1178 , n362 );
not ( n1180 , n362 );
and ( n1181 , n1177 , n552 );
not ( n1182 , n1181 );
nor ( n1183 , n1180 , n1182 );
nand ( n1184 , n1175 , n1183 );
nand ( n1185 , n1179 , n1184 );
nand ( n1186 , n742 , n219 );
and ( n1187 , n571 , n223 );
not ( n1188 , n652 );
and ( n1189 , n1188 , n225 );
nor ( n1190 , n1187 , n1189 );
buf ( n1191 , n553 );
nand ( n1192 , n1191 , n221 );
and ( n1193 , n1019 , n220 );
nor ( n1194 , n1193 , n719 );
nand ( n1195 , n1186 , n1190 , n1192 , n1194 );
not ( n1196 , n1027 );
nand ( n1197 , n1196 , n228 );
nand ( n1198 , n1197 , n596 );
nand ( n1199 , n1195 , n1198 );
and ( n1200 , n750 , n222 );
or ( n1201 , n671 , n719 );
not ( n1202 , n1201 );
and ( n1203 , n1202 , n224 );
nor ( n1204 , n1200 , n1203 );
nand ( n1205 , n635 , n229 );
nand ( n1206 , n605 , n231 );
nand ( n1207 , n611 , n230 );
nand ( n1208 , n1205 , n1206 , n1207 );
and ( n1209 , n1208 , n723 );
and ( n1210 , n871 , n227 );
nor ( n1211 , n1209 , n1210 );
nand ( n1212 , n1046 , n226 );
and ( n1213 , n1021 , n1212 );
nand ( n1214 , n1199 , n1204 , n1211 , n1213 );
not ( n1215 , n279 );
not ( n1216 , n1013 );
or ( n1217 , n1215 , n1216 );
nand ( n1218 , n1084 , n282 );
nand ( n1219 , n1217 , n1218 );
and ( n1220 , n752 , n280 );
nor ( n1221 , n1219 , n1220 );
not ( n1222 , n660 );
not ( n1223 , n1222 );
not ( n1224 , n281 );
not ( n1225 , n1224 );
and ( n1226 , n1223 , n1225 );
not ( n1227 , n278 );
not ( n1228 , n850 );
or ( n1229 , n1227 , n1228 );
nor ( n1230 , n16 , n283 );
not ( n1231 , n1230 );
nand ( n1232 , n1231 , n1019 );
nand ( n1233 , n1229 , n1232 );
and ( n1234 , n1233 , n597 );
nor ( n1235 , n1226 , n1234 );
nand ( n1236 , n622 , n285 );
nand ( n1237 , n605 , n286 );
nand ( n1238 , n635 , n287 );
nand ( n1239 , n611 , n288 );
nand ( n1240 , n1236 , n1237 , n1238 , n1239 );
and ( n1241 , n1240 , n723 );
and ( n1242 , n871 , n284 );
nor ( n1243 , n1241 , n1242 );
not ( n1244 , n1201 );
not ( n1245 , n159 );
not ( n1246 , n1245 );
and ( n1247 , n1244 , n1246 );
and ( n1248 , n1046 , n123 );
nor ( n1249 , n1247 , n1248 );
nand ( n1250 , n1221 , n1235 , n1243 , n1249 );
not ( n1251 , n1109 );
not ( n1252 , n16 );
not ( n1253 , n306 );
nand ( n1254 , n1252 , n1253 );
not ( n1255 , n1254 );
not ( n1256 , n1255 );
and ( n1257 , n1251 , n1256 );
and ( n1258 , n1046 , n60 );
nor ( n1259 , n1257 , n1258 );
nand ( n1260 , n850 , n300 );
not ( n1261 , n587 );
nand ( n1262 , n1261 , n304 );
nand ( n1263 , n577 , n302 );
nand ( n1264 , n303 , n852 );
nand ( n1265 , n1260 , n1262 , n1263 , n1264 );
nand ( n1266 , n1265 , n680 );
nand ( n1267 , n605 , n309 );
nand ( n1268 , n622 , n310 );
nand ( n1269 , n635 , n311 );
nand ( n1270 , n611 , n308 );
nand ( n1271 , n1267 , n1268 , n1269 , n1270 );
and ( n1272 , n1271 , n723 );
and ( n1273 , n871 , n307 );
nor ( n1274 , n1272 , n1273 );
and ( n1275 , n1013 , n301 );
not ( n1276 , n305 );
nor ( n1277 , n1276 , n1083 );
nor ( n1278 , n1275 , n1277 );
nand ( n1279 , n1259 , n1266 , n1274 , n1278 );
not ( n1280 , n328 );
nor ( n1281 , n587 , n1280 );
not ( n1282 , n325 );
not ( n1283 , n571 );
or ( n1284 , n1282 , n1283 );
nand ( n1285 , n327 , n651 );
nand ( n1286 , n1284 , n1285 );
or ( n1287 , n1281 , n1286 );
nand ( n1288 , n1287 , n681 );
and ( n1289 , n1021 , n1288 );
nand ( n1290 , n1009 , n329 );
nand ( n1291 , n730 , n861 );
and ( n1292 , n1044 , n869 );
nor ( n1293 , n1044 , n332 );
nor ( n1294 , n1292 , n1293 );
not ( n1295 , n861 );
not ( n1296 , n110 );
and ( n1297 , n1295 , n1296 );
nor ( n1298 , n1297 , n595 );
nand ( n1299 , n1291 , n1294 , n1298 );
nand ( n1300 , n1020 , n330 );
and ( n1301 , n1290 , n1299 , n1300 );
and ( n1302 , n750 , n324 );
and ( n1303 , n1202 , n326 );
nor ( n1304 , n1302 , n1303 );
nand ( n1305 , n635 , n333 );
nand ( n1306 , n605 , n335 );
nand ( n1307 , n611 , n334 );
nand ( n1308 , n1305 , n1306 , n1307 );
and ( n1309 , n1308 , n723 );
and ( n1310 , n871 , n331 );
nor ( n1311 , n1309 , n1310 );
nand ( n1312 , n1289 , n1301 , n1304 , n1311 );
and ( n1313 , n315 , n753 );
not ( n1314 , n16 );
not ( n1315 , n318 );
nand ( n1316 , n1314 , n1315 );
not ( n1317 , n1316 );
not ( n1318 , n1020 );
or ( n1319 , n1317 , n1318 );
nand ( n1320 , n1084 , n620 , n316 );
nand ( n1321 , n1319 , n1320 );
nor ( n1322 , n1313 , n1321 );
not ( n1323 , n1201 );
not ( n1324 , n314 );
not ( n1325 , n1324 );
and ( n1326 , n1323 , n1325 );
not ( n1327 , n863 );
and ( n1328 , n1327 , n84 );
nor ( n1329 , n1326 , n1328 );
and ( n1330 , n871 , n319 );
not ( n1331 , n313 );
nor ( n1332 , n1331 , n1012 );
nor ( n1333 , n1330 , n1332 );
nand ( n1334 , n605 , n323 );
nand ( n1335 , n622 , n320 );
nand ( n1336 , n635 , n321 );
nand ( n1337 , n611 , n322 );
nand ( n1338 , n1334 , n1335 , n1336 , n1337 );
and ( n1339 , n1338 , n723 );
nand ( n1340 , n312 , n850 );
nand ( n1341 , n1261 , n317 );
nand ( n1342 , n1340 , n1341 );
and ( n1343 , n1342 , n597 );
nor ( n1344 , n1339 , n1343 );
nand ( n1345 , n1322 , n1329 , n1333 , n1344 );
and ( n1346 , n250 , n753 );
nor ( n1347 , n16 , n245 );
not ( n1348 , n1347 );
not ( n1349 , n1348 );
not ( n1350 , n1020 );
or ( n1351 , n1349 , n1350 );
nand ( n1352 , n1084 , n552 , n246 );
nand ( n1353 , n1351 , n1352 );
nor ( n1354 , n1346 , n1353 );
not ( n1355 , n1201 );
not ( n1356 , n249 );
not ( n1357 , n1356 );
and ( n1358 , n1355 , n1357 );
and ( n1359 , n1327 , n96 );
nor ( n1360 , n1358 , n1359 );
and ( n1361 , n871 , n251 );
not ( n1362 , n248 );
nor ( n1363 , n1362 , n1012 );
nor ( n1364 , n1361 , n1363 );
nand ( n1365 , n605 , n255 );
nand ( n1366 , n622 , n252 );
nand ( n1367 , n635 , n253 );
nand ( n1368 , n611 , n254 );
nand ( n1369 , n1365 , n1366 , n1367 , n1368 );
and ( n1370 , n1369 , n723 );
not ( n1371 , n247 );
not ( n1372 , n850 );
or ( n1373 , n1371 , n1372 );
nand ( n1374 , n1261 , n244 );
nand ( n1375 , n1373 , n1374 );
and ( n1376 , n1375 , n680 );
nor ( n1377 , n1370 , n1376 );
nand ( n1378 , n1354 , n1360 , n1364 , n1377 );
not ( n1379 , n1222 );
and ( n1380 , n1379 , n9 );
and ( n1381 , n753 , n7 );
nor ( n1382 , n1380 , n1381 );
and ( n1383 , n1013 , n8 );
and ( n1384 , n1202 , n1 );
nor ( n1385 , n1383 , n1384 );
not ( n1386 , n28 );
not ( n1387 , n1028 );
or ( n1388 , n1386 , n1387 );
nand ( n1389 , n638 , n19 );
nand ( n1390 , n17 , n18 );
nand ( n1391 , n1389 , n646 , n1390 );
nand ( n1392 , n1388 , n1391 );
and ( n1393 , n1392 , n1029 );
and ( n1394 , n750 , n10 );
nor ( n1395 , n1393 , n1394 );
not ( n1396 , n680 );
not ( n1397 , n29 );
not ( n1398 , n605 );
or ( n1399 , n1397 , n1398 );
and ( n1400 , n635 , n27 );
and ( n1401 , n611 , n30 );
nor ( n1402 , n1400 , n1401 );
nand ( n1403 , n1399 , n1402 );
nand ( n1404 , n1396 , n1403 , n630 );
nand ( n1405 , n1382 , n1385 , n1395 , n1404 );
nor ( n1406 , n16 , n290 );
not ( n1407 , n1406 );
and ( n1408 , n1019 , n1407 );
and ( n1409 , n1082 , n291 );
nor ( n1410 , n1408 , n1409 );
nand ( n1411 , n744 , n294 );
nand ( n1412 , n1261 , n289 );
nand ( n1413 , n850 , n293 );
nand ( n1414 , n1410 , n1411 , n1412 , n1413 );
nand ( n1415 , n1414 , n597 );
not ( n1416 , n1201 );
not ( n1417 , n156 );
not ( n1418 , n1417 );
and ( n1419 , n1416 , n1418 );
and ( n1420 , n1327 , n48 );
nor ( n1421 , n1419 , n1420 );
nand ( n1422 , n605 , n297 );
nand ( n1423 , n622 , n296 );
nand ( n1424 , n298 , n635 );
nand ( n1425 , n611 , n299 );
nand ( n1426 , n1422 , n1423 , n1424 , n1425 );
and ( n1427 , n1426 , n723 );
and ( n1428 , n871 , n295 );
nor ( n1429 , n1427 , n1428 );
nand ( n1430 , n753 , n292 );
nand ( n1431 , n1415 , n1421 , n1429 , n1430 );
not ( n1432 , n40 );
not ( n1433 , n605 );
or ( n1434 , n1432 , n1433 );
nand ( n1435 , n611 , n39 );
nand ( n1436 , n1434 , n1435 );
and ( n1437 , n635 , n41 );
or ( n1438 , n1436 , n1437 );
nand ( n1439 , n1438 , n630 );
and ( n1440 , n1028 , n42 );
nor ( n1441 , n861 , n869 );
nand ( n1442 , n1441 , n37 );
not ( n1443 , n38 );
not ( n1444 , n641 );
or ( n1445 , n1443 , n1444 );
nand ( n1446 , n638 , n14 );
nand ( n1447 , n1445 , n1446 );
nand ( n1448 , n646 , n1447 );
nand ( n1449 , n1442 , n1448 , n659 );
nor ( n1450 , n1440 , n1449 );
and ( n1451 , n1439 , n1450 );
not ( n1452 , n36 );
not ( n1453 , n750 );
or ( n1454 , n1452 , n1453 );
nand ( n1455 , n620 , n1084 , n35 );
nand ( n1456 , n1454 , n1455 );
nor ( n1457 , n1451 , n1456 );
and ( n1458 , n742 , n106 );
and ( n1459 , n577 , n103 );
and ( n1460 , n744 , n105 );
nor ( n1461 , n1458 , n1459 , n1460 );
and ( n1462 , n1191 , n107 );
and ( n1463 , n850 , n108 );
nor ( n1464 , n1462 , n1463 );
not ( n1465 , n104 );
not ( n1466 , n1465 );
not ( n1467 , n597 );
or ( n1468 , n1466 , n1467 );
nand ( n1469 , n1468 , n653 );
and ( n1470 , n1461 , n1464 , n1469 );
nand ( n1471 , n605 , n114 );
nand ( n1472 , n622 , n111 );
nand ( n1473 , n1471 , n1472 , n630 );
not ( n1474 , n112 );
not ( n1475 , n635 );
or ( n1476 , n1474 , n1475 );
nand ( n1477 , n611 , n113 );
nand ( n1478 , n1476 , n1477 );
or ( n1479 , n1473 , n1478 );
and ( n1480 , n638 , n84 );
and ( n1481 , n641 , n110 );
and ( n1482 , n17 , n109 );
nor ( n1483 , n1480 , n1481 , n1482 );
nand ( n1484 , n1483 , n646 );
nand ( n1485 , n1479 , n1484 );
and ( n1486 , n1485 , n596 );
nor ( n1487 , n1470 , n1486 );
and ( n1488 , n1173 , n1177 , n365 );
and ( n1489 , n1181 , n366 );
nor ( n1490 , n1488 , n1489 );
not ( n1491 , n347 );
or ( n1492 , n1491 , n16 , n348 );
not ( n1493 , n353 );
nand ( n1494 , n1493 , n55 );
or ( n1495 , n1255 , n1494 );
not ( n1496 , n359 );
nand ( n1497 , n1496 , n67 );
or ( n1498 , n1497 , n1077 );
nand ( n1499 , n1495 , n1498 );
not ( n1500 , n1 );
and ( n1501 , n356 , n1500 );
not ( n1502 , n356 );
and ( n1503 , n1502 , n1 );
nor ( n1504 , n1501 , n1503 );
or ( n1505 , n1139 , n1504 );
and ( n1506 , n91 , n350 );
not ( n1507 , n91 );
not ( n1508 , n350 );
and ( n1509 , n1507 , n1508 );
or ( n1510 , n1506 , n1509 );
or ( n1511 , n1347 , n1510 );
nand ( n1512 , n1505 , n1511 );
nor ( n1513 , n1499 , n1512 );
not ( n1514 , n358 );
and ( n1515 , n357 , n1514 );
not ( n1516 , n357 );
and ( n1517 , n1516 , n358 );
nor ( n1518 , n1515 , n1517 );
or ( n1519 , n1114 , n1518 );
xnor ( n1520 , n351 , n43 );
or ( n1521 , n1520 , n1406 );
nand ( n1522 , n1519 , n1521 );
and ( n1523 , n79 , n352 );
not ( n1524 , n79 );
not ( n1525 , n352 );
and ( n1526 , n1524 , n1525 );
nor ( n1527 , n1523 , n1526 );
not ( n1528 , n1527 );
not ( n1529 , n1316 );
or ( n1530 , n1528 , n1529 );
nand ( n1531 , n1530 , n159 );
nor ( n1532 , n1522 , n1531 );
not ( n1533 , n355 );
and ( n1534 , n354 , n1533 );
not ( n1535 , n354 );
and ( n1536 , n1535 , n355 );
nor ( n1537 , n1534 , n1536 );
or ( n1538 , n1230 , n1537 );
not ( n1539 , n55 );
nand ( n1540 , n1539 , n353 );
or ( n1541 , n1255 , n1540 );
nand ( n1542 , n1538 , n1541 );
nor ( n1543 , n1077 , n1496 , n67 );
nor ( n1544 , n1542 , n1543 );
nand ( n1545 , n1513 , n1532 , n1544 );
nand ( n1546 , n163 , n349 );
nand ( n1547 , n1546 , n348 );
or ( n1548 , n1545 , n1547 );
nand ( n1549 , n1492 , n1548 );
or ( n1550 , n1172 , n1178 , n365 );
not ( n1551 , n365 );
nor ( n1552 , n1551 , n1182 );
nand ( n1553 , n1172 , n1552 );
nand ( n1554 , n1550 , n1553 );
not ( n1555 , n367 );
or ( n1556 , n1555 , n16 , n348 );
not ( n1557 , n1078 );
not ( n1558 , n71 );
nor ( n1559 , n1558 , n359 );
not ( n1560 , n1559 );
or ( n1561 , n1557 , n1560 );
not ( n1562 , n59 );
nand ( n1563 , n1562 , n1254 , n353 );
nand ( n1564 , n1561 , n1563 );
and ( n1565 , n83 , n352 );
not ( n1566 , n83 );
and ( n1567 , n1566 , n1525 );
nor ( n1568 , n1565 , n1567 );
not ( n1569 , n1568 );
not ( n1570 , n1316 );
or ( n1571 , n1569 , n1570 );
not ( n1572 , n1139 );
and ( n1573 , n10 , n356 );
not ( n1574 , n10 );
not ( n1575 , n356 );
and ( n1576 , n1574 , n1575 );
nor ( n1577 , n1573 , n1576 );
nand ( n1578 , n1572 , n1577 );
nand ( n1579 , n1571 , n1578 );
nor ( n1580 , n1564 , n1579 );
and ( n1581 , n95 , n350 );
not ( n1582 , n95 );
and ( n1583 , n1582 , n1508 );
nor ( n1584 , n1581 , n1583 );
not ( n1585 , n1584 );
not ( n1586 , n1348 );
or ( n1587 , n1585 , n1586 );
and ( n1588 , n357 , n369 );
not ( n1589 , n357 );
not ( n1590 , n369 );
and ( n1591 , n1589 , n1590 );
nor ( n1592 , n1588 , n1591 );
nand ( n1593 , n1113 , n1592 );
nand ( n1594 , n1587 , n1593 );
and ( n1595 , n351 , n47 );
not ( n1596 , n351 );
not ( n1597 , n47 );
and ( n1598 , n1596 , n1597 );
nor ( n1599 , n1595 , n1598 );
not ( n1600 , n1599 );
not ( n1601 , n1407 );
or ( n1602 , n1600 , n1601 );
nand ( n1603 , n1602 , n278 );
nor ( n1604 , n1594 , n1603 );
nand ( n1605 , n1078 , n1558 , n359 );
not ( n1606 , n59 );
nor ( n1607 , n1606 , n353 );
nand ( n1608 , n1254 , n1607 );
not ( n1609 , n1230 );
and ( n1610 , n354 , n368 );
not ( n1611 , n354 );
not ( n1612 , n368 );
and ( n1613 , n1611 , n1612 );
nor ( n1614 , n1610 , n1613 );
nand ( n1615 , n1609 , n1614 );
and ( n1616 , n1605 , n1608 , n1615 );
nand ( n1617 , n1580 , n1604 , n1616 );
nand ( n1618 , n161 , n349 );
nand ( n1619 , n1618 , n348 );
or ( n1620 , n1617 , n1619 );
nand ( n1621 , n1556 , n1620 );
nand ( n1622 , n1177 , n345 );
not ( n1623 , n1622 );
and ( n1624 , n1170 , n1623 );
and ( n1625 , n1181 , n364 );
nor ( n1626 , n1624 , n1625 );
nor ( n1627 , n1173 , n1626 );
nor ( n1628 , n1545 , n1546 );
not ( n1629 , n1167 );
not ( n1630 , n1169 );
or ( n1631 , n1629 , n1622 , n1630 );
not ( n1632 , n1170 );
or ( n1633 , n1632 , n1178 );
nand ( n1634 , n1631 , n1633 );
not ( n1635 , n337 );
not ( n1636 , n339 );
nor ( n1637 , n1636 , n338 );
nor ( n1638 , n340 , n341 );
not ( n1639 , n342 );
nand ( n1640 , n1637 , n1638 , n1639 , n153 );
nor ( n1641 , n16 , n343 );
not ( n1642 , n1641 );
nor ( n1643 , n1640 , n1642 );
not ( n1644 , n1643 );
or ( n1645 , n1635 , n1644 );
and ( n1646 , n1640 , n1641 );
and ( n1647 , n1646 , n247 );
and ( n1648 , n1642 , n317 );
nor ( n1649 , n1647 , n1648 );
nand ( n1650 , n1645 , n1649 );
not ( n1651 , n336 );
not ( n1652 , n1643 );
or ( n1653 , n1651 , n1652 );
and ( n1654 , n1646 , n312 );
and ( n1655 , n1642 , n289 );
nor ( n1656 , n1654 , n1655 );
nand ( n1657 , n1653 , n1656 );
not ( n1658 , n1646 );
not ( n1659 , n278 );
or ( n1660 , n1658 , n1659 );
nor ( n1661 , n289 , n317 );
or ( n1662 , n1661 , n1641 );
nand ( n1663 , n1643 , n160 );
nand ( n1664 , n1660 , n1662 , n1663 );
not ( n1665 , n152 );
not ( n1666 , n154 );
nand ( n1667 , n1665 , n1666 , n150 , n151 );
not ( n1668 , n155 );
nand ( n1669 , n1668 , n153 );
nor ( n1670 , n1667 , n1669 );
not ( n1671 , n1670 );
nor ( n1672 , n16 , n158 );
nand ( n1673 , n1671 , n1672 );
or ( n1674 , n1673 , n1417 );
and ( n1675 , n1670 , n1672 );
nand ( n1676 , n1675 , n157 );
nand ( n1677 , n1674 , n1676 );
or ( n1678 , n1673 , n1245 );
nand ( n1679 , n1675 , n160 );
nand ( n1680 , n1678 , n1679 );
or ( n1681 , n1673 , n1324 );
nand ( n1682 , n1675 , n336 );
nand ( n1683 , n1681 , n1682 );
or ( n1684 , n1356 , n1673 );
nand ( n1685 , n1675 , n337 );
nand ( n1686 , n1684 , n1685 );
not ( n1687 , n157 );
not ( n1688 , n1643 );
or ( n1689 , n1687 , n1688 );
nand ( n1690 , n1646 , n293 );
nand ( n1691 , n1689 , n1690 );
not ( n1692 , n1165 );
nand ( n1693 , n1692 , n360 );
not ( n1694 , n360 );
nand ( n1695 , n1694 , n345 , n344 );
and ( n1696 , n1693 , n1695 );
nor ( n1697 , n1696 , n1182 );
and ( n1698 , n1165 , n1177 , n360 );
and ( n1699 , n1181 , n361 );
nor ( n1700 , n1698 , n1699 );
nor ( n1701 , n1700 , n1629 );
not ( n1702 , n374 );
not ( n1703 , n1181 );
or ( n1704 , n1702 , n1703 );
nand ( n1705 , n1177 , n373 );
nand ( n1706 , n1704 , n1705 );
nor ( n1707 , n1622 , n1164 );
not ( n1708 , n371 );
and ( n1709 , n1708 , n391 );
and ( n1710 , n3 , n371 );
nor ( n1711 , n1709 , n1710 );
not ( n1712 , n1711 );
and ( n1713 , n1708 , n389 );
and ( n1714 , n351 , n371 );
nor ( n1715 , n1713 , n1714 );
not ( n1716 , n1715 );
and ( n1717 , n1708 , n390 );
and ( n1718 , n354 , n371 );
nor ( n1719 , n1717 , n1718 );
not ( n1720 , n1719 );
and ( n1721 , n1708 , n403 );
and ( n1722 , n2 , n371 );
nor ( n1723 , n1721 , n1722 );
not ( n1724 , n1723 );
and ( n1725 , n1708 , n394 );
and ( n1726 , n4 , n371 );
nor ( n1727 , n1725 , n1726 );
not ( n1728 , n1727 );
not ( n1729 , n379 );
not ( n1730 , n16 );
nand ( n1731 , n1730 , n378 );
nand ( n1732 , n1729 , n1731 );
nor ( n1733 , n376 , n377 );
nor ( n1734 , n1733 , n16 );
and ( n1735 , n371 , n402 );
not ( n1736 , n371 );
and ( n1737 , n1736 , n401 );
or ( n1738 , n1735 , n1737 );
and ( n1739 , n371 , n410 );
not ( n1740 , n371 );
and ( n1741 , n1740 , n409 );
or ( n1742 , n1739 , n1741 );
and ( n1743 , n371 , n348 , n370 );
and ( n1744 , n371 , n393 );
not ( n1745 , n371 );
and ( n1746 , n1745 , n392 );
or ( n1747 , n1744 , n1746 );
and ( n1748 , n371 , n398 );
not ( n1749 , n371 );
and ( n1750 , n1749 , n397 );
or ( n1751 , n1748 , n1750 );
and ( n1752 , n371 , n386 );
not ( n1753 , n371 );
and ( n1754 , n1753 , n385 );
or ( n1755 , n1752 , n1754 );
and ( n1756 , n371 , n388 );
not ( n1757 , n371 );
and ( n1758 , n1757 , n387 );
or ( n1759 , n1756 , n1758 );
and ( n1760 , n371 , n396 );
not ( n1761 , n371 );
and ( n1762 , n1761 , n395 );
or ( n1763 , n1760 , n1762 );
and ( n1764 , n371 , n400 );
not ( n1765 , n371 );
and ( n1766 , n1765 , n399 );
or ( n1767 , n1764 , n1766 );
and ( n1768 , n371 , n405 );
not ( n1769 , n371 );
and ( n1770 , n1769 , n404 );
or ( n1771 , n1768 , n1770 );
and ( n1772 , n371 , n407 );
not ( n1773 , n371 );
and ( n1774 , n1773 , n406 );
or ( n1775 , n1772 , n1774 );
and ( n1776 , n371 , n6 );
not ( n1777 , n371 );
and ( n1778 , n1777 , n408 );
or ( n1779 , n1776 , n1778 );
and ( n1780 , n371 , n5 );
not ( n1781 , n371 );
and ( n1782 , n1781 , n411 );
or ( n1783 , n1780 , n1782 );
or ( n1784 , n16 , n383 );
or ( n1785 , n16 , n382 );
not ( n1786 , n375 );
nor ( n1787 , n1786 , n16 );
nand ( n1788 , n370 , n372 );
or ( n1789 , n16 , n381 );
or ( n1790 , n16 , n380 );
or ( n1791 , n16 , n384 );
not ( n1792 , n16 );
not ( n1793 , n16 );
not ( n1794 , n1617 );
not ( n1795 , n1618 );
and ( n1796 , n1794 , n1795 );
nor ( n1797 , n1796 , n1628 );
and ( n1798 , n1743 , n1797 );
not ( n1799 , n1743 );
and ( n1800 , n1799 , n1788 );
nor ( n1801 , n1798 , n1800 );
not ( n1802 , n1175 );
nor ( n1803 , n1802 , n1490 );
endmodule
