module galois8MulOpt(
    input wire [7:0] in,
    output wire [7:0] out
);

  parameter constVal = 0;

  `define C(ind, val) assign tab[ind] = 8'd``val
  wire [7:0] tab [255:0];

  if (constVal == 8'h1) begin
    assign out = in;
  end if (constVal == 8'h94) begin
    `C(0, 0); `C(1, 148); `C(2, 235); `C(3, 127); `C(4, 21); `C(5, 129);
    `C(6, 254); `C(7, 106); `C(8, 42); `C(9, 190); `C(10, 193); `C(11, 85);
    `C(12, 63); `C(13, 171); `C(14, 212); `C(15, 64); `C(16, 84); `C(17, 192);
    `C(18, 191); `C(19, 43); `C(20, 65); `C(21, 213); `C(22, 170); `C(23, 62);
    `C(24, 126); `C(25, 234); `C(26, 149); `C(27, 1); `C(28, 107); `C(29, 255);
    `C(30, 128); `C(31, 20); `C(32, 168); `C(33, 60); `C(34, 67); `C(35, 215);
    `C(36, 189); `C(37, 41); `C(38, 86); `C(39, 194); `C(40, 130); `C(41, 22);
    `C(42, 105); `C(43, 253); `C(44, 151); `C(45, 3); `C(46, 124); `C(47, 232);
    `C(48, 252); `C(49, 104); `C(50, 23); `C(51, 131); `C(52, 233);
    `C(53, 125); `C(54, 2); `C(55, 150); `C(56, 214); `C(57, 66); `C(58, 61);
    `C(59, 169); `C(60, 195); `C(61, 87); `C(62, 40); `C(63, 188); `C(64, 147);
    `C(65, 7); `C(66, 120); `C(67, 236); `C(68, 134); `C(69, 18); `C(70, 109);
    `C(71, 249); `C(72, 185); `C(73, 45); `C(74, 82); `C(75, 198); `C(76, 172);
    `C(77, 56); `C(78, 71); `C(79, 211); `C(80, 199); `C(81, 83); `C(82, 44);
    `C(83, 184); `C(84, 210); `C(85, 70); `C(86, 57); `C(87, 173); `C(88, 237);
    `C(89, 121); `C(90, 6); `C(91, 146); `C(92, 248); `C(93, 108); `C(94, 19);
    `C(95, 135); `C(96, 59); `C(97, 175); `C(98, 208); `C(99, 68); `C(100, 46);
    `C(101, 186); `C(102, 197); `C(103, 81); `C(104, 17); `C(105, 133);
    `C(106, 250); `C(107, 110); `C(108, 4); `C(109, 144); `C(110, 239);
    `C(111, 123); `C(112, 111); `C(113, 251); `C(114, 132); `C(115, 16);
    `C(116, 122); `C(117, 238); `C(118, 145); `C(119, 5); `C(120, 69);
    `C(121, 209); `C(122, 174); `C(123, 58); `C(124, 80); `C(125, 196);
    `C(126, 187); `C(127, 47); `C(128, 229); `C(129, 113); `C(130, 14);
    `C(131, 154); `C(132, 240); `C(133, 100); `C(134, 27); `C(135, 143);
    `C(136, 207); `C(137, 91); `C(138, 36); `C(139, 176); `C(140, 218);
    `C(141, 78); `C(142, 49); `C(143, 165); `C(144, 177); `C(145, 37);
    `C(146, 90); `C(147, 206); `C(148, 164); `C(149, 48); `C(150, 79);
    `C(151, 219); `C(152, 155); `C(153, 15); `C(154, 112); `C(155, 228);
    `C(156, 142); `C(157, 26); `C(158, 101); `C(159, 241); `C(160, 77);
    `C(161, 217); `C(162, 166); `C(163, 50); `C(164, 88); `C(165, 204);
    `C(166, 179); `C(167, 39); `C(168, 103); `C(169, 243); `C(170, 140);
    `C(171, 24); `C(172, 114); `C(173, 230); `C(174, 153); `C(175, 13);
    `C(176, 25); `C(177, 141); `C(178, 242); `C(179, 102); `C(180, 12);
    `C(181, 152); `C(182, 231); `C(183, 115); `C(184, 51); `C(185, 167);
    `C(186, 216); `C(187, 76); `C(188, 38); `C(189, 178); `C(190, 205);
    `C(191, 89); `C(192, 118); `C(193, 226); `C(194, 157); `C(195, 9);
    `C(196, 99); `C(197, 247); `C(198, 136); `C(199, 28); `C(200, 92);
    `C(201, 200); `C(202, 183); `C(203, 35); `C(204, 73); `C(205, 221);
    `C(206, 162); `C(207, 54); `C(208, 34); `C(209, 182); `C(210, 201);
    `C(211, 93); `C(212, 55); `C(213, 163); `C(214, 220); `C(215, 72);
    `C(216, 8); `C(217, 156); `C(218, 227); `C(219, 119); `C(220, 29);
    `C(221, 137); `C(222, 246); `C(223, 98); `C(224, 222); `C(225, 74);
    `C(226, 53); `C(227, 161); `C(228, 203); `C(229, 95); `C(230, 32);
    `C(231, 180); `C(232, 244); `C(233, 96); `C(234, 31); `C(235, 139);
    `C(236, 225); `C(237, 117); `C(238, 10); `C(239, 158); `C(240, 138);
    `C(241, 30); `C(242, 97); `C(243, 245); `C(244, 159); `C(245, 11);
    `C(246, 116); `C(247, 224); `C(248, 160); `C(249, 52); `C(250, 75);
    `C(251, 223); `C(252, 181); `C(253, 33); `C(254, 94); `C(255, 202);
    assign out = tab[in];
  end if (constVal == 8'h20) begin
    `C(0, 0); `C(1, 32); `C(2, 64); `C(3, 96); `C(4, 128); `C(5, 160);
    `C(6, 192); `C(7, 224); `C(8, 195); `C(9, 227); `C(10, 131); `C(11, 163);
    `C(12, 67); `C(13, 99); `C(14, 3); `C(15, 35); `C(16, 69); `C(17, 101);
    `C(18, 5); `C(19, 37); `C(20, 197); `C(21, 229); `C(22, 133); `C(23, 165);
    `C(24, 134); `C(25, 166); `C(26, 198); `C(27, 230); `C(28, 6); `C(29, 38);
    `C(30, 70); `C(31, 102); `C(32, 138); `C(33, 170); `C(34, 202);
    `C(35, 234); `C(36, 10); `C(37, 42); `C(38, 74); `C(39, 106); `C(40, 73);
    `C(41, 105); `C(42, 9); `C(43, 41); `C(44, 201); `C(45, 233); `C(46, 137);
    `C(47, 169); `C(48, 207); `C(49, 239); `C(50, 143); `C(51, 175);
    `C(52, 79); `C(53, 111); `C(54, 15); `C(55, 47); `C(56, 12); `C(57, 44);
    `C(58, 76); `C(59, 108); `C(60, 140); `C(61, 172); `C(62, 204);
    `C(63, 236); `C(64, 215); `C(65, 247); `C(66, 151); `C(67, 183);
    `C(68, 87); `C(69, 119); `C(70, 23); `C(71, 55); `C(72, 20); `C(73, 52);
    `C(74, 84); `C(75, 116); `C(76, 148); `C(77, 180); `C(78, 212);
    `C(79, 244); `C(80, 146); `C(81, 178); `C(82, 210); `C(83, 242);
    `C(84, 18); `C(85, 50); `C(86, 82); `C(87, 114); `C(88, 81); `C(89, 113);
    `C(90, 17); `C(91, 49); `C(92, 209); `C(93, 241); `C(94, 145);
    `C(95, 177); `C(96, 93); `C(97, 125); `C(98, 29); `C(99, 61); `C(100, 221);
    `C(101, 253); `C(102, 157); `C(103, 189); `C(104, 158); `C(105, 190);
    `C(106, 222); `C(107, 254); `C(108, 30); `C(109, 62); `C(110, 94);
    `C(111, 126); `C(112, 24); `C(113, 56); `C(114, 88); `C(115, 120);
    `C(116, 152); `C(117, 184); `C(118, 216); `C(119, 248); `C(120, 219);
    `C(121, 251); `C(122, 155); `C(123, 187); `C(124, 91); `C(125, 123);
    `C(126, 27); `C(127, 59); `C(128, 109); `C(129, 77); `C(130, 45);
    `C(131, 13); `C(132, 237); `C(133, 205); `C(134, 173); `C(135, 141);
    `C(136, 174); `C(137, 142); `C(138, 238); `C(139, 206); `C(140, 46);
    `C(141, 14); `C(142, 110); `C(143, 78); `C(144, 40); `C(145, 8);
    `C(146, 104); `C(147, 72); `C(148, 168); `C(149, 136); `C(150, 232);
    `C(151, 200); `C(152, 235); `C(153, 203); `C(154, 171); `C(155, 139);
    `C(156, 107); `C(157, 75); `C(158, 43); `C(159, 11); `C(160, 231);
    `C(161, 199); `C(162, 167); `C(163, 135); `C(164, 103); `C(165, 71);
    `C(166, 39); `C(167, 7); `C(168, 36); `C(169, 4); `C(170, 100);
    `C(171, 68); `C(172, 164); `C(173, 132); `C(174, 228); `C(175, 196);
    `C(176, 162); `C(177, 130); `C(178, 226); `C(179, 194); `C(180, 34);
    `C(181, 2); `C(182, 98); `C(183, 66); `C(184, 97); `C(185, 65);
    `C(186, 33); `C(187, 1); `C(188, 225); `C(189, 193); `C(190, 161);
    `C(191, 129); `C(192, 186); `C(193, 154); `C(194, 250); `C(195, 218);
    `C(196, 58); `C(197, 26); `C(198, 122); `C(199, 90); `C(200, 121);
    `C(201, 89); `C(202, 57); `C(203, 25); `C(204, 249); `C(205, 217);
    `C(206, 185); `C(207, 153); `C(208, 255); `C(209, 223); `C(210, 191);
    `C(211, 159); `C(212, 127); `C(213, 95); `C(214, 63); `C(215, 31);
    `C(216, 60); `C(217, 28); `C(218, 124); `C(219, 92); `C(220, 188);
    `C(221, 156); `C(222, 252); `C(223, 220); `C(224, 48); `C(225, 16);
    `C(226, 112); `C(227, 80); `C(228, 176); `C(229, 144); `C(230, 240);
    `C(231, 208); `C(232, 243); `C(233, 211); `C(234, 179); `C(235, 147);
    `C(236, 115); `C(237, 83); `C(238, 51); `C(239, 19); `C(240, 117);
    `C(241, 85); `C(242, 53); `C(243, 21); `C(244, 245); `C(245, 213);
    `C(246, 181); `C(247, 149); `C(248, 182); `C(249, 150); `C(250, 246);
    `C(251, 214); `C(252, 54); `C(253, 22); `C(254, 118); `C(255, 86);
    assign out = tab[in];
  end if (constVal == 8'h85) begin
    `C(0, 0); `C(1, 133); `C(2, 201); `C(3, 76); `C(4, 81); `C(5, 212);
    `C(6, 152); `C(7, 29); `C(8, 162); `C(9, 39); `C(10, 107); `C(11, 238);
    `C(12, 243); `C(13, 118); `C(14, 58); `C(15, 191); `C(16, 135); `C(17, 2);
    `C(18, 78); `C(19, 203); `C(20, 214); `C(21, 83); `C(22, 31); `C(23, 154);
    `C(24, 37); `C(25, 160); `C(26, 236); `C(27, 105); `C(28, 116);
    `C(29, 241); `C(30, 189); `C(31, 56); `C(32, 205); `C(33, 72); `C(34, 4);
    `C(35, 129); `C(36, 156); `C(37, 25); `C(38, 85); `C(39, 208); `C(40, 111);
    `C(41, 234); `C(42, 166); `C(43, 35); `C(44, 62); `C(45, 187); `C(46, 247);
    `C(47, 114); `C(48, 74); `C(49, 207); `C(50, 131); `C(51, 6); `C(52, 27);
    `C(53, 158); `C(54, 210); `C(55, 87); `C(56, 232); `C(57, 109); `C(58, 33);
    `C(59, 164); `C(60, 185); `C(61, 60); `C(62, 112); `C(63, 245); `C(64, 89);
    `C(65, 220); `C(66, 144); `C(67, 21); `C(68, 8); `C(69, 141); `C(70, 193);
    `C(71, 68); `C(72, 251); `C(73, 126); `C(74, 50); `C(75, 183); `C(76, 170);
    `C(77, 47); `C(78, 99); `C(79, 230); `C(80, 222); `C(81, 91); `C(82, 23);
    `C(83, 146); `C(84, 143); `C(85, 10); `C(86, 70); `C(87, 195); `C(88, 124);
    `C(89, 249); `C(90, 181); `C(91, 48); `C(92, 45); `C(93, 168); `C(94, 228);
    `C(95, 97); `C(96, 148); `C(97, 17); `C(98, 93); `C(99, 216); `C(100, 197);
    `C(101, 64); `C(102, 12); `C(103, 137); `C(104, 54); `C(105, 179);
    `C(106, 255); `C(107, 122); `C(108, 103); `C(109, 226); `C(110, 174);
    `C(111, 43); `C(112, 19); `C(113, 150); `C(114, 218); `C(115, 95);
    `C(116, 66); `C(117, 199); `C(118, 139); `C(119, 14); `C(120, 177);
    `C(121, 52); `C(122, 120); `C(123, 253); `C(124, 224); `C(125, 101);
    `C(126, 41); `C(127, 172); `C(128, 178); `C(129, 55); `C(130, 123);
    `C(131, 254); `C(132, 227); `C(133, 102); `C(134, 42); `C(135, 175);
    `C(136, 16); `C(137, 149); `C(138, 217); `C(139, 92); `C(140, 65);
    `C(141, 196); `C(142, 136); `C(143, 13); `C(144, 53); `C(145, 176);
    `C(146, 252); `C(147, 121); `C(148, 100); `C(149, 225); `C(150, 173);
    `C(151, 40); `C(152, 151); `C(153, 18); `C(154, 94); `C(155, 219);
    `C(156, 198); `C(157, 67); `C(158, 15); `C(159, 138); `C(160, 127);
    `C(161, 250); `C(162, 182); `C(163, 51); `C(164, 46); `C(165, 171);
    `C(166, 231); `C(167, 98); `C(168, 221); `C(169, 88); `C(170, 20);
    `C(171, 145); `C(172, 140); `C(173, 9); `C(174, 69); `C(175, 192);
    `C(176, 248); `C(177, 125); `C(178, 49); `C(179, 180); `C(180, 169);
    `C(181, 44); `C(182, 96); `C(183, 229); `C(184, 90); `C(185, 223);
    `C(186, 147); `C(187, 22); `C(188, 11); `C(189, 142); `C(190, 194);
    `C(191, 71); `C(192, 235); `C(193, 110); `C(194, 34); `C(195, 167);
    `C(196, 186); `C(197, 63); `C(198, 115); `C(199, 246); `C(200, 73);
    `C(201, 204); `C(202, 128); `C(203, 5); `C(204, 24); `C(205, 157);
    `C(206, 209); `C(207, 84); `C(208, 108); `C(209, 233); `C(210, 165);
    `C(211, 32); `C(212, 61); `C(213, 184); `C(214, 244); `C(215, 113);
    `C(216, 206); `C(217, 75); `C(218, 7); `C(219, 130); `C(220, 159);
    `C(221, 26); `C(222, 86); `C(223, 211); `C(224, 38); `C(225, 163);
    `C(226, 239); `C(227, 106); `C(228, 119); `C(229, 242); `C(230, 190);
    `C(231, 59); `C(232, 132); `C(233, 1); `C(234, 77); `C(235, 200);
    `C(236, 213); `C(237, 80); `C(238, 28); `C(239, 153); `C(240, 161);
    `C(241, 36); `C(242, 104); `C(243, 237); `C(244, 240); `C(245, 117);
    `C(246, 57); `C(247, 188); `C(248, 3); `C(249, 134); `C(250, 202);
    `C(251, 79); `C(252, 82); `C(253, 215); `C(254, 155); `C(255, 30);
    assign out = tab[in];
  end if (constVal == 8'h10) begin
    `C(0, 0); `C(1, 16); `C(2, 32); `C(3, 48); `C(4, 64); `C(5, 80); `C(6, 96);
    `C(7, 112); `C(8, 128); `C(9, 144); `C(10, 160); `C(11, 176); `C(12, 192);
    `C(13, 208); `C(14, 224); `C(15, 240); `C(16, 195); `C(17, 211);
    `C(18, 227); `C(19, 243); `C(20, 131); `C(21, 147); `C(22, 163);
    `C(23, 179); `C(24, 67); `C(25, 83); `C(26, 99); `C(27, 115); `C(28, 3);
    `C(29, 19); `C(30, 35); `C(31, 51); `C(32, 69); `C(33, 85); `C(34, 101);
    `C(35, 117); `C(36, 5); `C(37, 21); `C(38, 37); `C(39, 53); `C(40, 197);
    `C(41, 213); `C(42, 229); `C(43, 245); `C(44, 133); `C(45, 149);
    `C(46, 165); `C(47, 181); `C(48, 134); `C(49, 150); `C(50, 166);
    `C(51, 182); `C(52, 198); `C(53, 214); `C(54, 230); `C(55, 246);
    `C(56, 6); `C(57, 22); `C(58, 38); `C(59, 54); `C(60, 70);
    `C(61, 86); `C(62, 102); `C(63, 118); `C(64, 138); `C(65, 154);
    `C(66, 170); `C(67, 186); `C(68, 202); `C(69, 218); `C(70, 234);
    `C(71, 250); `C(72, 10); `C(73, 26); `C(74, 42); `C(75, 58);
    `C(76, 74); `C(77, 90); `C(78, 106); `C(79, 122); `C(80, 73); `C(81, 89);
    `C(82, 105); `C(83, 121); `C(84, 9); `C(85, 25); `C(86, 41); `C(87, 57);
    `C(88, 201); `C(89, 217); `C(90, 233); `C(91, 249); `C(92, 137);
    `C(93, 153); `C(94, 169); `C(95, 185); `C(96, 207); `C(97, 223);
    `C(98, 239); `C(99, 255); `C(100, 143); `C(101, 159); `C(102, 175);
    `C(103, 191); `C(104, 79); `C(105, 95); `C(106, 111); `C(107, 127);
    `C(108, 15); `C(109, 31); `C(110, 47); `C(111, 63); `C(112, 12);
    `C(113, 28); `C(114, 44); `C(115, 60); `C(116, 76); `C(117, 92);
    `C(118, 108); `C(119, 124); `C(120, 140); `C(121, 156); `C(122, 172);
    `C(123, 188); `C(124, 204); `C(125, 220); `C(126, 236); `C(127, 252);
    `C(128, 215); `C(129, 199); `C(130, 247); `C(131, 231); `C(132, 151);
    `C(133, 135); `C(134, 183); `C(135, 167); `C(136, 87); `C(137, 71);
    `C(138, 119); `C(139, 103); `C(140, 23); `C(141, 7); `C(142, 55);
    `C(143, 39); `C(144, 20); `C(145, 4); `C(146, 52); `C(147, 36);
    `C(148, 84); `C(149, 68); `C(150, 116); `C(151, 100); `C(152, 148);
    `C(153, 132); `C(154, 180); `C(155, 164); `C(156, 212); `C(157, 196);
    `C(158, 244); `C(159, 228); `C(160, 146); `C(161, 130); `C(162, 178);
    `C(163, 162); `C(164, 210); `C(165, 194); `C(166, 242); `C(167, 226);
    `C(168, 18); `C(169, 2); `C(170, 50); `C(171, 34); `C(172, 82);
    `C(173, 66); `C(174, 114); `C(175, 98); `C(176, 81); `C(177, 65);
    `C(178, 113); `C(179, 97); `C(180, 17); `C(181, 1); `C(182, 49);
    `C(183, 33); `C(184, 209); `C(185, 193); `C(186, 241); `C(187, 225);
    `C(188, 145); `C(189, 129); `C(190, 177); `C(191, 161); `C(192, 93);
    `C(193, 77); `C(194, 125); `C(195, 109); `C(196, 29); `C(197, 13);
    `C(198, 61); `C(199, 45); `C(200, 221); `C(201, 205); `C(202, 253);
    `C(203, 237); `C(204, 157); `C(205, 141); `C(206, 189); `C(207, 173);
    `C(208, 158); `C(209, 142); `C(210, 190); `C(211, 174); `C(212, 222);
    `C(213, 206); `C(214, 254); `C(215, 238); `C(216, 30); `C(217, 14);
    `C(218, 62); `C(219, 46); `C(220, 94); `C(221, 78); `C(222, 126);
    `C(223, 110); `C(224, 24); `C(225, 8); `C(226, 56); `C(227, 40);
    `C(228, 88); `C(229, 72); `C(230, 120); `C(231, 104); `C(232, 152);
    `C(233, 136); `C(234, 184); `C(235, 168); `C(236, 216); `C(237, 200);
    `C(238, 248); `C(239, 232); `C(240, 219); `C(241, 203); `C(242, 251);
    `C(243, 235); `C(244, 155); `C(245, 139); `C(246, 187); `C(247, 171);
    `C(248, 91); `C(249, 75); `C(250, 123); `C(251, 107); `C(252, 27);
    `C(253, 11); `C(254, 59); `C(255, 43);
    assign out = tab[in];
  end if (constVal == 8'hC2) begin
    `C(0, 0); `C(1, 194); `C(2, 71); `C(3, 133); `C(4, 142); `C(5, 76);
    `C(6, 201); `C(7, 11); `C(8, 223); `C(9, 29); `C(10, 152); `C(11, 90);
    `C(12, 81); `C(13, 147); `C(14, 22); `C(15, 212); `C(16, 125); `C(17, 191);
    `C(18, 58); `C(19, 248); `C(20, 243); `C(21, 49); `C(22, 180); `C(23, 118);
    `C(24, 162); `C(25, 96); `C(26, 229); `C(27, 39); `C(28, 44); `C(29, 238);
    `C(30, 107); `C(31, 169); `C(32, 250); `C(33, 56); `C(34, 189);
    `C(35, 127); `C(36, 116); `C(37, 182); `C(38, 51); `C(39, 241); `C(40, 37);
    `C(41, 231); `C(42, 98); `C(43, 160); `C(44, 171); `C(45, 105);
    `C(46, 236); `C(47, 46); `C(48, 135); `C(49, 69); `C(50, 192); `C(51, 2);
    `C(52, 9); `C(53, 203); `C(54, 78); `C(55, 140); `C(56, 88); `C(57, 154);
    `C(58, 31); `C(59, 221); `C(60, 214); `C(61, 20); `C(62, 145); `C(63, 83);
    `C(64, 55); `C(65, 245); `C(66, 112); `C(67, 178); `C(68, 185);
    `C(69, 123); `C(70, 254); `C(71, 60); `C(72, 232); `C(73, 42); `C(74, 175);
    `C(75, 109); `C(76, 102); `C(77, 164); `C(78, 33); `C(79, 227); `C(80, 74);
    `C(81, 136); `C(82, 13); `C(83, 207); `C(84, 196); `C(85, 6); `C(86, 131);
    `C(87, 65); `C(88, 149); `C(89, 87); `C(90, 210); `C(91, 16); `C(92, 27);
    `C(93, 217); `C(94, 92); `C(95, 158); `C(96, 205); `C(97, 15); `C(98, 138);
    `C(99, 72); `C(100, 67); `C(101, 129); `C(102, 4); `C(103, 198);
    `C(104, 18); `C(105, 208); `C(106, 85); `C(107, 151); `C(108, 156);
    `C(109, 94); `C(110, 219); `C(111, 25); `C(112, 176); `C(113, 114);
    `C(114, 247); `C(115, 53); `C(116, 62); `C(117, 252); `C(118, 121);
    `C(119, 187); `C(120, 111); `C(121, 173); `C(122, 40); `C(123, 234);
    `C(124, 225); `C(125, 35); `C(126, 166); `C(127, 100); `C(128, 110);
    `C(129, 172); `C(130, 41); `C(131, 235); `C(132, 224); `C(133, 34);
    `C(134, 167); `C(135, 101); `C(136, 177); `C(137, 115); `C(138, 246);
    `C(139, 52); `C(140, 63); `C(141, 253); `C(142, 120); `C(143, 186);
    `C(144, 19); `C(145, 209); `C(146, 84); `C(147, 150); `C(148, 157);
    `C(149, 95); `C(150, 218); `C(151, 24); `C(152, 204); `C(153, 14);
    `C(154, 139); `C(155, 73); `C(156, 66); `C(157, 128); `C(158, 5);
    `C(159, 199); `C(160, 148); `C(161, 86); `C(162, 211); `C(163, 17);
    `C(164, 26); `C(165, 216); `C(166, 93); `C(167, 159); `C(168, 75);
    `C(169, 137); `C(170, 12); `C(171, 206); `C(172, 197); `C(173, 7);
    `C(174, 130); `C(175, 64); `C(176, 233); `C(177, 43); `C(178, 174);
    `C(179, 108); `C(180, 103); `C(181, 165); `C(182, 32); `C(183, 226);
    `C(184, 54); `C(185, 244); `C(186, 113); `C(187, 179); `C(188, 184);
    `C(189, 122); `C(190, 255); `C(191, 61); `C(192, 89); `C(193, 155);
    `C(194, 30); `C(195, 220); `C(196, 215); `C(197, 21); `C(198, 144);
    `C(199, 82); `C(200, 134); `C(201, 68); `C(202, 193); `C(203, 3);
    `C(204, 8); `C(205, 202); `C(206, 79); `C(207, 141); `C(208, 36);
    `C(209, 230); `C(210, 99); `C(211, 161); `C(212, 170); `C(213, 104);
    `C(214, 237); `C(215, 47); `C(216, 251); `C(217, 57); `C(218, 188);
    `C(219, 126); `C(220, 117); `C(221, 183); `C(222, 50); `C(223, 240);
    `C(224, 163); `C(225, 97); `C(226, 228); `C(227, 38); `C(228, 45);
    `C(229, 239); `C(230, 106); `C(231, 168); `C(232, 124); `C(233, 190);
    `C(234, 59); `C(235, 249); `C(236, 242); `C(237, 48); `C(238, 181);
    `C(239, 119); `C(240, 222); `C(241, 28); `C(242, 153); `C(243, 91);
    `C(244, 80); `C(245, 146); `C(246, 23); `C(247, 213); `C(248, 1);
    `C(249, 195); `C(250, 70); `C(251, 132); `C(252, 143); `C(253, 77);
    `C(254, 200); `C(255, 10);
    assign out = tab[in];
  end if (constVal == 8'hC0) begin
    `C(0, 0); `C(1, 192); `C(2, 67); `C(3, 131); `C(4, 134); `C(5, 70);
    `C(6, 197); `C(7, 5); `C(8, 207); `C(9, 15); `C(10, 140); `C(11, 76);
    `C(12, 73); `C(13, 137); `C(14, 10); `C(15, 202); `C(16, 93); `C(17, 157);
    `C(18, 30); `C(19, 222); `C(20, 219); `C(21, 27); `C(22, 152); `C(23, 88);
    `C(24, 146); `C(25, 82); `C(26, 209); `C(27, 17); `C(28, 20); `C(29, 212);
    `C(30, 87); `C(31, 151); `C(32, 186); `C(33, 122); `C(34, 249); `C(35, 57);
    `C(36, 60); `C(37, 252); `C(38, 127); `C(39, 191); `C(40, 117);
    `C(41, 181); `C(42, 54); `C(43, 246); `C(44, 243); `C(45, 51); `C(46, 176);
    `C(47, 112); `C(48, 231); `C(49, 39); `C(50, 164); `C(51, 100); `C(52, 97);
    `C(53, 161); `C(54, 34); `C(55, 226); `C(56, 40); `C(57, 232); `C(58, 107);
    `C(59, 171); `C(60, 174); `C(61, 110); `C(62, 237); `C(63, 45);
    `C(64, 183); `C(65, 119); `C(66, 244); `C(67, 52); `C(68, 49); `C(69, 241);
    `C(70, 114); `C(71, 178); `C(72, 120); `C(73, 184);
    `C(74, 59); `C(75, 251); `C(76, 254); `C(77, 62); `C(78, 189); `C(79, 125);
    `C(80, 234); `C(81, 42); `C(82, 169); `C(83, 105);
    `C(84, 108); `C(85, 172); `C(86, 47); `C(87, 239); `C(88, 37); `C(89, 229);
    `C(90, 102); `C(91, 166); `C(92, 163); `C(93, 99); `C(94, 224); `C(95, 32);
    `C(96, 13); `C(97, 205); `C(98, 78); `C(99, 142); `C(100, 139);
    `C(101, 75); `C(102, 200); `C(103, 8); `C(104, 194); `C(105, 2);
    `C(106, 129); `C(107, 65); `C(108, 68); `C(109, 132); `C(110, 7);
    `C(111, 199); `C(112, 80); `C(113, 144); `C(114, 19); `C(115, 211);
    `C(116, 214); `C(117, 22); `C(118, 149); `C(119, 85); `C(120, 159);
    `C(121, 95); `C(122, 220); `C(123, 28); `C(124, 25); `C(125, 217);
    `C(126, 90); `C(127, 154); `C(128, 173); `C(129, 109); `C(130, 238);
    `C(131, 46); `C(132, 43); `C(133, 235); `C(134, 104); `C(135, 168);
    `C(136, 98); `C(137, 162); `C(138, 33); `C(139, 225); `C(140, 228);
    `C(141, 36); `C(142, 167); `C(143, 103); `C(144, 240); `C(145, 48);
    `C(146, 179); `C(147, 115); `C(148, 118); `C(149, 182); `C(150, 53);
    `C(151, 245); `C(152, 63); `C(153, 255); `C(154, 124); `C(155, 188);
    `C(156, 185); `C(157, 121); `C(158, 250); `C(159, 58); `C(160, 23);
    `C(161, 215); `C(162, 84); `C(163, 148); `C(164, 145); `C(165, 81);
    `C(166, 210); `C(167, 18); `C(168, 216); `C(169, 24); `C(170, 155);
    `C(171, 91); `C(172, 94); `C(173, 158); `C(174, 29); `C(175, 221);
    `C(176, 74); `C(177, 138); `C(178, 9); `C(179, 201); `C(180, 204);
    `C(181, 12); `C(182, 143); `C(183, 79); `C(184, 133); `C(185, 69);
    `C(186, 198); `C(187, 6); `C(188, 3); `C(189, 195); `C(190, 64);
    `C(191, 128); `C(192, 26); `C(193, 218); `C(194, 89); `C(195, 153);
    `C(196, 156); `C(197, 92); `C(198, 223); `C(199, 31); `C(200, 213);
    `C(201, 21); `C(202, 150); `C(203, 86); `C(204, 83); `C(205, 147);
    `C(206, 16); `C(207, 208); `C(208, 71); `C(209, 135); `C(210, 4);
    `C(211, 196); `C(212, 193); `C(213, 1); `C(214, 130); `C(215, 66);
    `C(216, 136); `C(217, 72); `C(218, 203); `C(219, 11); `C(220, 14);
    `C(221, 206); `C(222, 77); `C(223, 141); `C(224, 160); `C(225, 96);
    `C(226, 227); `C(227, 35); `C(228, 38); `C(229, 230); `C(230, 101);
    `C(231, 165); `C(232, 111); `C(233, 175); `C(234, 44); `C(235, 236);
    `C(236, 233); `C(237, 41); `C(238, 170); `C(239, 106); `C(240, 253);
    `C(241, 61); `C(242, 190); `C(243, 126); `C(244, 123); `C(245, 187);
    `C(246, 56); `C(247, 248); `C(248, 50); `C(249, 242); `C(250, 113);
    `C(251, 177); `C(252, 180); `C(253, 116); `C(254, 247); `C(255, 55);
    assign out = tab[in];
  end if (constVal == 8'hFB) begin
    `C(0, 0); `C(1, 251); `C(2, 53); `C(3, 206); `C(4, 106); `C(5, 145);
    `C(6, 95); `C(7, 164); `C(8, 212); `C(9, 47); `C(10, 225); `C(11, 26);
    `C(12, 190); `C(13, 69); `C(14, 139); `C(15, 112); `C(16, 107);
    `C(17, 144); `C(18, 94); `C(19, 165); `C(20, 1); `C(21, 250); `C(22, 52);
    `C(23, 207); `C(24, 191); `C(25, 68); `C(26, 138); `C(27, 113);
    `C(28, 213); `C(29, 46); `C(30, 224); `C(31, 27); `C(32, 214); `C(33, 45);
    `C(34, 227); `C(35, 24); `C(36, 188); `C(37, 71); `C(38, 137); `C(39, 114);
    `C(40, 2); `C(41, 249); `C(42, 55); `C(43, 204); `C(44, 104); `C(45, 147);
    `C(46, 93); `C(47, 166); `C(48, 189); `C(49, 70); `C(50, 136); `C(51, 115);
    `C(52, 215); `C(53, 44); `C(54, 226); `C(55, 25); `C(56, 105); `C(57, 146);
    `C(58, 92); `C(59, 167); `C(60, 3); `C(61, 248); `C(62, 54); `C(63, 205);
    `C(64, 111); `C(65, 148); `C(66, 90); `C(67, 161); `C(68, 5); `C(69, 254);
    `C(70, 48); `C(71, 203); `C(72, 187); `C(73, 64); `C(74, 142); `C(75, 117);
    `C(76, 209); `C(77, 42); `C(78, 228); `C(79, 31); `C(80, 4); `C(81, 255);
    `C(82, 49); `C(83, 202); `C(84, 110); `C(85, 149); `C(86, 91); `C(87, 160);
    `C(88, 208); `C(89, 43); `C(90, 229); `C(91, 30); `C(92, 186); `C(93, 65);
    `C(94, 143); `C(95, 116); `C(96, 185); `C(97, 66); `C(98, 140);
    `C(99, 119); `C(100, 211); `C(101, 40); `C(102, 230); `C(103, 29);
    `C(104, 109); `C(105, 150); `C(106, 88); `C(107, 163); `C(108, 7);
    `C(109, 252); `C(110, 50); `C(111, 201); `C(112, 210); `C(113, 41);
    `C(114, 231); `C(115, 28); `C(116, 184); `C(117, 67); `C(118, 141);
    `C(119, 118); `C(120, 6); `C(121, 253); `C(122, 51); `C(123, 200);
    `C(124, 108); `C(125, 151); `C(126, 89); `C(127, 162); `C(128, 222);
    `C(129, 37); `C(130, 235); `C(131, 16); `C(132, 180); `C(133, 79);
    `C(134, 129); `C(135, 122); `C(136, 10); `C(137, 241); `C(138, 63);
    `C(139, 196); `C(140, 96); `C(141, 155); `C(142, 85); `C(143, 174);
    `C(144, 181); `C(145, 78); `C(146, 128); `C(147, 123); `C(148, 223);
    `C(149, 36); `C(150, 234); `C(151, 17); `C(152, 97); `C(153, 154);
    `C(154, 84); `C(155, 175); `C(156, 11); `C(157, 240); `C(158, 62);
    `C(159, 197); `C(160, 8); `C(161, 243); `C(162, 61); `C(163, 198);
    `C(164, 98); `C(165, 153); `C(166, 87); `C(167, 172); `C(168, 220);
    `C(169, 39); `C(170, 233); `C(171, 18); `C(172, 182); `C(173, 77);
    `C(174, 131); `C(175, 120); `C(176, 99); `C(177, 152); `C(178, 86);
    `C(179, 173); `C(180, 9); `C(181, 242); `C(182, 60); `C(183, 199);
    `C(184, 183); `C(185, 76); `C(186, 130); `C(187, 121); `C(188, 221);
    `C(189, 38); `C(190, 232); `C(191, 19); `C(192, 177); `C(193, 74);
    `C(194, 132); `C(195, 127); `C(196, 219); `C(197, 32); `C(198, 238);
    `C(199, 21); `C(200, 101); `C(201, 158); `C(202, 80); `C(203, 171);
    `C(204, 15); `C(205, 244); `C(206, 58); `C(207, 193); `C(208, 218);
    `C(209, 33); `C(210, 239); `C(211, 20); `C(212, 176); `C(213, 75);
    `C(214, 133); `C(215, 126); `C(216, 14); `C(217, 245); `C(218, 59);
    `C(219, 192); `C(220, 100); `C(221, 159); `C(222, 81); `C(223, 170);
    `C(224, 103); `C(225, 156); `C(226, 82); `C(227, 169); `C(228, 13);
    `C(229, 246); `C(230, 56); `C(231, 195); `C(232, 179); `C(233, 72);
    `C(234, 134); `C(235, 125); `C(236, 217); `C(237, 34); `C(238, 236);
    `C(239, 23); `C(240, 12); `C(241, 247); `C(242, 57); `C(243, 194);
    `C(244, 102); `C(245, 157); `C(246, 83); `C(247, 168); `C(248, 216);
    `C(249, 35); `C(250, 237); `C(251, 22); `C(252, 178); `C(253, 73);
    `C(254, 135); `C(255, 124);
    assign out = tab[in];
  end

endmodule
