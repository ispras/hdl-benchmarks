`timescale 1 ps / 1 ps

module lcell (gnd, marker_bep_outwire);
  input gnd;
  output marker_bep_outwire;
endmodule
