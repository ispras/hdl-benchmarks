module RAMB4_S4_S4 (CLKA, CLKB, RSTB, RSTA, DOA, ADDRA, DIA, ENA, WEA, DOB, ADDRB, DIB, ENB, WEB);
  input CLKA;
  input CLKB;
  input RSTB;
  input RSTA;
  output DOA;
  output ADDRA;
  input DIA;
  output ENA;
  input WEA;
  output DOB;
  output ADDRB;
  output DIB;
  output ENB;
  output WEB;
endmodule