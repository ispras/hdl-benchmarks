module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 ;
output n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
 n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
 n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
 n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
 n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
 n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
 n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
 n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
 n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
 n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
 n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
 n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
 n220 , n221 , n222 , n223 , n224 , n225 , n226 ;
wire n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , 
 n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , 
 n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , 
 n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , 
 n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , 
 n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , 
 n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , 
 n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , 
 n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , 
 n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , 
 n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , 
 n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , 
 n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , 
 n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , 
 n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , 
 n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , 
 n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , 
 n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , 
 n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , 
 n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , 
 n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , 
 n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , 
 n675 , n676 , n677 , n678 , n679 , n680 , n70358 , n70359 , n70360 , n70361 , 
 n70362 , n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , 
 n70372 , n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , 
 n70382 , n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , 
 n70392 , n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , 
 n70402 , n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , 
 n70412 , n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , 
 n70422 , n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , 
 n70432 , n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , 
 n70442 , n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , 
 n70452 , n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , 
 n70462 , n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , 
 n70472 , n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , 
 n70482 , n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , 
 n70492 , n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , 
 n70502 , n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , 
 n70512 , n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , 
 n70522 , n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , 
 n70532 , n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , 
 n70542 , n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , 
 n70552 , n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , 
 n70562 , n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , 
 n70572 , n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , 
 n70582 , n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , 
 n70592 , n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , 
 n70602 , n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , 
 n70612 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , 
 n70622 , n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , 
 n70632 , n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , 
 n70642 , n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , 
 n70652 , n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , 
 n70662 , n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , 
 n70672 , n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , 
 n70682 , n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , 
 n70692 , n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , 
 n70702 , n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , 
 n70712 , n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , 
 n682 , n70723 , n684 , n70725 , n686 , n687 , n70728 , n689 , n690 , n691 , 
 n692 , n693 , n70734 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , 
 n70742 , n703 , n70744 , n705 , n706 , n707 , n708 , n709 , n70750 , n711 , 
 n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , 
 n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , 
 n732 , n733 , n734 , n735 , n736 , n70777 , n741 , n70779 , n743 , n70781 , 
 n745 , n70783 , n747 , n748 , n70786 , n750 , n751 , n752 , n753 , n754 , 
 n758 , n70793 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n770 , 
 n70802 , n772 , n70804 , n774 , n775 , n776 , n777 , n778 , n782 , n70811 , 
 n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , 
 n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , 
 n804 , n805 , n806 , n807 , n808 , n809 , n70838 , n814 , n815 , n70841 , 
 n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n70851 , 
 n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , 
 n837 , n70863 , n839 , n843 , n70866 , n845 , n846 , n847 , n848 , n849 , 
 n850 , n851 , n852 , n853 , n70876 , n855 , n856 , n857 , n858 , n859 , 
 n860 , n861 , n862 , n863 , n864 , n70887 , n869 , n870 , n871 , n872 , 
 n873 , n874 , n70894 , n876 , n877 , n878 , n879 , n880 , n70900 , n882 , 
 n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , 
 n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , 
 n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n70930 , n912 , 
 n913 , n914 , n915 , n916 , n917 , n918 , n919 , n70939 , n921 , n922 , 
 n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , 
 n933 , n937 , n70954 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , 
 n946 , n947 , n948 , n949 , n950 , n951 , n70968 , n956 , n957 , n958 , 
 n959 , n960 , n961 , n962 , n963 , n70977 , n965 , n966 , n967 , n968 , 
 n969 , n970 , n971 , n972 , n973 , n70987 , n975 , n976 , n977 , n978 , 
 n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
 n989 , n990 , n991 , n992 , n993 , n71007 , n995 , n996 , n997 , n998 , 
 n999 , n1000 , n1001 , n1002 , n1003 , n1007 , n71018 , n1009 , n1010 , n1011 , 
 n1012 , n71023 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , 
 n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n71041 , 
 n1035 , n1036 , n71044 , n1038 , n1039 , n1040 , n1041 , n1042 , n71050 , n1044 , 
 n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , 
 n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , 
 n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , 
 n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , 
 n1085 , n1086 , n71094 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , 
 n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n71110 , n1104 , 
 n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , 
 n1115 , n1116 , n1117 , n1121 , n71126 , n1123 , n1124 , n1125 , n1126 , n1127 , 
 n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n71141 , 
 n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
 n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
 n1161 , n1162 , n71164 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
 n1171 , n1172 , n71174 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
 n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n71190 , n1190 , 
 n1191 , n1192 , n1193 , n71195 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
 n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1211 , n71210 , n1213 , 
 n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , 
 n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , 
 n1234 , n1235 , n1236 , n1237 , n71236 , n1242 , n1243 , n1244 , n1245 , n1246 , 
 n1247 , n1248 , n1249 , n71245 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , 
 n1257 , n1258 , n1259 , n71255 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , 
 n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , 
 n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , 
 n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , 
 n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n71299 , n1305 , n1306 , 
 n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , 
 n1317 , n1321 , n71314 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
 n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
 n1340 , n1341 , n71334 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
 n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
 n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n71360 , n1372 , 
 n1373 , n1374 , n1375 , n1376 , n1377 , n71367 , n1379 , n1380 , n1381 , n1382 , 
 n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , 
 n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , 
 n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n71398 , n1410 , n1411 , n1412 , 
 n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , 
 n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , 
 n1433 , n71423 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , 
 n1443 , n71433 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , 
 n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , 
 n1463 , n1467 , n71454 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , 
 n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , 
 n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n71480 , n1498 , 
 n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n71491 , 
 n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , 
 n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , 
 n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , 
 n71522 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , 
 n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , 
 n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , 
 n1569 , n71553 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , 
 n1579 , n1580 , n1581 , n1582 , n1583 , n71567 , n1585 , n1586 , n1587 , n1588 , 
 n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , 
 n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , 
 n1609 , n1610 , n1611 , n1612 , n1616 , n71597 , n1618 , n1619 , n1620 , n1621 , 
 n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , 
 n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n71621 , 
 n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , 
 n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , 
 n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n71648 , n1672 , n1673 , n1674 , 
 n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , 
 n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , 
 n1695 , n71673 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , 
 n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n71690 , n1714 , 
 n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n71699 , n1723 , n1724 , 
 n1725 , n1726 , n1730 , n71705 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , 
 n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , 
 n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , 
 n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , 
 n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , 
 n1778 , n1779 , n71754 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n71761 , 
 n1791 , n1792 , n1793 , n1794 , n1795 , n71767 , n1797 , n1798 , n1799 , n1800 , 
 n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
 n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
 n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
 n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
 n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
 n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
 n1861 , n1862 , n1863 , n1864 , n1865 , n71837 , n1867 , n1868 , n1869 , n1870 , 
 n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
 n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n71861 , 
 n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
 n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
 n1911 , n1912 , n1913 , n1917 , n71886 , n1919 , n1920 , n1921 , n1922 , n1923 , 
 n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , 
 n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , 
 n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n71918 , n1954 , n1955 , n1956 , 
 n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , 
 n1967 , n1968 , n71934 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , 
 n1977 , n1978 , n71944 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , 
 n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , 
 n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , 
 n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , 
 n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , 
 n2027 , n2028 , n2029 , n2030 , n2031 , n71997 , n2033 , n2034 , n2035 , n2036 , 
 n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , 
 n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , 
 n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , 
 n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , 
 n2077 , n2081 , n72044 , n2083 , n2084 , n2085 , n2086 , n72049 , n2088 , n2089 , 
 n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
 n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
 n2110 , n2111 , n72074 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , 
 n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , 
 n2133 , n72093 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , 
 n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , 
 n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , 
 n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , 
 n2173 , n72133 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , 
 n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , 
 n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , 
 n2203 , n2204 , n2205 , n2206 , n2207 , n72167 , n2209 , n2210 , n2211 , n2212 , 
 n2213 , n2217 , n72174 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , 
 n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , 
 n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n72199 , n2244 , n2245 , 
 n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , 
 n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , 
 n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , 
 n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , 
 n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , 
 n2296 , n2297 , n2298 , n2299 , n2300 , n72257 , n2305 , n2306 , n2307 , n2308 , 
 n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , 
 n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , 
 n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , 
 n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , 
 n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
 n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
 n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
 n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n72340 , n2388 , 
 n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
 n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , 
 n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , 
 n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , 
 n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , 
 n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , 
 n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , 
 n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n72420 , n2471 , 
 n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , 
 n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , 
 n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , 
 n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , 
 n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , 
 n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , 
 n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , 
 n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , 
 n2552 , n2553 , n2554 , n72505 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , 
 n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , 
 n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , 
 n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , 
 n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , 
 n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , 
 n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , 
 n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , 
 n72582 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , 
 n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , 
 n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , 
 n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , 
 n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , 
 n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , 
 n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , 
 n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , 
 n2715 , n2716 , n2717 , n2718 , n72666 , n2720 , n2721 , n2722 , n2723 , n2724 , 
 n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , 
 n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , 
 n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , 
 n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , 
 n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , 
 n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , 
 n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , 
 n2795 , n2796 , n2797 , n72745 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , 
 n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , 
 n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , 
 n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , 
 n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , 
 n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , 
 n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , 
 n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , 
 n2878 , n2879 , n2880 , n2881 , n72826 , n2883 , n2884 , n2885 , n2886 , n2887 , 
 n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , 
 n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , 
 n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , 
 n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , 
 n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , 
 n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , 
 n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n72901 , 
 n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
 n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
 n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
 n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
 n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
 n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
 n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
 n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n72978 , n3038 , n3039 , n3040 , 
 n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
 n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
 n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
 n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
 n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
 n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
 n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n73049 , n3112 , n3113 , 
 n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , 
 n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , 
 n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , 
 n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , 
 n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , 
 n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , 
 n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n73120 , n3183 , 
 n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , 
 n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , 
 n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , 
 n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , 
 n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , 
 n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , 
 n3244 , n3245 , n3246 , n73185 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , 
 n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , 
 n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , 
 n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , 
 n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , 
 n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , 
 n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , 
 n73252 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , 
 n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , 
 n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , 
 n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , 
 n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , 
 n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , 
 n3377 , n73313 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
 n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
 n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
 n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
 n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
 n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
 n3440 , n3441 , n73374 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
 n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
 n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
 n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
 n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
 n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n73431 , 
 n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
 n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , 
 n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
 n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
 n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
 n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n73488 , n3560 , n3561 , n3562 , 
 n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
 n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
 n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
 n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
 n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n73541 , 
 n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , 
 n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , 
 n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , 
 n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , 
 n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , 
 n73592 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , 
 n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , 
 n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , 
 n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , 
 n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n73640 , n3718 , 
 n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , 
 n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , 
 n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , 
 n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , 
 n3759 , n3760 , n3761 , n3762 , n3763 , n73687 , n3765 , n3766 , n3767 , n3768 , 
 n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , 
 n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , 
 n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , 
 n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n73731 , 
 n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , 
 n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , 
 n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , 
 n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , 
 n73772 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , 
 n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , 
 n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , 
 n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n73810 , n3894 , 
 n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , 
 n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , 
 n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , 
 n3925 , n3926 , n3927 , n3928 , n3929 , n73847 , n3931 , n3932 , n3933 , n3934 , 
 n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , 
 n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , 
 n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n73881 , 
 n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , 
 n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , 
 n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , 
 n73912 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , 
 n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , 
 n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4030 , n4031 , n4032 , 
 n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , 
 n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , 
 n4053 , n4054 , n4055 , n73965 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , 
 n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , 
 n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n73989 , n4084 , n4085 , 
 n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , 
 n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n74010 , n4105 , 
 n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , 
 n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n74028 , n4126 , n74030 , n74031 , 
 n4129 , n74033 , n74034 , n4132 , n74036 , n4134 , n4135 , n4136 , n74040 , n74041 , 
 n4139 , n74043 , n74044 , n4142 , n74046 , n74047 , n4145 , n4146 , n4147 , n74051 , 
 n74052 , n4150 , n74054 , n4152 , n74056 , n4154 , n4155 , n4156 , n4157 , n4158 , 
 n74062 , n4160 , n4161 , n4162 , n4163 , n74067 , n4165 , n74069 , n4167 , n74071 , 
 n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n74078 , n4176 , n4177 , n4178 , 
 n4179 , n4180 , n4181 , n4182 , n4183 , n74087 , n4185 , n74089 , n4187 , n4188 , 
 n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , 
 n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , 
 n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , 
 n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n74129 , n74130 , n4228 , 
 n74132 , n4230 , n74134 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , 
 n4239 , n4240 , n4241 , n74145 , n4243 , n4244 , n4245 , n4246 , n4247 , n74151 , 
 n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , 
 n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , 
 n4269 , n4270 , n4271 , n4272 , n74176 , n74177 , n4275 , n4276 , n4277 , n4278 , 
 n4279 , n74183 , n74184 , n4282 , n74186 , n4284 , n74188 , n4286 , n4287 , n4288 , 
 n4289 , n74193 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
 n4299 , n4300 , n74204 , n74205 , n4303 , n4304 , n4305 , n4306 , n4307 , n74211 , 
 n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
 n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n74230 , n74231 , 
 n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , 
 n4339 , n74243 , n74244 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , 
 n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , 
 n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , 
 n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
 n4379 , n4380 , n4381 , n4382 , n4383 , n74287 , n74288 , n4386 , n74290 , n4388 , 
 n74292 , n4390 , n4391 , n4392 , n4393 , n74297 , n4395 , n4396 , n4397 , n4398 , 
 n4399 , n4400 , n4401 , n4402 , n4403 , n74307 , n4405 , n4406 , n4407 , n4408 , 
 n4409 , n74313 , n4411 , n74315 , n4413 , n74317 , n4415 , n4416 , n4417 , n4418 , 
 n4419 , n74323 , n4421 , n4422 , n4423 , n4424 , n4425 , n74329 , n4427 , n74331 , 
 n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n74338 , n4436 , n4437 , n4438 , 
 n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
 n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
 n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
 n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
 n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
 n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n74400 , n4501 , 
 n74402 , n4503 , n74404 , n4505 , n4506 , n74407 , n4508 , n4509 , n4513 , n74411 , 
 n74412 , n4516 , n4517 , n4518 , n74416 , n74417 , n4521 , n4522 , n4523 , n4524 , 
 n4525 , n74423 , n4527 , n4528 , n4529 , n4530 , n4531 , n74429 , n74430 , n4534 , 
 n4535 , n4536 , n74434 , n74435 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , 
 n4545 , n74443 , n74444 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , 
 n74452 , n74453 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , 
 n4565 , n4566 , n74464 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , 
 n4575 , n4576 , n74474 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , 
 n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n74489 , n74490 , n4594 , 
 n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , 
 n4605 , n4606 , n4607 , n4608 , n74506 , n4610 , n4611 , n4612 , n4613 , n4614 , 
 n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n74521 , 
 n4625 , n4626 , n4627 , n4628 , n4629 , n74527 , n4631 , n4632 , n4633 , n4634 , 
 n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , 
 n4645 , n74543 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , 
 n4655 , n4656 , n74554 , n4661 , n74556 , n4663 , n4664 , n4665 , n74560 , n4670 , 
 n4671 , n4672 , n74564 , n74565 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
 n74572 , n74573 , n4683 , n4684 , n4685 , n4686 , n74578 , n4688 , n4689 , n4690 , 
 n4691 , n4692 , n4693 , n74585 , n74586 , n4696 , n4697 , n4698 , n4699 , n74591 , 
 n74592 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n74599 , n74600 , n4710 , 
 n4711 , n4712 , n4713 , n4714 , n4715 , n74607 , n4717 , n4718 , n4719 , n4720 , 
 n4721 , n4722 , n74614 , n4724 , n4725 , n4726 , n4727 , n4728 , n74620 , n4730 , 
 n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
 n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
 n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
 n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n74659 , n74660 , n4770 , 
 n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n74671 , 
 n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
 n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
 n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n74701 , 
 n4811 , n4812 , n4813 , n4814 , n4815 , n74707 , n4817 , n4818 , n4819 , n4820 , 
 n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n74718 , n4828 , n4829 , n4830 , 
 n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
 n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
 n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n74748 , n4861 , n74750 , n4863 , 
 n4864 , n74753 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n74761 , 
 n4877 , n4878 , n4879 , n74765 , n74766 , n4882 , n4883 , n4884 , n4885 , n4886 , 
 n4887 , n74773 , n74774 , n4890 , n4891 , n4892 , n4893 , n74779 , n4895 , n4896 , 
 n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , 
 n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n74799 , n74800 , n4916 , 
 n4917 , n4918 , n4919 , n4920 , n74806 , n74807 , n4923 , n4924 , n4925 , n4926 , 
 n4927 , n4928 , n74814 , n74815 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , 
 n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , 
 n4947 , n4948 , n74834 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , 
 n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n74849 , n4965 , n4966 , 
 n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n74859 , n4975 , n4976 , 
 n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , 
 n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , 
 n74882 , n74883 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , 
 n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , 
 n5017 , n5018 , n74904 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , 
 n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n74920 , n5036 , 
 n5037 , n5038 , n5039 , n5040 , n74926 , n5042 , n5043 , n5044 , n5045 , n5046 , 
 n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , 
 n5057 , n5058 , n5059 , n5060 , n5061 , n74947 , n5063 , n5064 , n5065 , n5066 , 
 n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , 
 n5077 , n74963 , n5082 , n74965 , n5084 , n5085 , n5086 , n5087 , n74970 , n5089 , 
 n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
 n74982 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n74990 , n74991 , 
 n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n74998 , n74999 , n5121 , n5122 , 
 n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n75009 , n5131 , n5132 , 
 n5133 , n5134 , n5135 , n5136 , n5137 , n75017 , n75018 , n5140 , n5141 , n5142 , 
 n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n75029 , n75030 , n5152 , 
 n5153 , n5154 , n5155 , n5156 , n5157 , n75037 , n75038 , n5160 , n5161 , n5162 , 
 n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n75048 , n5170 , n5171 , n5172 , 
 n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , 
 n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , 
 n5193 , n75073 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
 n5203 , n75083 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
 n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
 n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , 
 n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , 
 n5243 , n5244 , n75124 , n75125 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , 
 n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n75141 , 
 n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , 
 n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , 
 n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , 
 n75172 , n5294 , n5295 , n5296 , n5297 , n5298 , n75178 , n5300 , n5301 , n5302 , 
 n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , 
 n5313 , n5314 , n75194 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , 
 n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , 
 n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , 
 n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n75229 , n5354 , n75231 , 
 n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , 
 n75242 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n75250 , n75251 , 
 n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n75258 , n75259 , n5387 , n5388 , 
 n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n75270 , n5398 , 
 n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
 n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n75290 , n75291 , 
 n5419 , n5420 , n5421 , n5422 , n5423 , n75297 , n75298 , n5426 , n5427 , n5428 , 
 n5429 , n5430 , n5431 , n75305 , n75306 , n5434 , n5435 , n5436 , n5437 , n5438 , 
 n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
 n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
 n5459 , n5460 , n5461 , n75335 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
 n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
 n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n75359 , n5487 , n5488 , 
 n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
 n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
 n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n75390 , n5518 , 
 n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
 n5529 , n5530 , n5531 , n5532 , n75406 , n75407 , n5535 , n5536 , n5537 , n5538 , 
 n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
 n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
 n5559 , n5560 , n5561 , n5562 , n5563 , n75437 , n5565 , n5566 , n5567 , n5568 , 
 n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n75450 , n5578 , 
 n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n75460 , n5588 , 
 n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
 n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
 n5609 , n5610 , n5611 , n5612 , n5613 , n75487 , n5615 , n5616 , n5617 , n5618 , 
 n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
 n5629 , n75503 , n5634 , n75505 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , 
 n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n75521 , 
 n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n75529 , n75530 , n5664 , 
 n5665 , n5666 , n5667 , n5668 , n5669 , n75537 , n75538 , n5672 , n5673 , n5674 , 
 n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , 
 n5685 , n5686 , n75554 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , 
 n5695 , n5696 , n5697 , n75565 , n75566 , n5700 , n5701 , n5702 , n5703 , n5704 , 
 n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , 
 n5715 , n5716 , n5717 , n5718 , n75586 , n75587 , n5721 , n5722 , n5723 , n5724 , 
 n5725 , n5726 , n75594 , n75595 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , 
 n5735 , n5736 , n5737 , n5738 , n75606 , n5740 , n5741 , n5742 , n5743 , n5744 , 
 n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , 
 n5755 , n5756 , n5757 , n5758 , n75626 , n5760 , n5761 , n5762 , n5763 , n5764 , 
 n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , 
 n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , 
 n5785 , n5786 , n5787 , n5788 , n5789 , n75657 , n5791 , n5792 , n5793 , n5794 , 
 n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , 
 n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , 
 n5815 , n75683 , n75684 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , 
 n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , 
 n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n75709 , n5843 , n5844 , 
 n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , 
 n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , 
 n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , 
 n5875 , n5876 , n5877 , n75745 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , 
 n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n75759 , n5893 , n5894 , 
 n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , 
 n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n75781 , 
 n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , 
 n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , 
 n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , 
 n75812 , n5949 , n75814 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , 
 n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , 
 n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n75838 , n5978 , n5979 , n5980 , 
 n5981 , n5982 , n5983 , n5984 , n75846 , n75847 , n5987 , n5988 , n5989 , n5990 , 
 n5991 , n5992 , n75854 , n75855 , n5995 , n5996 , n5997 , n5998 , n5999 , n75861 , 
 n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
 n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
 n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
 n6031 , n6032 , n6033 , n6034 , n75896 , n75897 , n6037 , n6038 , n6039 , n6040 , 
 n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
 n75912 , n75913 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n75920 , n75921 , 
 n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
 n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
 n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n75951 , 
 n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
 n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
 n6111 , n6112 , n75974 , n6114 , n6115 , n6116 , n6117 , n6118 , n75980 , n6120 , 
 n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
 n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
 n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
 n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
 n6161 , n6162 , n6163 , n6164 , n6165 , n76027 , n76028 , n6168 , n6169 , n6170 , 
 n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
 n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
 n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
 n6201 , n6202 , n76064 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
 n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n76081 , 
 n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
 n6231 , n6232 , n6233 , n76095 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
 n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
 n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
 n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n76131 , 
 n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
 n6281 , n6282 , n76144 , n6287 , n76146 , n6289 , n6290 , n6291 , n6292 , n6293 , 
 n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , 
 n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n76170 , n6316 , 
 n6317 , n6318 , n6319 , n6320 , n76176 , n76177 , n6323 , n6324 , n6325 , n6326 , 
 n6327 , n6328 , n76184 , n76185 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , 
 n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n76198 , n76199 , n6345 , n6346 , 
 n6347 , n6348 , n6349 , n6350 , n76206 , n76207 , n6353 , n6354 , n6355 , n6356 , 
 n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , 
 n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , 
 n76232 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , 
 n6387 , n6388 , n76244 , n76245 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , 
 n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , 
 n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , 
 n6417 , n6418 , n6419 , n76275 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , 
 n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , 
 n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n76298 , n6444 , n6445 , n6446 , 
 n6447 , n6448 , n76304 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , 
 n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , 
 n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , 
 n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , 
 n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , 
 n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , 
 n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n76369 , n76370 , n6516 , 
 n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , 
 n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , 
 n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n76401 , 
 n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , 
 n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , 
 n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , 
 n6577 , n76433 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , 
 n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , 
 n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n76458 , n6604 , n6605 , n6606 , 
 n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , 
 n6617 , n6618 , n76474 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , 
 n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , 
 n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , 
 n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n76510 , n6659 , 
 n76512 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
 n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
 n6680 , n6681 , n6682 , n6683 , n76536 , n6688 , n6689 , n6690 , n6691 , n6692 , 
 n6693 , n76543 , n76544 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n76551 , 
 n76552 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , 
 n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , 
 n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , 
 n6733 , n6734 , n6735 , n6736 , n6737 , n76587 , n76588 , n6740 , n6741 , n6742 , 
 n6743 , n6744 , n6745 , n76595 , n76596 , n6748 , n6749 , n6750 , n6751 , n6752 , 
 n76602 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , 
 n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , 
 n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , 
 n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , 
 n6793 , n76643 , n76644 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , 
 n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , 
 n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n76668 , n6820 , n6821 , n6822 , 
 n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , 
 n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , 
 n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n76701 , 
 n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n76711 , 
 n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , 
 n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , 
 n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , 
 n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , 
 n6903 , n6904 , n76754 , n76755 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , 
 n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , 
 n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , 
 n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , 
 n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n76800 , n6952 , 
 n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , 
 n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n76818 , n6970 , n6971 , n6972 , 
 n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
 n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , 
 n6993 , n76843 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , 
 n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , 
 n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , 
 n7023 , n76873 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , 
 n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n76891 , 
 n7046 , n76893 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , 
 n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , 
 n7066 , n7067 , n7068 , n7069 , n7070 , n76917 , n7075 , n7076 , n7077 , n7078 , 
 n7079 , n7080 , n7081 , n76925 , n76926 , n7084 , n7085 , n7086 , n7087 , n7088 , 
 n7089 , n76933 , n76934 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
 n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n76948 , n7106 , n7107 , n7108 , 
 n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
 n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
 n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
 n7139 , n7140 , n7141 , n7142 , n7143 , n76987 , n76988 , n7146 , n7147 , n7148 , 
 n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
 n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
 n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n77020 , n77021 , 
 n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n77028 , n77029 , n7187 , n7188 , 
 n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
 n7199 , n7200 , n7201 , n7202 , n77046 , n7204 , n7205 , n7206 , n7207 , n7208 , 
 n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
 n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
 n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
 n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
 n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
 n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
 n7269 , n7270 , n7271 , n7272 , n77116 , n7274 , n7275 , n7276 , n7277 , n7278 , 
 n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
 n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n77141 , 
 n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
 n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
 n7319 , n7320 , n7321 , n77165 , n77166 , n7324 , n7325 , n7326 , n7327 , n7328 , 
 n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
 n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n77191 , 
 n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
 n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
 n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
 n7379 , n7380 , n77224 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
 n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
 n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
 n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n77259 , n7417 , n7418 , 
 n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
 n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n77279 , n7437 , n7438 , 
 n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
 n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
 n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n77311 , 
 n7472 , n77313 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , 
 n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , 
 n7492 , n7493 , n7494 , n7495 , n7496 , n77337 , n7501 , n7502 , n7503 , n7504 , 
 n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , 
 n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n77358 , n77359 , n7523 , n7524 , 
 n7525 , n7526 , n7527 , n7528 , n77366 , n77367 , n7531 , n7532 , n7533 , n7534 , 
 n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , 
 n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n77388 , n7552 , n7553 , n7554 , 
 n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , 
 n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , 
 n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , 
 n77422 , n77423 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , 
 n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , 
 n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n77450 , n77451 , 
 n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n77458 , n77459 , n7623 , n7624 , 
 n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , 
 n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , 
 n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , 
 n7655 , n7656 , n7657 , n77495 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , 
 n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , 
 n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , 
 n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , 
 n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , 
 n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , 
 n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , 
 n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , 
 n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , 
 n7745 , n7746 , n7747 , n7748 , n7749 , n77587 , n77588 , n7752 , n7753 , n7754 , 
 n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , 
 n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , 
 n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , 
 n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , 
 n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , 
 n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , 
 n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n77658 , n7822 , n7823 , n7824 , 
 n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , 
 n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , 
 n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , 
 n7855 , n77693 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , 
 n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , 
 n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , 
 n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , 
 n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n77738 , n7905 , n77740 , n7907 , 
 n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , 
 n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , 
 n7928 , n7929 , n77764 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
 n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
 n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n77790 , n77791 , 
 n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n77798 , n77799 , n7969 , n7970 , 
 n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
 n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
 n77822 , n77823 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n77830 , n77831 , 
 n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
 n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
 n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
 n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n77871 , 
 n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
 n8051 , n8052 , n8053 , n8054 , n77886 , n77887 , n8057 , n8058 , n8059 , n8060 , 
 n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
 n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
 n8081 , n8082 , n77914 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
 n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
 n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
 n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
 n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
 n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
 n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
 n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
 n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
 n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n78008 , n78009 , n8179 , n8180 , 
 n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
 n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
 n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
 n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
 n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
 n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
 n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
 n78082 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
 n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
 n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
 n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
 n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
 n8301 , n78133 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
 n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
 n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
 n8331 , n8332 , n8333 , n78165 , n8338 , n78167 , n8340 , n8341 , n8342 , n8343 , 
 n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , 
 n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n78191 , 
 n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n78199 , n8375 , n8376 , 
 n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , 
 n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , 
 n8397 , n8398 , n78224 , n78225 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , 
 n78232 , n78233 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , 
 n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , 
 n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , 
 n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , 
 n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , 
 n8457 , n8458 , n8459 , n78285 , n78286 , n8462 , n8463 , n8464 , n8465 , n8466 , 
 n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , 
 n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n78310 , n78311 , 
 n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n78318 , n78319 , n8495 , n8496 , 
 n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , 
 n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , 
 n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , 
 n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , 
 n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n78369 , n8545 , n8546 , 
 n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , 
 n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , 
 n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , 
 n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , 
 n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , 
 n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , 
 n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , 
 n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , 
 n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , 
 n8637 , n78463 , n78464 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , 
 n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , 
 n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , 
 n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , 
 n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , 
 n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , 
 n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , 
 n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n78541 , 
 n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , 
 n78552 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , 
 n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , 
 n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , 
 n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , 
 n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , 
 n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , 
 n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , 
 n8797 , n8798 , n78624 , n8803 , n78626 , n8805 , n8806 , n8807 , n8808 , n8809 , 
 n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
 n8820 , n8821 , n8822 , n78645 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , 
 n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , 
 n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , 
 n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n78680 , n78681 , 
 n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n78688 , n78689 , n8871 , n8872 , 
 n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , 
 n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n78709 , n78710 , n8892 , 
 n8893 , n8894 , n8895 , n8896 , n8897 , n78717 , n78718 , n8900 , n8901 , n8902 , 
 n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , 
 n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , 
 n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , 
 n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , 
 n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , 
 n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , 
 n8963 , n8964 , n8965 , n78785 , n78786 , n8968 , n8969 , n8970 , n8971 , n8972 , 
 n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , 
 n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , 
 n78812 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , 
 n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , 
 n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , 
 n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , 
 n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , 
 n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , 
 n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , 
 n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , 
 n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , 
 n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , 
 n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9102 , n9103 , 
 n9104 , n9105 , n9106 , n9107 , n78926 , n78927 , n9110 , n9111 , n9112 , n9113 , 
 n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , 
 n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , 
 n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , 
 n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , 
 n9154 , n9155 , n9156 , n78975 , n9158 , n9159 , n9160 , n9161 , n9162 , n78981 , 
 n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , 
 n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , 
 n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , 
 n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , 
 n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , 
 n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , 
 n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , 
 n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n79061 , 
 n9247 , n79063 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , 
 n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , 
 n9267 , n9268 , n9269 , n9270 , n9271 , n79087 , n9276 , n9277 , n9278 , n9279 , 
 n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n79099 , n79100 , n9289 , 
 n9290 , n9291 , n9292 , n9293 , n9294 , n79107 , n79108 , n9297 , n9298 , n9299 , 
 n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
 n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
 n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
 n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
 n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
 n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
 n9360 , n9361 , n9362 , n9363 , n9364 , n79177 , n79178 , n9367 , n9368 , n9369 , 
 n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
 n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
 n79202 , n79203 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n79210 , n79211 , 
 n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
 n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
 n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
 n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
 n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
 n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
 n9460 , n79273 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
 n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
 n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
 n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
 n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
 n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
 n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
 n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
 n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
 n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
 n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
 n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
 n9580 , n79393 , n79394 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
 n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
 n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
 n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
 n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n79438 , n9627 , n79440 , n9629 , 
 n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
 n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
 n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
 n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
 n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
 n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
 n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
 n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
 n9710 , n9711 , n79524 , n9716 , n79526 , n9718 , n9719 , n9720 , n9721 , n9722 , 
 n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , 
 n9733 , n9734 , n9735 , n79545 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , 
 n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , 
 n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , 
 n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , 
 n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , 
 n9786 , n9787 , n79594 , n79595 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , 
 n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , 
 n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , 
 n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , 
 n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , 
 n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , 
 n79652 , n79653 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , 
 n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , 
 n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , 
 n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n79689 , n79690 , n9885 , 
 n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , 
 n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , 
 n9906 , n9907 , n9908 , n9909 , n79716 , n9911 , n9912 , n9913 , n9914 , n9915 , 
 n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , 
 n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , 
 n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , 
 n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , 
 n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , 
 n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , 
 n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , 
 n9986 , n79793 , n79794 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , 
 n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , 
 n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , 
 n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , 
 n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , 
 n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , 
 n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , 
 n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n79871 , 
 n10066 , n10067 , n10068 , n10069 , n10070 , n79877 , n10072 , n10073 , n10074 , n10075 , 
 n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , 
 n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , 
 n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , 
 n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , 
 n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , 
 n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , 
 n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , 
 n10146 , n10147 , n10148 , n10149 , n79956 , n10154 , n79958 , n10156 , n10157 , n10158 , 
 n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
 n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
 n79982 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , 
 n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , 
 n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , 
 n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , 
 n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , 
 n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , 
 n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , 
 n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , 
 n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , 
 n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , 
 n10282 , n10283 , n10284 , n80085 , n80086 , n10287 , n10288 , n10289 , n10290 , n10291 , 
 n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , 
 n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , 
 n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , 
 n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , 
 n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , 
 n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n80148 , n10349 , n10350 , n10351 , 
 n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , 
 n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , 
 n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , 
 n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , 
 n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , 
 n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , 
 n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , 
 n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , 
 n10432 , n10433 , n10434 , n80235 , n80236 , n10437 , n10438 , n10439 , n10440 , n10441 , 
 n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , 
 n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , 
 n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , 
 n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , 
 n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , 
 n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , 
 n10502 , n10503 , n80304 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , 
 n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , 
 n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , 
 n10532 , n80333 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , 
 n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , 
 n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , 
 n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , 
 n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , 
 n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n80391 , 
 n10595 , n80393 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , 
 n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , 
 n80412 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , 
 n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , 
 n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , 
 n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , 
 n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , 
 n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , 
 n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , 
 n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , 
 n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n80498 , n80499 , n10706 , n10707 , 
 n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , 
 n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , 
 n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , 
 n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , 
 n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , 
 n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , 
 n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , 
 n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n80578 , n10785 , n10786 , n10787 , 
 n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , 
 n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , 
 n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , 
 n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , 
 n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , 
 n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , 
 n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n80649 , n80650 , n10857 , 
 n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , 
 n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , 
 n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , 
 n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , 
 n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , 
 n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , 
 n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , 
 n10928 , n80723 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , 
 n10938 , n80733 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , 
 n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , 
 n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , 
 n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , 
 n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , 
 n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , 
 n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , 
 n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , 
 n11018 , n80813 , n11023 , n80815 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , 
 n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , 
 n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n80839 , n11052 , n11053 , 
 n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , 
 n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , 
 n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , 
 n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , 
 n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , 
 n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , 
 n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , 
 n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , 
 n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , 
 n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , 
 n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n80949 , n80950 , n11163 , 
 n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , 
 n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , 
 n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , 
 n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , 
 n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n81000 , n11213 , 
 n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , 
 n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , 
 n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , 
 n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , 
 n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , 
 n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , 
 n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , 
 n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n81081 , 
 n81082 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , 
 n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , 
 n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , 
 n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , 
 n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , 
 n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , 
 n11354 , n11355 , n11356 , n11357 , n81146 , n11359 , n11360 , n11361 , n11362 , n11363 , 
 n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , 
 n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , 
 n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , 
 n11394 , n11395 , n11396 , n81185 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , 
 n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , 
 n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , 
 n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , 
 n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , 
 n11444 , n11445 , n81234 , n11450 , n81236 , n11452 , n11453 , n11454 , n11455 , n11456 , 
 n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , 
 n11467 , n11468 , n11469 , n11470 , n81256 , n11475 , n11476 , n11477 , n11478 , n11479 , 
 n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
 n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
 n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
 n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
 n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
 n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
 n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
 n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
 n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n81349 , n81350 , n11569 , 
 n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
 n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
 n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
 n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
 n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
 n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
 n11630 , n11631 , n81414 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
 n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
 n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
 n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
 n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
 n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
 n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
 n81482 , n81483 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
 n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
 n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
 n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
 n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
 n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
 n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n81550 , n11769 , 
 n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
 n11780 , n11781 , n11782 , n81565 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
 n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
 n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
 n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
 n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
 n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
 n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
 n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n81638 , n11860 , n81640 , n11862 , 
 n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , 
 n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , 
 n11883 , n11884 , n81664 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , 
 n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , 
 n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , 
 n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , 
 n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , 
 n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , 
 n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , 
 n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , 
 n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , 
 n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , 
 n11986 , n81763 , n81764 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , 
 n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , 
 n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , 
 n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , 
 n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , 
 n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n81818 , n12043 , n12044 , n12045 , 
 n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , 
 n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , 
 n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , 
 n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , 
 n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , 
 n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , 
 n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n81890 , n81891 , 
 n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , 
 n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , 
 n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , 
 n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , 
 n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , 
 n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , 
 n12176 , n12177 , n12178 , n12179 , n12180 , n81957 , n12182 , n12183 , n12184 , n12185 , 
 n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , 
 n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , 
 n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , 
 n81992 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , 
 n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , 
 n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , 
 n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , 
 n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , 
 n12266 , n12267 , n12268 , n82045 , n12273 , n82047 , n12275 , n12276 , n12277 , n12278 , 
 n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
 n12289 , n12290 , n12291 , n12292 , n12293 , n82067 , n12298 , n12299 , n12300 , n12301 , 
 n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , 
 n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , 
 n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , 
 n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , 
 n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , 
 n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , 
 n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , 
 n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , 
 n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n82160 , n82161 , 
 n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , 
 n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , 
 n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , 
 n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , 
 n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , 
 n12442 , n12443 , n12444 , n82215 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , 
 n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , 
 n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , 
 n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , 
 n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , 
 n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , 
 n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , 
 n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , 
 n12522 , n12523 , n12524 , n82295 , n82296 , n12527 , n12528 , n12529 , n12530 , n12531 , 
 n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , 
 n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , 
 n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , 
 n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , 
 n82342 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , 
 n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , 
 n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , 
 n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n82381 , 
 n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , 
 n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , 
 n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , 
 n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , 
 n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n82430 , n12664 , 
 n82432 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , 
 n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , 
 n12685 , n12686 , n12687 , n12688 , n82456 , n12693 , n12694 , n12695 , n12696 , n12697 , 
 n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , 
 n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , 
 n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , 
 n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , 
 n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , 
 n12748 , n12749 , n12750 , n12751 , n82516 , n82517 , n12754 , n12755 , n12756 , n12757 , 
 n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , 
 n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , 
 n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , 
 n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , 
 n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , 
 n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , 
 n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , 
 n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n82600 , n12837 , 
 n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , 
 n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , 
 n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , 
 n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , 
 n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , 
 n12888 , n12889 , n12890 , n12891 , n12892 , n82657 , n82658 , n12895 , n12896 , n12897 , 
 n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , 
 n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , 
 n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , 
 n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , 
 n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , 
 n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , 
 n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n82728 , n12965 , n12966 , n12967 , 
 n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n82739 , n12976 , n12977 , 
 n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , 
 n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , 
 n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , 
 n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , 
 n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , 
 n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , 
 n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , 
 n13048 , n13049 , n13050 , n13051 , n82816 , n13056 , n82818 , n13058 , n13059 , n13060 , 
 n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , 
 n13071 , n13072 , n13073 , n13074 , n13075 , n82837 , n13080 , n13081 , n13082 , n13083 , 
 n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , 
 n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , 
 n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , 
 n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , 
 n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , 
 n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n82900 , n82901 , 
 n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , 
 n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , 
 n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , 
 n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , 
 n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , 
 n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , 
 n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , 
 n13214 , n13215 , n13216 , n82975 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , 
 n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , 
 n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , 
 n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , 
 n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , 
 n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , 
 n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , 
 n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , 
 n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , 
 n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n83069 , n83070 , n13313 , 
 n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , 
 n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , 
 n83092 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , 
 n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , 
 n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , 
 n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , 
 n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , 
 n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , 
 n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , 
 n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , 
 n13414 , n13415 , n13416 , n13417 , n83176 , n13422 , n83178 , n13424 , n13425 , n13426 , 
 n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , 
 n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , 
 n83202 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
 n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
 n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
 n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
 n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
 n13500 , n13501 , n13502 , n13503 , n83256 , n83257 , n13506 , n13507 , n13508 , n13509 , 
 n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
 n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
 n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
 n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
 n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
 n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
 n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
 n13580 , n13581 , n13582 , n83335 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
 n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
 n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
 n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
 n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
 n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
 n13640 , n13641 , n13642 , n13643 , n13644 , n83397 , n83398 , n13647 , n13648 , n13649 , 
 n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
 n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
 n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
 n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
 n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
 n13700 , n83453 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
 n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
 n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
 n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
 n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
 n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
 n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
 n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , 
 n13780 , n13781 , n13782 , n83535 , n13787 , n83537 , n13789 , n13790 , n13791 , n13792 , 
 n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , 
 n13803 , n13804 , n13805 , n13806 , n83556 , n13811 , n13812 , n13813 , n13814 , n13815 , 
 n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , 
 n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , 
 n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , 
 n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , 
 n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n83609 , n83610 , n13865 , 
 n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , 
 n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , 
 n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , 
 n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , 
 n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , 
 n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , 
 n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , 
 n13936 , n13937 , n13938 , n13939 , n83686 , n13941 , n13942 , n13943 , n13944 , n13945 , 
 n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , 
 n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , 
 n13966 , n13967 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , 
 n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , 
 n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , 
 n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , 
 n14007 , n14008 , n14009 , n14010 , n83756 , n83757 , n14013 , n14014 , n14015 , n14016 , 
 n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , 
 n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , 
 n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , 
 n14047 , n14048 , n83794 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , 
 n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , 
 n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , 
 n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , 
 n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , 
 n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , 
 n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , 
 n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , 
 n14127 , n14128 , n83874 , n14133 , n83876 , n14135 , n14136 , n14137 , n14138 , n14139 , 
 n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , 
 n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n83900 , n14162 , 
 n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , 
 n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , 
 n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , 
 n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , 
 n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n83949 , n83950 , n14212 , 
 n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , 
 n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , 
 n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , 
 n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , 
 n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , 
 n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , 
 n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , 
 n14283 , n14284 , n14285 , n14286 , n84026 , n14288 , n14289 , n14290 , n14291 , n14292 , 
 n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , 
 n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , 
 n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , 
 n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , 
 n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , 
 n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , 
 n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , 
 n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , 
 n14373 , n14374 , n84114 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , 
 n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , 
 n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , 
 n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , 
 n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , 
 n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , 
 n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , 
 n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , 
 n14453 , n14454 , n84194 , n14459 , n84196 , n14461 , n14462 , n14463 , n14464 , n14465 , 
 n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , 
 n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , 
 n84222 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , 
 n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , 
 n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
 n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , 
 n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , 
 n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , 
 n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n84289 , n84290 , n14558 , 
 n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , 
 n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , 
 n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , 
 n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , 
 n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , 
 n84342 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , 
 n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , 
 n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , 
 n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , 
 n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , 
 n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , 
 n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , 
 n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , 
 n14689 , n14690 , n14691 , n84425 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , 
 n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , 
 n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , 
 n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , 
 n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , 
 n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , 
 n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , 
 n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n84501 , 
 n14772 , n84503 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , 
 n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , 
 n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n84531 , 
 n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , 
 n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , 
 n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , 
 n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , 
 n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , 
 n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n84590 , n84591 , 
 n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , 
 n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , 
 n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , 
 n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , 
 n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , 
 n14915 , n14916 , n14917 , n14918 , n14919 , n84647 , n14921 , n14922 , n14923 , n14924 , 
 n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , 
 n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14942 , n14943 , n14944 , n14945 , 
 n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , 
 n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , 
 n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , 
 n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , 
 n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , 
 n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , 
 n15006 , n15007 , n84734 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , 
 n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , 
 n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , 
 n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , 
 n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , 
 n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , 
 n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n84801 , 
 n15080 , n84803 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , 
 n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , 
 n15100 , n15101 , n15102 , n84825 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , 
 n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , 
 n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , 
 n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , 
 n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , 
 n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n84878 , n84879 , n15161 , n15162 , 
 n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , 
 n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , 
 n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , 
 n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , 
 n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , 
 n15213 , n15214 , n15215 , n84935 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , 
 n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , 
 n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , 
 n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , 
 n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , 
 n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , 
 n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , 
 n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , 
 n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n85018 , n15300 , n15301 , n15302 , 
 n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , 
 n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , 
 n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , 
 n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , 
 n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , 
 n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , 
 n85082 , n15367 , n85084 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , 
 n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , 
 n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n85109 , n15397 , n15398 , 
 n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , 
 n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , 
 n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , 
 n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , 
 n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , 
 n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , 
 n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , 
 n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , 
 n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n85198 , n15486 , n15487 , n15488 , 
 n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , 
 n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , 
 n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , 
 n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , 
 n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , 
 n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , 
 n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , 
 n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n85281 , 
 n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , 
 n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , 
 n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , 
 n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , 
 n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , 
 n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n85339 , n15630 , n85341 , 
 n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , 
 n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n85360 , n15654 , 
 n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , 
 n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , 
 n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , 
 n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , 
 n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , 
 n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , 
 n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , 
 n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , 
 n15735 , n15736 , n15737 , n15738 , n15739 , n85447 , n15741 , n15742 , n15743 , n15744 , 
 n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , 
 n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , 
 n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , 
 n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , 
 n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , 
 n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , 
 n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n85519 , n15813 , n15814 , 
 n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , 
 n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , 
 n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , 
 n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , 
 n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , 
 n15865 , n85573 , n15870 , n85575 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , 
 n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , 
 n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n85599 , n15899 , n15900 , 
 n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , 
 n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , 
 n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , 
 n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , 
 n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , 
 n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , 
 n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , 
 n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n85681 , 
 n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , 
 n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , 
 n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , 
 n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , 
 n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , 
 n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , 
 n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n85748 , n16048 , n16049 , n16050 , 
 n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , 
 n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , 
 n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , 
 n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , 
 n16091 , n16092 , n16093 , n16094 , n85796 , n16099 , n85798 , n16101 , n16102 , n16103 , 
 n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , 
 n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , 
 n16124 , n16125 , n85824 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , 
 n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , 
 n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , 
 n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , 
 n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , 
 n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , 
 n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , 
 n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , 
 n16207 , n16208 , n16209 , n16210 , n85906 , n16212 , n16213 , n16214 , n16215 , n16216 , 
 n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , 
 n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , 
 n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , 
 n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , 
 n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , 
 n16267 , n16268 , n16269 , n85965 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , 
 n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , 
 n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , 
 n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , 
 n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n86009 , n16318 , n86011 , 
 n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , 
 n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , 
 n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n86039 , n16351 , n16352 , 
 n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , 
 n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , 
 n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , 
 n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , 
 n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , 
 n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , 
 n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , 
 n16423 , n16424 , n16425 , n16426 , n16427 , n86117 , n16429 , n16430 , n16431 , n16432 , 
 n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , 
 n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , 
 n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , 
 n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , 
 n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , 
 n16483 , n16484 , n86174 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , 
 n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , 
 n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , 
 n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , 
 n86212 , n16527 , n86214 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , 
 n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , 
 n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n86240 , n16558 , 
 n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , 
 n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , 
 n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , 
 n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , 
 n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , 
 n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , 
 n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , 
 n16629 , n86313 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , 
 n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , 
 n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , 
 n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , 
 n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , 
 n16679 , n16680 , n16681 , n16682 , n16683 , n86367 , n16685 , n16686 , n16687 , n16688 , 
 n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , 
 n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , 
 n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n86401 , 
 n16722 , n86403 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , 
 n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , 
 n16742 , n16743 , n16744 , n16745 , n16746 , n86427 , n16751 , n16752 , n16753 , n16754 , 
 n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , 
 n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , 
 n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , 
 n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , 
 n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , 
 n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , 
 n16815 , n16816 , n16817 , n86495 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , 
 n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , 
 n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , 
 n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , 
 n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , 
 n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n86549 , n16873 , n16874 , 
 n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , 
 n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , 
 n16895 , n16896 , n16897 , n16898 , n16899 , n86577 , n16904 , n86579 , n16906 , n16907 , 
 n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , 
 n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n86599 , n16929 , n16930 , 
 n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , 
 n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , 
 n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , 
 n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , 
 n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , 
 n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n86661 , 
 n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , 
 n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , 
 n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , 
 n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , 
 n17031 , n86703 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , 
 n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , 
 n17051 , n17052 , n17053 , n17054 , n17055 , n86727 , n17060 , n86729 , n17062 , n17063 , 
 n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , 
 n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , 
 n17084 , n86753 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , 
 n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , 
 n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , 
 n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , 
 n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , 
 n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n86809 , n17145 , n17146 , 
 n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , 
 n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , 
 n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , 
 n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , 
 n86852 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , 
 n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n86870 , n17209 , 
 n86872 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , 
 n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n86891 , 
 n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , 
 n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , 
 n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , 
 n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , 
 n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , 
 n17283 , n17284 , n86944 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , 
 n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , 
 n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , 
 n17313 , n17314 , n17315 , n86975 , n17320 , n86977 , n17322 , n17323 , n17324 , n17325 , 
 n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , 
 n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , 
 n17346 , n87003 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , 
 n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , 
 n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , 
 n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , 
 n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n87051 , 
 n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , 
 n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , 
 n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , 
 n17429 , n17430 , n17431 , n17432 , n87086 , n17437 , n87088 , n17439 , n17440 , n17441 , 
 n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , 
 n17452 , n17453 , n17454 , n17455 , n17456 , n87107 , n17461 , n17462 , n17463 , n17464 , 
 n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , 
 n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , 
 n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , 
 n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n87149 , n17503 , n17504 , 
 n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , 
 n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , 
 n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n87181 , 
 n17538 , n87183 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , 
 n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n87200 , n17560 , 
 n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , 
 n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , 
 n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , 
 n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n87238 , n17598 , n17599 , n17600 , 
 n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , 
 n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , 
 n17621 , n17622 , n87264 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , 
 n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , 
 n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , 
 n17654 , n17655 , n17656 , n17657 , n87296 , n17659 , n17660 , n17661 , n17662 , n17663 , 
 n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , 
 n17674 , n17675 , n17676 , n17677 , n87316 , n17682 , n17683 , n17684 , n17685 , n17686 , 
 n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , 
 n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , 
 n87342 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , 
 n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n87358 , n17727 , n17728 , n17729 , 
 n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , 
 n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n87381 , 
 n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n87390 , n17762 , 
 n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , 
 n17773 , n17774 , n17775 , n17776 , n87406 , n17781 , n87408 , n87409 , n87410 , n87411 , 
 n87412 , n87413 , n87414 , n87415 , n87416 , n87417 , n87418 , n87419 , n87420 , n87421 , 
 n87422 , n87423 , n87424 , n87425 , n87426 , n87427 , n87428 , n87429 , n87430 , n87431 , 
 n87432 , n87433 , n87434 , n87435 , n87436 , n87437 , n87438 , n87439 , n87440 , n87441 , 
 n87442 , n87443 , n87444 , n87445 , n87446 , n87447 , n87448 , n87449 , n87450 , n87451 , 
 n87452 , n87453 , n87454 , n87455 , n87456 , n87457 , n87458 , n87459 , n87460 , n87461 , 
 n87462 , n87463 , n87464 , n87465 , n87466 , n87467 , n87468 , n87469 , n87470 , n87471 , 
 n87472 , n87473 , n87474 , n87475 , n87476 , n87477 , n87478 , n87479 , n87480 , n87481 , 
 n87482 , n87483 , n87484 , n87485 , n87486 , n87487 , n87488 , n87489 , n87490 , n87491 , 
 n87492 , n87493 , n87494 , n87495 , n87496 , n87497 , n87498 , n87499 , n87500 , n87501 , 
 n87502 , n87503 , n87504 , n87505 , n87506 , n87507 , n87508 , n87509 , n87510 , n87511 , 
 n87512 , n87513 , n87514 , n87515 , n87516 , n87517 , n87518 , n87519 , n87520 , n87521 , 
 n87522 , n87523 , n87524 , n87525 , n87526 , n87527 , n87528 , n87529 , n87530 , n87531 , 
 n87532 , n87533 , n87534 , n87535 , n87536 , n87537 , n87538 , n87539 , n87540 , n87541 , 
 n87542 , n87543 , n87544 , n87545 , n87546 , n87547 , n87548 , n87549 , n87550 , n87551 , 
 n87552 , n87553 , n87554 , n87555 , n87556 , n87557 , n87558 , n87559 , n87560 , n87561 , 
 n87562 , n87563 , n87564 , n87565 , n87566 , n87567 , n87568 , n87569 , n87570 , n87571 , 
 n87572 , n87573 , n87574 , n87575 , n87576 , n87577 , n87578 , n87579 , n87580 , n87581 , 
 n87582 , n87583 , n87584 , n87585 , n87586 , n87587 , n87588 , n87589 , n87590 , n87591 , 
 n87592 , n87593 , n87594 , n87595 , n87596 , n87597 , n87598 , n87599 , n87600 , n87601 , 
 n87602 , n87603 , n87604 , n87605 , n87606 , n87607 , n87608 , n87609 , n87610 , n87611 , 
 n87612 , n87613 , n87614 , n87615 , n87616 , n87617 , n87618 , n87619 , n87620 , n87621 , 
 n87622 , n87623 , n87624 , n87625 , n87626 , n87627 , n87628 , n87629 , n87630 , n87631 , 
 n87632 , n87633 , n87634 , n87635 , n87636 , n87637 , n87638 , n87639 , n87640 , n87641 , 
 n87642 , n87643 , n87644 , n87645 , n87646 , n87647 , n87648 , n87649 , n87650 , n87651 , 
 n87652 , n87653 , n87654 , n87655 , n87656 , n87657 , n87658 , n87659 , n87660 , n87661 , 
 n87662 , n87663 , n87664 , n87665 , n87666 , n87667 , n87668 , n87669 , n87670 , n87671 , 
 n87672 , n87673 , n87674 , n87675 , n87676 , n87677 , n87678 , n87679 , n87680 , n87681 , 
 n87682 , n87683 , n87684 , n87685 , n87686 , n87687 , n87688 , n87689 , n87690 , n87691 , 
 n87692 , n87693 , n87694 , n87695 , n87696 , n87697 , n87698 , n87699 , n87700 , n87701 , 
 n87702 , n87703 , n87704 , n87705 , n87706 , n87707 , n87708 , n87709 , n87710 , n87711 , 
 n87712 , n87713 , n87714 , n87715 , n87716 , n87717 , n87718 , n87719 , n87720 , n87721 , 
 n87722 , n87723 , n87724 , n87725 , n87726 , n87727 , n87728 , n87729 , n87730 , n87731 , 
 n87732 , n87733 , n87734 , n87735 , n87736 , n87737 , n87738 , n87739 , n87740 , n87741 , 
 n87742 , n87743 , n87744 , n87745 , n87746 , n87747 , n87748 , n87749 , n87750 , n87751 , 
 n87752 , n87753 , n87754 , n87755 , n87756 , n87757 , n87758 , n87759 , n87760 , n87761 , 
 n87762 , n87763 , n87764 , n87765 , n87766 , n87767 , n87768 , n87769 , n87770 , n87771 , 
 n87772 , n87773 , n87774 , n87775 , n87776 , n87777 , n87778 , n87779 , n87780 , n87781 , 
 n87782 , n87783 , n87784 , n87785 , n87786 , n87787 , n87788 , n87789 , n87790 , n87791 , 
 n87792 , n87793 , n87794 , n87795 , n87796 , n87797 , n87798 , n87799 , n87800 , n87801 , 
 n87802 , n87803 , n87804 , n87805 , n87806 , n87807 , n87808 , n87809 , n87810 , n87811 , 
 n87812 , n87813 , n87814 , n87815 , n87816 , n87817 , n87818 , n87819 , n87820 , n87821 , 
 n87822 , n87823 , n87824 , n87825 , n87826 , n87827 , n87828 , n87829 , n87830 , n87831 , 
 n87832 , n87833 , n87834 , n87835 , n87836 , n87837 , n87838 , n87839 , n87840 , n87841 , 
 n87842 , n87843 , n87844 , n87845 , n87846 , n87847 , n87848 , n87849 , n87850 , n87851 , 
 n87852 , n87853 , n87854 , n87855 , n87856 , n87857 , n87858 , n87859 , n87860 , n87861 , 
 n87862 , n87863 , n87864 , n87865 , n87866 , n87867 , n87868 , n87869 , n87870 , n87871 , 
 n87872 , n87873 , n87874 , n87875 , n87876 , n87877 , n87878 , n87879 , n87880 , n87881 , 
 n87882 , n87883 , n87884 , n87885 , n87886 , n87887 , n87888 , n87889 , n87890 , n87891 , 
 n87892 , n87893 , n87894 , n87895 , n87896 , n87897 , n87898 , n87899 , n87900 , n87901 , 
 n87902 , n87903 , n87904 , n87905 , n87906 , n87907 , n87908 , n87909 , n87910 , n87911 , 
 n87912 , n87913 , n87914 , n87915 , n87916 , n87917 , n87918 , n87919 , n87920 , n87921 , 
 n87922 , n87923 , n87924 , n87925 , n87926 , n87927 , n87928 , n87929 , n87930 , n87931 , 
 n87932 , n87933 , n87934 , n87935 , n87936 , n87937 , n87938 , n87939 , n87940 , n87941 , 
 n87942 , n87943 , n87944 , n87945 , n87946 , n87947 , n87948 , n87949 , n87950 , n87951 , 
 n87952 , n87953 , n87954 , n87955 , n87956 , n87957 , n87958 , n87959 , n87960 , n87961 , 
 n87962 , n87963 , n87964 , n87965 , n87966 , n87967 , n87968 , n87969 , n87970 , n87971 , 
 n87972 , n87973 , n87974 , n87975 , n87976 , n87977 , n87978 , n87979 , n87980 , n87981 , 
 n87982 , n87983 , n87984 , n87985 , n87986 , n87987 , n87988 , n87989 , n87990 , n87991 , 
 n87992 , n87993 , n87994 , n87995 , n87996 , n87997 , n87998 , n87999 , n88000 , n88001 , 
 n88002 , n88003 , n88004 , n88005 , n88006 , n88007 , n88008 , n88009 , n88010 , n88011 , 
 n88012 , n88013 , n88014 , n88015 , n88016 , n88017 , n88018 , n88019 , n88020 , n88021 , 
 n88022 , n88023 , n88024 , n88025 , n88026 , n88027 , n88028 , n88029 , n88030 , n88031 , 
 n88032 , n88033 , n88034 , n88035 , n88036 , n88037 , n88038 , n88039 , n88040 , n88041 , 
 n88042 , n88043 , n88044 , n88045 , n88046 , n88047 , n88048 , n88049 , n88050 , n88051 , 
 n88052 , n88053 , n88054 , n88055 , n88056 , n88057 , n88058 , n88059 , n88060 , n88061 , 
 n88062 , n88063 , n88064 , n88065 , n88066 , n88067 , n88068 , n88069 , n88070 , n88071 , 
 n88072 , n88073 , n88074 , n88075 , n88076 , n88077 , n88078 , n88079 , n88080 , n88081 , 
 n88082 , n88083 , n88084 , n88085 , n88086 , n88087 , n88088 , n88089 , n88090 , n88091 , 
 n88092 , n88093 , n88094 , n88095 , n88096 , n88097 , n88098 , n88099 , n88100 , n88101 , 
 n88102 , n88103 , n88104 , n88105 , n88106 , n88107 , n88108 , n88109 , n88110 , n88111 , 
 n88112 , n88113 , n88114 , n88115 , n88116 , n88117 , n88118 , n88119 , n88120 , n88121 , 
 n88122 , n88123 , n88124 , n88125 , n88126 , n88127 , n88128 , n88129 , n88130 , n88131 , 
 n88132 , n88133 , n88134 , n88135 , n88136 , n88137 , n88138 , n88139 , n88140 , n88141 , 
 n88142 , n88143 , n88144 , n88145 , n88146 , n88147 , n88148 , n88149 , n88150 , n88151 , 
 n88152 , n88153 , n88154 , n88155 , n88156 , n88157 , n88158 , n88159 , n88160 , n88161 , 
 n88162 , n88163 , n88164 , n88165 , n88166 , n88167 , n88168 , n88169 , n88170 , n17782 , 
 n88172 , n17784 , n88174 , n17789 , n17790 , n88177 , n17792 , n88179 , n17797 , n17798 , 
 n88182 , n17800 , n88184 , n17805 , n17806 , n88187 , n17808 , n88189 , n17813 , n17814 , 
 n88192 , n17816 , n88194 , n17821 , n88196 , n88197 , n88198 , n88199 , n88200 , n88201 , 
 n88202 , n88203 , n88204 , n88205 , n88206 , n88207 , n88208 , n88209 , n88210 , n88211 , 
 n88212 , n88213 , n88214 , n88215 , n88216 , n88217 , n88218 , n88219 , n88220 , n88221 , 
 n88222 , n88223 , n88224 , n88225 , n88226 , n88227 , n88228 , n88229 , n88230 , n88231 , 
 n88232 , n88233 , n88234 , n88235 , n88236 , n88237 , n88238 , n88239 , n88240 , n88241 , 
 n88242 , n88243 , n88244 , n88245 , n88246 , n88247 , n88248 , n88249 , n88250 , n88251 , 
 n88252 , n88253 , n88254 , n88255 , n88256 , n88257 , n88258 , n88259 , n88260 , n88261 , 
 n88262 , n88263 , n88264 , n88265 , n88266 , n88267 , n88268 , n88269 , n88270 , n88271 , 
 n88272 , n88273 , n88274 , n88275 , n88276 , n88277 , n88278 , n88279 , n88280 , n88281 , 
 n88282 , n88283 , n88284 , n88285 , n88286 , n88287 , n88288 , n88289 , n88290 , n88291 , 
 n88292 , n88293 , n88294 , n88295 , n88296 , n88297 , n88298 , n88299 , n88300 , n88301 , 
 n88302 , n88303 , n88304 , n88305 , n88306 , n88307 , n88308 , n88309 , n88310 , n88311 , 
 n88312 , n88313 , n88314 , n88315 , n88316 , n88317 , n88318 , n88319 , n88320 , n88321 , 
 n88322 , n88323 , n88324 , n88325 , n88326 , n88327 , n88328 , n88329 , n88330 , n88331 , 
 n88332 , n88333 , n88334 , n88335 , n88336 , n88337 , n88338 , n88339 , n88340 , n88341 , 
 n88342 , n88343 , n88344 , n88345 , n88346 , n88347 , n88348 , n88349 , n88350 , n88351 , 
 n88352 , n88353 , n88354 , n88355 , n88356 , n88357 , n88358 , n88359 , n88360 , n88361 , 
 n88362 , n88363 , n88364 , n88365 , n88366 , n88367 , n88368 , n88369 , n88370 , n88371 , 
 n88372 , n88373 , n88374 , n88375 , n88376 , n88377 , n88378 , n88379 , n88380 , n88381 , 
 n88382 , n88383 , n88384 , n88385 , n88386 , n88387 , n88388 , n88389 , n88390 , n88391 , 
 n88392 , n88393 , n88394 , n88395 , n88396 , n88397 , n88398 , n88399 , n88400 , n88401 , 
 n88402 , n88403 , n88404 , n88405 , n88406 , n88407 , n88408 , n88409 , n88410 , n88411 , 
 n88412 , n88413 , n88414 , n88415 , n88416 , n88417 , n88418 , n88419 , n88420 , n88421 , 
 n88422 , n88423 , n88424 , n88425 , n88426 , n88427 , n88428 , n88429 , n88430 , n88431 , 
 n88432 , n88433 , n88434 , n88435 , n88436 , n88437 , n88438 , n88439 , n88440 , n88441 , 
 n88442 , n88443 , n88444 , n88445 , n88446 , n88447 , n88448 , n88449 , n88450 , n88451 , 
 n88452 , n88453 , n88454 , n88455 , n88456 , n88457 , n88458 , n88459 , n88460 , n88461 , 
 n88462 , n88463 , n88464 , n88465 , n88466 , n88467 , n88468 , n88469 , n88470 , n88471 , 
 n88472 , n88473 , n88474 , n88475 , n88476 , n88477 , n88478 , n88479 , n88480 , n88481 , 
 n88482 , n88483 , n88484 , n88485 , n88486 , n88487 , n88488 , n88489 , n88490 , n88491 , 
 n88492 , n88493 , n88494 , n88495 , n88496 , n88497 , n88498 , n88499 , n88500 , n88501 , 
 n88502 , n88503 , n88504 , n88505 , n88506 , n88507 , n88508 , n88509 , n88510 , n88511 , 
 n88512 , n88513 , n88514 , n88515 , n88516 , n88517 , n88518 , n88519 , n88520 , n88521 , 
 n88522 , n88523 , n88524 , n88525 , n88526 , n88527 , n88528 , n88529 , n88530 , n88531 , 
 n88532 , n88533 , n88534 , n88535 , n88536 , n88537 , n88538 , n88539 , n88540 , n88541 , 
 n88542 , n88543 , n88544 , n88545 , n88546 , n88547 , n88548 , n88549 , n88550 , n88551 , 
 n88552 , n88553 , n88554 , n88555 , n88556 , n88557 , n88558 , n88559 , n88560 , n88561 , 
 n88562 , n88563 , n88564 , n88565 , n88566 , n88567 , n88568 , n88569 , n88570 , n88571 , 
 n88572 , n88573 , n88574 , n88575 , n88576 , n88577 , n88578 , n88579 , n88580 , n88581 , 
 n88582 , n88583 , n88584 , n88585 , n88586 , n88587 , n88588 , n88589 , n88590 , n88591 , 
 n88592 , n88593 , n88594 , n88595 , n88596 , n88597 , n88598 , n88599 , n88600 , n88601 , 
 n88602 , n88603 , n88604 , n88605 , n88606 , n88607 , n88608 , n88609 , n88610 , n88611 , 
 n88612 , n88613 , n88614 , n88615 , n88616 , n88617 , n88618 , n88619 , n88620 , n88621 , 
 n88622 , n88623 , n88624 , n88625 , n88626 , n88627 , n88628 , n88629 , n88630 , n88631 , 
 n88632 , n88633 , n88634 , n88635 , n88636 , n88637 , n88638 , n88639 , n88640 , n88641 , 
 n88642 , n88643 , n88644 , n88645 , n88646 , n88647 , n88648 , n88649 , n88650 , n88651 , 
 n88652 , n88653 , n88654 , n88655 , n88656 , n88657 , n88658 , n88659 , n88660 , n88661 , 
 n88662 , n88663 , n88664 , n88665 , n88666 , n88667 , n88668 , n88669 , n88670 , n88671 , 
 n88672 , n88673 , n88674 , n88675 , n88676 , n88677 , n88678 , n88679 , n88680 , n88681 , 
 n88682 , n88683 , n88684 , n88685 , n88686 , n88687 , n88688 , n88689 , n88690 , n88691 , 
 n88692 , n88693 , n88694 , n88695 , n88696 , n88697 , n88698 , n88699 , n88700 , n88701 , 
 n88702 , n88703 , n88704 , n88705 , n88706 , n88707 , n88708 , n88709 , n88710 , n88711 , 
 n88712 , n88713 , n88714 , n88715 , n88716 , n88717 , n88718 , n88719 , n88720 , n88721 , 
 n88722 , n88723 , n88724 , n88725 , n88726 , n88727 , n88728 , n88729 , n88730 , n88731 , 
 n88732 , n88733 , n88734 , n88735 , n88736 , n88737 , n88738 , n88739 , n88740 , n88741 , 
 n88742 , n88743 , n88744 , n88745 , n88746 , n88747 , n88748 , n88749 , n88750 , n88751 , 
 n88752 , n88753 , n88754 , n88755 , n88756 , n88757 , n88758 , n88759 , n88760 , n88761 , 
 n88762 , n88763 , n88764 , n88765 , n88766 , n88767 , n88768 , n88769 , n88770 , n88771 , 
 n88772 , n88773 , n88774 , n88775 , n88776 , n88777 , n88778 , n88779 , n88780 , n88781 , 
 n88782 , n88783 , n88784 , n88785 , n88786 , n88787 , n88788 , n88789 , n88790 , n88791 , 
 n88792 , n88793 , n88794 , n88795 , n88796 , n88797 , n88798 , n88799 , n88800 , n88801 , 
 n88802 , n88803 , n88804 , n88805 , n88806 , n88807 , n88808 , n88809 , n88810 , n88811 , 
 n88812 , n88813 , n88814 , n88815 , n88816 , n88817 , n88818 , n88819 , n88820 , n88821 , 
 n88822 , n88823 , n88824 , n88825 , n88826 , n88827 , n88828 , n88829 , n88830 , n88831 , 
 n88832 , n88833 , n88834 , n88835 , n88836 , n88837 , n88838 , n88839 , n88840 , n88841 , 
 n88842 , n88843 , n88844 , n88845 , n88846 , n88847 , n88848 , n88849 , n88850 , n88851 , 
 n88852 , n88853 , n88854 , n88855 , n88856 , n88857 , n88858 , n88859 , n88860 , n88861 , 
 n88862 , n88863 , n88864 , n88865 , n88866 , n88867 , n88868 , n88869 , n88870 , n88871 , 
 n88872 , n88873 , n88874 , n88875 , n88876 , n88877 , n88878 , n88879 , n88880 , n88881 , 
 n88882 , n88883 , n88884 , n88885 , n88886 , n88887 , n88888 , n88889 , n88890 , n88891 , 
 n88892 , n88893 , n88894 , n88895 , n88896 , n88897 , n88898 , n88899 , n88900 , n88901 , 
 n88902 , n88903 , n88904 , n88905 , n88906 , n88907 , n88908 , n88909 , n88910 , n88911 , 
 n88912 , n88913 , n88914 , n88915 , n88916 , n88917 , n88918 , n88919 , n88920 , n88921 , 
 n88922 , n88923 , n88924 , n88925 , n88926 , n88927 , n88928 , n88929 , n88930 , n88931 , 
 n88932 , n88933 , n88934 , n88935 , n88936 , n88937 , n88938 , n88939 , n88940 , n88941 , 
 n88942 , n88943 , n88944 , n88945 , n88946 , n88947 , n88948 , n88949 , n88950 , n88951 , 
 n88952 , n88953 , n88954 , n88955 , n88956 , n88957 , n88958 , n88959 , n88960 , n88961 , 
 n88962 , n88963 , n88964 , n88965 , n88966 , n88967 , n88968 , n88969 , n88970 , n88971 , 
 n88972 , n88973 , n88974 , n88975 , n88976 , n88977 , n88978 , n88979 , n88980 , n88981 , 
 n88982 , n88983 , n88984 , n88985 , n88986 , n88987 , n88988 , n88989 , n88990 , n88991 , 
 n88992 , n88993 , n88994 , n88995 , n88996 , n88997 , n88998 , n88999 , n89000 , n89001 , 
 n89002 , n89003 , n89004 , n89005 , n89006 , n89007 , n89008 , n89009 , n89010 , n89011 , 
 n89012 , n89013 , n89014 , n89015 , n89016 , n89017 , n89018 , n89019 , n89020 , n89021 , 
 n89022 , n89023 , n89024 , n89025 , n89026 , n89027 , n89028 , n89029 , n89030 , n89031 , 
 n89032 , n89033 , n89034 , n89035 , n89036 , n89037 , n89038 , n89039 , n89040 , n89041 , 
 n89042 , n89043 , n89044 , n89045 , n89046 , n89047 , n89048 , n89049 , n89050 , n89051 , 
 n89052 , n89053 , n89054 , n89055 , n89056 , n89057 , n89058 , n89059 , n89060 , n89061 , 
 n89062 , n89063 , n89064 , n89065 , n89066 , n89067 , n89068 , n89069 , n89070 , n89071 , 
 n89072 , n89073 , n89074 , n89075 , n89076 , n89077 , n89078 , n89079 , n89080 , n89081 , 
 n89082 , n89083 , n89084 , n89085 , n89086 , n89087 , n89088 , n89089 , n89090 , n89091 , 
 n89092 , n89093 , n89094 , n89095 , n89096 , n89097 , n89098 , n89099 , n89100 , n89101 , 
 n89102 , n89103 , n89104 , n89105 , n89106 , n89107 , n89108 , n89109 , n89110 , n89111 , 
 n89112 , n89113 , n89114 , n89115 , n89116 , n89117 , n89118 , n89119 , n89120 , n89121 , 
 n89122 , n89123 , n89124 , n89125 , n89126 , n89127 , n89128 , n89129 , n89130 , n89131 , 
 n89132 , n89133 , n89134 , n89135 , n89136 , n89137 , n89138 , n89139 , n89140 , n89141 , 
 n89142 , n89143 , n89144 , n89145 , n89146 , n89147 , n89148 , n89149 , n89150 , n89151 , 
 n89152 , n89153 , n89154 , n89155 , n89156 , n89157 , n89158 , n89159 , n89160 , n89161 , 
 n89162 , n89163 , n89164 , n89165 , n89166 , n89167 , n89168 , n89169 , n89170 , n89171 , 
 n89172 , n89173 , n89174 , n89175 , n89176 , n89177 , n89178 , n89179 , n89180 , n89181 , 
 n89182 , n89183 , n89184 , n89185 , n89186 , n89187 , n89188 , n89189 , n89190 , n89191 , 
 n89192 , n89193 , n89194 , n89195 , n89196 , n89197 , n89198 , n89199 , n89200 , n89201 , 
 n89202 , n89203 , n89204 , n89205 , n89206 , n89207 , n89208 , n89209 , n89210 , n89211 , 
 n89212 , n89213 , n89214 , n89215 , n89216 , n89217 , n89218 , n89219 , n89220 , n89221 , 
 n89222 , n89223 , n89224 , n89225 , n89226 , n89227 , n89228 , n89229 , n89230 , n89231 , 
 n89232 , n89233 , n89234 , n89235 , n89236 , n89237 , n89238 , n89239 , n89240 , n89241 , 
 n89242 , n89243 , n89244 , n89245 , n89246 , n89247 , n89248 , n89249 , n89250 , n89251 , 
 n89252 , n89253 , n89254 , n89255 , n89256 , n89257 , n89258 , n89259 , n89260 , n89261 , 
 n89262 , n89263 , n89264 , n89265 , n89266 , n89267 , n89268 , n89269 , n89270 , n89271 , 
 n89272 , n89273 , n89274 , n89275 , n89276 , n89277 , n89278 , n89279 , n89280 , n89281 , 
 n89282 , n89283 , n89284 , n89285 , n89286 , n89287 , n89288 , n89289 , n89290 , n89291 , 
 n89292 , n89293 , n89294 , n89295 , n89296 , n89297 , n89298 , n89299 , n89300 , n89301 , 
 n89302 , n89303 , n89304 , n89305 , n89306 , n89307 , n89308 , n89309 , n89310 , n89311 , 
 n89312 , n89313 , n89314 , n89315 , n89316 , n89317 , n89318 , n89319 , n89320 , n89321 , 
 n89322 , n89323 , n89324 , n89325 , n89326 , n89327 , n89328 , n89329 , n89330 , n89331 , 
 n89332 , n89333 , n89334 , n89335 , n89336 , n89337 , n89338 , n89339 , n89340 , n89341 , 
 n89342 , n89343 , n89344 , n89345 , n89346 , n89347 , n89348 , n89349 , n89350 , n89351 , 
 n89352 , n89353 , n89354 , n89355 , n89356 , n89357 , n89358 , n89359 , n89360 , n89361 , 
 n89362 , n89363 , n89364 , n89365 , n89366 , n89367 , n89368 , n89369 , n89370 , n89371 , 
 n89372 , n89373 , n89374 , n89375 , n89376 , n89377 , n89378 , n89379 , n89380 , n89381 , 
 n89382 , n89383 , n89384 , n89385 , n89386 , n89387 , n89388 , n89389 , n89390 , n89391 , 
 n89392 , n89393 , n89394 , n89395 , n89396 , n89397 , n89398 , n89399 , n89400 , n89401 , 
 n89402 , n89403 , n89404 , n89405 , n89406 , n89407 , n89408 , n89409 , n89410 , n89411 , 
 n89412 , n89413 , n89414 , n89415 , n89416 , n89417 , n89418 , n89419 , n89420 , n89421 , 
 n89422 , n89423 , n89424 , n89425 , n89426 , n89427 , n89428 , n89429 , n89430 , n89431 , 
 n89432 , n89433 , n89434 , n89435 , n89436 , n89437 , n89438 , n89439 , n89440 , n89441 , 
 n89442 , n89443 , n89444 , n89445 , n89446 , n89447 , n89448 , n89449 , n89450 , n89451 , 
 n89452 , n89453 , n89454 , n89455 , n89456 , n89457 , n89458 , n89459 , n89460 , n89461 , 
 n89462 , n89463 , n89464 , n89465 , n89466 , n89467 , n89468 , n89469 , n89470 , n89471 , 
 n89472 , n89473 , n89474 , n89475 , n89476 , n89477 , n89478 , n89479 , n89480 , n89481 , 
 n89482 , n89483 , n89484 , n89485 , n89486 , n89487 , n89488 , n89489 , n89490 , n89491 , 
 n89492 , n89493 , n89494 , n89495 , n89496 , n89497 , n89498 , n89499 , n89500 , n89501 , 
 n89502 , n89503 , n89504 , n89505 , n89506 , n89507 , n89508 , n89509 , n89510 , n89511 , 
 n89512 , n89513 , n89514 , n89515 , n89516 , n89517 , n89518 , n89519 , n89520 , n89521 , 
 n89522 , n89523 , n89524 , n89525 , n89526 , n89527 , n89528 , n89529 , n89530 , n89531 , 
 n89532 , n89533 , n89534 , n89535 , n89536 , n89537 , n89538 , n89539 , n89540 , n89541 , 
 n89542 , n89543 , n89544 , n89545 , n89546 , n89547 , n89548 , n89549 , n89550 , n89551 , 
 n89552 , n89553 , n89554 , n89555 , n89556 , n89557 , n89558 , n89559 , n89560 , n89561 , 
 n89562 , n89563 , n89564 , n89565 , n89566 , n89567 , n89568 , n89569 , n89570 , n89571 , 
 n89572 , n89573 , n89574 , n89575 , n89576 , n89577 , n89578 , n89579 , n89580 , n89581 , 
 n89582 , n89583 , n89584 , n89585 , n89586 , n89587 , n89588 , n89589 , n89590 , n89591 , 
 n89592 , n89593 , n89594 , n89595 , n89596 , n89597 , n89598 , n89599 , n89600 , n89601 , 
 n89602 , n89603 , n89604 , n89605 , n89606 , n89607 , n89608 , n89609 , n89610 , n89611 , 
 n89612 , n89613 , n89614 , n89615 , n89616 , n89617 , n89618 , n89619 , n89620 , n89621 , 
 n89622 , n89623 , n89624 , n89625 , n89626 , n89627 , n89628 , n89629 , n89630 , n89631 , 
 n89632 , n89633 , n89634 , n89635 , n89636 , n89637 , n89638 , n89639 , n89640 , n89641 , 
 n89642 , n89643 , n89644 , n89645 , n89646 , n89647 , n89648 , n89649 , n89650 , n89651 , 
 n89652 , n89653 , n89654 , n89655 , n89656 , n89657 , n89658 , n89659 , n89660 , n89661 , 
 n89662 , n89663 , n89664 , n89665 , n89666 , n89667 , n89668 , n89669 , n89670 , n89671 , 
 n89672 , n89673 , n89674 , n89675 , n89676 , n89677 , n89678 , n89679 , n89680 , n89681 , 
 n89682 , n89683 , n89684 , n89685 , n89686 , n89687 , n89688 , n89689 , n89690 , n89691 , 
 n89692 , n89693 , n89694 , n89695 , n89696 , n89697 , n89698 , n89699 , n89700 , n89701 , 
 n89702 , n89703 , n89704 , n89705 , n89706 , n89707 , n89708 , n89709 , n89710 , n89711 , 
 n89712 , n89713 , n89714 , n89715 , n89716 , n89717 , n89718 , n89719 , n89720 , n89721 , 
 n89722 , n89723 , n89724 , n89725 , n89726 , n89727 , n89728 , n89729 , n89730 , n89731 , 
 n89732 , n89733 , n89734 , n89735 , n89736 , n89737 , n89738 , n89739 , n89740 , n89741 , 
 n89742 , n89743 , n89744 , n89745 , n89746 , n89747 , n89748 , n89749 , n89750 , n89751 , 
 n89752 , n89753 , n89754 , n89755 , n89756 , n89757 , n89758 , n89759 , n89760 , n89761 , 
 n89762 , n89763 , n89764 , n89765 , n89766 , n89767 , n89768 , n89769 , n89770 , n89771 , 
 n89772 , n89773 , n89774 , n89775 , n89776 , n89777 , n89778 , n89779 , n89780 , n89781 , 
 n89782 , n89783 , n89784 , n89785 , n89786 , n89787 , n89788 , n89789 , n89790 , n89791 , 
 n89792 , n89793 , n89794 , n89795 , n89796 , n89797 , n89798 , n89799 , n89800 , n89801 , 
 n89802 , n89803 , n89804 , n89805 , n89806 , n89807 , n89808 , n89809 , n89810 , n89811 , 
 n89812 , n89813 , n89814 , n89815 , n89816 , n89817 , n89818 , n89819 , n89820 , n89821 , 
 n89822 , n89823 , n89824 , n89825 , n89826 , n89827 , n89828 , n89829 , n89830 , n89831 , 
 n89832 , n89833 , n89834 , n89835 , n89836 , n89837 , n89838 , n89839 , n89840 , n89841 , 
 n89842 , n89843 , n89844 , n89845 , n89846 , n89847 , n89848 , n89849 , n89850 , n89851 , 
 n89852 , n89853 , n89854 , n89855 , n89856 , n89857 , n89858 , n89859 , n89860 , n89861 , 
 n89862 , n89863 , n89864 , n89865 , n89866 , n89867 , n89868 , n89869 , n89870 , n89871 , 
 n89872 , n89873 , n89874 , n89875 , n89876 , n89877 , n89878 , n89879 , n89880 , n89881 , 
 n89882 , n89883 , n89884 , n89885 , n89886 , n89887 , n89888 , n89889 , n89890 , n89891 , 
 n89892 , n89893 , n89894 , n89895 , n89896 , n89897 , n89898 , n89899 , n89900 , n89901 , 
 n89902 , n89903 , n89904 , n89905 , n89906 , n89907 , n89908 , n89909 , n89910 , n89911 , 
 n89912 , n89913 , n89914 , n89915 , n89916 , n89917 , n89918 , n89919 , n89920 , n89921 , 
 n89922 , n89923 , n89924 , n89925 , n89926 , n89927 , n89928 , n89929 , n89930 , n89931 , 
 n89932 , n89933 , n89934 , n89935 , n89936 , n89937 , n89938 , n89939 , n89940 , n89941 , 
 n89942 , n89943 , n89944 , n89945 , n89946 , n89947 , n89948 , n89949 , n89950 , n89951 , 
 n89952 , n89953 , n89954 , n89955 , n89956 , n89957 , n89958 , n89959 , n89960 , n89961 , 
 n89962 , n89963 , n89964 , n89965 , n89966 , n89967 , n89968 , n89969 , n89970 , n89971 , 
 n89972 , n89973 , n89974 , n89975 , n89976 , n89977 , n89978 , n89979 , n89980 , n89981 , 
 n89982 , n89983 , n89984 , n89985 , n89986 , n89987 , n89988 , n89989 , n89990 , n89991 , 
 n89992 , n89993 , n89994 , n89995 , n89996 , n89997 , n89998 , n89999 , n90000 , n90001 , 
 n90002 , n90003 , n90004 , n90005 , n90006 , n90007 , n90008 , n90009 , n90010 , n90011 , 
 n90012 , n90013 , n90014 , n90015 , n90016 , n90017 , n90018 , n90019 , n90020 , n90021 , 
 n90022 , n90023 , n90024 , n90025 , n90026 , n90027 , n90028 , n90029 , n90030 , n90031 , 
 n90032 , n90033 , n90034 , n90035 , n90036 , n90037 , n90038 , n90039 , n90040 , n90041 , 
 n90042 , n90043 , n90044 , n90045 , n90046 , n90047 , n90048 , n90049 , n90050 , n90051 , 
 n90052 , n90053 , n90054 , n90055 , n90056 , n90057 , n90058 , n90059 , n90060 , n90061 , 
 n90062 , n90063 , n90064 , n90065 , n90066 , n90067 , n90068 , n90069 , n90070 , n90071 , 
 n90072 , n90073 , n90074 , n90075 , n90076 , n90077 , n90078 , n90079 , n90080 , n90081 , 
 n90082 , n90083 , n90084 , n90085 , n90086 , n90087 , n90088 , n90089 , n90090 , n90091 , 
 n90092 , n90093 , n90094 , n90095 , n90096 , n90097 , n90098 , n90099 , n90100 , n90101 , 
 n90102 , n90103 , n90104 , n90105 , n90106 , n90107 , n90108 , n90109 , n90110 , n90111 , 
 n90112 , n90113 , n90114 , n90115 , n90116 , n90117 , n90118 , n90119 , n90120 , n90121 , 
 n90122 , n90123 , n90124 , n90125 , n90126 , n90127 , n90128 , n90129 , n90130 , n90131 , 
 n90132 , n90133 , n90134 , n90135 , n90136 , n90137 , n90138 , n90139 , n90140 , n90141 , 
 n90142 , n90143 , n90144 , n90145 , n90146 , n90147 , n90148 , n90149 , n90150 , n90151 , 
 n90152 , n90153 , n90154 , n90155 , n90156 , n90157 , n90158 , n90159 , n90160 , n90161 , 
 n90162 , n90163 , n90164 , n90165 , n90166 , n90167 , n90168 , n90169 , n90170 , n90171 , 
 n90172 , n90173 , n90174 , n90175 , n90176 , n90177 , n90178 , n90179 , n90180 , n90181 , 
 n90182 , n90183 , n90184 , n90185 , n90186 , n90187 , n90188 , n90189 , n90190 , n90191 , 
 n90192 , n90193 , n90194 , n90195 , n90196 , n90197 , n90198 , n90199 , n90200 , n90201 , 
 n90202 , n90203 , n90204 , n90205 , n90206 , n90207 , n90208 , n90209 , n90210 , n90211 , 
 n90212 , n90213 , n90214 , n90215 , n90216 , n90217 , n90218 , n90219 , n90220 , n90221 , 
 n90222 , n90223 , n90224 , n90225 , n90226 , n90227 , n90228 , n90229 , n90230 , n90231 , 
 n90232 , n90233 , n90234 , n90235 , n90236 , n90237 , n90238 , n90239 , n90240 , n90241 , 
 n90242 , n90243 , n90244 , n90245 , n90246 , n90247 , n90248 , n90249 , n90250 , n90251 , 
 n90252 , n90253 , n90254 , n90255 , n90256 , n90257 , n90258 , n90259 , n90260 , n90261 , 
 n90262 , n90263 , n90264 , n90265 , n90266 , n90267 , n90268 , n90269 , n90270 , n90271 , 
 n90272 , n90273 , n90274 , n90275 , n90276 , n90277 , n90278 , n90279 , n90280 , n90281 , 
 n90282 , n90283 , n90284 , n90285 , n90286 , n90287 , n90288 , n90289 , n90290 , n90291 , 
 n90292 , n90293 , n90294 , n90295 , n90296 , n90297 , n90298 , n90299 , n90300 , n90301 , 
 n90302 , n90303 , n90304 , n90305 , n90306 , n90307 , n90308 , n90309 , n90310 , n90311 , 
 n90312 , n90313 , n90314 , n90315 , n90316 , n90317 , n90318 , n90319 , n90320 , n90321 , 
 n90322 , n90323 , n90324 , n90325 , n90326 , n90327 , n90328 , n90329 , n90330 , n90331 , 
 n90332 , n90333 , n90334 , n90335 , n90336 , n90337 , n90338 , n90339 , n90340 , n90341 , 
 n90342 , n90343 , n90344 , n90345 , n90346 , n90347 , n90348 , n90349 , n90350 , n90351 , 
 n90352 , n90353 , n90354 , n90355 , n90356 , n90357 , n90358 , n90359 , n90360 , n90361 , 
 n90362 , n90363 , n90364 , n90365 , n90366 , n90367 , n90368 , n90369 , n90370 , n90371 , 
 n90372 , n90373 , n90374 , n90375 , n90376 , n90377 , n90378 , n90379 , n90380 , n90381 , 
 n90382 , n90383 , n90384 , n90385 , n90386 , n90387 , n90388 , n90389 , n90390 , n90391 , 
 n90392 , n90393 , n90394 , n90395 , n90396 , n90397 , n90398 , n90399 , n90400 , n90401 , 
 n90402 , n90403 , n90404 , n90405 , n90406 , n90407 , n90408 , n90409 , n90410 , n90411 , 
 n90412 , n90413 , n90414 , n90415 , n90416 , n90417 , n90418 , n90419 , n90420 , n90421 , 
 n90422 , n90423 , n90424 , n90425 , n90426 , n90427 , n90428 , n90429 , n90430 , n90431 , 
 n90432 , n90433 , n90434 , n90435 , n90436 , n90437 , n90438 , n90439 , n90440 , n90441 , 
 n90442 , n90443 , n90444 , n90445 , n90446 , n90447 , n90448 , n90449 , n90450 , n90451 , 
 n90452 , n90453 , n90454 , n90455 , n90456 , n90457 , n90458 , n90459 , n90460 , n90461 , 
 n90462 , n90463 , n90464 , n90465 , n90466 , n90467 , n90468 , n90469 , n90470 , n90471 , 
 n90472 , n90473 , n90474 , n90475 , n90476 , n90477 , n90478 , n90479 , n90480 , n90481 , 
 n90482 , n90483 , n90484 , n90485 , n90486 , n90487 , n90488 , n90489 , n90490 , n90491 , 
 n90492 , n90493 , n90494 , n90495 , n90496 , n90497 , n90498 , n90499 , n90500 , n90501 , 
 n90502 , n90503 , n90504 , n90505 , n90506 , n90507 , n90508 , n90509 , n90510 , n90511 , 
 n90512 , n90513 , n90514 , n90515 , n90516 , n90517 , n90518 , n90519 , n90520 , n90521 , 
 n90522 , n90523 , n90524 , n90525 , n90526 , n90527 , n90528 , n90529 , n90530 , n90531 , 
 n90532 , n90533 , n90534 , n90535 , n90536 , n90537 , n90538 , n90539 , n90540 , n90541 , 
 n90542 , n90543 , n90544 , n90545 , n90546 , n90547 , n90548 , n90549 , n90550 , n90551 , 
 n90552 , n90553 , n90554 , n90555 , n90556 , n90557 , n90558 , n90559 , n90560 , n90561 , 
 n90562 , n90563 , n90564 , n90565 , n90566 , n90567 , n90568 , n90569 , n90570 , n90571 , 
 n90572 , n90573 , n90574 , n90575 , n90576 , n90577 , n90578 , n90579 , n90580 , n90581 , 
 n90582 , n90583 , n90584 , n90585 , n90586 , n90587 , n90588 , n90589 , n90590 , n90591 , 
 n90592 , n90593 , n90594 , n90595 , n90596 , n90597 , n90598 , n90599 , n90600 , n90601 , 
 n90602 , n90603 , n90604 , n90605 , n90606 , n90607 , n90608 , n90609 , n90610 , n90611 , 
 n90612 , n90613 , n90614 , n90615 , n90616 , n90617 , n90618 , n90619 , n90620 , n90621 , 
 n90622 , n90623 , n90624 , n90625 , n90626 , n90627 , n90628 , n90629 , n90630 , n90631 , 
 n90632 , n90633 , n90634 , n90635 , n90636 , n90637 , n90638 , n90639 , n90640 , n90641 , 
 n90642 , n90643 , n90644 , n90645 , n90646 , n90647 , n90648 , n90649 , n90650 , n90651 , 
 n90652 , n90653 , n90654 , n90655 , n90656 , n90657 , n90658 , n90659 , n90660 , n90661 , 
 n90662 , n90663 , n90664 , n90665 , n90666 , n90667 , n90668 , n90669 , n90670 , n90671 , 
 n90672 , n90673 , n90674 , n90675 , n90676 , n90677 , n90678 , n90679 , n90680 , n90681 , 
 n90682 , n90683 , n90684 , n90685 , n90686 , n90687 , n90688 , n90689 , n90690 , n90691 , 
 n90692 , n90693 , n90694 , n90695 , n90696 , n90697 , n90698 , n90699 , n90700 , n90701 , 
 n90702 , n90703 , n90704 , n90705 , n90706 , n90707 , n90708 , n90709 , n90710 , n90711 , 
 n90712 , n90713 , n90714 , n90715 , n90716 , n90717 , n90718 , n90719 , n90720 , n90721 , 
 n90722 , n90723 , n90724 , n90725 , n90726 , n90727 , n90728 , n90729 , n90730 , n90731 , 
 n90732 , n90733 , n90734 , n90735 , n90736 , n90737 , n90738 , n90739 , n90740 , n90741 , 
 n90742 , n90743 , n90744 , n90745 , n90746 , n90747 , n90748 , n90749 , n90750 , n90751 , 
 n90752 , n90753 , n90754 , n90755 , n90756 , n90757 , n90758 , n90759 , n90760 , n90761 , 
 n90762 , n90763 , n90764 , n90765 , n90766 , n90767 , n90768 , n90769 , n90770 , n90771 , 
 n90772 , n90773 , n90774 , n90775 , n90776 , n90777 , n90778 , n90779 , n90780 , n90781 , 
 n90782 , n90783 , n90784 , n90785 , n90786 , n90787 , n90788 , n90789 , n90790 , n90791 , 
 n90792 , n90793 , n90794 , n90795 , n90796 , n90797 , n90798 , n90799 , n90800 , n90801 , 
 n90802 , n90803 , n90804 , n90805 , n90806 , n90807 , n90808 , n90809 , n90810 , n90811 , 
 n90812 , n90813 , n90814 , n90815 , n90816 , n90817 , n90818 , n90819 , n90820 , n90821 , 
 n90822 , n90823 , n90824 , n90825 , n90826 , n90827 , n90828 , n90829 , n90830 , n90831 , 
 n90832 , n90833 , n90834 , n90835 , n90836 , n90837 , n90838 , n90839 , n90840 , n90841 , 
 n90842 , n90843 , n90844 , n90845 , n90846 , n90847 , n90848 , n90849 , n90850 , n90851 , 
 n90852 , n90853 , n90854 , n90855 , n90856 , n90857 , n90858 , n90859 , n90860 , n90861 , 
 n90862 , n90863 , n90864 , n90865 , n90866 , n90867 , n90868 , n90869 , n90870 , n90871 , 
 n90872 , n90873 , n90874 , n90875 , n90876 , n90877 , n90878 , n90879 , n90880 , n90881 , 
 n90882 , n90883 , n90884 , n90885 , n90886 , n90887 , n90888 , n90889 , n90890 , n90891 , 
 n90892 , n90893 , n90894 , n90895 , n90896 , n90897 , n90898 , n90899 , n90900 , n90901 , 
 n90902 , n90903 , n90904 , n90905 , n90906 , n90907 , n90908 , n90909 , n90910 , n90911 , 
 n90912 , n90913 , n90914 , n90915 , n90916 , n90917 , n90918 , n90919 , n90920 , n90921 , 
 n90922 , n90923 , n90924 , n90925 , n90926 , n90927 , n90928 , n90929 , n90930 , n90931 , 
 n90932 , n90933 , n90934 , n90935 , n90936 , n90937 , n90938 , n90939 , n90940 , n90941 , 
 n90942 , n90943 , n90944 , n90945 , n90946 , n90947 , n90948 , n90949 , n90950 , n90951 , 
 n90952 , n90953 , n90954 , n90955 , n90956 , n90957 , n90958 , n90959 , n90960 , n90961 , 
 n90962 , n90963 , n90964 , n90965 , n90966 , n90967 , n90968 , n90969 , n90970 , n90971 , 
 n90972 , n90973 , n90974 , n90975 , n90976 , n90977 , n90978 , n90979 , n90980 , n90981 , 
 n90982 , n90983 , n90984 , n90985 , n90986 , n90987 , n90988 , n90989 , n90990 , n90991 , 
 n90992 , n90993 , n90994 , n90995 , n90996 , n90997 , n90998 , n90999 , n91000 , n91001 , 
 n91002 , n91003 , n91004 , n91005 , n91006 , n91007 , n91008 , n91009 , n91010 , n91011 , 
 n91012 , n91013 , n91014 , n91015 , n91016 , n91017 , n91018 , n91019 , n91020 , n91021 , 
 n91022 , n91023 , n91024 , n91025 , n91026 , n91027 , n91028 , n91029 , n91030 , n91031 , 
 n91032 , n91033 , n91034 , n91035 , n91036 , n91037 , n91038 , n91039 , n91040 , n91041 , 
 n91042 , n91043 , n91044 , n91045 , n91046 , n91047 , n91048 , n91049 , n91050 , n91051 , 
 n91052 , n91053 , n91054 , n91055 , n91056 , n91057 , n91058 , n91059 , n91060 , n91061 , 
 n91062 , n91063 , n91064 , n91065 , n91066 , n91067 , n91068 , n91069 , n91070 , n91071 , 
 n91072 , n91073 , n91074 , n91075 , n91076 , n91077 , n91078 , n91079 , n91080 , n91081 , 
 n91082 , n91083 , n91084 , n91085 , n91086 , n91087 , n91088 , n91089 , n91090 , n91091 , 
 n91092 , n91093 , n91094 , n91095 , n91096 , n91097 , n91098 , n91099 , n91100 , n91101 , 
 n91102 , n91103 , n91104 , n91105 , n91106 , n91107 , n91108 , n91109 , n91110 , n91111 , 
 n91112 , n91113 , n91114 , n91115 , n91116 , n91117 , n91118 , n91119 , n91120 , n91121 , 
 n91122 , n91123 , n91124 , n91125 , n91126 , n91127 , n91128 , n91129 , n91130 , n91131 , 
 n91132 , n91133 , n91134 , n91135 , n91136 , n91137 , n91138 , n91139 , n91140 , n91141 , 
 n91142 , n91143 , n91144 , n91145 , n91146 , n91147 , n91148 , n91149 , n91150 , n91151 , 
 n91152 , n91153 , n91154 , n91155 , n91156 , n91157 , n91158 , n91159 , n91160 , n91161 , 
 n91162 , n91163 , n91164 , n91165 , n91166 , n91167 , n91168 , n91169 , n91170 , n91171 , 
 n91172 , n91173 , n91174 , n91175 , n91176 , n91177 , n91178 , n91179 , n91180 , n91181 , 
 n91182 , n91183 , n91184 , n91185 , n91186 , n91187 , n91188 , n91189 , n91190 , n91191 , 
 n91192 , n91193 , n91194 , n91195 , n91196 , n91197 , n91198 , n91199 , n91200 , n91201 , 
 n91202 , n91203 , n91204 , n91205 , n91206 , n91207 , n91208 , n91209 , n91210 , n91211 , 
 n91212 , n91213 , n91214 , n91215 , n91216 , n91217 , n91218 , n91219 , n91220 , n91221 , 
 n91222 , n91223 , n91224 , n91225 , n91226 , n91227 , n91228 , n91229 , n91230 , n91231 , 
 n91232 , n91233 , n91234 , n91235 , n91236 , n91237 , n91238 , n91239 , n91240 , n91241 , 
 n91242 , n91243 , n91244 , n91245 , n91246 , n91247 , n91248 , n91249 , n91250 , n91251 , 
 n91252 , n91253 , n91254 , n91255 , n91256 , n91257 , n91258 , n91259 , n91260 , n91261 , 
 n91262 , n91263 , n91264 , n91265 , n91266 , n91267 , n91268 , n91269 , n91270 , n91271 , 
 n91272 , n91273 , n91274 , n91275 , n91276 , n91277 , n91278 , n91279 , n91280 , n91281 , 
 n91282 , n91283 , n91284 , n91285 , n91286 , n91287 , n91288 , n91289 , n91290 , n91291 , 
 n91292 , n91293 , n91294 , n91295 , n91296 , n91297 , n91298 , n91299 , n91300 , n91301 , 
 n91302 , n91303 , n91304 , n91305 , n91306 , n91307 , n91308 , n91309 , n91310 , n91311 , 
 n91312 , n91313 , n91314 , n91315 , n91316 , n91317 , n91318 , n91319 , n91320 , n91321 , 
 n91322 , n91323 , n91324 , n91325 , n91326 , n91327 , n91328 , n91329 , n91330 , n91331 , 
 n91332 , n91333 , n91334 , n91335 , n91336 , n91337 , n91338 , n91339 , n91340 , n91341 , 
 n91342 , n91343 , n91344 , n91345 , n91346 , n91347 , n91348 , n91349 , n91350 , n91351 , 
 n91352 , n91353 , n91354 , n91355 , n91356 , n91357 , n91358 , n91359 , n91360 , n91361 , 
 n91362 , n91363 , n91364 , n91365 , n91366 , n91367 , n91368 , n91369 , n91370 , n91371 , 
 n91372 , n91373 , n91374 , n91375 , n91376 , n91377 , n91378 , n91379 , n91380 , n91381 , 
 n91382 , n91383 , n91384 , n91385 , n91386 , n91387 , n91388 , n91389 , n91390 , n91391 , 
 n91392 , n91393 , n91394 , n91395 , n91396 , n91397 , n91398 , n91399 , n91400 , n91401 , 
 n91402 , n91403 , n91404 , n91405 , n91406 , n91407 , n91408 , n91409 , n91410 , n91411 , 
 n91412 , n91413 , n91414 , n91415 , n91416 , n91417 , n91418 , n91419 , n91420 , n91421 , 
 n91422 , n91423 , n91424 , n91425 , n91426 , n91427 , n91428 , n91429 , n91430 , n91431 , 
 n91432 , n91433 , n91434 , n91435 , n91436 , n91437 , n91438 , n91439 , n91440 , n91441 , 
 n91442 , n91443 , n91444 , n91445 , n91446 , n91447 , n91448 , n91449 , n91450 , n91451 , 
 n91452 , n91453 , n91454 , n91455 , n91456 , n91457 , n91458 , n91459 , n91460 , n91461 , 
 n91462 , n91463 , n91464 , n91465 , n91466 , n91467 , n91468 , n91469 , n91470 , n91471 , 
 n91472 , n91473 , n91474 , n91475 , n91476 , n91477 , n91478 , n91479 , n91480 , n91481 , 
 n91482 , n91483 , n91484 , n91485 , n91486 , n91487 , n91488 , n91489 , n91490 , n91491 , 
 n91492 , n91493 , n91494 , n91495 , n91496 , n91497 , n91498 , n91499 , n91500 , n91501 , 
 n91502 , n91503 , n91504 , n91505 , n91506 , n91507 , n91508 , n91509 , n91510 , n91511 , 
 n91512 , n91513 , n91514 , n91515 , n91516 , n91517 , n91518 , n91519 , n91520 , n91521 , 
 n91522 , n91523 , n91524 , n91525 , n91526 , n91527 , n91528 , n91529 , n91530 , n91531 , 
 n91532 , n91533 , n91534 , n91535 , n91536 , n91537 , n91538 , n91539 , n91540 , n91541 , 
 n91542 , n91543 , n91544 , n91545 , n91546 , n91547 , n91548 , n91549 , n91550 , n91551 , 
 n91552 , n91553 , n91554 , n91555 , n91556 , n91557 , n91558 , n91559 , n91560 , n91561 , 
 n91562 , n91563 , n91564 , n91565 , n91566 , n91567 , n91568 , n91569 , n91570 , n91571 , 
 n91572 , n91573 , n91574 , n91575 , n91576 , n91577 , n91578 , n91579 , n91580 , n91581 , 
 n91582 , n91583 , n91584 , n91585 , n91586 , n91587 , n91588 , n91589 , n91590 , n91591 , 
 n91592 , n91593 , n91594 , n91595 , n91596 , n91597 , n91598 , n91599 , n91600 , n91601 , 
 n91602 , n91603 , n91604 , n91605 , n91606 , n91607 , n91608 , n91609 , n91610 , n91611 , 
 n91612 , n91613 , n91614 , n91615 , n91616 , n91617 , n91618 , n91619 , n91620 , n91621 , 
 n91622 , n91623 , n91624 , n91625 , n91626 , n91627 , n91628 , n91629 , n91630 , n91631 , 
 n91632 , n91633 , n91634 , n91635 , n91636 , n91637 , n91638 , n91639 , n91640 , n91641 , 
 n91642 , n91643 , n91644 , n91645 , n91646 , n91647 , n91648 , n91649 , n91650 , n91651 , 
 n91652 , n91653 , n91654 , n91655 , n91656 , n91657 , n91658 , n91659 , n91660 , n91661 , 
 n91662 , n91663 , n91664 , n91665 , n91666 , n91667 , n91668 , n91669 , n91670 , n91671 , 
 n91672 , n91673 , n91674 , n91675 , n91676 , n91677 , n91678 , n91679 , n91680 , n91681 , 
 n91682 , n91683 , n91684 , n91685 , n91686 , n91687 , n91688 , n91689 , n91690 , n91691 , 
 n91692 , n91693 , n91694 , n91695 , n91696 , n91697 , n91698 , n91699 , n91700 , n91701 , 
 n91702 , n91703 , n91704 , n91705 , n91706 , n91707 , n91708 , n91709 , n91710 , n91711 , 
 n91712 , n91713 , n91714 , n91715 , n91716 , n91717 , n91718 , n91719 , n91720 , n91721 , 
 n91722 , n91723 , n91724 , n91725 , n91726 , n91727 , n91728 , n91729 , n91730 , n91731 , 
 n91732 , n91733 , n91734 , n91735 , n91736 , n91737 , n91738 , n91739 , n91740 , n91741 , 
 n91742 , n91743 , n91744 , n91745 , n91746 , n91747 , n91748 , n91749 , n91750 , n91751 , 
 n91752 , n91753 , n91754 , n91755 , n91756 , n91757 , n91758 , n91759 , n91760 , n91761 , 
 n91762 , n91763 , n91764 , n91765 , n91766 , n91767 , n91768 , n91769 , n91770 , n91771 , 
 n91772 , n91773 , n91774 , n91775 , n91776 , n91777 , n91778 , n91779 , n91780 , n91781 , 
 n91782 , n91783 , n91784 , n91785 , n91786 , n91787 , n91788 , n91789 , n91790 , n91791 , 
 n91792 , n91793 , n91794 , n91795 , n91796 , n91797 , n91798 , n91799 , n91800 , n91801 , 
 n91802 , n91803 , n91804 , n91805 , n91806 , n91807 , n91808 , n91809 , n91810 , n91811 , 
 n91812 , n91813 , n91814 , n91815 , n91816 , n91817 , n91818 , n91819 , n91820 , n91821 , 
 n91822 , n91823 , n91824 , n91825 , n91826 , n91827 , n91828 , n91829 , n91830 , n91831 , 
 n91832 , n91833 , n91834 , n91835 , n91836 , n91837 , n91838 , n91839 , n91840 , n91841 , 
 n91842 , n91843 , n91844 , n91845 , n91846 , n91847 , n91848 , n91849 , n91850 , n91851 , 
 n91852 , n91853 , n91854 , n91855 , n91856 , n91857 , n91858 , n91859 , n91860 , n91861 , 
 n91862 , n91863 , n91864 , n91865 , n91866 , n91867 , n91868 , n91869 , n91870 , n91871 , 
 n91872 , n91873 , n91874 , n91875 , n91876 , n91877 , n91878 , n91879 , n91880 , n91881 , 
 n91882 , n91883 , n91884 , n91885 , n91886 , n91887 , n91888 , n91889 , n91890 , n91891 , 
 n91892 , n91893 , n91894 , n91895 , n91896 , n91897 , n91898 , n91899 , n91900 , n91901 , 
 n91902 , n91903 , n91904 , n91905 , n91906 , n91907 , n91908 , n91909 , n91910 , n91911 , 
 n91912 , n91913 , n91914 , n91915 , n91916 , n91917 , n91918 , n91919 , n91920 , n91921 , 
 n91922 , n91923 , n91924 , n91925 , n91926 , n91927 , n91928 , n91929 , n91930 , n91931 , 
 n91932 , n91933 , n91934 , n91935 , n91936 , n91937 , n91938 , n91939 , n91940 , n91941 , 
 n91942 , n91943 , n91944 , n91945 , n91946 , n91947 , n91948 , n91949 , n91950 , n91951 , 
 n91952 , n91953 , n91954 , n91955 , n91956 , n91957 , n91958 , n91959 , n91960 , n91961 , 
 n91962 , n91963 , n91964 , n91965 , n91966 , n91967 , n91968 , n91969 , n91970 , n91971 , 
 n91972 , n91973 , n91974 , n91975 , n91976 , n91977 , n91978 , n91979 , n91980 , n91981 , 
 n91982 , n91983 , n91984 , n91985 , n91986 , n91987 , n91988 , n91989 , n91990 , n91991 , 
 n91992 , n91993 , n91994 , n91995 , n91996 , n91997 , n91998 , n91999 , n92000 , n92001 , 
 n92002 , n92003 , n92004 , n92005 , n92006 , n92007 , n92008 , n92009 , n92010 , n92011 , 
 n92012 , n92013 , n92014 , n92015 , n92016 , n92017 , n92018 , n92019 , n92020 , n92021 , 
 n92022 , n92023 , n92024 , n92025 , n92026 , n92027 , n92028 , n92029 , n92030 , n92031 , 
 n92032 , n92033 , n92034 , n92035 , n92036 , n92037 , n92038 , n92039 , n92040 , n92041 , 
 n92042 , n92043 , n92044 , n92045 , n92046 , n92047 , n92048 , n92049 , n92050 , n92051 , 
 n92052 , n92053 , n92054 , n92055 , n92056 , n92057 , n92058 , n92059 , n92060 , n92061 , 
 n92062 , n92063 , n92064 , n92065 , n92066 , n92067 , n92068 , n92069 , n92070 , n92071 , 
 n92072 , n92073 , n92074 , n92075 , n92076 , n92077 , n92078 , n92079 , n92080 , n92081 , 
 n92082 , n92083 , n92084 , n92085 , n92086 , n92087 , n92088 , n92089 , n92090 , n92091 , 
 n92092 , n92093 , n92094 , n92095 , n92096 , n92097 , n92098 , n92099 , n92100 , n92101 , 
 n92102 , n92103 , n92104 , n92105 , n92106 , n92107 , n92108 , n92109 , n92110 , n92111 , 
 n92112 , n92113 , n92114 , n92115 , n92116 , n92117 , n92118 , n92119 , n92120 , n92121 , 
 n92122 , n92123 , n92124 , n92125 , n92126 , n92127 , n92128 , n92129 , n92130 , n92131 , 
 n92132 , n92133 , n92134 , n92135 , n92136 , n92137 , n92138 , n92139 , n92140 , n92141 , 
 n92142 , n92143 , n92144 , n92145 , n92146 , n92147 , n92148 , n92149 , n92150 , n92151 , 
 n92152 , n92153 , n92154 , n92155 , n92156 , n92157 , n92158 , n92159 , n92160 , n92161 , 
 n92162 , n92163 , n92164 , n92165 , n92166 , n92167 , n92168 , n92169 , n92170 , n92171 , 
 n92172 , n92173 , n92174 , n92175 , n92176 , n92177 , n92178 , n92179 , n92180 , n92181 , 
 n92182 , n92183 , n92184 , n92185 , n92186 , n92187 , n92188 , n92189 , n92190 , n92191 , 
 n92192 , n92193 , n92194 , n92195 , n92196 , n92197 , n92198 , n92199 , n92200 , n92201 , 
 n92202 , n92203 , n92204 , n92205 , n92206 , n92207 , n92208 , n92209 , n92210 , n92211 , 
 n92212 , n92213 , n92214 , n92215 , n92216 , n92217 , n92218 , n92219 , n92220 , n92221 , 
 n92222 , n92223 , n92224 , n92225 , n92226 , n92227 , n92228 , n92229 , n92230 , n92231 , 
 n92232 , n92233 , n92234 , n92235 , n92236 , n92237 , n92238 , n92239 , n92240 , n92241 , 
 n92242 , n92243 , n92244 , n92245 , n92246 , n92247 , n92248 , n92249 , n92250 , n92251 , 
 n92252 , n92253 , n92254 , n92255 , n92256 , n92257 , n92258 , n92259 , n92260 , n92261 , 
 n92262 , n92263 , n92264 , n92265 , n92266 , n92267 , n92268 , n92269 , n92270 , n92271 , 
 n92272 , n92273 , n92274 , n92275 , n92276 , n92277 , n92278 , n92279 , n92280 , n92281 , 
 n92282 , n92283 , n92284 , n92285 , n92286 , n92287 , n92288 , n92289 , n92290 , n92291 , 
 n92292 , n92293 , n92294 , n92295 , n92296 , n92297 , n92298 , n92299 , n92300 , n92301 , 
 n92302 , n92303 , n92304 , n92305 , n92306 , n92307 , n92308 , n92309 , n92310 , n92311 , 
 n92312 , n92313 , n92314 , n92315 , n92316 , n92317 , n92318 , n92319 , n92320 , n92321 , 
 n92322 , n92323 , n92324 , n92325 , n92326 , n92327 , n92328 , n92329 , n92330 , n92331 , 
 n92332 , n92333 , n92334 , n92335 , n92336 , n92337 , n92338 , n92339 , n92340 , n92341 , 
 n92342 , n92343 , n92344 , n92345 , n92346 , n92347 , n92348 , n92349 , n92350 , n92351 , 
 n92352 , n92353 , n92354 , n92355 , n92356 , n92357 , n92358 , n92359 , n92360 , n92361 , 
 n92362 , n92363 , n92364 , n92365 , n92366 , n92367 , n92368 , n92369 , n92370 , n92371 , 
 n92372 , n92373 , n92374 , n92375 , n92376 , n92377 , n92378 , n92379 , n92380 , n92381 , 
 n92382 , n92383 , n92384 , n92385 , n92386 , n92387 , n92388 , n92389 , n92390 , n92391 , 
 n92392 , n92393 , n92394 , n92395 , n92396 , n92397 , n92398 , n92399 , n92400 , n92401 , 
 n92402 , n92403 , n92404 , n92405 , n92406 , n92407 , n92408 , n92409 , n92410 , n92411 , 
 n92412 , n92413 , n92414 , n92415 , n92416 , n92417 , n92418 , n92419 , n92420 , n92421 , 
 n92422 , n92423 , n92424 , n92425 , n92426 , n92427 , n92428 , n92429 , n92430 , n92431 , 
 n92432 , n92433 , n92434 , n92435 , n92436 , n92437 , n92438 , n92439 , n92440 , n92441 , 
 n92442 , n92443 , n92444 , n92445 , n92446 , n92447 , n92448 , n92449 , n92450 , n92451 , 
 n92452 , n92453 , n92454 , n92455 , n92456 , n92457 , n92458 , n92459 , n92460 , n92461 , 
 n92462 , n92463 , n92464 , n92465 , n92466 , n92467 , n92468 , n92469 , n92470 , n92471 , 
 n92472 , n92473 , n92474 , n92475 , n92476 , n92477 , n92478 , n92479 , n92480 , n92481 , 
 n92482 , n92483 , n92484 , n92485 , n92486 , n92487 , n92488 , n92489 , n92490 , n92491 , 
 n92492 , n92493 , n92494 , n92495 , n92496 , n92497 , n92498 , n92499 , n92500 , n92501 , 
 n92502 , n92503 , n92504 , n92505 , n92506 , n92507 , n92508 , n92509 , n92510 , n92511 , 
 n92512 , n92513 , n92514 , n92515 , n92516 , n92517 , n92518 , n92519 , n92520 , n92521 , 
 n92522 , n92523 , n92524 , n92525 , n92526 , n92527 , n92528 , n92529 , n92530 , n92531 , 
 n92532 , n92533 , n92534 , n92535 , n92536 , n92537 , n92538 , n92539 , n92540 , n92541 , 
 n92542 , n92543 , n92544 , n92545 , n92546 , n92547 , n92548 , n92549 , n92550 , n92551 , 
 n92552 , n92553 , n92554 , n92555 , n92556 , n92557 , n92558 , n92559 , n92560 , n92561 , 
 n92562 , n92563 , n92564 , n92565 , n92566 , n92567 , n92568 , n92569 , n92570 , n92571 , 
 n92572 , n92573 , n92574 , n92575 , n92576 , n92577 , n92578 , n92579 , n92580 , n92581 , 
 n92582 , n92583 , n92584 , n92585 , n92586 , n92587 , n92588 , n92589 , n92590 , n92591 , 
 n92592 , n92593 , n92594 , n92595 , n92596 , n92597 , n92598 , n92599 , n92600 , n92601 , 
 n92602 , n92603 , n92604 , n92605 , n92606 , n92607 , n92608 , n92609 , n92610 , n92611 , 
 n92612 , n92613 , n92614 , n92615 , n92616 , n92617 , n92618 , n92619 , n92620 , n92621 , 
 n92622 , n92623 , n92624 , n92625 , n92626 , n92627 , n92628 , n92629 , n92630 , n92631 , 
 n92632 , n92633 , n92634 , n92635 , n92636 , n92637 , n92638 , n92639 , n92640 , n92641 , 
 n92642 , n92643 , n92644 , n92645 , n92646 , n92647 , n92648 , n92649 , n92650 , n92651 , 
 n92652 , n92653 , n92654 , n92655 , n92656 , n92657 , n92658 , n92659 , n92660 , n92661 , 
 n92662 , n92663 , n92664 , n92665 , n92666 , n92667 , n92668 , n92669 , n92670 , n92671 , 
 n92672 , n92673 , n92674 , n92675 , n92676 , n92677 , n92678 , n92679 , n92680 , n92681 , 
 n92682 , n92683 , n92684 , n92685 , n92686 , n92687 , n92688 , n92689 , n92690 , n92691 , 
 n92692 , n92693 , n92694 , n92695 , n92696 , n92697 , n92698 , n92699 , n92700 , n92701 , 
 n92702 , n92703 , n92704 , n92705 , n92706 , n92707 , n92708 , n92709 , n92710 , n92711 , 
 n92712 , n92713 , n92714 , n92715 , n92716 , n92717 , n92718 , n92719 , n92720 , n92721 , 
 n92722 , n92723 , n92724 , n92725 , n92726 , n92727 , n92728 , n92729 , n92730 , n92731 , 
 n92732 , n92733 , n92734 , n92735 , n92736 , n92737 , n92738 , n92739 , n92740 , n92741 , 
 n92742 , n92743 , n92744 , n92745 , n92746 , n92747 , n92748 , n92749 , n92750 , n92751 , 
 n92752 , n92753 , n92754 , n92755 , n92756 , n92757 , n92758 , n92759 , n92760 , n92761 , 
 n92762 , n92763 , n92764 , n92765 , n92766 , n92767 , n92768 , n92769 , n92770 , n92771 , 
 n92772 , n92773 , n92774 , n92775 , n92776 , n92777 , n92778 , n92779 , n92780 , n92781 , 
 n92782 , n92783 , n92784 , n92785 , n92786 , n92787 , n92788 , n92789 , n92790 , n92791 , 
 n92792 , n92793 , n92794 , n92795 , n92796 , n92797 , n92798 , n92799 , n92800 , n92801 , 
 n92802 , n92803 , n92804 , n92805 , n92806 , n92807 , n92808 , n92809 , n92810 , n92811 , 
 n92812 , n92813 , n92814 , n92815 , n92816 , n92817 , n92818 , n92819 , n92820 , n92821 , 
 n92822 , n92823 , n92824 , n92825 , n92826 , n92827 , n92828 , n92829 , n92830 , n92831 , 
 n92832 , n92833 , n92834 , n92835 , n92836 , n92837 , n92838 , n92839 , n92840 , n92841 , 
 n92842 , n92843 , n92844 , n92845 , n92846 , n92847 , n92848 , n92849 , n92850 , n92851 , 
 n92852 , n92853 , n92854 , n92855 , n92856 , n92857 , n92858 , n92859 , n92860 , n92861 , 
 n92862 , n92863 , n92864 , n92865 , n92866 , n92867 , n92868 , n92869 , n92870 , n92871 , 
 n92872 , n92873 , n92874 , n92875 , n92876 , n92877 , n92878 , n92879 , n92880 , n92881 , 
 n92882 , n92883 , n92884 , n92885 , n92886 , n92887 , n92888 , n92889 , n92890 , n92891 , 
 n92892 , n92893 , n92894 , n92895 , n92896 , n92897 , n92898 , n92899 , n92900 , n92901 , 
 n92902 , n92903 , n92904 , n92905 , n92906 , n92907 , n92908 , n92909 , n92910 , n92911 , 
 n92912 , n92913 , n92914 , n92915 , n92916 , n92917 , n92918 , n92919 , n92920 , n92921 , 
 n92922 , n92923 , n92924 , n92925 , n92926 , n92927 , n92928 , n92929 , n92930 , n92931 , 
 n92932 , n92933 , n92934 , n92935 , n92936 , n92937 , n92938 , n92939 , n92940 , n92941 , 
 n92942 , n92943 , n92944 , n92945 , n92946 , n92947 , n92948 , n92949 , n92950 , n92951 , 
 n92952 , n92953 , n92954 , n92955 , n92956 , n92957 , n92958 , n92959 , n92960 , n92961 , 
 n92962 , n92963 , n92964 , n92965 , n92966 , n92967 , n92968 , n92969 , n92970 , n92971 , 
 n92972 , n92973 , n92974 , n92975 , n92976 , n92977 , n92978 , n92979 , n92980 , n92981 , 
 n92982 , n92983 , n92984 , n92985 , n92986 , n92987 , n92988 , n92989 , n92990 , n92991 , 
 n92992 , n92993 , n92994 , n92995 , n92996 , n92997 , n92998 , n92999 , n93000 , n93001 , 
 n93002 , n93003 , n93004 , n93005 , n93006 , n93007 , n93008 , n93009 , n93010 , n93011 , 
 n93012 , n93013 , n93014 , n93015 , n93016 , n93017 , n93018 , n93019 , n93020 , n93021 , 
 n93022 , n93023 , n93024 , n93025 , n93026 , n93027 , n93028 , n93029 , n93030 , n93031 , 
 n93032 , n93033 , n93034 , n93035 , n93036 , n93037 , n93038 , n93039 , n93040 , n93041 , 
 n93042 , n93043 , n93044 , n93045 , n93046 , n93047 , n93048 , n93049 , n93050 , n93051 , 
 n93052 , n93053 , n93054 , n93055 , n93056 , n93057 , n93058 , n93059 , n93060 , n93061 , 
 n93062 , n93063 , n93064 , n93065 , n93066 , n93067 , n93068 , n93069 , n93070 , n93071 , 
 n93072 , n93073 , n93074 , n93075 , n93076 , n93077 , n93078 , n93079 , n93080 , n93081 , 
 n93082 , n93083 , n93084 , n93085 , n93086 , n93087 , n93088 , n93089 , n93090 , n93091 , 
 n93092 , n93093 , n93094 , n93095 , n93096 , n93097 , n93098 , n93099 , n93100 , n93101 , 
 n93102 , n93103 , n93104 , n93105 , n93106 , n93107 , n93108 , n93109 , n93110 , n93111 , 
 n93112 , n93113 , n93114 , n93115 , n93116 , n93117 , n93118 , n93119 , n93120 , n93121 , 
 n93122 , n93123 , n93124 , n93125 , n93126 , n93127 , n93128 , n93129 , n93130 , n93131 , 
 n93132 , n93133 , n93134 , n93135 , n93136 , n93137 , n93138 , n93139 , n93140 , n93141 , 
 n93142 , n93143 , n93144 , n93145 , n93146 , n93147 , n93148 , n93149 , n93150 , n93151 , 
 n93152 , n93153 , n93154 , n93155 , n93156 , n93157 , n93158 , n93159 , n93160 , n93161 , 
 n93162 , n93163 , n93164 , n93165 , n93166 , n93167 , n93168 , n93169 , n93170 , n93171 , 
 n93172 , n93173 , n93174 , n93175 , n93176 , n93177 , n93178 , n93179 , n93180 , n93181 , 
 n93182 , n93183 , n93184 , n93185 , n93186 , n93187 , n93188 , n93189 , n93190 , n93191 , 
 n93192 , n93193 , n93194 , n93195 , n93196 , n93197 , n93198 , n93199 , n93200 , n93201 , 
 n93202 , n93203 , n93204 , n93205 , n93206 , n93207 , n93208 , n93209 , n93210 , n93211 , 
 n93212 , n93213 , n93214 , n93215 , n93216 , n93217 , n93218 , n93219 , n93220 , n93221 , 
 n93222 , n93223 , n93224 , n93225 , n93226 , n93227 , n93228 , n93229 , n93230 , n93231 , 
 n93232 , n93233 , n93234 , n93235 , n93236 , n93237 , n93238 , n93239 , n93240 , n93241 , 
 n93242 , n93243 , n93244 , n93245 , n93246 , n93247 , n93248 , n93249 , n93250 , n93251 , 
 n93252 , n93253 , n93254 , n93255 , n93256 , n93257 , n93258 , n93259 , n93260 , n93261 , 
 n93262 , n93263 , n93264 , n93265 , n93266 , n93267 , n93268 , n93269 , n93270 , n93271 , 
 n93272 , n93273 , n93274 , n93275 , n93276 , n93277 , n93278 , n93279 , n93280 , n93281 , 
 n93282 , n93283 , n93284 , n93285 , n93286 , n93287 , n93288 , n93289 , n93290 , n93291 , 
 n93292 , n93293 , n93294 , n93295 , n93296 , n93297 , n93298 , n93299 , n93300 , n93301 , 
 n93302 , n93303 , n93304 , n93305 , n93306 , n93307 , n93308 , n93309 , n93310 , n93311 , 
 n93312 , n93313 , n93314 , n93315 , n93316 , n93317 , n93318 , n93319 , n93320 , n93321 , 
 n93322 , n93323 , n93324 , n93325 , n93326 , n93327 , n93328 , n93329 , n93330 , n93331 , 
 n93332 , n93333 , n93334 , n93335 , n93336 , n93337 , n93338 , n93339 , n93340 , n93341 , 
 n93342 , n93343 , n93344 , n93345 , n93346 , n93347 , n93348 , n93349 , n93350 , n93351 , 
 n93352 , n93353 , n93354 , n93355 , n93356 , n93357 , n93358 , n93359 , n93360 , n93361 , 
 n93362 , n93363 , n93364 , n93365 , n93366 , n93367 , n93368 , n93369 , n93370 , n93371 , 
 n93372 , n93373 , n93374 , n93375 , n93376 , n93377 , n93378 , n93379 , n93380 , n93381 , 
 n93382 , n93383 , n93384 , n93385 , n93386 , n93387 , n93388 , n93389 , n93390 , n93391 , 
 n93392 , n93393 , n93394 , n93395 , n93396 , n93397 , n93398 , n93399 , n93400 , n93401 , 
 n93402 , n93403 , n93404 , n93405 , n93406 , n93407 , n93408 , n93409 , n93410 , n93411 , 
 n93412 , n93413 , n93414 , n93415 , n93416 , n93417 , n93418 , n93419 , n93420 , n93421 , 
 n93422 , n93423 , n93424 , n93425 , n93426 , n93427 , n93428 , n93429 , n93430 , n93431 , 
 n93432 , n93433 , n93434 , n93435 , n93436 , n93437 , n93438 , n93439 , n93440 , n93441 , 
 n93442 , n93443 , n93444 , n93445 , n93446 , n93447 , n93448 , n93449 , n93450 , n93451 , 
 n93452 , n93453 , n93454 , n93455 , n93456 , n93457 , n93458 , n93459 , n93460 , n93461 , 
 n93462 , n93463 , n93464 , n93465 , n93466 , n93467 , n93468 , n93469 , n93470 , n93471 , 
 n93472 , n93473 , n93474 , n93475 , n93476 , n93477 , n93478 , n93479 , n93480 , n93481 , 
 n93482 , n93483 , n93484 , n93485 , n93486 , n93487 , n93488 , n93489 , n93490 , n93491 , 
 n93492 , n93493 , n93494 , n93495 , n93496 , n93497 , n93498 , n93499 , n93500 , n93501 , 
 n93502 , n93503 , n93504 , n93505 , n93506 , n93507 , n93508 , n93509 , n93510 , n93511 , 
 n93512 , n93513 , n93514 , n93515 , n93516 , n93517 , n93518 , n93519 , n93520 , n93521 , 
 n93522 , n93523 , n93524 , n93525 , n93526 , n93527 , n93528 , n93529 , n93530 , n93531 , 
 n93532 , n93533 , n93534 , n93535 , n93536 , n93537 , n93538 , n93539 , n93540 , n93541 , 
 n93542 , n93543 , n93544 , n93545 , n93546 , n93547 , n93548 , n93549 , n93550 , n93551 , 
 n93552 , n93553 , n93554 , n93555 , n93556 , n93557 , n93558 , n93559 , n93560 , n93561 , 
 n93562 , n93563 , n93564 , n93565 , n93566 , n93567 , n93568 , n93569 , n93570 , n93571 , 
 n93572 , n93573 , n93574 , n93575 , n93576 , n93577 , n93578 , n93579 , n93580 , n93581 , 
 n93582 , n93583 , n93584 , n93585 , n93586 , n93587 , n93588 , n93589 , n93590 , n93591 , 
 n93592 , n93593 , n93594 , n93595 , n93596 , n93597 , n93598 , n93599 , n93600 , n93601 , 
 n93602 , n93603 , n93604 , n93605 , n93606 , n93607 , n93608 , n93609 , n93610 , n93611 , 
 n93612 , n93613 , n93614 , n93615 , n93616 , n93617 , n93618 , n93619 , n93620 , n93621 , 
 n93622 , n93623 , n93624 , n93625 , n93626 , n93627 , n93628 , n93629 , n93630 , n93631 , 
 n93632 , n93633 , n93634 , n93635 , n93636 , n93637 , n93638 , n93639 , n93640 , n93641 , 
 n93642 , n93643 , n93644 , n93645 , n93646 , n93647 , n93648 , n93649 , n93650 , n93651 , 
 n93652 , n93653 , n93654 , n93655 , n93656 , n93657 , n93658 , n93659 , n93660 , n93661 , 
 n93662 , n93663 , n93664 , n93665 , n93666 , n93667 , n93668 , n93669 , n93670 , n93671 , 
 n93672 , n93673 , n93674 , n93675 , n93676 , n93677 , n93678 , n93679 , n93680 , n93681 , 
 n93682 , n93683 , n93684 , n93685 , n93686 , n93687 , n93688 , n93689 , n93690 , n93691 , 
 n93692 , n93693 , n93694 , n93695 , n93696 , n93697 , n93698 , n93699 , n93700 , n93701 , 
 n93702 , n93703 , n93704 , n93705 , n93706 , n93707 , n93708 , n93709 , n93710 , n93711 , 
 n93712 , n93713 , n93714 , n93715 , n93716 , n93717 , n93718 , n93719 , n93720 , n93721 , 
 n93722 , n93723 , n93724 , n93725 , n93726 , n93727 , n93728 , n93729 , n93730 , n93731 , 
 n93732 , n93733 , n93734 , n93735 , n93736 , n93737 , n93738 , n93739 , n93740 , n93741 , 
 n93742 , n93743 , n93744 , n93745 , n93746 , n93747 , n93748 , n93749 , n93750 , n93751 , 
 n93752 , n93753 , n93754 , n93755 , n93756 , n93757 , n93758 , n93759 , n93760 , n93761 , 
 n93762 , n93763 , n93764 , n93765 , n93766 , n93767 , n93768 , n93769 , n93770 , n93771 , 
 n93772 , n93773 , n93774 , n93775 , n93776 , n93777 , n93778 , n93779 , n93780 , n93781 , 
 n93782 , n93783 , n93784 , n93785 , n93786 , n93787 , n93788 , n93789 , n93790 , n93791 , 
 n93792 , n93793 , n93794 , n93795 , n93796 , n93797 , n93798 , n93799 , n93800 , n93801 , 
 n93802 , n93803 , n93804 , n93805 , n93806 , n93807 , n93808 , n93809 , n93810 , n93811 , 
 n93812 , n93813 , n93814 , n93815 , n93816 , n93817 , n93818 , n93819 , n93820 , n93821 , 
 n93822 , n93823 , n93824 , n93825 , n93826 , n93827 , n93828 , n93829 , n93830 , n93831 , 
 n93832 , n93833 , n93834 , n93835 , n93836 , n93837 , n93838 , n93839 , n93840 , n93841 , 
 n93842 , n93843 , n93844 , n93845 , n93846 , n93847 , n93848 , n93849 , n93850 , n93851 , 
 n93852 , n93853 , n93854 , n93855 , n93856 , n93857 , n93858 , n93859 , n93860 , n93861 , 
 n93862 , n93863 , n93864 , n93865 , n93866 , n93867 , n93868 , n93869 , n93870 , n93871 , 
 n93872 , n93873 , n93874 , n93875 , n93876 , n93877 , n93878 , n93879 , n93880 , n93881 , 
 n93882 , n93883 , n93884 , n93885 , n93886 , n93887 , n93888 , n93889 , n93890 , n93891 , 
 n93892 , n93893 , n93894 , n93895 , n93896 , n93897 , n93898 , n93899 , n93900 , n93901 , 
 n93902 , n93903 , n93904 , n93905 , n93906 , n93907 , n93908 , n93909 , n93910 , n93911 , 
 n93912 , n93913 , n93914 , n93915 , n93916 , n93917 , n93918 , n93919 , n93920 , n93921 , 
 n93922 , n93923 , n93924 , n93925 , n93926 , n93927 , n93928 , n93929 , n93930 , n93931 , 
 n93932 , n93933 , n93934 , n93935 , n93936 , n93937 , n93938 , n93939 , n93940 , n93941 , 
 n93942 , n93943 , n93944 , n93945 , n93946 , n93947 , n93948 , n93949 , n93950 , n93951 , 
 n93952 , n93953 , n93954 , n93955 , n93956 , n93957 , n93958 , n93959 , n93960 , n93961 , 
 n93962 , n93963 , n93964 , n93965 , n93966 , n93967 , n93968 , n93969 , n93970 , n93971 , 
 n93972 , n93973 , n93974 , n93975 , n93976 , n93977 , n93978 , n93979 , n93980 , n93981 , 
 n93982 , n93983 , n93984 , n93985 , n93986 , n93987 , n93988 , n93989 , n93990 , n93991 , 
 n93992 , n93993 , n93994 , n93995 , n93996 , n93997 , n93998 , n93999 , n94000 , n94001 , 
 n94002 , n94003 , n94004 , n94005 , n94006 , n94007 , n94008 , n94009 , n94010 , n94011 , 
 n94012 , n94013 , n94014 , n94015 , n94016 , n94017 , n94018 , n94019 , n94020 , n94021 , 
 n94022 , n94023 , n94024 , n94025 , n94026 , n94027 , n94028 , n94029 , n94030 , n94031 , 
 n94032 , n94033 , n94034 , n94035 , n94036 , n94037 , n94038 , n94039 , n94040 , n94041 , 
 n94042 , n94043 , n94044 , n94045 , n94046 , n94047 , n94048 , n94049 , n94050 , n94051 , 
 n94052 , n94053 , n94054 , n94055 , n94056 , n94057 , n94058 , n94059 , n94060 , n94061 , 
 n94062 , n94063 , n94064 , n94065 , n94066 , n94067 , n94068 , n94069 , n94070 , n94071 , 
 n94072 , n94073 , n94074 , n94075 , n94076 , n94077 , n94078 , n94079 , n94080 , n94081 , 
 n94082 , n94083 , n94084 , n94085 , n94086 , n94087 , n94088 , n94089 , n94090 , n94091 , 
 n94092 , n94093 , n94094 , n94095 , n94096 , n94097 , n94098 , n94099 , n94100 , n94101 , 
 n94102 , n94103 , n94104 , n94105 , n94106 , n94107 , n94108 , n94109 , n94110 , n94111 , 
 n94112 , n94113 , n94114 , n94115 , n94116 , n94117 , n94118 , n94119 , n94120 , n94121 , 
 n94122 , n94123 , n94124 , n94125 , n94126 , n94127 , n94128 , n94129 , n94130 , n94131 , 
 n94132 , n94133 , n94134 , n94135 , n94136 , n94137 , n94138 , n94139 , n94140 , n94141 , 
 n94142 , n94143 , n94144 , n94145 , n94146 , n94147 , n94148 , n94149 , n94150 , n94151 , 
 n94152 , n94153 , n94154 , n94155 , n94156 , n94157 , n94158 , n94159 , n94160 , n94161 , 
 n94162 , n94163 , n94164 , n94165 , n94166 , n94167 , n94168 , n94169 , n94170 , n94171 , 
 n94172 , n94173 , n94174 , n94175 , n94176 , n94177 , n94178 , n94179 , n94180 , n94181 , 
 n94182 , n94183 , n94184 , n94185 , n94186 , n94187 , n94188 , n94189 , n94190 , n94191 , 
 n94192 , n94193 , n94194 , n94195 , n94196 , n94197 , n94198 , n94199 , n94200 , n94201 , 
 n94202 , n94203 , n94204 , n94205 , n94206 , n94207 , n94208 , n94209 , n94210 , n94211 , 
 n94212 , n94213 , n94214 , n94215 , n94216 , n94217 , n94218 , n94219 , n94220 , n94221 , 
 n94222 , n94223 , n94224 , n94225 , n94226 , n94227 , n94228 , n94229 , n94230 , n94231 , 
 n94232 , n94233 , n94234 , n94235 , n94236 , n94237 , n94238 , n94239 , n94240 , n94241 , 
 n94242 , n94243 , n94244 , n94245 , n94246 , n94247 , n94248 , n94249 , n94250 , n94251 , 
 n94252 , n94253 , n94254 , n94255 , n94256 , n94257 , n94258 , n94259 , n94260 , n94261 , 
 n94262 , n94263 , n94264 , n94265 , n94266 , n94267 , n94268 , n94269 , n94270 , n94271 , 
 n94272 , n94273 , n94274 , n94275 , n94276 , n94277 , n94278 , n94279 , n94280 , n94281 , 
 n94282 , n94283 , n94284 , n94285 , n94286 , n94287 , n94288 , n94289 , n94290 , n94291 , 
 n94292 , n94293 , n94294 , n94295 , n94296 , n94297 , n94298 , n94299 , n94300 , n94301 , 
 n94302 , n94303 , n94304 , n94305 , n94306 , n94307 , n94308 , n94309 , n94310 , n94311 , 
 n94312 , n94313 , n94314 , n94315 , n94316 , n94317 , n94318 , n94319 , n94320 , n94321 , 
 n94322 , n94323 , n94324 , n94325 , n94326 , n94327 , n94328 , n94329 , n94330 , n94331 , 
 n94332 , n94333 , n94334 , n94335 , n94336 , n94337 , n94338 , n94339 , n94340 , n94341 , 
 n94342 , n94343 , n94344 , n94345 , n94346 , n94347 , n94348 , n94349 , n94350 , n94351 , 
 n94352 , n94353 , n94354 , n94355 , n94356 , n94357 , n94358 , n94359 , n94360 , n94361 , 
 n94362 , n94363 , n94364 , n94365 , n94366 , n94367 , n94368 , n94369 , n94370 , n94371 , 
 n94372 , n94373 , n94374 , n94375 , n94376 , n94377 , n94378 , n94379 , n94380 , n94381 , 
 n94382 , n94383 , n94384 , n94385 , n94386 , n94387 , n94388 , n94389 , n94390 , n94391 , 
 n94392 , n94393 , n94394 , n94395 , n94396 , n94397 , n94398 , n94399 , n94400 , n94401 , 
 n94402 , n94403 , n94404 , n94405 , n94406 , n94407 , n94408 , n94409 , n94410 , n94411 , 
 n94412 , n94413 , n94414 , n94415 , n94416 , n94417 , n94418 , n94419 , n94420 , n94421 , 
 n94422 , n94423 , n94424 , n94425 , n94426 , n94427 , n94428 , n94429 , n94430 , n94431 , 
 n94432 , n94433 , n94434 , n94435 , n94436 , n94437 , n94438 , n94439 , n94440 , n94441 , 
 n94442 , n94443 , n94444 , n94445 , n94446 , n94447 , n94448 , n94449 , n94450 , n94451 , 
 n94452 , n94453 , n94454 , n94455 , n94456 , n94457 , n94458 , n94459 , n94460 , n94461 , 
 n94462 , n94463 , n94464 , n94465 , n94466 , n94467 , n94468 , n94469 , n94470 , n94471 , 
 n94472 , n94473 , n94474 , n94475 , n94476 , n94477 , n94478 , n94479 , n94480 , n94481 , 
 n94482 , n94483 , n94484 , n94485 , n94486 , n94487 , n94488 , n94489 , n94490 , n94491 , 
 n94492 , n94493 , n94494 , n94495 , n94496 , n94497 , n94498 , n94499 , n94500 , n94501 , 
 n94502 , n94503 , n94504 , n94505 , n94506 , n94507 , n94508 , n94509 , n94510 , n94511 , 
 n94512 , n94513 , n94514 , n94515 , n94516 , n94517 , n94518 , n94519 , n94520 , n94521 , 
 n94522 , n94523 , n94524 , n94525 , n94526 , n94527 , n94528 , n94529 , n94530 , n94531 , 
 n94532 , n94533 , n94534 , n94535 , n94536 , n94537 , n94538 , n94539 , n94540 , n94541 , 
 n94542 , n94543 , n94544 , n94545 , n94546 , n94547 , n94548 , n94549 , n94550 , n94551 , 
 n94552 , n94553 , n94554 , n94555 , n94556 , n94557 , n94558 , n94559 , n94560 , n94561 , 
 n94562 , n94563 , n94564 , n94565 , n94566 , n94567 , n94568 , n94569 , n94570 , n94571 , 
 n94572 , n94573 , n94574 , n94575 , n94576 , n94577 , n94578 , n94579 , n94580 , n94581 , 
 n94582 , n94583 , n94584 , n94585 , n94586 , n94587 , n94588 , n94589 , n94590 , n94591 , 
 n94592 , n94593 , n94594 , n94595 , n94596 , n94597 , n94598 , n94599 , n94600 , n94601 , 
 n94602 , n94603 , n94604 , n94605 , n94606 , n94607 , n94608 , n94609 , n94610 , n94611 , 
 n94612 , n94613 , n94614 , n94615 , n94616 , n94617 , n94618 , n94619 , n94620 , n94621 , 
 n94622 , n94623 , n94624 , n94625 , n94626 , n94627 , n94628 , n94629 , n94630 , n94631 , 
 n94632 , n94633 , n94634 , n94635 , n94636 , n94637 , n94638 , n94639 , n94640 , n94641 , 
 n94642 , n94643 , n94644 , n94645 , n94646 , n94647 , n94648 , n94649 , n94650 , n94651 , 
 n94652 , n94653 , n94654 , n94655 , n94656 , n94657 , n94658 , n94659 , n94660 , n94661 , 
 n94662 , n94663 , n94664 , n94665 , n94666 , n94667 , n94668 , n94669 , n94670 , n94671 , 
 n94672 , n94673 , n94674 , n94675 , n94676 , n94677 , n94678 , n94679 , n94680 , n94681 , 
 n94682 , n94683 , n94684 , n94685 , n94686 , n94687 , n94688 , n94689 , n94690 , n94691 , 
 n94692 , n94693 , n94694 , n94695 , n94696 , n94697 , n94698 , n94699 , n94700 , n94701 , 
 n94702 , n94703 , n94704 , n94705 , n94706 , n94707 , n94708 , n94709 , n94710 , n94711 , 
 n94712 , n94713 , n94714 , n94715 , n94716 , n94717 , n94718 , n94719 , n94720 , n94721 , 
 n94722 , n94723 , n94724 , n94725 , n94726 , n94727 , n94728 , n94729 , n94730 , n94731 , 
 n94732 , n94733 , n94734 , n94735 , n94736 , n94737 , n94738 , n94739 , n94740 , n94741 , 
 n94742 , n94743 , n94744 , n94745 , n94746 , n94747 , n94748 , n94749 , n94750 , n94751 , 
 n94752 , n94753 , n94754 , n94755 , n94756 , n94757 , n94758 , n94759 , n94760 , n94761 , 
 n94762 , n94763 , n94764 , n94765 , n94766 , n94767 , n94768 , n94769 , n94770 , n94771 , 
 n94772 , n94773 , n94774 , n94775 , n94776 , n94777 , n94778 , n94779 , n94780 , n94781 , 
 n94782 , n94783 , n94784 , n94785 , n94786 , n94787 , n94788 , n94789 , n94790 , n94791 , 
 n94792 , n94793 , n94794 , n94795 , n94796 , n94797 , n94798 , n94799 , n94800 , n94801 , 
 n94802 , n94803 , n94804 , n94805 , n94806 , n94807 , n94808 , n94809 , n94810 , n94811 , 
 n94812 , n94813 , n94814 , n94815 , n94816 , n94817 , n94818 , n94819 , n94820 , n94821 , 
 n94822 , n94823 , n94824 , n94825 , n94826 , n94827 , n94828 , n94829 , n94830 , n94831 , 
 n94832 , n94833 , n94834 , n94835 , n94836 , n94837 , n94838 , n94839 , n94840 , n94841 , 
 n94842 , n94843 , n94844 , n94845 , n94846 , n94847 , n94848 , n94849 , n94850 , n94851 , 
 n94852 , n94853 , n94854 , n94855 , n94856 , n94857 , n94858 , n94859 , n94860 , n94861 , 
 n94862 , n94863 , n94864 , n94865 , n94866 , n94867 , n94868 , n94869 , n94870 , n94871 , 
 n94872 , n94873 , n94874 , n94875 , n94876 , n94877 , n94878 , n94879 , n94880 , n94881 , 
 n94882 , n94883 , n94884 , n94885 , n94886 , n94887 , n94888 , n94889 , n94890 , n94891 , 
 n94892 , n94893 , n94894 , n94895 , n94896 , n94897 , n94898 , n94899 , n94900 , n94901 , 
 n94902 , n94903 , n94904 , n94905 , n94906 , n94907 , n94908 , n94909 , n94910 , n94911 , 
 n94912 , n94913 , n94914 , n94915 , n94916 , n94917 , n94918 , n94919 , n94920 , n94921 , 
 n94922 , n94923 , n94924 , n94925 , n94926 , n94927 , n94928 , n94929 , n94930 , n94931 , 
 n94932 , n94933 , n94934 , n94935 , n94936 , n94937 , n94938 , n94939 , n94940 , n94941 , 
 n94942 , n94943 , n94944 , n94945 , n94946 , n94947 , n94948 , n94949 , n94950 , n94951 , 
 n94952 , n94953 , n94954 , n94955 , n94956 , n94957 , n94958 , n94959 , n94960 , n94961 , 
 n94962 , n94963 , n94964 , n94965 , n94966 , n94967 , n94968 , n94969 , n94970 , n94971 , 
 n94972 , n94973 , n94974 , n94975 , n94976 , n94977 , n94978 , n94979 , n94980 , n94981 , 
 n94982 , n94983 , n94984 , n94985 , n94986 , n94987 , n94988 , n94989 , n94990 , n94991 , 
 n94992 , n94993 , n94994 , n94995 , n94996 , n94997 , n94998 , n94999 , n95000 , n95001 , 
 n95002 , n95003 , n95004 , n95005 , n95006 , n95007 , n95008 , n95009 , n95010 , n95011 , 
 n95012 , n95013 , n95014 , n95015 , n95016 , n95017 , n95018 , n95019 , n95020 , n95021 , 
 n95022 , n95023 , n95024 , n95025 , n95026 , n95027 , n95028 , n95029 , n95030 , n95031 , 
 n95032 , n95033 , n95034 , n95035 , n95036 , n95037 , n95038 , n95039 , n95040 , n95041 , 
 n95042 , n95043 , n95044 , n95045 , n95046 , n95047 , n95048 , n95049 , n95050 , n95051 , 
 n95052 , n95053 , n95054 , n95055 , n95056 , n95057 , n95058 , n95059 , n95060 , n95061 , 
 n95062 , n95063 , n95064 , n95065 , n95066 , n95067 , n95068 , n95069 , n95070 , n95071 , 
 n95072 , n95073 , n95074 , n95075 , n95076 , n95077 , n95078 , n95079 , n95080 , n95081 , 
 n95082 , n95083 , n95084 , n95085 , n95086 , n95087 , n95088 , n95089 , n95090 , n95091 , 
 n95092 , n95093 , n95094 , n95095 , n95096 , n95097 , n95098 , n95099 , n95100 , n95101 , 
 n95102 , n95103 , n95104 , n95105 , n95106 , n95107 , n95108 , n95109 , n95110 , n95111 , 
 n95112 , n95113 , n95114 , n95115 , n95116 , n95117 , n95118 , n95119 , n95120 , n95121 , 
 n95122 , n95123 , n95124 , n95125 , n95126 , n95127 , n95128 , n95129 , n95130 , n95131 , 
 n95132 , n95133 , n95134 , n95135 , n95136 , n95137 , n95138 , n95139 , n95140 , n95141 , 
 n95142 , n95143 , n95144 , n95145 , n95146 , n95147 , n95148 , n95149 , n95150 , n95151 , 
 n95152 , n95153 , n95154 , n95155 , n95156 , n95157 , n95158 , n95159 , n95160 , n95161 , 
 n95162 , n95163 , n95164 , n95165 , n95166 , n95167 , n95168 , n95169 , n95170 , n95171 , 
 n95172 , n95173 , n95174 , n95175 , n95176 , n95177 , n95178 , n95179 , n95180 , n95181 , 
 n95182 , n95183 , n95184 , n95185 , n95186 , n95187 , n95188 , n95189 , n95190 , n95191 , 
 n95192 , n95193 , n95194 , n95195 , n95196 , n95197 , n95198 , n95199 , n95200 , n95201 , 
 n95202 , n95203 , n95204 , n95205 , n95206 , n95207 , n95208 , n95209 , n95210 , n95211 , 
 n95212 , n95213 , n95214 , n95215 , n95216 , n95217 , n95218 , n95219 , n95220 , n95221 , 
 n95222 , n95223 , n95224 , n95225 , n95226 , n95227 , n95228 , n95229 , n95230 , n95231 , 
 n95232 , n95233 , n95234 , n95235 , n95236 , n95237 , n95238 , n95239 , n95240 , n95241 , 
 n95242 , n95243 , n95244 , n95245 , n95246 , n95247 , n95248 , n95249 , n95250 , n95251 , 
 n95252 , n95253 , n95254 , n95255 , n95256 , n95257 , n95258 , n95259 , n95260 , n95261 , 
 n95262 , n95263 , n95264 , n95265 , n95266 , n95267 , n95268 , n95269 , n95270 , n95271 , 
 n95272 , n95273 , n95274 , n95275 , n95276 , n95277 , n95278 , n95279 , n95280 , n95281 , 
 n95282 , n95283 , n95284 , n95285 , n95286 , n95287 , n95288 , n95289 , n95290 , n95291 , 
 n95292 , n95293 , n95294 , n95295 , n95296 , n95297 , n95298 , n95299 , n95300 , n95301 , 
 n95302 , n95303 , n95304 , n95305 , n95306 , n95307 , n95308 , n95309 , n95310 , n95311 , 
 n95312 , n95313 , n95314 , n95315 , n95316 , n95317 , n95318 , n95319 , n95320 , n95321 , 
 n95322 , n95323 , n95324 , n95325 , n95326 , n95327 , n95328 , n95329 , n95330 , n95331 , 
 n95332 , n95333 , n95334 , n95335 , n95336 , n95337 , n95338 , n95339 , n95340 , n95341 , 
 n95342 , n95343 , n95344 , n95345 , n95346 , n95347 , n95348 , n95349 , n95350 , n95351 , 
 n95352 , n95353 , n95354 , n95355 , n95356 , n95357 , n95358 , n95359 , n95360 , n95361 , 
 n95362 , n95363 , n95364 , n95365 , n95366 , n95367 , n95368 , n95369 , n95370 , n95371 , 
 n95372 , n95373 , n95374 , n95375 , n95376 , n95377 , n95378 , n95379 , n95380 , n95381 , 
 n95382 , n95383 , n95384 , n95385 , n95386 , n95387 , n95388 , n95389 , n95390 , n95391 , 
 n95392 , n95393 , n95394 , n95395 , n95396 , n95397 , n95398 , n95399 , n95400 , n95401 , 
 n95402 , n95403 , n95404 , n95405 , n95406 , n95407 , n95408 , n95409 , n95410 , n95411 , 
 n95412 , n95413 , n95414 , n95415 , n95416 , n95417 , n95418 , n95419 , n95420 , n95421 , 
 n95422 , n95423 , n95424 , n95425 , n95426 , n95427 , n95428 , n95429 , n95430 , n95431 , 
 n95432 , n95433 , n95434 , n95435 , n95436 , n95437 , n95438 , n95439 , n95440 , n95441 , 
 n95442 , n95443 , n95444 , n95445 , n95446 , n95447 , n95448 , n95449 , n95450 , n95451 , 
 n95452 , n95453 , n95454 , n95455 , n95456 , n95457 , n95458 , n95459 , n95460 , n95461 , 
 n95462 , n95463 , n95464 , n95465 , n95466 , n95467 , n95468 , n95469 , n95470 , n95471 , 
 n95472 , n95473 , n95474 , n95475 , n95476 , n95477 , n95478 , n95479 , n95480 , n95481 , 
 n95482 , n95483 , n95484 , n95485 , n95486 , n95487 , n95488 , n95489 , n95490 , n95491 , 
 n95492 , n95493 , n95494 , n95495 , n95496 , n95497 , n95498 , n95499 , n95500 , n95501 , 
 n95502 , n95503 , n95504 , n95505 , n95506 , n95507 , n95508 , n95509 , n95510 , n95511 , 
 n95512 , n95513 , n95514 , n95515 , n95516 , n95517 , n95518 , n95519 , n95520 , n95521 , 
 n95522 , n95523 , n95524 , n95525 , n95526 , n95527 , n95528 , n95529 , n95530 , n95531 , 
 n95532 , n95533 , n95534 , n95535 , n95536 , n95537 , n95538 , n95539 , n95540 , n95541 , 
 n95542 , n95543 , n95544 , n95545 , n95546 , n95547 , n95548 , n95549 , n95550 , n95551 , 
 n95552 , n95553 , n95554 , n95555 , n95556 , n95557 , n95558 , n95559 , n95560 , n95561 , 
 n95562 , n95563 , n95564 , n95565 , n95566 , n95567 , n95568 , n95569 , n95570 , n95571 , 
 n95572 , n95573 , n95574 , n95575 , n95576 , n95577 , n95578 , n95579 , n95580 , n95581 , 
 n95582 , n95583 , n95584 , n95585 , n95586 , n95587 , n95588 , n95589 , n95590 , n95591 , 
 n95592 , n95593 , n95594 , n95595 , n95596 , n95597 , n95598 , n95599 , n95600 , n95601 , 
 n95602 , n95603 , n95604 , n95605 , n95606 , n95607 , n95608 , n95609 , n95610 , n95611 , 
 n95612 , n95613 , n95614 , n95615 , n95616 , n95617 , n95618 , n95619 , n95620 , n95621 , 
 n95622 , n95623 , n95624 , n95625 , n95626 , n95627 , n95628 , n95629 , n95630 , n95631 , 
 n95632 , n95633 , n95634 , n95635 , n95636 , n95637 , n95638 , n95639 , n95640 , n95641 , 
 n95642 , n95643 , n95644 , n95645 , n95646 , n95647 , n95648 , n95649 , n95650 , n95651 , 
 n95652 , n95653 , n95654 , n95655 , n95656 , n95657 , n95658 , n95659 , n95660 , n95661 , 
 n95662 , n95663 , n95664 , n95665 , n95666 , n95667 , n95668 , n95669 , n95670 , n95671 , 
 n95672 , n95673 , n95674 , n95675 , n95676 , n95677 , n95678 , n95679 , n95680 , n95681 , 
 n95682 , n95683 , n95684 , n95685 , n95686 , n95687 , n95688 , n95689 , n95690 , n95691 , 
 n95692 , n95693 , n95694 , n95695 , n95696 , n95697 , n95698 , n95699 , n95700 , n95701 , 
 n95702 , n95703 , n95704 , n95705 , n95706 , n95707 , n95708 , n95709 , n95710 , n95711 , 
 n95712 , n95713 , n95714 , n95715 , n95716 , n95717 , n95718 , n95719 , n95720 , n95721 , 
 n95722 , n95723 , n95724 , n95725 , n95726 , n95727 , n95728 , n95729 , n95730 , n95731 , 
 n95732 , n95733 , n95734 , n95735 , n95736 , n95737 , n95738 , n95739 , n95740 , n95741 , 
 n95742 , n95743 , n95744 , n95745 , n95746 , n95747 , n95748 , n95749 , n95750 , n95751 , 
 n95752 , n95753 , n95754 , n95755 , n95756 , n95757 , n95758 , n95759 , n95760 , n95761 , 
 n95762 , n95763 , n95764 , n95765 , n95766 , n95767 , n95768 , n95769 , n95770 , n95771 , 
 n95772 , n95773 , n95774 , n95775 , n95776 , n95777 , n95778 , n95779 , n95780 , n95781 , 
 n95782 , n95783 , n95784 , n95785 , n95786 , n95787 , n95788 , n95789 , n95790 , n95791 , 
 n95792 , n95793 , n95794 , n95795 , n95796 , n95797 , n95798 , n95799 , n95800 , n95801 , 
 n95802 , n95803 , n95804 , n95805 , n95806 , n95807 , n95808 , n95809 , n95810 , n95811 , 
 n95812 , n95813 , n95814 , n95815 , n95816 , n95817 , n95818 , n95819 , n95820 , n95821 , 
 n95822 , n95823 , n95824 , n95825 , n95826 , n95827 , n95828 , n95829 , n95830 , n95831 , 
 n95832 , n95833 , n95834 , n95835 , n95836 , n95837 , n95838 , n95839 , n95840 , n95841 , 
 n95842 , n95843 , n95844 , n95845 , n95846 , n95847 , n95848 , n95849 , n95850 , n95851 , 
 n95852 , n95853 , n95854 , n95855 , n95856 , n95857 , n95858 , n95859 , n95860 , n95861 , 
 n95862 , n95863 , n95864 , n95865 , n95866 , n95867 , n95868 , n95869 , n95870 , n95871 , 
 n95872 , n95873 , n95874 , n95875 , n95876 , n95877 , n95878 , n95879 , n95880 , n95881 , 
 n95882 , n95883 , n95884 , n95885 , n95886 , n95887 , n95888 , n95889 , n95890 , n95891 , 
 n95892 , n95893 , n95894 , n95895 , n95896 , n95897 , n95898 , n95899 , n95900 , n95901 , 
 n95902 , n95903 , n95904 , n95905 , n95906 , n95907 , n95908 , n95909 , n95910 , n95911 , 
 n95912 , n95913 , n95914 , n95915 , n95916 , n95917 , n95918 , n95919 , n95920 , n95921 , 
 n95922 , n95923 , n95924 , n95925 , n95926 , n95927 , n95928 , n95929 , n95930 , n95931 , 
 n95932 , n95933 , n95934 , n95935 , n95936 , n95937 , n95938 , n95939 , n95940 , n95941 , 
 n95942 , n95943 , n95944 , n95945 , n95946 , n95947 , n95948 , n95949 , n95950 , n95951 , 
 n95952 , n95953 , n95954 , n95955 , n95956 , n95957 , n95958 , n95959 , n95960 , n95961 , 
 n95962 , n95963 , n95964 , n95965 , n95966 , n95967 , n95968 , n95969 , n95970 , n95971 , 
 n95972 , n95973 , n95974 , n95975 , n95976 , n95977 , n95978 , n95979 , n95980 , n95981 , 
 n95982 , n95983 , n95984 , n95985 , n95986 , n95987 , n95988 , n95989 , n95990 , n95991 , 
 n95992 , n95993 , n95994 , n95995 , n95996 , n95997 , n95998 , n95999 , n96000 , n96001 , 
 n96002 , n96003 , n96004 , n96005 , n96006 , n96007 , n96008 , n96009 , n96010 , n96011 , 
 n96012 , n96013 , n96014 , n96015 , n96016 , n96017 , n96018 , n96019 , n96020 , n96021 , 
 n96022 , n96023 , n96024 , n96025 , n96026 , n96027 , n96028 , n96029 , n96030 , n96031 , 
 n96032 , n96033 , n96034 , n96035 , n96036 , n96037 , n96038 , n96039 , n96040 , n96041 , 
 n96042 , n96043 , n96044 , n96045 , n96046 , n96047 , n96048 , n96049 , n96050 , n96051 , 
 n96052 , n96053 , n96054 , n96055 , n96056 , n96057 , n96058 , n96059 , n96060 , n96061 , 
 n96062 , n96063 , n96064 , n96065 , n96066 , n96067 , n96068 , n96069 , n96070 , n96071 , 
 n96072 , n96073 , n96074 , n96075 , n96076 , n96077 , n96078 , n96079 , n96080 , n96081 , 
 n96082 , n96083 , n96084 , n96085 , n96086 , n96087 , n96088 , n96089 , n96090 , n96091 , 
 n96092 , n96093 , n96094 , n96095 , n96096 , n96097 , n96098 , n96099 , n96100 , n96101 , 
 n96102 , n96103 , n96104 , n96105 , n96106 , n96107 , n96108 , n96109 , n96110 , n96111 , 
 n96112 , n96113 , n96114 , n96115 , n96116 , n96117 , n96118 , n96119 , n96120 , n96121 , 
 n96122 , n96123 , n96124 , n96125 , n96126 , n96127 , n96128 , n96129 , n96130 , n96131 , 
 n96132 , n96133 , n96134 , n96135 , n96136 , n96137 , n96138 , n96139 , n96140 , n96141 , 
 n96142 , n96143 , n96144 , n96145 , n96146 , n96147 , n96148 , n96149 , n96150 , n96151 , 
 n96152 , n96153 , n96154 , n96155 , n96156 , n96157 , n96158 , n96159 , n96160 , n96161 , 
 n96162 , n96163 , n96164 , n96165 , n96166 , n96167 , n96168 , n96169 , n96170 , n96171 , 
 n96172 , n96173 , n96174 , n96175 , n96176 , n96177 , n96178 , n96179 , n96180 , n96181 , 
 n96182 , n96183 , n96184 , n96185 , n96186 , n96187 , n96188 , n96189 , n96190 , n96191 , 
 n96192 , n96193 , n96194 , n96195 , n96196 , n96197 , n96198 , n96199 , n96200 , n96201 , 
 n96202 , n96203 , n96204 , n96205 , n96206 , n96207 , n96208 , n96209 , n96210 , n96211 , 
 n96212 , n96213 , n96214 , n96215 , n96216 , n96217 , n96218 , n96219 , n96220 , n96221 , 
 n96222 , n96223 , n96224 , n96225 , n96226 , n96227 , n96228 , n96229 , n96230 , n96231 , 
 n96232 , n96233 , n96234 , n96235 , n96236 , n96237 , n96238 , n96239 , n96240 , n96241 , 
 n96242 , n96243 , n96244 , n96245 , n96246 , n96247 , n96248 , n96249 , n96250 , n96251 , 
 n96252 , n96253 , n96254 , n96255 , n96256 , n96257 , n96258 , n96259 , n96260 , n96261 , 
 n96262 , n96263 , n96264 , n96265 , n96266 , n96267 , n96268 , n96269 , n96270 , n96271 , 
 n96272 , n96273 , n96274 , n96275 , n96276 , n96277 , n96278 , n96279 , n96280 , n96281 , 
 n96282 , n96283 , n96284 , n96285 , n96286 , n96287 , n96288 , n96289 , n96290 , n96291 , 
 n96292 , n96293 , n96294 , n96295 , n96296 , n96297 , n96298 , n96299 , n96300 , n96301 , 
 n96302 , n96303 , n96304 , n96305 , n96306 , n96307 , n96308 , n96309 , n96310 , n96311 , 
 n96312 , n96313 , n96314 , n96315 , n96316 , n96317 , n96318 , n96319 , n96320 , n96321 , 
 n96322 , n96323 , n96324 , n96325 , n96326 , n96327 , n96328 , n96329 , n96330 , n96331 , 
 n96332 , n96333 , n96334 , n96335 , n96336 , n96337 , n96338 , n96339 , n96340 , n96341 , 
 n96342 , n96343 , n96344 , n96345 , n96346 , n96347 , n96348 , n96349 , n96350 , n96351 , 
 n96352 , n96353 , n96354 , n96355 , n96356 , n96357 , n96358 , n96359 , n96360 , n96361 , 
 n96362 , n96363 , n96364 , n96365 , n96366 , n96367 , n96368 , n96369 , n96370 , n96371 , 
 n96372 , n96373 , n96374 , n96375 , n96376 , n96377 , n96378 , n96379 , n96380 , n96381 , 
 n96382 , n96383 , n96384 , n96385 , n96386 , n96387 , n96388 , n96389 , n96390 , n96391 , 
 n96392 , n96393 , n96394 , n96395 , n96396 , n96397 , n96398 , n96399 , n96400 , n96401 , 
 n96402 , n96403 , n96404 , n96405 , n96406 , n96407 , n96408 , n96409 , n96410 , n96411 , 
 n96412 , n96413 , n96414 , n96415 , n96416 , n96417 , n96418 , n96419 , n96420 , n96421 , 
 n96422 , n96423 , n96424 , n96425 , n96426 , n96427 , n96428 , n96429 , n96430 , n96431 , 
 n96432 , n96433 , n96434 , n96435 , n96436 , n96437 , n96438 , n96439 , n96440 , n96441 , 
 n96442 , n96443 , n96444 , n96445 , n96446 , n96447 , n96448 , n96449 , n96450 , n96451 , 
 n96452 , n96453 , n96454 , n96455 , n96456 , n96457 , n96458 , n96459 , n96460 , n96461 , 
 n96462 , n96463 , n96464 , n96465 , n96466 , n96467 , n96468 , n96469 , n96470 , n96471 , 
 n96472 , n96473 , n96474 , n96475 , n96476 , n96477 , n96478 , n96479 , n96480 , n96481 , 
 n96482 , n96483 , n96484 , n96485 , n96486 , n96487 , n96488 , n96489 , n96490 , n96491 , 
 n96492 , n96493 , n96494 , n96495 , n96496 , n96497 , n96498 , n96499 , n96500 , n96501 , 
 n96502 , n96503 , n96504 , n96505 , n96506 , n96507 , n96508 , n96509 , n96510 , n96511 , 
 n96512 , n96513 , n96514 , n96515 , n96516 , n96517 , n96518 , n96519 , n96520 , n96521 , 
 n96522 , n96523 , n96524 , n96525 , n96526 , n96527 , n96528 , n96529 , n96530 , n96531 , 
 n96532 , n96533 , n96534 , n96535 , n96536 , n96537 , n96538 , n96539 , n96540 , n96541 , 
 n96542 , n96543 , n96544 , n96545 , n96546 , n96547 , n96548 , n96549 , n96550 , n96551 , 
 n96552 , n96553 , n96554 , n96555 , n96556 , n96557 , n96558 , n96559 , n96560 , n96561 , 
 n96562 , n96563 , n96564 , n96565 , n96566 , n96567 , n96568 , n96569 , n96570 , n96571 , 
 n96572 , n96573 , n96574 , n96575 , n96576 , n96577 , n96578 , n96579 , n96580 , n96581 , 
 n96582 , n96583 , n96584 , n96585 , n96586 , n96587 , n96588 , n96589 , n96590 , n96591 , 
 n96592 , n96593 , n96594 , n96595 , n96596 , n96597 , n96598 , n96599 , n96600 , n96601 , 
 n96602 , n96603 , n96604 , n96605 , n96606 , n96607 , n96608 , n96609 , n96610 , n96611 , 
 n96612 , n96613 , n96614 , n96615 , n96616 , n96617 , n96618 , n96619 , n96620 , n96621 , 
 n96622 , n96623 , n96624 , n96625 , n96626 , n96627 , n96628 , n96629 , n96630 , n96631 , 
 n96632 , n96633 , n96634 , n96635 , n96636 , n96637 , n96638 , n96639 , n96640 , n96641 , 
 n96642 , n96643 , n96644 , n96645 , n96646 , n96647 , n96648 , n96649 , n96650 , n96651 , 
 n96652 , n96653 , n96654 , n96655 , n96656 , n96657 , n96658 , n96659 , n96660 , n96661 , 
 n96662 , n96663 , n96664 , n96665 , n96666 , n96667 , n96668 , n96669 , n96670 , n96671 , 
 n96672 , n96673 , n96674 , n96675 , n96676 , n96677 , n96678 , n96679 , n96680 , n96681 , 
 n96682 , n96683 , n96684 , n96685 , n96686 , n96687 , n96688 , n96689 , n96690 , n96691 , 
 n96692 , n96693 , n96694 , n96695 , n96696 , n96697 , n96698 , n96699 , n96700 , n96701 , 
 n96702 , n96703 , n96704 , n96705 , n96706 , n96707 , n96708 , n96709 , n96710 , n96711 , 
 n96712 , n96713 , n96714 , n96715 , n96716 , n96717 , n96718 , n96719 , n96720 , n96721 , 
 n96722 , n96723 , n96724 , n96725 , n96726 , n96727 , n96728 , n96729 , n96730 , n96731 , 
 n96732 , n96733 , n96734 , n96735 , n96736 , n96737 , n96738 , n96739 , n96740 , n96741 , 
 n96742 , n96743 , n96744 , n96745 , n96746 , n96747 , n96748 , n96749 , n96750 , n96751 , 
 n96752 , n96753 , n96754 , n96755 , n96756 , n96757 , n96758 , n96759 , n96760 , n96761 , 
 n96762 , n96763 , n96764 , n96765 , n96766 , n96767 , n96768 , n96769 , n96770 , n96771 , 
 n96772 , n96773 , n96774 , n96775 , n96776 , n96777 , n96778 , n96779 , n96780 , n96781 , 
 n96782 , n96783 , n96784 , n96785 , n96786 , n96787 , n96788 , n96789 , n96790 , n96791 , 
 n96792 , n96793 , n96794 , n96795 , n96796 , n96797 , n96798 , n96799 , n96800 , n96801 , 
 n96802 , n96803 , n96804 , n96805 , n96806 , n96807 , n96808 , n96809 , n96810 , n96811 , 
 n96812 , n96813 , n96814 , n96815 , n96816 , n96817 , n96818 , n96819 , n96820 , n96821 , 
 n96822 , n96823 , n96824 , n96825 , n96826 , n96827 , n96828 , n96829 , n96830 , n96831 , 
 n96832 , n96833 , n96834 , n96835 , n96836 , n96837 , n96838 , n96839 , n96840 , n96841 , 
 n96842 , n96843 , n96844 , n96845 , n96846 , n96847 , n96848 , n96849 , n96850 , n96851 , 
 n96852 , n96853 , n96854 , n96855 , n96856 , n96857 , n96858 , n96859 , n96860 , n96861 , 
 n96862 , n96863 , n96864 , n96865 , n96866 , n96867 , n96868 , n96869 , n96870 , n96871 , 
 n96872 , n96873 , n96874 , n96875 , n96876 , n96877 , n96878 , n96879 , n96880 , n96881 , 
 n96882 , n96883 , n96884 , n96885 , n96886 , n96887 , n96888 , n96889 , n96890 , n96891 , 
 n96892 , n96893 , n96894 , n96895 , n96896 , n96897 , n96898 , n96899 , n96900 , n96901 , 
 n96902 , n96903 , n96904 , n96905 , n96906 , n96907 , n96908 , n96909 , n96910 , n96911 , 
 n96912 , n96913 , n96914 , n96915 , n96916 , n96917 , n96918 , n96919 , n96920 , n96921 , 
 n96922 , n96923 , n96924 , n96925 , n96926 , n96927 , n96928 , n96929 , n96930 , n96931 , 
 n96932 , n96933 , n96934 , n96935 , n96936 , n96937 , n96938 , n96939 , n96940 , n96941 , 
 n96942 , n96943 , n96944 , n96945 , n96946 , n96947 , n96948 , n96949 , n96950 , n96951 , 
 n96952 , n96953 , n96954 , n96955 , n96956 , n96957 , n96958 , n96959 , n96960 , n96961 , 
 n96962 , n96963 , n96964 , n96965 , n96966 , n96967 , n96968 , n96969 , n96970 , n96971 , 
 n96972 , n96973 , n96974 , n96975 , n96976 , n96977 , n96978 , n96979 , n96980 , n96981 , 
 n96982 , n96983 , n96984 , n96985 , n96986 , n96987 , n96988 , n96989 , n96990 , n96991 , 
 n96992 , n96993 , n96994 , n96995 , n96996 , n96997 , n96998 , n96999 , n97000 , n97001 , 
 n97002 , n97003 , n97004 , n97005 , n97006 , n97007 , n97008 , n97009 , n97010 , n97011 , 
 n97012 , n97013 , n97014 , n97015 , n97016 , n97017 , n97018 , n97019 , n97020 , n97021 , 
 n97022 , n97023 , n97024 , n97025 , n97026 , n97027 , n97028 , n97029 , n97030 , n97031 , 
 n97032 , n97033 , n97034 , n97035 , n97036 , n97037 , n97038 , n97039 , n97040 , n97041 , 
 n97042 , n97043 , n97044 , n97045 , n97046 , n97047 , n97048 , n97049 , n97050 , n97051 , 
 n97052 , n97053 , n97054 , n97055 , n97056 , n97057 , n97058 , n97059 , n97060 , n97061 , 
 n97062 , n97063 , n97064 , n97065 , n97066 , n97067 , n97068 , n97069 , n97070 , n97071 , 
 n97072 , n97073 , n97074 , n97075 , n97076 , n97077 , n97078 , n97079 , n97080 , n97081 , 
 n97082 , n97083 , n97084 , n97085 , n97086 , n97087 , n97088 , n97089 , n97090 , n97091 , 
 n97092 , n97093 , n97094 , n97095 , n97096 , n97097 , n97098 , n97099 , n97100 , n97101 , 
 n97102 , n97103 , n97104 , n97105 , n97106 , n97107 , n97108 , n97109 , n97110 , n97111 , 
 n97112 , n97113 , n97114 , n97115 , n97116 , n97117 , n97118 , n97119 , n97120 , n97121 , 
 n97122 , n97123 , n97124 , n97125 , n97126 , n97127 , n97128 , n97129 , n97130 , n97131 , 
 n97132 , n97133 , n97134 , n97135 , n97136 , n97137 , n97138 , n97139 , n97140 , n97141 , 
 n97142 , n97143 , n97144 , n97145 , n97146 , n97147 , n97148 , n97149 , n97150 , n97151 , 
 n97152 , n97153 , n97154 , n97155 , n97156 , n97157 , n97158 , n97159 , n97160 , n97161 , 
 n97162 , n97163 , n97164 , n97165 , n97166 , n97167 , n97168 , n97169 , n97170 , n97171 , 
 n97172 , n97173 , n97174 , n97175 , n97176 , n97177 , n97178 , n97179 , n97180 , n97181 , 
 n97182 , n97183 , n97184 , n97185 , n97186 , n97187 , n97188 , n97189 , n97190 , n97191 , 
 n97192 , n97193 , n97194 , n97195 , n97196 , n97197 , n97198 , n97199 , n97200 , n97201 , 
 n97202 , n97203 , n97204 , n97205 , n97206 , n97207 , n97208 , n97209 , n97210 , n97211 , 
 n97212 , n97213 , n97214 , n97215 , n97216 , n97217 , n97218 , n97219 , n97220 , n97221 , 
 n97222 , n97223 , n97224 , n97225 , n97226 , n97227 , n97228 , n97229 , n97230 , n97231 , 
 n97232 , n97233 , n97234 , n97235 , n97236 , n97237 , n97238 , n97239 , n97240 , n97241 , 
 n97242 , n97243 , n97244 , n97245 , n97246 , n97247 , n97248 , n97249 , n97250 , n97251 , 
 n97252 , n97253 , n97254 , n97255 , n97256 , n97257 , n97258 , n97259 , n97260 , n97261 , 
 n97262 , n97263 , n97264 , n97265 , n97266 , n97267 , n97268 , n97269 , n97270 , n97271 , 
 n97272 , n97273 , n97274 , n97275 , n97276 , n97277 , n97278 , n97279 , n97280 , n97281 , 
 n97282 , n97283 , n97284 , n97285 , n97286 , n97287 , n97288 , n97289 , n97290 , n97291 , 
 n97292 , n97293 , n97294 , n97295 , n97296 , n97297 , n97298 , n97299 , n97300 , n97301 , 
 n97302 , n97303 , n97304 , n97305 , n97306 , n97307 , n97308 , n97309 , n97310 , n97311 , 
 n97312 , n97313 , n97314 , n97315 , n97316 , n97317 , n97318 , n97319 , n97320 , n97321 , 
 n97322 , n97323 , n97324 , n97325 , n97326 , n97327 , n97328 , n97329 , n97330 , n97331 , 
 n97332 , n97333 , n97334 , n97335 , n97336 , n97337 , n97338 , n97339 , n97340 , n97341 , 
 n97342 , n97343 , n97344 , n97345 , n97346 , n97347 , n97348 , n97349 , n97350 , n97351 , 
 n97352 , n97353 , n97354 , n97355 , n97356 , n97357 , n97358 , n97359 , n97360 , n97361 , 
 n97362 , n97363 , n97364 , n97365 , n97366 , n97367 , n97368 , n97369 , n97370 , n97371 , 
 n97372 , n97373 , n97374 , n97375 , n97376 , n97377 , n97378 , n97379 , n97380 , n97381 , 
 n97382 , n97383 , n97384 , n97385 , n97386 , n97387 , n97388 , n97389 , n97390 , n97391 , 
 n97392 , n97393 , n97394 , n97395 , n97396 , n97397 , n97398 , n97399 , n97400 , n97401 , 
 n97402 , n97403 , n97404 , n97405 , n97406 , n97407 , n97408 , n97409 , n97410 , n97411 , 
 n97412 , n97413 , n97414 , n97415 , n97416 , n97417 , n97418 , n97419 , n97420 , n97421 , 
 n97422 , n97423 , n97424 , n97425 , n97426 , n97427 , n97428 , n97429 , n97430 , n97431 , 
 n97432 , n97433 , n97434 , n97435 , n97436 , n97437 , n97438 , n97439 , n97440 , n97441 , 
 n97442 , n97443 , n97444 , n97445 , n97446 , n97447 , n97448 , n97449 , n97450 , n97451 , 
 n97452 , n97453 , n97454 , n97455 , n97456 , n97457 , n97458 , n97459 , n97460 , n97461 , 
 n97462 , n97463 , n97464 , n97465 , n97466 , n97467 , n97468 , n97469 , n97470 , n97471 , 
 n97472 , n97473 , n97474 , n97475 , n97476 , n97477 , n97478 , n97479 , n97480 , n97481 , 
 n97482 , n97483 , n97484 , n97485 , n97486 , n97487 , n97488 , n97489 , n97490 , n97491 , 
 n97492 , n97493 , n97494 , n97495 , n97496 , n97497 , n97498 , n97499 , n97500 , n97501 , 
 n97502 , n97503 , n97504 , n97505 , n97506 , n97507 , n97508 , n97509 , n97510 , n97511 , 
 n97512 , n97513 , n97514 , n97515 , n97516 , n97517 , n97518 , n97519 , n97520 , n97521 , 
 n97522 , n97523 , n97524 , n97525 , n97526 , n97527 , n97528 , n97529 , n97530 , n97531 , 
 n97532 , n97533 , n97534 , n97535 , n97536 , n97537 , n97538 , n97539 , n97540 , n97541 , 
 n97542 , n97543 , n97544 , n97545 , n97546 , n97547 , n97548 , n97549 , n97550 , n97551 , 
 n97552 , n97553 , n97554 , n97555 , n97556 , n97557 , n97558 , n97559 , n97560 , n97561 , 
 n97562 , n97563 , n97564 , n97565 , n97566 , n97567 , n97568 , n97569 , n97570 , n97571 , 
 n97572 , n97573 , n97574 , n97575 , n97576 , n97577 , n97578 , n97579 , n97580 , n97581 , 
 n97582 , n97583 , n97584 , n97585 , n97586 , n97587 , n97588 , n97589 , n97590 , n97591 , 
 n97592 , n97593 , n97594 , n97595 , n97596 , n97597 , n97598 , n97599 , n97600 , n97601 , 
 n97602 , n97603 , n97604 , n97605 , n97606 , n97607 , n97608 , n97609 , n97610 , n97611 , 
 n97612 , n97613 , n97614 , n97615 , n97616 , n97617 , n97618 , n97619 , n97620 , n97621 , 
 n97622 , n97623 , n97624 , n97625 , n97626 , n97627 , n97628 , n97629 , n97630 , n97631 , 
 n97632 , n97633 , n97634 , n97635 , n97636 , n97637 , n97638 , n97639 , n97640 , n97641 , 
 n97642 , n97643 , n97644 , n97645 , n97646 , n97647 , n97648 , n97649 , n97650 , n97651 , 
 n97652 , n97653 , n97654 , n97655 , n97656 , n97657 , n97658 , n97659 , n97660 , n97661 , 
 n97662 , n97663 , n97664 , n97665 , n97666 , n97667 , n97668 , n97669 , n97670 , n97671 , 
 n97672 , n97673 , n97674 , n97675 , n97676 , n97677 , n97678 , n97679 , n97680 , n97681 , 
 n97682 , n97683 , n97684 , n97685 , n97686 , n97687 , n97688 , n97689 , n97690 , n97691 , 
 n97692 , n97693 , n97694 , n97695 , n97696 , n97697 , n97698 , n97699 , n97700 , n97701 , 
 n97702 , n97703 , n97704 , n97705 , n97706 , n97707 , n97708 , n97709 , n97710 , n97711 , 
 n97712 , n97713 , n97714 , n97715 , n97716 , n97717 , n97718 , n97719 , n97720 , n97721 , 
 n97722 , n97723 , n97724 , n97725 , n97726 , n97727 , n97728 , n97729 , n97730 , n97731 , 
 n97732 , n97733 , n97734 , n97735 , n97736 , n97737 , n97738 , n97739 , n97740 , n97741 , 
 n97742 , n97743 , n97744 , n97745 , n97746 , n97747 , n97748 , n97749 , n97750 , n97751 , 
 n97752 , n97753 , n97754 , n97755 , n97756 , n97757 , n97758 , n97759 , n97760 , n97761 , 
 n97762 , n97763 , n97764 , n97765 , n97766 , n97767 , n97768 , n97769 , n97770 , n97771 , 
 n97772 , n97773 , n97774 , n97775 , n97776 , n97777 , n97778 , n97779 , n97780 , n97781 , 
 n97782 , n97783 , n97784 , n97785 , n97786 , n97787 , n97788 , n97789 , n97790 , n97791 , 
 n97792 , n97793 , n97794 , n97795 , n97796 , n97797 , n97798 , n97799 , n97800 , n97801 , 
 n97802 , n97803 , n97804 , n97805 , n97806 , n97807 , n97808 , n97809 , n97810 , n97811 , 
 n97812 , n97813 , n97814 , n97815 , n97816 , n97817 , n97818 , n97819 , n97820 , n97821 , 
 n97822 , n97823 , n97824 , n97825 , n97826 , n97827 , n97828 , n97829 , n97830 , n97831 , 
 n97832 , n97833 , n97834 , n97835 , n97836 , n97837 , n97838 , n97839 , n97840 , n97841 , 
 n97842 , n97843 , n97844 , n97845 , n97846 , n97847 , n97848 , n97849 , n97850 , n97851 , 
 n97852 , n97853 , n97854 , n97855 , n97856 , n97857 , n97858 , n97859 , n97860 , n97861 , 
 n97862 , n97863 , n97864 , n97865 , n97866 , n97867 , n97868 , n97869 , n97870 , n97871 , 
 n97872 , n97873 , n97874 , n97875 , n97876 , n97877 , n97878 , n97879 , n97880 , n97881 , 
 n97882 , n97883 , n97884 , n97885 , n97886 , n97887 , n97888 , n97889 , n97890 , n97891 , 
 n97892 , n97893 , n97894 , n97895 , n97896 , n97897 , n97898 , n97899 , n97900 , n97901 , 
 n97902 , n97903 , n97904 , n97905 , n97906 , n97907 , n97908 , n97909 , n97910 , n97911 , 
 n97912 , n97913 , n97914 , n97915 , n97916 , n97917 , n97918 , n97919 , n97920 , n97921 , 
 n97922 , n97923 , n97924 , n97925 , n97926 , n97927 , n97928 , n97929 , n97930 , n97931 , 
 n97932 , n97933 , n97934 , n97935 , n97936 , n97937 , n97938 , n97939 , n97940 , n97941 , 
 n97942 , n97943 , n97944 , n97945 , n97946 , n97947 , n97948 , n97949 , n97950 , n97951 , 
 n97952 , n97953 , n97954 , n97955 , n97956 , n97957 , n97958 , n97959 , n97960 , n97961 , 
 n97962 , n97963 , n97964 , n97965 , n97966 , n97967 , n97968 , n97969 , n97970 , n97971 , 
 n97972 , n97973 , n97974 , n97975 , n97976 , n97977 , n97978 , n97979 , n97980 , n97981 , 
 n97982 , n97983 , n97984 , n97985 , n97986 , n97987 , n97988 , n97989 , n97990 , n97991 , 
 n97992 , n97993 , n97994 , n97995 , n97996 , n97997 , n97998 , n97999 , n98000 , n98001 , 
 n98002 , n98003 , n98004 , n98005 , n98006 , n98007 , n98008 , n98009 , n98010 , n98011 , 
 n98012 , n98013 , n98014 , n98015 , n98016 , n98017 , n98018 , n98019 , n98020 , n98021 , 
 n98022 , n98023 , n98024 , n98025 , n98026 , n98027 , n98028 , n98029 , n98030 , n98031 , 
 n98032 , n98033 , n98034 , n98035 , n98036 , n98037 , n98038 , n98039 , n98040 , n98041 , 
 n98042 , n98043 , n98044 , n98045 , n98046 , n98047 , n98048 , n98049 , n98050 , n98051 , 
 n98052 , n98053 , n98054 , n98055 , n98056 , n98057 , n98058 , n98059 , n98060 , n98061 , 
 n98062 , n98063 , n98064 , n98065 , n98066 , n98067 , n98068 , n98069 , n98070 , n98071 , 
 n98072 , n98073 , n98074 , n98075 , n98076 , n98077 , n98078 , n98079 , n98080 , n98081 , 
 n98082 , n98083 , n98084 , n98085 , n98086 , n98087 , n98088 , n98089 , n98090 , n98091 , 
 n98092 , n98093 , n98094 , n98095 , n98096 , n98097 , n98098 , n98099 , n98100 , n98101 , 
 n98102 , n98103 , n98104 , n98105 , n98106 , n98107 , n98108 , n98109 , n98110 , n98111 , 
 n98112 , n98113 , n98114 , n98115 , n98116 , n98117 , n98118 , n98119 , n98120 , n98121 , 
 n98122 , n98123 , n98124 , n98125 , n98126 , n98127 , n98128 , n98129 , n98130 , n98131 , 
 n98132 , n98133 , n98134 , n98135 , n98136 , n98137 , n98138 , n98139 , n98140 , n98141 , 
 n98142 , n98143 , n98144 , n98145 , n98146 , n98147 , n98148 , n98149 , n98150 , n98151 , 
 n98152 , n98153 , n98154 , n98155 , n98156 , n98157 , n98158 , n98159 , n98160 , n98161 , 
 n98162 , n98163 , n98164 , n98165 , n98166 , n98167 , n98168 , n98169 , n98170 , n98171 , 
 n98172 , n98173 , n98174 , n98175 , n98176 , n98177 , n98178 , n98179 , n98180 , n98181 , 
 n98182 , n98183 , n98184 , n98185 , n98186 , n98187 , n98188 , n98189 , n98190 , n98191 , 
 n98192 , n98193 , n98194 , n98195 , n98196 , n98197 , n98198 , n98199 , n98200 , n98201 , 
 n98202 , n98203 , n98204 , n98205 , n98206 , n98207 , n98208 , n98209 , n98210 , n98211 , 
 n98212 , n98213 , n98214 , n98215 , n98216 , n98217 , n98218 , n98219 , n98220 , n98221 , 
 n98222 , n98223 , n98224 , n98225 , n98226 , n98227 , n98228 , n98229 , n98230 , n98231 , 
 n98232 , n98233 , n98234 , n98235 , n98236 , n98237 , n98238 , n98239 , n98240 , n98241 , 
 n98242 , n98243 , n98244 , n98245 , n98246 , n98247 , n98248 , n98249 , n98250 , n98251 , 
 n98252 , n98253 , n98254 , n98255 , n98256 , n98257 , n98258 , n98259 , n98260 , n98261 , 
 n98262 , n98263 , n98264 , n98265 , n98266 , n98267 , n98268 , n98269 , n98270 , n98271 , 
 n98272 , n98273 , n98274 , n98275 , n98276 , n98277 , n98278 , n98279 , n98280 , n98281 , 
 n98282 , n98283 , n98284 , n98285 , n98286 , n98287 , n98288 , n98289 , n98290 , n98291 , 
 n98292 , n98293 , n98294 , n98295 , n98296 , n98297 , n98298 , n98299 , n98300 , n98301 , 
 n98302 , n98303 , n98304 , n98305 , n98306 , n98307 , n98308 , n98309 , n98310 , n98311 , 
 n98312 , n98313 , n98314 , n98315 , n98316 , n98317 , n98318 , n98319 , n98320 , n98321 , 
 n98322 , n98323 , n98324 , n98325 , n98326 , n98327 , n98328 , n98329 , n98330 , n98331 , 
 n98332 , n98333 , n98334 , n98335 , n98336 , n98337 , n98338 , n98339 , n98340 , n98341 , 
 n98342 , n98343 , n98344 , n98345 , n98346 , n98347 , n98348 , n98349 , n98350 , n98351 , 
 n98352 , n98353 , n98354 , n98355 , n98356 , n98357 , n98358 , n98359 , n98360 , n98361 , 
 n98362 , n98363 , n98364 , n98365 , n98366 , n98367 , n98368 , n98369 , n98370 , n98371 , 
 n98372 , n98373 , n98374 , n98375 , n98376 , n98377 , n98378 , n98379 , n98380 , n98381 , 
 n98382 , n98383 , n98384 , n98385 , n98386 , n98387 , n98388 , n98389 , n98390 , n98391 , 
 n98392 , n98393 , n98394 , n98395 , n98396 , n98397 , n98398 , n98399 , n98400 , n98401 , 
 n98402 , n98403 , n98404 , n98405 , n98406 , n98407 , n98408 , n98409 , n98410 , n98411 , 
 n98412 , n98413 , n98414 , n98415 , n98416 , n98417 , n98418 , n98419 , n98420 , n98421 , 
 n98422 , n98423 , n98424 , n98425 , n98426 , n98427 , n98428 , n98429 , n98430 , n98431 , 
 n98432 , n98433 , n98434 , n98435 , n98436 , n98437 , n98438 , n98439 , n98440 , n98441 , 
 n98442 , n98443 , n98444 , n98445 , n98446 , n98447 , n98448 , n98449 , n98450 , n98451 , 
 n98452 , n98453 , n98454 , n98455 , n98456 , n98457 , n98458 , n98459 , n98460 , n98461 , 
 n98462 , n98463 , n98464 , n98465 , n98466 , n98467 , n98468 , n98469 , n98470 , n98471 , 
 n98472 , n98473 , n98474 , n98475 , n98476 , n98477 , n98478 , n98479 , n98480 , n98481 , 
 n98482 , n98483 , n98484 , n98485 , n98486 , n98487 , n98488 , n98489 , n98490 , n98491 , 
 n98492 , n98493 , n98494 , n98495 , n98496 , n98497 , n98498 , n98499 , n98500 , n98501 , 
 n98502 , n98503 , n98504 , n98505 , n98506 , n98507 , n98508 , n98509 , n98510 , n98511 , 
 n98512 , n98513 , n98514 , n98515 , n98516 , n98517 , n98518 , n98519 , n98520 , n98521 , 
 n98522 , n98523 , n98524 , n98525 , n98526 , n98527 , n98528 , n98529 , n98530 , n98531 , 
 n98532 , n98533 , n98534 , n98535 , n98536 , n98537 , n98538 , n98539 , n98540 , n98541 , 
 n98542 , n98543 , n98544 , n98545 , n98546 , n98547 , n98548 , n98549 , n98550 , n98551 , 
 n98552 , n98553 , n98554 , n98555 , n98556 , n98557 , n98558 , n98559 , n98560 , n98561 , 
 n98562 , n98563 , n98564 , n98565 , n98566 , n98567 , n98568 , n98569 , n98570 , n98571 , 
 n98572 , n98573 , n98574 , n98575 , n98576 , n98577 , n98578 , n98579 , n98580 , n98581 , 
 n98582 , n98583 , n98584 , n98585 , n98586 , n98587 , n98588 , n98589 , n98590 , n98591 , 
 n98592 , n98593 , n98594 , n98595 , n98596 , n98597 , n98598 , n98599 , n98600 , n98601 , 
 n98602 , n98603 , n98604 , n98605 , n98606 , n98607 , n98608 , n98609 , n98610 , n98611 , 
 n98612 , n98613 , n98614 , n98615 , n98616 , n98617 , n98618 , n98619 , n98620 , n98621 , 
 n98622 , n98623 , n98624 , n98625 , n98626 , n98627 , n98628 , n98629 , n98630 , n98631 , 
 n98632 , n98633 , n98634 , n98635 , n98636 , n98637 , n98638 , n98639 , n98640 , n98641 , 
 n98642 , n98643 , n98644 , n98645 , n98646 , n98647 , n98648 , n98649 , n98650 , n98651 , 
 n98652 , n98653 , n98654 , n98655 , n98656 , n98657 , n98658 , n98659 , n98660 , n98661 , 
 n98662 , n98663 , n98664 , n98665 , n98666 , n98667 , n98668 , n98669 , n98670 , n98671 , 
 n98672 , n98673 , n98674 , n98675 , n98676 , n98677 , n98678 , n98679 , n98680 , n98681 , 
 n98682 , n98683 , n98684 , n98685 , n98686 , n98687 , n98688 , n98689 , n98690 , n98691 , 
 n98692 , n98693 , n98694 , n98695 , n98696 , n98697 , n98698 , n98699 , n98700 , n98701 , 
 n98702 , n98703 , n98704 , n98705 , n98706 , n98707 , n98708 , n98709 , n98710 , n98711 , 
 n98712 , n98713 , n98714 , n98715 , n98716 , n98717 , n98718 , n98719 , n98720 , n98721 , 
 n98722 , n98723 , n98724 , n98725 , n98726 , n98727 , n98728 , n98729 , n98730 , n98731 , 
 n98732 , n98733 , n98734 , n98735 , n98736 , n98737 , n98738 , n98739 , n98740 , n98741 , 
 n98742 , n98743 , n98744 , n98745 , n98746 , n98747 , n98748 , n98749 , n98750 , n98751 , 
 n98752 , n98753 , n98754 , n98755 , n98756 , n98757 , n98758 , n98759 , n98760 , n98761 , 
 n98762 , n98763 , n98764 , n98765 , n98766 , n98767 , n98768 , n98769 , n98770 , n98771 , 
 n98772 , n98773 , n98774 , n98775 , n98776 , n98777 , n98778 , n98779 , n98780 , n98781 , 
 n98782 , n98783 , n98784 , n98785 , n98786 , n98787 , n98788 , n98789 , n98790 , n98791 , 
 n98792 , n98793 , n98794 , n98795 , n98796 , n98797 , n98798 , n98799 , n98800 , n98801 , 
 n98802 , n98803 , n98804 , n98805 , n98806 , n98807 , n98808 , n98809 , n98810 , n98811 , 
 n98812 , n98813 , n98814 , n98815 , n98816 , n98817 , n98818 , n98819 , n98820 , n98821 , 
 n98822 , n98823 , n98824 , n98825 , n98826 , n98827 , n98828 , n98829 , n98830 , n98831 , 
 n98832 , n98833 , n98834 , n98835 , n98836 , n98837 , n98838 , n98839 , n98840 , n98841 , 
 n98842 , n98843 , n98844 , n98845 , n98846 , n98847 , n98848 , n98849 , n98850 , n98851 , 
 n98852 , n98853 , n98854 , n98855 , n98856 , n98857 , n98858 , n98859 , n98860 , n98861 , 
 n98862 , n98863 , n98864 , n98865 , n98866 , n98867 , n98868 , n98869 , n98870 , n98871 , 
 n98872 , n98873 , n98874 , n98875 , n98876 , n98877 , n98878 , n98879 , n98880 , n98881 , 
 n98882 , n98883 , n98884 , n98885 , n98886 , n98887 , n98888 , n98889 , n98890 , n98891 , 
 n98892 , n98893 , n98894 , n98895 , n98896 , n98897 , n98898 , n98899 , n98900 , n98901 , 
 n98902 , n98903 , n98904 , n98905 , n98906 , n98907 , n98908 , n98909 , n98910 , n98911 , 
 n98912 , n98913 , n98914 , n98915 , n98916 , n98917 , n98918 , n98919 , n98920 , n98921 , 
 n98922 , n98923 , n98924 , n98925 , n98926 , n98927 , n98928 , n98929 , n98930 , n98931 , 
 n98932 , n98933 , n98934 , n98935 , n98936 , n98937 , n98938 , n98939 , n98940 , n98941 , 
 n98942 , n98943 , n98944 , n98945 , n98946 , n98947 , n98948 , n98949 , n98950 , n98951 , 
 n98952 , n98953 , n98954 , n98955 , n98956 , n98957 , n98958 , n98959 , n98960 , n98961 , 
 n98962 , n98963 , n98964 , n98965 , n98966 , n98967 , n98968 , n98969 , n98970 , n98971 , 
 n98972 , n98973 , n98974 , n98975 , n98976 , n98977 , n98978 , n98979 , n98980 , n98981 , 
 n98982 , n98983 , n98984 , n98985 , n98986 , n98987 , n98988 , n98989 , n98990 , n98991 , 
 C0n , C0 , C1n , C1 ;
buf ( n454 , n0 );
buf ( n455 , n1 );
buf ( n456 , n2 );
buf ( n457 , n3 );
buf ( n458 , n4 );
buf ( n459 , n5 );
buf ( n460 , n6 );
buf ( n461 , n7 );
buf ( n462 , n8 );
buf ( n463 , n9 );
buf ( n464 , n10 );
buf ( n465 , n11 );
buf ( n466 , n12 );
buf ( n467 , n13 );
buf ( n468 , n14 );
buf ( n469 , n15 );
buf ( n470 , n16 );
buf ( n471 , n17 );
buf ( n472 , n18 );
buf ( n473 , n19 );
buf ( n474 , n20 );
buf ( n475 , n21 );
buf ( n476 , n22 );
buf ( n477 , n23 );
buf ( n478 , n24 );
buf ( n479 , n25 );
buf ( n480 , n26 );
buf ( n481 , n27 );
buf ( n482 , n28 );
buf ( n483 , n29 );
buf ( n484 , n30 );
buf ( n485 , n31 );
buf ( n486 , n32 );
buf ( n487 , n33 );
buf ( n488 , n34 );
buf ( n489 , n35 );
buf ( n490 , n36 );
buf ( n491 , n37 );
buf ( n492 , n38 );
buf ( n493 , n39 );
buf ( n494 , n40 );
buf ( n495 , n41 );
buf ( n496 , n42 );
buf ( n497 , n43 );
buf ( n498 , n44 );
buf ( n499 , n45 );
buf ( n500 , n46 );
buf ( n501 , n47 );
buf ( n502 , n48 );
buf ( n503 , n49 );
buf ( n504 , n50 );
buf ( n505 , n51 );
buf ( n506 , n52 );
buf ( n507 , n53 );
buf ( n508 , n54 );
buf ( n509 , n55 );
buf ( n510 , n56 );
buf ( n511 , n57 );
buf ( n512 , n58 );
buf ( n513 , n59 );
buf ( n514 , n60 );
buf ( n515 , n61 );
buf ( n516 , n62 );
buf ( n517 , n63 );
buf ( n518 , n64 );
buf ( n519 , n65 );
buf ( n520 , n66 );
buf ( n521 , n67 );
buf ( n522 , n68 );
buf ( n523 , n69 );
buf ( n524 , n70 );
buf ( n525 , n71 );
buf ( n526 , n72 );
buf ( n527 , n73 );
buf ( n528 , n74 );
buf ( n529 , n75 );
buf ( n530 , n76 );
buf ( n531 , n77 );
buf ( n532 , n78 );
buf ( n533 , n79 );
buf ( n534 , n80 );
buf ( n535 , n81 );
buf ( n536 , n82 );
buf ( n537 , n83 );
buf ( n538 , n84 );
buf ( n539 , n85 );
buf ( n540 , n86 );
buf ( n541 , n87 );
buf ( n542 , n88 );
buf ( n543 , n89 );
buf ( n544 , n90 );
buf ( n545 , n91 );
buf ( n546 , n92 );
buf ( n547 , n93 );
buf ( n548 , n94 );
buf ( n549 , n95 );
buf ( n550 , n96 );
buf ( n551 , n97 );
buf ( n552 , n98 );
buf ( n99 , n553 );
buf ( n100 , n554 );
buf ( n101 , n555 );
buf ( n102 , n556 );
buf ( n103 , n557 );
buf ( n104 , n558 );
buf ( n105 , n559 );
buf ( n106 , n560 );
buf ( n107 , n561 );
buf ( n108 , n562 );
buf ( n109 , n563 );
buf ( n110 , n564 );
buf ( n111 , n565 );
buf ( n112 , n566 );
buf ( n113 , n567 );
buf ( n114 , n568 );
buf ( n115 , n569 );
buf ( n116 , n570 );
buf ( n117 , n571 );
buf ( n118 , n572 );
buf ( n119 , n573 );
buf ( n120 , n574 );
buf ( n121 , n575 );
buf ( n122 , n576 );
buf ( n123 , n577 );
buf ( n124 , n578 );
buf ( n125 , n579 );
buf ( n126 , n580 );
buf ( n127 , n581 );
buf ( n128 , n582 );
buf ( n129 , n583 );
buf ( n130 , n584 );
buf ( n131 , n585 );
buf ( n132 , n586 );
buf ( n133 , n587 );
buf ( n134 , n588 );
buf ( n135 , n589 );
buf ( n136 , n590 );
buf ( n137 , n591 );
buf ( n138 , n592 );
buf ( n139 , n593 );
buf ( n140 , n594 );
buf ( n141 , n595 );
buf ( n142 , n596 );
buf ( n143 , n597 );
buf ( n144 , n598 );
buf ( n145 , n599 );
buf ( n146 , n600 );
buf ( n147 , n601 );
buf ( n148 , n602 );
buf ( n149 , n603 );
buf ( n150 , n604 );
buf ( n151 , n605 );
buf ( n152 , n606 );
buf ( n153 , n607 );
buf ( n154 , n608 );
buf ( n155 , n609 );
buf ( n156 , n610 );
buf ( n157 , n611 );
buf ( n158 , n612 );
buf ( n159 , n613 );
buf ( n160 , n614 );
buf ( n161 , n615 );
buf ( n162 , n616 );
buf ( n163 , n617 );
buf ( n164 , n618 );
buf ( n165 , n619 );
buf ( n166 , n620 );
buf ( n167 , n621 );
buf ( n168 , n622 );
buf ( n169 , n623 );
buf ( n170 , n624 );
buf ( n171 , n625 );
buf ( n172 , n626 );
buf ( n173 , n627 );
buf ( n174 , n628 );
buf ( n175 , n629 );
buf ( n176 , n630 );
buf ( n177 , n631 );
buf ( n178 , n632 );
buf ( n179 , n633 );
buf ( n180 , n634 );
buf ( n181 , n635 );
buf ( n182 , n636 );
buf ( n183 , n637 );
buf ( n184 , n638 );
buf ( n185 , n639 );
buf ( n186 , n640 );
buf ( n187 , n641 );
buf ( n188 , n642 );
buf ( n189 , n643 );
buf ( n190 , n644 );
buf ( n191 , n645 );
buf ( n192 , n646 );
buf ( n193 , n647 );
buf ( n194 , n648 );
buf ( n195 , n649 );
buf ( n196 , n650 );
buf ( n197 , n651 );
buf ( n198 , n652 );
buf ( n199 , n653 );
buf ( n200 , n654 );
buf ( n201 , n655 );
buf ( n202 , n656 );
buf ( n203 , n657 );
buf ( n204 , n658 );
buf ( n205 , n659 );
buf ( n206 , n660 );
buf ( n207 , n661 );
buf ( n208 , n662 );
buf ( n209 , n663 );
buf ( n210 , n664 );
buf ( n211 , n665 );
buf ( n212 , n666 );
buf ( n213 , n667 );
buf ( n214 , n668 );
buf ( n215 , n669 );
buf ( n216 , n670 );
buf ( n217 , n671 );
buf ( n218 , n672 );
buf ( n219 , n673 );
buf ( n220 , n674 );
buf ( n221 , n675 );
buf ( n222 , n676 );
buf ( n223 , n677 );
buf ( n224 , n678 );
buf ( n225 , n679 );
buf ( n226 , n680 );
buf ( n553 , C0 );
buf ( n554 , C0 );
buf ( n555 , C0 );
buf ( n556 , C0 );
buf ( n557 , C0 );
buf ( n558 , C0 );
buf ( n559 , C0 );
buf ( n560 , C0 );
buf ( n561 , C0 );
buf ( n562 , C0 );
buf ( n563 , C0 );
buf ( n564 , C0 );
buf ( n565 , C0 );
buf ( n566 , C0 );
buf ( n567 , C0 );
buf ( n568 , C0 );
buf ( n569 , n98439 );
buf ( n570 , n98451 );
buf ( n571 , n98441 );
buf ( n572 , n98308 );
buf ( n573 , n97286 );
buf ( n574 , n98226 );
buf ( n575 , n98173 );
buf ( n576 , n98134 );
buf ( n577 , n94938 );
buf ( n578 , n95072 );
buf ( n579 , n95113 );
buf ( n580 , n94973 );
buf ( n581 , n95146 );
buf ( n582 , n95142 );
buf ( n583 , n95175 );
buf ( n584 , n98991 );
buf ( n585 , n16704 );
buf ( n586 , n16712 );
buf ( n587 , n15958 );
buf ( n588 , n16033 );
buf ( n589 , n16048 );
buf ( n590 , n15995 );
buf ( n591 , n16758 );
buf ( n592 , n17504 );
buf ( n593 , n17477 );
buf ( n594 , n17483 );
buf ( n595 , n17514 );
buf ( n596 , n16880 );
buf ( n597 , n16786 );
buf ( n598 , n16835 );
buf ( n599 , n16846 );
buf ( n600 , n16817 );
buf ( n601 , n16895 );
buf ( n602 , n16942 );
buf ( n603 , n16983 );
buf ( n604 , n17020 );
buf ( n605 , n17055 );
buf ( n606 , n17098 );
buf ( n607 , n17135 );
buf ( n608 , n17173 );
buf ( n609 , n17211 );
buf ( n610 , n17246 );
buf ( n611 , n17265 );
buf ( n612 , n98863 );
buf ( n613 , n98873 );
buf ( n614 , n98975 );
buf ( n615 , n98877 );
buf ( n616 , n96987 );
buf ( n617 , C0 );
buf ( n618 , C0 );
buf ( n619 , C0 );
buf ( n620 , C0 );
buf ( n621 , C0 );
buf ( n622 , C0 );
buf ( n623 , C0 );
buf ( n624 , C0 );
buf ( n625 , C0 );
buf ( n626 , C0 );
buf ( n627 , C0 );
buf ( n628 , C0 );
buf ( n629 , C0 );
buf ( n630 , C0 );
buf ( n631 , C0 );
buf ( n632 , C0 );
buf ( n633 , n98918 );
buf ( n634 , n98748 );
buf ( n635 , n98739 );
buf ( n636 , n98794 );
buf ( n637 , n98960 );
buf ( n638 , n98727 );
buf ( n639 , n98841 );
buf ( n640 , n98791 );
buf ( n641 , n98765 );
buf ( n642 , n98810 );
buf ( n643 , n98705 );
buf ( n644 , n98828 );
buf ( n645 , n96699 );
buf ( n646 , n98663 );
buf ( n647 , n96760 );
buf ( n648 , n98680 );
buf ( n649 , n98653 );
buf ( n650 , n96827 );
buf ( n651 , n98636 );
buf ( n652 , n96859 );
buf ( n653 , n93516 );
buf ( n654 , n98969 );
buf ( n655 , n98990 );
buf ( n656 , n93560 );
buf ( n657 , n93571 );
buf ( n658 , n93583 );
buf ( n659 , n98911 );
buf ( n660 , n93610 );
buf ( n661 , n98901 );
buf ( n662 , n93627 );
buf ( n663 , n96717 );
buf ( n664 , n96724 );
buf ( n665 , n96743 );
buf ( n666 , n96772 );
buf ( n667 , n98943 );
buf ( n668 , n96786 );
buf ( n669 , n98857 );
buf ( n670 , n98923 );
buf ( n671 , n96798 );
buf ( n672 , n96809 );
buf ( n673 , n96834 );
buf ( n674 , n98928 );
buf ( n675 , n97002 );
buf ( n676 , n98986 );
buf ( n677 , n98882 );
buf ( n678 , n98948 );
buf ( n679 , n98974 );
buf ( n680 , n98869 );
not ( n70358 , n504 );
nand ( n70359 , n70358 , n503 );
not ( n70360 , n70359 );
xor ( n70361 , n503 , n520 );
and ( n70362 , n70360 , n70361 );
not ( n70363 , n70362 );
not ( n70364 , n502 );
not ( n70365 , n503 );
not ( n70366 , n70365 );
or ( n70367 , n70364 , n70366 );
not ( n70368 , n502 );
nand ( n70369 , n70368 , n503 );
nand ( n70370 , n70367 , n70369 );
buf ( n70371 , n70370 );
nand ( n70372 , n520 , n70371 );
nand ( n70373 , n70363 , n70372 );
xor ( n70374 , n503 , n519 );
not ( n70375 , n70374 );
nand ( n70376 , n503 , n504 );
nor ( n70377 , n70375 , n70376 , n520 );
or ( n70378 , n70373 , n70377 );
not ( n70379 , n70374 );
not ( n70380 , n70360 );
or ( n70381 , n70379 , n70380 );
xor ( n70382 , n518 , n503 );
nand ( n70383 , n70382 , n504 );
nand ( n70384 , n70381 , n70383 );
nand ( n70385 , n70378 , n70384 );
nand ( n70386 , C1 , n70385 );
not ( n70387 , n70386 );
not ( n70388 , n504 );
xor ( n70389 , n503 , n517 );
not ( n70390 , n70389 );
or ( n70391 , n70388 , n70390 );
nand ( n70392 , n70382 , n70360 );
nand ( n70393 , n70391 , n70392 );
or ( n70394 , n520 , n502 );
nand ( n70395 , n70394 , n503 );
nand ( n70396 , n520 , n502 );
and ( n70397 , n70395 , n70396 , n501 );
and ( n70398 , n70393 , n70397 );
not ( n70399 , n70393 );
not ( n70400 , n70397 );
and ( n70401 , n70399 , n70400 );
nor ( n70402 , n70398 , n70401 );
xor ( n70403 , n501 , n520 );
not ( n70404 , n70403 );
and ( n70405 , n502 , n503 );
not ( n70406 , n502 );
not ( n70407 , n503 );
and ( n70408 , n70406 , n70407 );
nor ( n70409 , n70405 , n70408 );
not ( n70410 , n70409 );
xor ( n70411 , n501 , n502 );
nand ( n70412 , n70410 , n70411 );
not ( n70413 , n70412 );
not ( n70414 , n70413 );
or ( n70415 , n70404 , n70414 );
xor ( n70416 , n519 , n501 );
nand ( n70417 , n70416 , n70371 );
nand ( n70418 , n70415 , n70417 );
nor ( n70419 , n70402 , n70418 );
not ( n70420 , n70419 );
not ( n70421 , n70420 );
or ( n70422 , n70387 , n70421 );
nand ( n70423 , n70418 , n70402 );
nand ( n70424 , n70422 , n70423 );
not ( n70425 , n70424 );
xor ( n70426 , n500 , n501 );
and ( n70427 , n70426 , n520 );
not ( n70428 , n70427 );
nand ( n70429 , n70411 , n70416 );
or ( n70430 , n70429 , n70371 );
not ( n70431 , n518 );
not ( n70432 , n501 );
not ( n70433 , n70432 );
or ( n70434 , n70431 , n70433 );
not ( n70435 , n518 );
nand ( n70436 , n70435 , n501 );
nand ( n70437 , n70434 , n70436 );
xor ( n70438 , n502 , n503 );
nand ( n70439 , n70437 , n70438 );
nand ( n70440 , n70430 , n70439 );
not ( n70441 , n70440 );
not ( n70442 , n70441 );
or ( n70443 , n70428 , n70442 );
not ( n70444 , n70427 );
nand ( n70445 , n70444 , n70440 );
nand ( n70446 , n70443 , n70445 );
not ( n70447 , n504 );
xor ( n70448 , n503 , n516 );
not ( n70449 , n70448 );
or ( n70450 , n70447 , n70449 );
nand ( n70451 , n70389 , n70360 );
nand ( n70452 , n70450 , n70451 );
not ( n70453 , n70452 );
and ( n70454 , n70446 , n70453 );
not ( n70455 , n70446 );
and ( n70456 , n70455 , n70452 );
nor ( n70457 , n70454 , n70456 );
and ( n70458 , n70393 , n70397 );
and ( n70459 , n70457 , n70458 );
nand ( n70460 , n70425 , n70459 );
not ( n70461 , n70458 );
nand ( n70462 , n70457 , n70461 );
not ( n70463 , n70462 );
nor ( n70464 , n70457 , n70461 );
or ( n70465 , n70463 , n70464 );
nand ( n70466 , n70465 , n70424 );
nor ( n70467 , n70457 , n70458 );
nand ( n70468 , n70425 , n70467 );
nand ( n70469 , n70460 , n70466 , n70468 );
not ( n70470 , n455 );
nand ( n70471 , n70469 , n70470 );
not ( n70472 , n70438 );
xor ( n70473 , n513 , n501 );
not ( n70474 , n70473 );
or ( n70475 , n70472 , n70474 );
xor ( n70476 , n501 , n514 );
not ( n70477 , n503 );
nand ( n70478 , n70477 , n502 );
nand ( n70479 , n503 , n70368 );
nand ( n70480 , n70411 , n70476 , n70478 , n70479 );
nand ( n70481 , n70475 , n70480 );
not ( n70482 , n497 );
or ( n70483 , n520 , n496 );
not ( n70484 , n70483 );
or ( n70485 , n70482 , n70484 );
nand ( n70486 , n520 , n496 );
and ( n70487 , n70486 , n495 );
nand ( n70488 , n70485 , n70487 );
not ( n70489 , n70488 );
and ( n70490 , n70481 , n70489 );
xor ( n70491 , n494 , n495 );
nand ( n70492 , n70491 , n520 );
and ( n70493 , n517 , n497 );
not ( n70494 , n517 );
not ( n70495 , n497 );
and ( n70496 , n70494 , n70495 );
nor ( n70497 , n70493 , n70496 );
not ( n70498 , n70497 );
xor ( n70499 , n498 , n499 );
not ( n70500 , n70499 );
not ( n70501 , n497 );
not ( n70502 , n498 );
not ( n70503 , n70502 );
or ( n70504 , n70501 , n70503 );
not ( n70505 , n497 );
nand ( n70506 , n70505 , n498 );
nand ( n70507 , n70504 , n70506 );
nand ( n70508 , n70500 , n70507 );
not ( n70509 , n70508 );
not ( n70510 , n70509 );
or ( n70511 , n70498 , n70510 );
xor ( n70512 , n516 , n497 );
buf ( n70513 , n70499 );
nand ( n70514 , n70512 , n70513 );
nand ( n70515 , n70511 , n70514 );
xor ( n70516 , n70492 , n70515 );
and ( n70517 , n70473 , n70411 );
not ( n70518 , n70517 );
not ( n70519 , n70371 );
not ( n70520 , n70519 );
or ( n70521 , n70518 , n70520 );
not ( n70522 , n70410 );
xor ( n70523 , n512 , n501 );
nand ( n70524 , n70522 , n70523 );
nand ( n70525 , n70521 , n70524 );
xnor ( n70526 , n70516 , n70525 );
xor ( n70527 , n70490 , n70526 );
xor ( n70528 , n520 , n495 );
not ( n70529 , n70528 );
not ( n70530 , n497 );
nor ( n70531 , n70530 , n496 );
not ( n70532 , n70531 );
nand ( n70533 , n70495 , n496 );
xor ( n70534 , n496 , n495 );
nand ( n70535 , n70532 , n70533 , n70534 );
not ( n70536 , n70535 );
not ( n70537 , n70536 );
or ( n70538 , n70529 , n70537 );
and ( n70539 , n496 , n497 );
not ( n70540 , n496 );
not ( n70541 , n497 );
and ( n70542 , n70540 , n70541 );
nor ( n70543 , n70539 , n70542 );
buf ( n70544 , n70543 );
xor ( n70545 , n519 , n495 );
nand ( n70546 , n70544 , n70545 );
nand ( n70547 , n70538 , n70546 );
not ( n70548 , n70547 );
and ( n70549 , n503 , n512 );
not ( n70550 , n503 );
not ( n70551 , n512 );
and ( n70552 , n70550 , n70551 );
nor ( n70553 , n70549 , n70552 );
not ( n70554 , n70553 );
not ( n70555 , n70360 );
or ( n70556 , n70554 , n70555 );
xor ( n70557 , n511 , n503 );
nand ( n70558 , n70557 , n504 );
nand ( n70559 , n70556 , n70558 );
not ( n70560 , n70559 );
or ( n70561 , n70548 , n70560 );
nor ( n70562 , n70559 , n70547 );
xor ( n70563 , n518 , n497 );
not ( n70564 , n70563 );
and ( n70565 , n70500 , n70507 );
not ( n70566 , n70565 );
or ( n70567 , n70564 , n70566 );
nand ( n70568 , n70513 , n70497 );
nand ( n70569 , n70567 , n70568 );
not ( n70570 , n70569 );
or ( n70571 , n70562 , n70570 );
nand ( n70572 , n70561 , n70571 );
xor ( n70573 , n70527 , n70572 );
not ( n70574 , n504 );
xor ( n70575 , n503 , n510 );
not ( n70576 , n70575 );
or ( n70577 , n70574 , n70576 );
nand ( n70578 , n70557 , n70360 );
nand ( n70579 , n70577 , n70578 );
not ( n70580 , n70579 );
not ( n70581 , n70580 );
not ( n70582 , n70545 );
not ( n70583 , n70505 );
not ( n70584 , n496 );
not ( n70585 , n70584 );
or ( n70586 , n70583 , n70585 );
nand ( n70587 , n496 , n497 );
nand ( n70588 , n70586 , n70587 );
and ( n70589 , n70588 , n70534 );
not ( n70590 , n70589 );
or ( n70591 , n70582 , n70590 );
and ( n70592 , n518 , n495 );
not ( n70593 , n518 );
not ( n70594 , n495 );
and ( n70595 , n70593 , n70594 );
nor ( n70596 , n70592 , n70595 );
nand ( n70597 , n70543 , n70596 );
nand ( n70598 , n70591 , n70597 );
not ( n70599 , n70598 );
or ( n70600 , n70581 , n70599 );
not ( n70601 , n70598 );
nand ( n70602 , n70601 , n70579 );
nand ( n70603 , n70600 , n70602 );
xor ( n70604 , n499 , n515 );
not ( n70605 , n70604 );
and ( n70606 , n500 , n501 );
not ( n70607 , n500 );
not ( n70608 , n501 );
and ( n70609 , n70607 , n70608 );
nor ( n70610 , n70606 , n70609 );
not ( n70611 , n70610 );
not ( n70612 , n500 );
not ( n70613 , n499 );
nand ( n70614 , n70612 , n70613 );
nand ( n70615 , n500 , n499 );
and ( n70616 , n70611 , n70614 , n70615 );
not ( n70617 , n70616 );
or ( n70618 , n70605 , n70617 );
xor ( n70619 , n514 , n499 );
nand ( n70620 , n70426 , n70619 );
nand ( n70621 , n70618 , n70620 );
xnor ( n70622 , n70603 , n70621 );
not ( n70623 , n70360 );
xor ( n70624 , n513 , n503 );
not ( n70625 , n70624 );
or ( n70626 , n70623 , n70625 );
nand ( n70627 , n70553 , n504 );
nand ( n70628 , n70626 , n70627 );
not ( n70629 , n70628 );
nand ( n70630 , n70544 , n520 );
not ( n70631 , n70630 );
not ( n70632 , n70631 );
or ( n70633 , n70629 , n70632 );
not ( n70634 , n70630 );
not ( n70635 , n70628 );
not ( n70636 , n70635 );
or ( n70637 , n70634 , n70636 );
xor ( n70638 , n519 , n497 );
not ( n70639 , n70638 );
buf ( n70640 , n70509 );
not ( n70641 , n70640 );
or ( n70642 , n70639 , n70641 );
nand ( n70643 , n70513 , n70563 );
nand ( n70644 , n70642 , n70643 );
nand ( n70645 , n70637 , n70644 );
nand ( n70646 , n70633 , n70645 );
not ( n70647 , n70646 );
xor ( n70648 , n516 , n499 );
not ( n70649 , n70648 );
xor ( n70650 , n500 , n499 );
nand ( n70651 , n70611 , n70650 );
not ( n70652 , n70651 );
not ( n70653 , n70652 );
or ( n70654 , n70649 , n70653 );
xor ( n70655 , n500 , n501 );
nand ( n70656 , n70655 , n70604 );
nand ( n70657 , n70654 , n70656 );
not ( n70658 , n70657 );
not ( n70659 , n70489 );
not ( n70660 , n70481 );
or ( n70661 , n70659 , n70660 );
or ( n70662 , n70481 , n70489 );
nand ( n70663 , n70661 , n70662 );
nand ( n70664 , n70658 , n70663 );
not ( n70665 , n70664 );
or ( n70666 , n70647 , n70665 );
not ( n70667 , n70663 );
nand ( n70668 , n70667 , n70657 );
nand ( n70669 , n70666 , n70668 );
or ( n70670 , n70622 , n70669 );
nand ( n70671 , n70622 , n70669 );
nand ( n70672 , n70670 , n70671 );
not ( n70673 , n70672 );
and ( n70674 , n70573 , n70673 );
not ( n70675 , n70573 );
and ( n70676 , n70675 , n70672 );
nor ( n70677 , n70674 , n70676 );
not ( n70678 , n70646 );
not ( n70679 , n70678 );
and ( n70680 , n70657 , n70663 );
not ( n70681 , n70657 );
and ( n70682 , n70481 , n70488 );
not ( n70683 , n70481 );
and ( n70684 , n70683 , n70489 );
or ( n70685 , n70682 , n70684 );
and ( n70686 , n70681 , n70685 );
nor ( n70687 , n70680 , n70686 );
not ( n70688 , n70687 );
not ( n70689 , n70688 );
or ( n70690 , n70679 , n70689 );
nand ( n70691 , n70687 , n70646 );
nand ( n70692 , n70690 , n70691 );
xor ( n70693 , n515 , n501 );
not ( n70694 , n70693 );
not ( n70695 , n70413 );
or ( n70696 , n70694 , n70695 );
nand ( n70697 , n70371 , n70476 );
nand ( n70698 , n70696 , n70697 );
not ( n70699 , n70698 );
xor ( n70700 , n517 , n499 );
not ( n70701 , n70700 );
not ( n70702 , n70652 );
or ( n70703 , n70701 , n70702 );
xor ( n70704 , n500 , n501 );
nand ( n70705 , n70704 , n70648 );
nand ( n70706 , n70703 , n70705 );
not ( n70707 , n70706 );
nand ( n70708 , n520 , n498 );
or ( n70709 , n520 , n498 );
nand ( n70710 , n70709 , n499 );
nand ( n70711 , n70708 , n70710 , n497 );
not ( n70712 , n70711 );
xor ( n70713 , n514 , n503 );
not ( n70714 , n70713 );
not ( n70715 , n70360 );
or ( n70716 , n70714 , n70715 );
nand ( n70717 , n70624 , n504 );
nand ( n70718 , n70716 , n70717 );
nand ( n70719 , n70712 , n70718 );
nand ( n70720 , n70707 , n70719 );
not ( n70721 , n70720 );
or ( n682 , n70699 , n70721 );
not ( n70723 , n70719 );
nand ( n684 , n70723 , n70706 );
nand ( n70725 , n682 , n684 );
buf ( n686 , n70725 );
or ( n687 , n70692 , n686 );
not ( n70728 , n70547 );
not ( n689 , n70559 );
xor ( n690 , n689 , n70569 );
xnor ( n691 , n70728 , n690 );
not ( n692 , n691 );
nand ( n693 , n687 , n692 );
nand ( n70734 , n70692 , n686 );
nand ( n695 , n70677 , n693 , n70734 );
not ( n696 , n695 );
xor ( n697 , n520 , n499 );
not ( n698 , n697 );
not ( n699 , n70651 );
not ( n700 , n699 );
or ( n701 , n698 , n700 );
xor ( n70742 , n519 , n499 );
nand ( n703 , n70655 , n70742 );
nand ( n70744 , n701 , n703 );
not ( n705 , n70744 );
not ( n706 , n70448 );
not ( n707 , n70360 );
or ( n708 , n706 , n707 );
xor ( n709 , n515 , n503 );
nand ( n70750 , n709 , n504 );
nand ( n711 , n708 , n70750 );
or ( n712 , n520 , n500 );
nand ( n713 , n712 , n501 );
nand ( n714 , n520 , n500 );
nand ( n715 , n713 , n714 , n499 );
and ( n716 , n711 , n715 );
not ( n717 , n711 );
not ( n718 , n715 );
and ( n719 , n717 , n718 );
nor ( n720 , n716 , n719 );
not ( n721 , n720 );
or ( n722 , n705 , n721 );
or ( n723 , n720 , n70744 );
nand ( n724 , n722 , n723 );
xor ( n725 , n517 , n501 );
and ( n726 , n725 , n70371 );
not ( n727 , n70437 );
nand ( n728 , n70410 , n70411 );
nor ( n729 , n727 , n728 );
nor ( n730 , n726 , n729 );
not ( n731 , n730 );
and ( n732 , n724 , n731 );
not ( n733 , n724 );
and ( n734 , n733 , n730 );
nor ( n735 , n732 , n734 );
not ( n736 , n70427 );
nand ( n70777 , n736 , n70453 );
buf ( n741 , n70440 );
nand ( n70779 , n70777 , n741 );
nand ( n743 , n70427 , n70452 );
nand ( n70781 , n70779 , n743 );
nand ( n745 , n735 , n70781 );
not ( n70783 , n745 );
not ( n747 , n70462 );
not ( n748 , n70424 );
or ( n70786 , n747 , n748 );
not ( n750 , n70464 );
nand ( n751 , n70786 , n750 );
nor ( n752 , n70783 , n751 );
not ( n753 , n735 );
not ( n754 , n741 );
not ( n758 , n70777 );
or ( n70793 , n754 , n758 );
nand ( n760 , n70793 , n743 );
not ( n761 , n760 );
nand ( n762 , n753 , n761 );
nand ( n763 , n711 , n718 );
not ( n764 , n763 );
not ( n765 , n764 );
not ( n766 , n70742 );
not ( n770 , n699 );
or ( n70802 , n766 , n770 );
xor ( n772 , n518 , n499 );
nand ( n70804 , n70704 , n772 );
nand ( n774 , n70802 , n70804 );
not ( n775 , n774 );
not ( n776 , n775 );
or ( n777 , n765 , n776 );
nand ( n778 , n774 , n763 );
nand ( n782 , n777 , n778 );
not ( n70811 , n70360 );
not ( n784 , n709 );
or ( n785 , n70811 , n784 );
nand ( n786 , n70713 , n504 );
nand ( n787 , n785 , n786 );
not ( n788 , n787 );
nand ( n789 , n70513 , n520 );
not ( n790 , n789 );
not ( n791 , n790 );
or ( n792 , n788 , n791 );
not ( n793 , n787 );
nand ( n794 , n793 , n789 );
nand ( n795 , n792 , n794 );
not ( n796 , n725 );
not ( n797 , n70413 );
or ( n798 , n796 , n797 );
xor ( n799 , n516 , n501 );
nand ( n800 , n70371 , n799 );
nand ( n801 , n798 , n800 );
not ( n802 , n801 );
and ( n803 , n795 , n802 );
not ( n804 , n795 );
and ( n805 , n804 , n801 );
nor ( n806 , n803 , n805 );
not ( n807 , n806 );
and ( n808 , n782 , n807 );
not ( n809 , n782 );
and ( n70838 , n809 , n806 );
nor ( n814 , n808 , n70838 );
nand ( n815 , n70744 , n731 );
not ( n70841 , n730 );
not ( n817 , n70744 );
not ( n818 , n817 );
or ( n819 , n70841 , n818 );
not ( n820 , n720 );
nand ( n821 , n819 , n820 );
nand ( n822 , n814 , n815 , n821 );
nand ( n823 , n762 , n822 );
nor ( n824 , n752 , n823 );
not ( n825 , n824 );
not ( n70851 , n774 );
not ( n827 , n764 );
or ( n828 , n70851 , n827 );
nand ( n829 , n763 , n775 );
nand ( n830 , n829 , n806 );
nand ( n831 , n828 , n830 );
not ( n832 , n831 );
not ( n833 , n789 );
not ( n834 , n793 );
or ( n835 , n833 , n834 );
nand ( n836 , n835 , n801 );
nand ( n837 , n787 , n790 );
nand ( n70863 , n836 , n837 );
not ( n839 , n70863 );
not ( n843 , n70718 );
not ( n70866 , n70711 );
and ( n845 , n843 , n70866 );
and ( n846 , n70718 , n70711 );
nor ( n847 , n845 , n846 );
not ( n848 , n847 );
and ( n849 , n839 , n848 );
and ( n850 , n70863 , n847 );
nor ( n851 , n849 , n850 );
not ( n852 , n772 );
not ( n853 , n70616 );
or ( n70876 , n852 , n853 );
nand ( n855 , n70700 , n70426 );
nand ( n856 , n70876 , n855 );
not ( n857 , n856 );
not ( n858 , n799 );
not ( n859 , n70413 );
or ( n860 , n858 , n859 );
nand ( n861 , n70371 , n70693 );
nand ( n862 , n860 , n861 );
not ( n863 , n862 );
not ( n864 , n863 );
or ( n70887 , n857 , n864 );
not ( n869 , n856 );
nand ( n870 , n862 , n869 );
nand ( n871 , n70887 , n870 );
xor ( n872 , n520 , n497 );
not ( n873 , n872 );
not ( n874 , n70640 );
or ( n70894 , n873 , n874 );
nand ( n876 , n70513 , n70638 );
nand ( n877 , n70894 , n876 );
and ( n878 , n871 , n877 );
not ( n879 , n871 );
not ( n880 , n877 );
and ( n70900 , n879 , n880 );
nor ( n882 , n878 , n70900 );
not ( n883 , n882 );
and ( n884 , n851 , n883 );
not ( n885 , n851 );
and ( n886 , n885 , n882 );
nor ( n887 , n884 , n886 );
not ( n888 , n887 );
nand ( n889 , n832 , n888 );
not ( n890 , n889 );
or ( n891 , n825 , n890 );
not ( n892 , n763 );
nand ( n893 , n892 , n774 );
not ( n894 , n893 );
not ( n895 , n830 );
or ( n896 , n894 , n895 );
nand ( n897 , n896 , n887 );
not ( n898 , n897 );
not ( n899 , n814 );
nand ( n900 , n815 , n821 );
nand ( n901 , n899 , n900 );
not ( n902 , n901 );
or ( n903 , n898 , n902 );
nand ( n904 , n903 , n889 );
nand ( n905 , n891 , n904 );
not ( n906 , n905 );
and ( n907 , n70628 , n70630 );
not ( n908 , n70628 );
and ( n909 , n70544 , n520 );
and ( n910 , n908 , n909 );
nor ( n70930 , n907 , n910 );
and ( n912 , n70930 , n70644 );
not ( n913 , n70930 );
not ( n914 , n70644 );
and ( n915 , n913 , n914 );
nor ( n916 , n912 , n915 );
not ( n917 , n869 );
not ( n918 , n863 );
or ( n919 , n917 , n918 );
nand ( n70939 , n919 , n877 );
nand ( n921 , n862 , n856 );
nand ( n922 , n916 , n70939 , n921 );
not ( n923 , n922 );
nand ( n924 , n684 , n70720 );
xnor ( n925 , n924 , n70698 );
not ( n926 , n925 );
or ( n927 , n923 , n926 );
not ( n928 , n916 );
nand ( n929 , n70939 , n921 );
nand ( n930 , n928 , n929 );
nand ( n931 , n927 , n930 );
not ( n932 , n931 );
not ( n933 , n691 );
not ( n937 , n70725 );
and ( n70954 , n933 , n937 );
and ( n939 , n70725 , n691 );
nor ( n940 , n70954 , n939 );
xor ( n941 , n70692 , n940 );
nand ( n942 , n932 , n941 );
not ( n943 , n916 );
not ( n944 , n943 );
not ( n945 , n929 );
not ( n946 , n945 );
or ( n947 , n944 , n946 );
nand ( n948 , n929 , n916 );
nand ( n949 , n947 , n948 );
not ( n950 , n925 );
and ( n951 , n949 , n950 );
not ( n70968 , n949 );
and ( n956 , n70968 , n925 );
nor ( n957 , n951 , n956 );
not ( n958 , n883 );
not ( n959 , n70863 );
nand ( n960 , n959 , n847 );
and ( n961 , n958 , n960 );
not ( n962 , n70863 );
nor ( n963 , n962 , n847 );
nor ( n70977 , n961 , n963 );
nand ( n965 , n957 , n70977 );
and ( n966 , n942 , n965 );
not ( n967 , n966 );
or ( n968 , n906 , n967 );
not ( n969 , n941 );
nand ( n970 , n969 , n931 );
not ( n971 , n970 );
not ( n972 , n957 );
not ( n973 , n70977 );
nand ( n70987 , n972 , n973 );
not ( n975 , n70987 );
or ( n976 , n971 , n975 );
buf ( n977 , n942 );
nand ( n978 , n976 , n977 );
nand ( n979 , n968 , n978 );
not ( n980 , n979 );
or ( n981 , n696 , n980 );
nand ( n982 , n70734 , n693 );
not ( n983 , n70673 );
buf ( n984 , n70573 );
not ( n985 , n984 );
or ( n986 , n983 , n985 );
or ( n987 , n984 , n70673 );
nand ( n988 , n986 , n987 );
nand ( n989 , n982 , n988 );
nand ( n990 , n981 , n989 );
not ( n991 , n70491 );
not ( n992 , n991 );
and ( n993 , n520 , n992 );
not ( n71007 , n993 );
not ( n995 , n70515 );
or ( n996 , n71007 , n995 );
nand ( n997 , n992 , n520 );
not ( n998 , n997 );
not ( n999 , n70515 );
not ( n1000 , n999 );
or ( n1001 , n998 , n1000 );
nand ( n1002 , n1001 , n70525 );
nand ( n1003 , n996 , n1002 );
not ( n1007 , n1003 );
or ( n71018 , n70598 , n70579 );
nand ( n1009 , n71018 , n70621 );
nand ( n1010 , n70598 , n70579 );
nand ( n1011 , n1009 , n1010 );
not ( n1012 , n1011 );
nand ( n71023 , n1007 , n1012 );
not ( n1014 , n71023 );
not ( n1015 , n70575 );
not ( n1016 , n70360 );
or ( n1017 , n1015 , n1016 );
xor ( n1018 , n503 , n509 );
nand ( n1019 , n504 , n1018 );
nand ( n1020 , n1017 , n1019 );
not ( n1021 , n70596 );
and ( n1022 , n497 , n496 );
not ( n1023 , n497 );
not ( n1024 , n496 );
and ( n1025 , n1023 , n1024 );
nor ( n1026 , n1022 , n1025 );
not ( n1027 , n1026 );
nand ( n1028 , n1027 , n70534 );
not ( n1029 , n1028 );
not ( n1030 , n1029 );
or ( n71041 , n1021 , n1030 );
xor ( n1035 , n495 , n517 );
nand ( n1036 , n1035 , n1026 );
nand ( n71044 , n71041 , n1036 );
xor ( n1038 , n1020 , n71044 );
not ( n1039 , n516 );
xnor ( n1040 , n1039 , n497 );
not ( n1041 , n1040 );
not ( n1042 , n70640 );
or ( n71050 , n1041 , n1042 );
xor ( n1044 , n515 , n497 );
nand ( n1045 , n70513 , n1044 );
nand ( n1046 , n71050 , n1045 );
xor ( n1047 , n1038 , n1046 );
not ( n1048 , n1047 );
or ( n1049 , n1014 , n1048 );
nand ( n1050 , n1003 , n1011 );
nand ( n1051 , n1049 , n1050 );
xor ( n1052 , n1020 , n71044 );
and ( n1053 , n1052 , n1046 );
and ( n1054 , n1020 , n71044 );
or ( n1055 , n1053 , n1054 );
not ( n1056 , n1055 );
not ( n1057 , n728 );
not ( n1058 , n1057 );
not ( n1059 , n70523 );
or ( n1060 , n1058 , n1059 );
xor ( n1061 , n511 , n501 );
nand ( n1062 , n70371 , n1061 );
nand ( n1063 , n1060 , n1062 );
nand ( n1064 , n520 , n494 );
or ( n1065 , n520 , n494 );
nand ( n1066 , n1065 , n495 );
nand ( n1067 , n1064 , n493 , n1066 );
not ( n1068 , n1067 );
nand ( n1069 , n1063 , n1068 );
not ( n1070 , n1069 );
not ( n1071 , n1070 );
xor ( n1072 , n513 , n499 );
not ( n1073 , n1072 );
not ( n1074 , n699 );
or ( n1075 , n1073 , n1074 );
not ( n1076 , n512 );
not ( n1077 , n499 );
not ( n1078 , n1077 );
or ( n1079 , n1076 , n1078 );
nand ( n1080 , n70551 , n499 );
nand ( n1081 , n1079 , n1080 );
nand ( n1082 , n70655 , n1081 );
nand ( n1083 , n1075 , n1082 );
not ( n1084 , n1083 );
not ( n1085 , n1084 );
and ( n1086 , n1071 , n1085 );
and ( n71094 , n1070 , n1084 );
nor ( n1088 , n1086 , n71094 );
not ( n1089 , n1088 );
or ( n1090 , n1056 , n1089 );
or ( n1091 , n1088 , n1055 );
nand ( n1092 , n1090 , n1091 );
not ( n1093 , n1092 );
and ( n1094 , n1051 , n1093 );
not ( n1095 , n1051 );
and ( n1096 , n1095 , n1092 );
nor ( n1097 , n1094 , n1096 );
not ( n1098 , n503 );
nor ( n1099 , n1098 , n504 );
not ( n1100 , n1099 );
not ( n1101 , n1018 );
or ( n1102 , n1100 , n1101 );
xor ( n71110 , n503 , n508 );
nand ( n1104 , n71110 , n504 );
nand ( n1105 , n1102 , n1104 );
not ( n1106 , n1035 );
not ( n1107 , n70589 );
or ( n1108 , n1106 , n1107 );
not ( n1109 , n1027 );
xor ( n1110 , n495 , n516 );
nand ( n1111 , n1109 , n1110 );
nand ( n1112 , n1108 , n1111 );
xor ( n1113 , n1105 , n1112 );
xor ( n1114 , n519 , n493 );
not ( n1115 , n1114 );
xor ( n1116 , n494 , n495 );
xor ( n1117 , n493 , n494 );
not ( n1121 , n1117 );
nor ( n71126 , n1116 , n1121 );
not ( n1123 , n71126 );
or ( n1124 , n1115 , n1123 );
xor ( n1125 , n518 , n493 );
nand ( n1126 , n70491 , n1125 );
nand ( n1127 , n1124 , n1126 );
xor ( n1128 , n1113 , n1127 );
xor ( n1129 , n492 , n493 );
and ( n1130 , n1129 , n520 );
not ( n1131 , n1061 );
not ( n1132 , n70413 );
or ( n1133 , n1131 , n1132 );
xor ( n1134 , n510 , n501 );
nand ( n1135 , n70371 , n1134 );
nand ( n1136 , n1133 , n1135 );
xor ( n71141 , n1130 , n1136 );
not ( n1141 , n1044 );
not ( n1142 , n70509 );
or ( n1143 , n1141 , n1142 );
xor ( n1144 , n514 , n497 );
nand ( n1145 , n70513 , n1144 );
nand ( n1146 , n1143 , n1145 );
xor ( n1147 , n71141 , n1146 );
xor ( n1148 , n1128 , n1147 );
not ( n1149 , n70619 );
not ( n1150 , n70616 );
or ( n1151 , n1149 , n1150 );
nand ( n1152 , n70426 , n1072 );
nand ( n1153 , n1151 , n1152 );
xor ( n1154 , n520 , n493 );
not ( n1155 , n1154 );
not ( n1156 , n1116 );
and ( n1157 , n1156 , n1117 );
not ( n1158 , n1157 );
or ( n1159 , n1155 , n1158 );
nand ( n1160 , n70491 , n1114 );
nand ( n1161 , n1159 , n1160 );
or ( n1162 , n1153 , n1161 );
not ( n71164 , n1162 );
and ( n1164 , n1063 , n1067 );
not ( n1165 , n1063 );
and ( n1166 , n1165 , n1068 );
or ( n1167 , n1164 , n1166 );
not ( n1168 , n1167 );
or ( n1169 , n71164 , n1168 );
nand ( n1170 , n1153 , n1161 );
nand ( n1171 , n1169 , n1170 );
not ( n1172 , n1171 );
xor ( n71174 , n1148 , n1172 );
not ( n1174 , n71174 );
and ( n1175 , n1097 , n1174 );
not ( n1176 , n1097 );
and ( n1177 , n1176 , n71174 );
nor ( n1178 , n1175 , n1177 );
xor ( n1179 , n70490 , n70526 );
and ( n1180 , n1179 , n70572 );
and ( n1181 , n70490 , n70526 );
or ( n1182 , n1180 , n1181 );
not ( n1183 , n1182 );
xor ( n1184 , n1153 , n1161 );
not ( n1185 , n1167 );
xor ( n1186 , n1184 , n1185 );
and ( n1187 , n1003 , n1012 );
not ( n1188 , n1003 );
and ( n71190 , n1188 , n1011 );
nor ( n1190 , n1187 , n71190 );
and ( n1191 , n1190 , n1047 );
not ( n1192 , n1190 );
not ( n1193 , n1047 );
and ( n71195 , n1192 , n1193 );
nor ( n1195 , n1191 , n71195 );
nand ( n1196 , n1186 , n1195 );
not ( n1197 , n1196 );
or ( n1198 , n1183 , n1197 );
not ( n1199 , n1195 );
not ( n1200 , n1186 );
nand ( n1201 , n1199 , n1200 );
nand ( n1202 , n1198 , n1201 );
not ( n1203 , n1202 );
nand ( n1204 , n1178 , n1203 );
not ( n1205 , n70669 );
nand ( n1206 , n1205 , n70622 );
not ( n1207 , n1206 );
not ( n1211 , n70573 );
or ( n71210 , n1207 , n1211 );
not ( n1213 , n70622 );
nand ( n1214 , n1213 , n70669 );
nand ( n1215 , n71210 , n1214 );
not ( n1216 , n1215 );
and ( n1217 , n1195 , n1200 );
not ( n1218 , n1195 );
and ( n1219 , n1218 , n1186 );
nor ( n1220 , n1217 , n1219 );
xor ( n1221 , n1182 , n1220 );
nand ( n1222 , n1216 , n1221 );
and ( n1223 , n1204 , n1222 );
not ( n1224 , n1174 );
xnor ( n1225 , n1055 , n1088 );
not ( n1226 , n1225 );
or ( n1227 , n1224 , n1226 );
not ( n1228 , n1093 );
not ( n1229 , n71174 );
or ( n1230 , n1228 , n1229 );
nand ( n1231 , n1230 , n1051 );
nand ( n1232 , n1227 , n1231 );
not ( n1233 , n1232 );
not ( n1234 , n1055 );
nand ( n1235 , n1084 , n1069 );
not ( n1236 , n1235 );
or ( n1237 , n1234 , n1236 );
not ( n71236 , n1084 );
nand ( n1242 , n71236 , n1070 );
nand ( n1243 , n1237 , n1242 );
xor ( n1244 , n520 , n491 );
not ( n1245 , n1244 );
xnor ( n1246 , n491 , n492 );
xor ( n1247 , n492 , n493 );
nor ( n1248 , n1246 , n1247 );
not ( n1249 , n1248 );
or ( n71245 , n1245 , n1249 );
xor ( n1251 , n491 , n519 );
nand ( n1252 , n1129 , n1251 );
nand ( n1253 , n71245 , n1252 );
not ( n1254 , n1081 );
not ( n1255 , n70652 );
or ( n1256 , n1254 , n1255 );
not ( n1257 , n511 );
not ( n1258 , n499 );
not ( n1259 , n1258 );
or ( n71255 , n1257 , n1259 );
not ( n1261 , n511 );
nand ( n1262 , n1261 , n499 );
nand ( n1263 , n71255 , n1262 );
nand ( n1264 , n70704 , n1263 );
nand ( n1265 , n1256 , n1264 );
xor ( n1266 , n1253 , n1265 );
not ( n1267 , n1125 );
and ( n1268 , n1156 , n1117 );
not ( n1269 , n1268 );
or ( n1270 , n1267 , n1269 );
xor ( n1271 , n517 , n493 );
nand ( n1272 , n70491 , n1271 );
nand ( n1273 , n1270 , n1272 );
xor ( n1274 , n1266 , n1273 );
not ( n1275 , n1134 );
not ( n1276 , n1057 );
or ( n1277 , n1275 , n1276 );
and ( n1278 , n509 , n70432 );
not ( n1279 , n509 );
and ( n1280 , n1279 , n501 );
or ( n1281 , n1278 , n1280 );
nand ( n1282 , n70371 , n1281 );
nand ( n1283 , n1277 , n1282 );
not ( n1284 , n1144 );
not ( n1285 , n70565 );
or ( n1286 , n1284 , n1285 );
and ( n1287 , n513 , n497 );
not ( n1288 , n513 );
and ( n1289 , n1288 , n70495 );
nor ( n1290 , n1287 , n1289 );
nand ( n1291 , n70513 , n1290 );
nand ( n1292 , n1286 , n1291 );
xor ( n1293 , n1283 , n1292 );
not ( n1294 , n1110 );
not ( n1295 , n1029 );
or ( n1296 , n1294 , n1295 );
not ( n1297 , n1027 );
xor ( n1298 , n515 , n495 );
nand ( n1299 , n1297 , n1298 );
nand ( n1300 , n1296 , n1299 );
not ( n1301 , n1300 );
and ( n1302 , n1293 , n1301 );
not ( n1303 , n1293 );
and ( n71299 , n1303 , n1300 );
nor ( n1305 , n1302 , n71299 );
xor ( n1306 , n1274 , n1305 );
xor ( n1307 , n1243 , n1306 );
not ( n1308 , n1307 );
nand ( n1309 , n520 , n492 );
or ( n1310 , n520 , n492 );
nand ( n1311 , n1310 , n493 );
and ( n1312 , n1309 , n1311 , n491 );
not ( n1313 , n1312 );
not ( n1314 , n1099 );
not ( n1315 , n71110 );
or ( n1316 , n1314 , n1315 );
xor ( n1317 , n503 , n507 );
nand ( n1321 , n1317 , n504 );
nand ( n71314 , n1316 , n1321 );
not ( n1323 , n71314 );
or ( n1324 , n1313 , n1323 );
or ( n1325 , n1312 , n71314 );
nand ( n1326 , n1324 , n1325 );
not ( n1327 , n1105 );
not ( n1328 , n1112 );
or ( n1329 , n1327 , n1328 );
not ( n1330 , n1035 );
not ( n1331 , n70589 );
or ( n1332 , n1330 , n1331 );
nand ( n1333 , n1332 , n1111 );
or ( n1334 , n1105 , n1333 );
nand ( n1335 , n1334 , n1127 );
nand ( n1336 , n1329 , n1335 );
xor ( n1337 , n1326 , n1336 );
xor ( n1338 , n1130 , n1136 );
and ( n1339 , n1338 , n1146 );
and ( n1340 , n1130 , n1136 );
or ( n1341 , n1339 , n1340 );
xor ( n71334 , n1337 , n1341 );
not ( n1343 , n71334 );
not ( n1344 , n1343 );
not ( n1345 , n1128 );
not ( n1346 , n1345 );
not ( n1347 , n1346 );
not ( n1348 , n1147 );
or ( n1349 , n1347 , n1348 );
not ( n1350 , n1345 );
not ( n1351 , n1147 );
not ( n1352 , n1351 );
or ( n1353 , n1350 , n1352 );
nand ( n1354 , n1353 , n1171 );
nand ( n1355 , n1349 , n1354 );
not ( n1356 , n1355 );
not ( n1357 , n1356 );
or ( n1358 , n1344 , n1357 );
nand ( n1359 , n71334 , n1355 );
nand ( n1360 , n1358 , n1359 );
not ( n1361 , n1360 );
not ( n1362 , n1361 );
or ( n1363 , n1308 , n1362 );
not ( n1364 , n1307 );
nand ( n1365 , n1360 , n1364 );
nand ( n1366 , n1363 , n1365 );
nand ( n1367 , n1233 , n1366 );
not ( n71360 , n1263 );
xor ( n1372 , n500 , n499 );
and ( n1373 , n1372 , n70611 );
not ( n1374 , n1373 );
or ( n1375 , n71360 , n1374 );
not ( n1376 , n70704 );
not ( n1377 , n1376 );
and ( n71367 , n510 , n499 );
not ( n1379 , n510 );
not ( n1380 , n499 );
and ( n1381 , n1379 , n1380 );
nor ( n1382 , n71367 , n1381 );
nand ( n1383 , n1377 , n1382 );
nand ( n1384 , n1375 , n1383 );
not ( n1385 , n1290 );
not ( n1386 , n70565 );
or ( n1387 , n1385 , n1386 );
xor ( n1388 , n512 , n497 );
nand ( n1389 , n70513 , n1388 );
nand ( n1390 , n1387 , n1389 );
xor ( n1391 , n1384 , n1390 );
not ( n1392 , n1298 );
not ( n1393 , n70589 );
or ( n1394 , n1392 , n1393 );
xor ( n1395 , n514 , n495 );
nand ( n1396 , n70544 , n1395 );
nand ( n1397 , n1394 , n1396 );
xor ( n1398 , n1391 , n1397 );
not ( n1399 , n1251 );
not ( n1400 , n1248 );
or ( n1401 , n1399 , n1400 );
xor ( n1402 , n491 , n518 );
nand ( n1403 , n1129 , n1402 );
nand ( n1404 , n1401 , n1403 );
not ( n1405 , n1404 );
nand ( n1406 , n71314 , n1312 );
xor ( n1407 , n1405 , n1406 );
not ( n1408 , n1156 );
nand ( n71398 , n1271 , n1117 );
not ( n1410 , n71398 );
or ( n1411 , n1408 , n1410 );
xnor ( n1412 , n516 , n493 );
nand ( n1413 , n1412 , n1116 );
nand ( n1414 , n1411 , n1413 );
xor ( n1415 , n1407 , n1414 );
and ( n1416 , n1398 , n1415 );
not ( n1417 , n1398 );
not ( n1418 , n1415 );
and ( n1419 , n1417 , n1418 );
nor ( n1420 , n1416 , n1419 );
not ( n1421 , n1336 );
nand ( n1422 , n1421 , n1326 );
not ( n1423 , n1422 );
not ( n1424 , n1341 );
or ( n1425 , n1423 , n1424 );
not ( n1426 , n1326 );
nand ( n1427 , n1426 , n1336 );
nand ( n1428 , n1425 , n1427 );
xor ( n1429 , n1420 , n1428 );
not ( n1430 , n1265 );
not ( n1431 , n1273 );
or ( n1432 , n1430 , n1431 );
not ( n1433 , n1081 );
not ( n71423 , n70652 );
or ( n1435 , n1433 , n71423 );
nand ( n1436 , n70426 , n1263 );
nand ( n1437 , n1435 , n1436 );
or ( n1438 , n1273 , n1437 );
nand ( n1439 , n1438 , n1253 );
nand ( n1440 , n1432 , n1439 );
not ( n1441 , n1300 );
not ( n1442 , n1283 );
or ( n1443 , n1441 , n1442 );
or ( n71433 , n1283 , n1300 );
nand ( n1445 , n71433 , n1292 );
nand ( n1446 , n1443 , n1445 );
xor ( n1447 , n1440 , n1446 );
xor ( n1448 , n490 , n491 );
and ( n1449 , n1448 , n520 );
not ( n1450 , n1449 );
not ( n1451 , n1450 );
not ( n1452 , n1317 );
not ( n1453 , n70360 );
or ( n1454 , n1452 , n1453 );
and ( n1455 , n503 , n506 );
not ( n1456 , n503 );
not ( n1457 , n506 );
and ( n1458 , n1456 , n1457 );
nor ( n1459 , n1455 , n1458 );
nand ( n1460 , n1459 , n504 );
nand ( n1461 , n1454 , n1460 );
not ( n1462 , n1461 );
or ( n1463 , n1451 , n1462 );
not ( n1467 , n1461 );
nand ( n71454 , n1467 , n1449 );
nand ( n1469 , n1463 , n71454 );
xor ( n1470 , n508 , n501 );
nand ( n1471 , n1470 , n70371 );
nand ( n1472 , n70413 , n1281 );
nand ( n1473 , n1471 , n1472 );
xor ( n1474 , n1469 , n1473 );
xor ( n1475 , n1447 , n1474 );
or ( n1476 , n1429 , n1475 );
nand ( n1477 , n1429 , n1475 );
nand ( n1478 , n1476 , n1477 );
buf ( n1479 , n1305 );
not ( n1480 , n1274 );
nand ( n1481 , n1479 , n1480 );
not ( n1482 , n1481 );
not ( n1483 , n1243 );
or ( n1484 , n1482 , n1483 );
or ( n1485 , n1479 , n1480 );
nand ( n1486 , n1484 , n1485 );
not ( n1487 , n1486 );
and ( n1488 , n1478 , n1487 );
not ( n1489 , n1478 );
and ( n1490 , n1489 , n1486 );
nor ( n1491 , n1488 , n1490 );
not ( n1492 , n1364 );
not ( n1493 , n1343 );
or ( n71480 , n1492 , n1493 );
not ( n1498 , n71334 );
not ( n1499 , n1307 );
or ( n1500 , n1498 , n1499 );
nand ( n1501 , n1500 , n1355 );
nand ( n1502 , n71480 , n1501 );
not ( n1503 , n1502 );
nand ( n1504 , n1491 , n1503 );
nand ( n1505 , n990 , n1223 , n1367 , n1504 );
not ( n1506 , n1204 );
nor ( n1507 , n1216 , n1221 );
not ( n71491 , n1507 );
or ( n1509 , n1506 , n71491 );
not ( n1510 , n1178 );
nand ( n1511 , n1510 , n1202 );
nand ( n1512 , n1509 , n1511 );
nand ( n1513 , n1512 , n1367 , n1504 );
not ( n1514 , n1503 );
not ( n1515 , n1491 );
or ( n1516 , n1514 , n1515 );
not ( n1517 , n1232 );
nor ( n1518 , n1366 , n1517 );
nand ( n1519 , n1516 , n1518 );
not ( n1520 , n1491 );
nand ( n1521 , n1520 , n1502 );
nand ( n1522 , n1505 , n1513 , n1519 , n1521 );
xor ( n1523 , n1384 , n1390 );
and ( n1524 , n1523 , n1397 );
and ( n1525 , n1384 , n1390 );
or ( n1526 , n1524 , n1525 );
not ( n1527 , n1388 );
not ( n1528 , n70509 );
or ( n1529 , n1527 , n1528 );
xor ( n1530 , n511 , n497 );
nand ( n1531 , n70513 , n1530 );
nand ( n1532 , n1529 , n1531 );
not ( n1533 , n1532 );
not ( n1534 , n1470 );
not ( n1535 , n1057 );
or ( n1536 , n1534 , n1535 );
and ( n1537 , n507 , n501 );
not ( n1538 , n507 );
not ( n71522 , n501 );
and ( n1540 , n1538 , n71522 );
nor ( n1541 , n1537 , n1540 );
nand ( n1542 , n70371 , n1541 );
nand ( n1543 , n1536 , n1542 );
not ( n1544 , n1543 );
not ( n1545 , n1544 );
or ( n1546 , n1533 , n1545 );
not ( n1547 , n1532 );
nand ( n1548 , n1543 , n1547 );
nand ( n1549 , n1546 , n1548 );
xor ( n1550 , n489 , n490 );
xor ( n1551 , n520 , n489 );
nand ( n1552 , n1550 , n1551 );
buf ( n1553 , n1448 );
or ( n1554 , n1552 , n1553 );
xor ( n1555 , n519 , n489 );
nand ( n1556 , n1553 , n1555 );
nand ( n1557 , n1554 , n1556 );
not ( n1558 , n1557 );
not ( n1559 , n1558 );
and ( n1560 , n1549 , n1559 );
not ( n1561 , n1549 );
and ( n1562 , n1561 , n1558 );
nor ( n1563 , n1560 , n1562 );
xor ( n1564 , n1526 , n1563 );
and ( n1565 , n493 , n1039 );
not ( n1566 , n493 );
and ( n1567 , n1566 , n516 );
nor ( n1568 , n1565 , n1567 );
nor ( n1569 , n1121 , n1568 );
not ( n71553 , n1569 );
not ( n1571 , n1156 );
or ( n1572 , n71553 , n1571 );
xor ( n1573 , n515 , n493 );
nand ( n1574 , n70491 , n1573 );
nand ( n1575 , n1572 , n1574 );
not ( n1576 , n1395 );
not ( n1577 , n1029 );
or ( n1578 , n1576 , n1577 );
xor ( n1579 , n513 , n495 );
and ( n1580 , n496 , n497 );
not ( n1581 , n496 );
and ( n1582 , n1581 , n70530 );
nor ( n1583 , n1580 , n1582 );
nand ( n71567 , n1579 , n1583 );
nand ( n1585 , n1578 , n71567 );
xor ( n1586 , n1575 , n1585 );
not ( n1587 , n1382 );
not ( n1588 , n699 );
or ( n1589 , n1587 , n1588 );
and ( n1590 , n509 , n499 );
not ( n1591 , n509 );
and ( n1592 , n1591 , n1380 );
nor ( n1593 , n1590 , n1592 );
nand ( n1594 , n70655 , n1593 );
nand ( n1595 , n1589 , n1594 );
xor ( n1596 , n1586 , n1595 );
xor ( n1597 , n1564 , n1596 );
not ( n1598 , n1341 );
not ( n1599 , n1422 );
or ( n1600 , n1598 , n1599 );
nand ( n1601 , n1600 , n1427 );
or ( n1602 , n1418 , n1601 );
buf ( n1603 , n1398 );
nand ( n1604 , n1602 , n1603 );
nand ( n1605 , n1601 , n1418 );
nand ( n1606 , n1604 , n1605 );
not ( n1607 , n1606 );
and ( n1608 , n1597 , n1607 );
not ( n1609 , n1597 );
and ( n1610 , n1609 , n1606 );
nor ( n1611 , n1608 , n1610 );
xor ( n1612 , n1405 , n1406 );
and ( n1616 , n1612 , n1414 );
and ( n71597 , n1405 , n1406 );
or ( n1618 , n1616 , n71597 );
nand ( n1619 , n1467 , n1450 );
not ( n1620 , n1619 );
not ( n1621 , n1473 );
or ( n1622 , n1620 , n1621 );
nand ( n1623 , n1449 , n1461 );
nand ( n1624 , n1622 , n1623 );
not ( n1625 , n1402 );
xnor ( n1626 , n491 , n492 );
nor ( n1627 , n1626 , n1247 );
not ( n1628 , n1627 );
or ( n1629 , n1625 , n1628 );
buf ( n1630 , n1129 );
xor ( n1631 , n517 , n491 );
nand ( n1632 , n1630 , n1631 );
nand ( n1633 , n1629 , n1632 );
not ( n1634 , n1633 );
not ( n1635 , n1459 );
not ( n1636 , n504 );
and ( n1637 , n1636 , n503 );
not ( n1638 , n1637 );
or ( n1639 , n1635 , n1638 );
xor ( n1640 , n503 , n505 );
nand ( n71621 , n1640 , n504 );
nand ( n1645 , n1639 , n71621 );
or ( n1646 , n520 , n490 );
nand ( n1647 , n1646 , n491 );
and ( n1648 , n520 , n490 );
not ( n1649 , n489 );
nor ( n1650 , n1648 , n1649 );
and ( n1651 , n1647 , n1650 );
nor ( n1652 , n1645 , n1651 );
not ( n1653 , n1652 );
nand ( n1654 , n1651 , n1645 );
nand ( n1655 , n1653 , n1654 );
or ( n1656 , n1634 , n1655 );
nand ( n1657 , n1655 , n1634 );
nand ( n1658 , n1656 , n1657 );
xor ( n1659 , n1624 , n1658 );
xor ( n1660 , n1618 , n1659 );
xor ( n1661 , n1440 , n1446 );
and ( n1662 , n1661 , n1474 );
and ( n1663 , n1440 , n1446 );
or ( n1664 , n1662 , n1663 );
xnor ( n1665 , n1660 , n1664 );
and ( n1666 , n1611 , n1665 );
not ( n1667 , n1611 );
not ( n1668 , n1665 );
and ( n1669 , n1667 , n1668 );
nor ( n1670 , n1666 , n1669 );
not ( n71648 , n1475 );
not ( n1672 , n1486 );
or ( n1673 , n71648 , n1672 );
or ( n1674 , n1486 , n1475 );
not ( n1675 , n1429 );
nand ( n1676 , n1674 , n1675 );
nand ( n1677 , n1673 , n1676 );
nand ( n1678 , n1670 , n1677 );
buf ( n1679 , n1678 );
not ( n1680 , n1677 );
not ( n1681 , n1670 );
nand ( n1682 , n1680 , n1681 );
nand ( n1683 , n1679 , n1682 );
xnor ( n1684 , n1522 , n1683 );
nand ( n1685 , n1684 , n70470 );
and ( n1686 , n492 , n493 );
not ( n1687 , n492 );
not ( n1688 , n493 );
and ( n1689 , n1687 , n1688 );
nor ( n1690 , n1686 , n1689 );
not ( n1691 , n1690 );
not ( n1692 , n492 );
not ( n1693 , n491 );
not ( n1694 , n1693 );
or ( n1695 , n1692 , n1694 );
not ( n71673 , n492 );
nand ( n1697 , n71673 , n491 );
nand ( n1698 , n1695 , n1697 );
nand ( n1699 , n1691 , n1698 );
not ( n1700 , n1699 );
not ( n1701 , n1700 );
not ( n1702 , n491 );
and ( n1703 , n456 , n464 );
not ( n1704 , n456 );
and ( n1705 , n1704 , n480 );
nor ( n1706 , n1703 , n1705 );
not ( n1707 , n1706 );
or ( n1708 , n1702 , n1707 );
not ( n1709 , n464 );
and ( n1710 , n456 , n1709 );
not ( n1711 , n456 );
not ( n1712 , n480 );
and ( n71690 , n1711 , n1712 );
nor ( n1714 , n1710 , n71690 );
not ( n1715 , n491 );
nand ( n1716 , n1714 , n1715 );
nand ( n1717 , n1708 , n1716 );
not ( n1718 , n1717 );
or ( n1719 , n1701 , n1718 );
not ( n1720 , n1715 );
not ( n1721 , n479 );
not ( n71699 , n456 );
not ( n1723 , n71699 );
or ( n1724 , n1721 , n1723 );
nand ( n1725 , n456 , n463 );
nand ( n1726 , n1724 , n1725 );
not ( n1730 , n1726 );
or ( n71705 , n1720 , n1730 );
and ( n1732 , n456 , n463 );
not ( n1733 , n456 );
and ( n1734 , n1733 , n479 );
nor ( n1735 , n1732 , n1734 );
nand ( n1736 , n1735 , n491 );
nand ( n1737 , n71705 , n1736 );
not ( n1738 , n1690 );
not ( n1739 , n1738 );
nand ( n1740 , n1737 , n1739 );
nand ( n1741 , n1719 , n1740 );
not ( n1742 , n495 );
and ( n1743 , n456 , n460 );
not ( n1744 , n456 );
and ( n1745 , n1744 , n476 );
nor ( n1746 , n1743 , n1745 );
not ( n1747 , n1746 );
or ( n1748 , n1742 , n1747 );
not ( n1749 , n495 );
and ( n1750 , n456 , n460 );
not ( n1751 , n456 );
and ( n1752 , n1751 , n476 );
nor ( n1753 , n1750 , n1752 );
not ( n1754 , n1753 );
nand ( n1755 , n1749 , n1754 );
nand ( n1756 , n1748 , n1755 );
not ( n1757 , n1756 );
not ( n1758 , n495 );
nand ( n1759 , n1758 , n497 , n496 );
not ( n1760 , n497 );
nand ( n1761 , n70584 , n1760 , n495 );
nand ( n1762 , n1759 , n1761 );
buf ( n1763 , n1762 );
not ( n1764 , n1763 );
or ( n1765 , n1757 , n1764 );
and ( n1766 , n456 , n459 );
not ( n1767 , n456 );
and ( n1768 , n1767 , n475 );
nor ( n1769 , n1766 , n1768 );
buf ( n1770 , n1769 );
and ( n1771 , n495 , n1770 );
not ( n1772 , n495 );
not ( n1773 , n459 );
and ( n1774 , n456 , n1773 );
not ( n1775 , n456 );
not ( n1776 , n475 );
and ( n1777 , n1775 , n1776 );
nor ( n1778 , n1774 , n1777 );
and ( n1779 , n1772 , n1778 );
or ( n71754 , n1771 , n1779 );
xor ( n1784 , n497 , n496 );
nand ( n1785 , n71754 , n1784 );
nand ( n1786 , n1765 , n1785 );
xor ( n1787 , n1741 , n1786 );
xor ( n1788 , n491 , n490 );
not ( n1789 , n1788 );
not ( n71761 , n1789 );
not ( n1791 , n71761 );
and ( n1792 , n456 , n465 );
not ( n1793 , n456 );
and ( n1794 , n1793 , n481 );
nor ( n1795 , n1792 , n1794 );
not ( n71767 , n1795 );
not ( n1797 , n71767 );
not ( n1798 , n1649 );
or ( n1799 , n1797 , n1798 );
not ( n1800 , n465 );
nand ( n1801 , n1800 , n456 );
not ( n1802 , n1801 );
or ( n1803 , n456 , n481 );
not ( n1804 , n1803 );
or ( n1805 , n1802 , n1804 );
nand ( n1806 , n1805 , n489 );
nand ( n1807 , n1799 , n1806 );
not ( n1808 , n1807 );
or ( n1809 , n1791 , n1808 );
not ( n1810 , n1649 );
and ( n1811 , n456 , n466 );
not ( n1812 , n456 );
and ( n1813 , n1812 , n482 );
nor ( n1814 , n1811 , n1813 );
not ( n1815 , n1814 );
not ( n1816 , n1815 );
or ( n1817 , n1810 , n1816 );
or ( n1818 , n1815 , n1649 );
nand ( n1819 , n1817 , n1818 );
not ( n1820 , n489 );
nor ( n1821 , n490 , n491 );
not ( n1822 , n1821 );
or ( n1823 , n1820 , n1822 );
not ( n1824 , n489 );
nand ( n1825 , n1824 , n491 , n490 );
nand ( n1826 , n1823 , n1825 );
not ( n1827 , n1826 );
not ( n1828 , n1827 );
nand ( n1829 , n1819 , n1828 );
nand ( n1830 , n1809 , n1829 );
and ( n1831 , n1787 , n1830 );
and ( n1832 , n1741 , n1786 );
or ( n1833 , n1831 , n1832 );
xor ( n1834 , n500 , n501 );
not ( n1835 , n499 );
nor ( n1836 , n500 , n501 );
not ( n1837 , n1836 );
or ( n1838 , n1835 , n1837 );
nand ( n1839 , n1258 , n501 , n500 );
nand ( n1840 , n1838 , n1839 );
or ( n1841 , n1834 , n1840 );
nand ( n1842 , n1841 , n499 );
not ( n1843 , n498 );
not ( n1844 , n1077 );
or ( n1845 , n1843 , n1844 );
nand ( n1846 , n70502 , n499 );
nand ( n1847 , n1845 , n1846 );
buf ( n1848 , n1847 );
not ( n1849 , n1848 );
and ( n1850 , n456 , n457 );
not ( n1851 , n456 );
and ( n1852 , n1851 , n473 );
nor ( n1853 , n1850 , n1852 );
not ( n1854 , n1853 );
not ( n1855 , n1854 );
and ( n1856 , n497 , n1855 );
not ( n1857 , n497 );
not ( n1858 , n1855 );
and ( n1859 , n1857 , n1858 );
or ( n1860 , n1856 , n1859 );
not ( n1861 , n1860 );
or ( n1862 , n1849 , n1861 );
not ( n1863 , n498 );
not ( n1864 , n499 );
nand ( n1865 , n1863 , n1864 , n497 );
not ( n71837 , n497 );
nand ( n1867 , n71837 , n498 , n499 );
nand ( n1868 , n1865 , n1867 );
buf ( n1869 , n1868 );
buf ( n1870 , n1869 );
and ( n1871 , n456 , n458 );
not ( n1872 , n456 );
and ( n1873 , n1872 , n474 );
nor ( n1874 , n1871 , n1873 );
and ( n1875 , n497 , n1874 );
not ( n1876 , n497 );
and ( n1877 , n456 , n458 );
not ( n1878 , n456 );
and ( n1879 , n1878 , n474 );
nor ( n1880 , n1877 , n1879 );
not ( n1881 , n1880 );
and ( n1882 , n1876 , n1881 );
or ( n1883 , n1875 , n1882 );
nand ( n1884 , n1870 , n1883 );
nand ( n1885 , n1862 , n1884 );
xor ( n1886 , n1842 , n1885 );
and ( n1887 , n70594 , n494 );
not ( n1888 , n494 );
and ( n1889 , n1888 , n495 );
nor ( n71861 , n1887 , n1889 );
not ( n1891 , n71861 );
not ( n1892 , n1891 );
and ( n1893 , n456 , n461 );
not ( n1894 , n456 );
and ( n1895 , n1894 , n477 );
nor ( n1896 , n1893 , n1895 );
and ( n1897 , n493 , n1896 );
not ( n1898 , n493 );
not ( n1899 , n1896 );
and ( n1900 , n1898 , n1899 );
or ( n1901 , n1897 , n1900 );
not ( n1902 , n1901 );
or ( n1903 , n1892 , n1902 );
nor ( n1904 , n494 , n495 );
nand ( n1905 , n1904 , n493 );
not ( n1906 , n493 );
nand ( n1907 , n1906 , n495 , n494 );
nand ( n1908 , n1905 , n1907 );
buf ( n1909 , n1908 );
not ( n1910 , n493 );
and ( n1911 , n456 , n462 );
not ( n1912 , n456 );
and ( n1913 , n1912 , n478 );
nor ( n1917 , n1911 , n1913 );
not ( n71886 , n1917 );
or ( n1919 , n1910 , n71886 );
or ( n1920 , n1917 , n493 );
nand ( n1921 , n1919 , n1920 );
nand ( n1922 , n1909 , n1921 );
nand ( n1923 , n1903 , n1922 );
and ( n1924 , n1886 , n1923 );
and ( n1925 , n1842 , n1885 );
or ( n1926 , n1924 , n1925 );
xor ( n1927 , n1833 , n1926 );
xor ( n1928 , n493 , n492 );
not ( n1929 , n1928 );
not ( n1930 , n491 );
not ( n1931 , n1917 );
or ( n1932 , n1930 , n1931 );
not ( n1933 , n462 );
and ( n1934 , n1933 , n456 );
nor ( n1935 , n456 , n478 );
nor ( n1936 , n1934 , n1935 );
nand ( n1937 , n1936 , n1715 );
nand ( n1938 , n1932 , n1937 );
not ( n1939 , n1938 );
or ( n1940 , n1929 , n1939 );
and ( n1941 , n1738 , n1698 );
nand ( n1942 , n1737 , n1941 );
nand ( n1943 , n1940 , n1942 );
not ( n1944 , n1807 );
not ( n1945 , n1828 );
or ( n1946 , n1944 , n1945 );
not ( n1947 , n489 );
not ( n1948 , n1706 );
or ( n1949 , n1947 , n1948 );
nand ( n71918 , n1714 , n1649 );
nand ( n1954 , n1949 , n71918 );
buf ( n1955 , n1788 );
nand ( n1956 , n1954 , n1955 );
nand ( n1957 , n1946 , n1956 );
xor ( n1958 , n1943 , n1957 );
not ( n1959 , n1870 );
not ( n1960 , n1860 );
or ( n1961 , n1959 , n1960 );
buf ( n1962 , n1848 );
nand ( n1963 , n1962 , n497 );
nand ( n1964 , n1961 , n1963 );
xor ( n1965 , n1958 , n1964 );
xor ( n1966 , n1927 , n1965 );
and ( n1967 , n456 , n466 );
not ( n1968 , n456 );
and ( n71934 , n1968 , n482 );
nor ( n1970 , n1967 , n71934 );
not ( n1971 , n1970 );
and ( n1972 , n1971 , n489 );
not ( n1973 , n1909 );
not ( n1974 , n1901 );
or ( n1975 , n1973 , n1974 );
not ( n1976 , n493 );
not ( n1977 , n1976 );
and ( n1978 , n456 , n460 );
not ( n71944 , n456 );
and ( n1980 , n71944 , n476 );
nor ( n1981 , n1978 , n1980 );
not ( n1982 , n1981 );
not ( n1983 , n1982 );
or ( n1984 , n1977 , n1983 );
or ( n1985 , n1982 , n1976 );
nand ( n1986 , n1984 , n1985 );
nand ( n1987 , n1986 , n1891 );
nand ( n1988 , n1975 , n1987 );
xor ( n1989 , n1972 , n1988 );
not ( n1990 , n1763 );
not ( n1991 , n71754 );
or ( n1992 , n1990 , n1991 );
and ( n1993 , n495 , n1874 );
not ( n1994 , n495 );
not ( n1995 , n1874 );
and ( n1996 , n1994 , n1995 );
or ( n1997 , n1993 , n1996 );
nand ( n1998 , n1997 , n1784 );
nand ( n1999 , n1992 , n1998 );
not ( n2000 , n1999 );
xor ( n2001 , n1989 , n2000 );
and ( n2002 , n456 , n467 );
not ( n2003 , n456 );
and ( n2004 , n2003 , n483 );
nor ( n2005 , n2002 , n2004 );
not ( n2006 , n2005 );
and ( n2007 , n2006 , n489 );
buf ( n2008 , n1840 );
not ( n2009 , n473 );
nor ( n2010 , n2009 , n456 );
not ( n2011 , n2010 );
nand ( n2012 , n456 , n457 );
nand ( n2013 , n2011 , n2012 );
or ( n2014 , n2013 , n70613 );
nand ( n2015 , n1854 , n70613 );
nand ( n2016 , n2014 , n2015 );
and ( n2017 , n2008 , n2016 );
xor ( n2018 , n500 , n501 );
and ( n2019 , n2018 , n499 );
nor ( n2020 , n2017 , n2019 );
not ( n2021 , n2020 );
xor ( n2022 , n2007 , n2021 );
not ( n2023 , n1869 );
and ( n2024 , n456 , n459 );
not ( n2025 , n456 );
and ( n2026 , n2025 , n475 );
or ( n2027 , n2024 , n2026 );
not ( n2028 , n2027 );
not ( n2029 , n1760 );
or ( n2030 , n2028 , n2029 );
nand ( n2031 , n497 , n1769 );
nand ( n71997 , n2030 , n2031 );
not ( n2033 , n71997 );
or ( n2034 , n2023 , n2033 );
nand ( n2035 , n1883 , n1848 );
nand ( n2036 , n2034 , n2035 );
nand ( n2037 , n1888 , n495 );
nand ( n2038 , n70594 , n494 );
nand ( n2039 , n2037 , n2038 );
not ( n2040 , n2039 );
not ( n2041 , n1921 );
or ( n2042 , n2040 , n2041 );
not ( n2043 , n1726 );
not ( n2044 , n1976 );
or ( n2045 , n2043 , n2044 );
nand ( n2046 , n1735 , n493 );
nand ( n2047 , n2045 , n2046 );
nand ( n2048 , n2047 , n1908 );
nand ( n2049 , n2042 , n2048 );
xor ( n2050 , n2036 , n2049 );
not ( n2051 , n1928 );
not ( n2052 , n1717 );
or ( n2053 , n2051 , n2052 );
not ( n2054 , n491 );
and ( n2055 , n456 , n465 );
not ( n2056 , n456 );
and ( n2057 , n2056 , n481 );
nor ( n2058 , n2055 , n2057 );
not ( n2059 , n2058 );
or ( n2060 , n2054 , n2059 );
and ( n2061 , n456 , n465 );
not ( n2062 , n456 );
and ( n2063 , n2062 , n481 );
nor ( n2064 , n2061 , n2063 );
not ( n2065 , n2064 );
nand ( n2066 , n2065 , n1715 );
nand ( n2067 , n2060 , n2066 );
nand ( n2068 , n2067 , n1700 );
nand ( n2069 , n2053 , n2068 );
and ( n2070 , n2050 , n2069 );
and ( n2071 , n2036 , n2049 );
or ( n2072 , n2070 , n2071 );
and ( n2073 , n2022 , n2072 );
and ( n2074 , n2007 , n2021 );
or ( n2075 , n2073 , n2074 );
xor ( n2076 , n2001 , n2075 );
not ( n2077 , n1763 );
and ( n2081 , n495 , n1896 );
not ( n72044 , n495 );
not ( n2083 , n461 );
not ( n2084 , n456 );
or ( n2085 , n2083 , n2084 );
not ( n2086 , n456 );
nand ( n72049 , n2086 , n477 );
nand ( n2088 , n2085 , n72049 );
and ( n2089 , n72044 , n2088 );
or ( n2090 , n2081 , n2089 );
not ( n2091 , n2090 );
or ( n2092 , n2077 , n2091 );
nand ( n2093 , n1756 , n1784 );
nand ( n2094 , n2092 , n2093 );
not ( n2095 , n1826 );
not ( n2096 , n1649 );
not ( n2097 , n467 );
and ( n2098 , n456 , n2097 );
not ( n2099 , n456 );
not ( n2100 , n483 );
and ( n2101 , n2099 , n2100 );
nor ( n2102 , n2098 , n2101 );
not ( n2103 , n2102 );
or ( n2104 , n2096 , n2103 );
nand ( n2105 , n2005 , n489 );
nand ( n2106 , n2104 , n2105 );
not ( n2107 , n2106 );
or ( n2108 , n2095 , n2107 );
nand ( n2109 , n1819 , n1788 );
nand ( n2110 , n2108 , n2109 );
xor ( n2111 , n2094 , n2110 );
and ( n72074 , n456 , n468 );
not ( n2116 , n456 );
and ( n2117 , n2116 , n484 );
nor ( n2118 , n72074 , n2117 );
not ( n2119 , n2118 );
and ( n2120 , n489 , n2119 );
and ( n2121 , n2111 , n2120 );
and ( n2122 , n2094 , n2110 );
or ( n2123 , n2121 , n2122 );
xor ( n2124 , n1741 , n1786 );
xor ( n2125 , n2124 , n1830 );
xor ( n2126 , n2123 , n2125 );
xor ( n2127 , n1842 , n1885 );
xor ( n2128 , n2127 , n1923 );
and ( n2129 , n2126 , n2128 );
and ( n2130 , n2123 , n2125 );
or ( n2131 , n2129 , n2130 );
xor ( n2132 , n2076 , n2131 );
xor ( n2133 , n1966 , n2132 );
xor ( n72093 , n2007 , n2021 );
xor ( n2135 , n72093 , n2072 );
not ( n2136 , n502 );
not ( n2137 , n503 );
not ( n2138 , n2137 );
or ( n2139 , n2136 , n2138 );
not ( n2140 , n502 );
nand ( n2141 , n2140 , n503 );
nand ( n2142 , n2139 , n2141 );
not ( n2143 , n2142 );
not ( n2144 , n2143 );
not ( n2145 , n501 );
nand ( n2146 , n2145 , n503 , n502 );
not ( n2147 , n502 );
not ( n2148 , n503 );
nand ( n2149 , n2147 , n2148 , n501 );
and ( n2150 , n2146 , n2149 );
not ( n2151 , n2150 );
or ( n2152 , n2144 , n2151 );
nand ( n2153 , n2152 , n501 );
not ( n2154 , n1834 );
not ( n2155 , n2016 );
or ( n2156 , n2154 , n2155 );
not ( n2157 , n499 );
not ( n2158 , n1874 );
or ( n2159 , n2157 , n2158 );
not ( n2160 , n499 );
nand ( n2161 , n2160 , n1881 );
nand ( n2162 , n2159 , n2161 );
not ( n2163 , n499 );
nor ( n2164 , n500 , n501 );
not ( n2165 , n2164 );
or ( n2166 , n2163 , n2165 );
nand ( n2167 , n2166 , n1839 );
nand ( n2168 , n2162 , n2167 );
nand ( n2169 , n2156 , n2168 );
xor ( n2170 , n2153 , n2169 );
not ( n2171 , n1763 );
not ( n2172 , n495 );
and ( n2173 , n456 , n462 );
not ( n72133 , n456 );
and ( n2175 , n72133 , n478 );
nor ( n2176 , n2173 , n2175 );
not ( n2177 , n2176 );
or ( n2178 , n2172 , n2177 );
or ( n2179 , n2176 , n495 );
nand ( n2180 , n2178 , n2179 );
not ( n2181 , n2180 );
or ( n2182 , n2171 , n2181 );
nand ( n2183 , n2090 , n1784 );
nand ( n2184 , n2182 , n2183 );
and ( n2185 , n2170 , n2184 );
and ( n2186 , n2153 , n2169 );
or ( n2187 , n2185 , n2186 );
xor ( n2188 , n2020 , n2187 );
and ( n2189 , n456 , n469 );
not ( n2190 , n456 );
and ( n2191 , n2190 , n485 );
nor ( n2192 , n2189 , n2191 );
nor ( n2193 , n2192 , n1824 );
not ( n2194 , n2039 );
not ( n2195 , n2047 );
or ( n2196 , n2194 , n2195 );
or ( n2197 , n1712 , n456 );
nand ( n2198 , n456 , n464 );
nand ( n2199 , n2197 , n2198 );
and ( n2200 , n493 , n2199 );
not ( n2201 , n493 );
not ( n2202 , n456 );
and ( n2203 , n2202 , n480 );
not ( n2204 , n2202 );
and ( n2205 , n2204 , n464 );
nor ( n2206 , n2203 , n2205 );
and ( n2207 , n2201 , n2206 );
nor ( n72167 , n2200 , n2207 );
nand ( n2209 , n1908 , n72167 );
nand ( n2210 , n2196 , n2209 );
xor ( n2211 , n2193 , n2210 );
not ( n2212 , n1869 );
not ( n2213 , n497 );
not ( n2217 , n2213 );
not ( n72174 , n1754 );
or ( n2219 , n2217 , n72174 );
or ( n2220 , n1754 , n2213 );
nand ( n2221 , n2219 , n2220 );
not ( n2222 , n2221 );
or ( n2223 , n2212 , n2222 );
nand ( n2224 , n71997 , n1848 );
nand ( n2225 , n2223 , n2224 );
and ( n2226 , n2211 , n2225 );
and ( n2227 , n2193 , n2210 );
or ( n2228 , n2226 , n2227 );
and ( n2229 , n2188 , n2228 );
and ( n2230 , n2020 , n2187 );
or ( n2231 , n2229 , n2230 );
xor ( n2232 , n2135 , n2231 );
xor ( n2233 , n2094 , n2110 );
xor ( n2234 , n2233 , n2120 );
xor ( n2235 , n2036 , n2049 );
xor ( n2236 , n2235 , n2069 );
xor ( n2237 , n2234 , n2236 );
not ( n2238 , n1928 );
not ( n2239 , n2067 );
or ( n2240 , n2238 , n2239 );
and ( n2241 , n493 , n1693 , n492 );
and ( n2242 , n1971 , n2241 );
not ( n72199 , n1971 );
not ( n2244 , n492 );
nand ( n2245 , n2244 , n1688 , n491 );
not ( n2246 , n2245 );
and ( n2247 , n72199 , n2246 );
nor ( n2248 , n2242 , n2247 );
nand ( n2249 , n2240 , n2248 );
not ( n2250 , n71761 );
not ( n2251 , n2106 );
or ( n2252 , n2250 , n2251 );
xor ( n2253 , n489 , n2119 );
nand ( n2254 , n2253 , n1826 );
nand ( n2255 , n2252 , n2254 );
xor ( n2256 , n2249 , n2255 );
nand ( n2257 , n2147 , n2148 , n501 );
nand ( n2258 , n2145 , n503 , n502 );
nand ( n2259 , n2257 , n2258 );
not ( n2260 , n2259 );
not ( n2261 , n501 );
nand ( n2262 , n1854 , n2261 );
nand ( n2263 , n1855 , n501 );
nand ( n2264 , n2262 , n2263 );
not ( n2265 , n2264 );
or ( n2266 , n2260 , n2265 );
and ( n2267 , n502 , n503 );
not ( n2268 , n502 );
not ( n2269 , n503 );
and ( n2270 , n2268 , n2269 );
nor ( n2271 , n2267 , n2270 );
buf ( n2272 , n2271 );
nand ( n2273 , n2272 , n501 );
nand ( n2274 , n2266 , n2273 );
and ( n2275 , n2256 , n2274 );
and ( n2276 , n2249 , n2255 );
or ( n2277 , n2275 , n2276 );
and ( n2278 , n2237 , n2277 );
and ( n2279 , n2234 , n2236 );
or ( n2280 , n2278 , n2279 );
and ( n2281 , n2232 , n2280 );
and ( n2282 , n2135 , n2231 );
or ( n2283 , n2281 , n2282 );
xor ( n2284 , n2133 , n2283 );
xor ( n2285 , n2123 , n2125 );
xor ( n2286 , n2285 , n2128 );
xor ( n2287 , n2135 , n2231 );
xor ( n2288 , n2287 , n2280 );
xor ( n2289 , n2286 , n2288 );
xor ( n2290 , n2020 , n2187 );
xor ( n2291 , n2290 , n2228 );
not ( n2292 , n2039 );
not ( n2293 , n72167 );
or ( n2294 , n2292 , n2293 );
not ( n2295 , n2064 );
not ( n2296 , n493 );
nand ( n2297 , n2296 , n495 , n494 );
not ( n2298 , n2297 );
and ( n2299 , n2295 , n2298 );
not ( n2300 , n1905 );
and ( n72257 , n2300 , n2058 );
nor ( n2305 , n2299 , n72257 );
nand ( n2306 , n2294 , n2305 );
not ( n2307 , n1869 );
not ( n2308 , n70505 );
not ( n2309 , n2088 );
or ( n2310 , n2308 , n2309 );
nand ( n2311 , n456 , n461 );
nand ( n2312 , n2086 , n477 );
nand ( n2313 , n2311 , n2312 , n497 );
nand ( n2314 , n2310 , n2313 );
not ( n2315 , n2314 );
or ( n2316 , n2307 , n2315 );
nand ( n2317 , n2221 , n1848 );
nand ( n2318 , n2316 , n2317 );
xor ( n2319 , n2306 , n2318 );
not ( n2320 , n1700 );
not ( n2321 , n1715 );
not ( n2322 , n2006 );
or ( n2323 , n2321 , n2322 );
or ( n2324 , n2006 , n1715 );
nand ( n2325 , n2323 , n2324 );
not ( n2326 , n2325 );
or ( n2327 , n2320 , n2326 );
not ( n2328 , n491 );
not ( n2329 , n1970 );
or ( n2330 , n2328 , n2329 );
nand ( n2331 , n1971 , n1715 );
nand ( n2332 , n2330 , n2331 );
nand ( n2333 , n2332 , n1739 );
nand ( n2334 , n2327 , n2333 );
and ( n2335 , n2319 , n2334 );
and ( n2336 , n2306 , n2318 );
or ( n2337 , n2335 , n2336 );
not ( n2338 , n2018 );
not ( n2339 , n2162 );
or ( n2340 , n2338 , n2339 );
not ( n2341 , n1077 );
and ( n2342 , n456 , n1773 );
not ( n2343 , n456 );
and ( n2344 , n2343 , n1776 );
nor ( n2345 , n2342 , n2344 );
not ( n2346 , n2345 );
or ( n2347 , n2341 , n2346 );
not ( n2348 , n459 );
nand ( n2349 , n2348 , n456 );
not ( n2350 , n2349 );
not ( n2351 , n456 );
nand ( n2352 , n2351 , n1776 );
not ( n2353 , n2352 );
or ( n2354 , n2350 , n2353 );
nand ( n2355 , n2354 , n499 );
nand ( n2356 , n2347 , n2355 );
nand ( n2357 , n1840 , n2356 );
nand ( n2358 , n2340 , n2357 );
not ( n2359 , n470 );
and ( n2360 , n456 , n2359 );
not ( n2361 , n456 );
not ( n2362 , n486 );
and ( n2363 , n2361 , n2362 );
nor ( n2364 , n2360 , n2363 );
and ( n2365 , n2364 , n489 );
xor ( n2366 , n2358 , n2365 );
not ( n2367 , n1784 );
not ( n2368 , n2180 );
or ( n2369 , n2367 , n2368 );
not ( n2370 , n495 );
not ( n2371 , n1735 );
or ( n2372 , n2370 , n2371 );
not ( n2373 , n456 );
not ( n2374 , n463 );
not ( n2375 , n2374 );
or ( n2376 , n2373 , n2375 );
nor ( n2377 , n456 , n479 );
nor ( n2378 , n2377 , n495 );
nand ( n2379 , n2376 , n2378 );
nand ( n2380 , n2372 , n2379 );
nand ( n2381 , n2380 , n1763 );
nand ( n2382 , n2369 , n2381 );
and ( n2383 , n2366 , n2382 );
and ( n2384 , n2358 , n2365 );
or ( n2385 , n2383 , n2384 );
xor ( n2386 , n2337 , n2385 );
xor ( n72340 , n2153 , n2169 );
xor ( n2388 , n72340 , n2184 );
and ( n2389 , n2386 , n2388 );
and ( n2390 , n2337 , n2385 );
or ( n2391 , n2389 , n2390 );
xor ( n2392 , n2291 , n2391 );
xor ( n2393 , n2193 , n2210 );
xor ( n2394 , n2393 , n2225 );
xor ( n2395 , n2249 , n2255 );
xor ( n2396 , n2395 , n2274 );
xor ( n2397 , n2394 , n2396 );
not ( n2398 , n71761 );
not ( n2399 , n2253 );
or ( n2400 , n2398 , n2399 );
and ( n2401 , n456 , n469 );
not ( n2402 , n456 );
and ( n2403 , n2402 , n485 );
nor ( n2404 , n2401 , n2403 );
not ( n2405 , n2404 );
not ( n2406 , n489 );
or ( n2407 , n2405 , n2406 );
and ( n2408 , n456 , n469 );
not ( n2409 , n456 );
and ( n2410 , n2409 , n485 );
nor ( n2411 , n2408 , n2410 );
not ( n2412 , n2411 );
nand ( n2413 , n2412 , n1649 );
nand ( n2414 , n2407 , n2413 );
nand ( n2415 , n2414 , n1828 );
nand ( n2416 , n2400 , n2415 );
not ( n2417 , n2274 );
xor ( n2418 , n2416 , n2417 );
not ( n2419 , n504 );
nand ( n2420 , n2419 , n503 );
not ( n2421 , n2420 );
not ( n2422 , n2421 );
nand ( n2423 , n503 , n504 );
nand ( n2424 , n2422 , n2423 );
not ( n2425 , n2424 );
and ( n2426 , n2418 , n2425 );
and ( n2427 , n2416 , n2417 );
or ( n2428 , n2426 , n2427 );
and ( n2429 , n2397 , n2428 );
and ( n2430 , n2394 , n2396 );
or ( n2431 , n2429 , n2430 );
and ( n2432 , n2392 , n2431 );
and ( n2433 , n2291 , n2391 );
or ( n2434 , n2432 , n2433 );
and ( n2435 , n2289 , n2434 );
and ( n2436 , n2286 , n2288 );
or ( n2437 , n2435 , n2436 );
or ( n2438 , n2284 , n2437 );
nand ( n2439 , n2284 , n2437 );
and ( n2440 , n2438 , n2439 );
xor ( n2441 , n2234 , n2236 );
xor ( n2442 , n2441 , n2277 );
xor ( n2443 , n2291 , n2391 );
xor ( n2444 , n2443 , n2431 );
xor ( n2445 , n2442 , n2444 );
xor ( n2446 , n2337 , n2385 );
xor ( n2447 , n2446 , n2388 );
not ( n2448 , n1848 );
not ( n2449 , n2314 );
or ( n2450 , n2448 , n2449 );
not ( n2451 , n497 );
not ( n2452 , n1917 );
or ( n2453 , n2451 , n2452 );
not ( n2454 , n497 );
and ( n2455 , n456 , n462 );
not ( n2456 , n456 );
and ( n2457 , n2456 , n478 );
or ( n2458 , n2455 , n2457 );
nand ( n2459 , n2454 , n2458 );
nand ( n2460 , n2453 , n2459 );
nand ( n2461 , n1869 , n2460 );
nand ( n2462 , n2450 , n2461 );
not ( n2463 , n2414 );
not ( n2464 , n1955 );
or ( n2465 , n2463 , n2464 );
not ( n2466 , n1649 );
and ( n72420 , n456 , n470 );
not ( n2471 , n456 );
and ( n2472 , n2471 , n486 );
or ( n2473 , n72420 , n2472 );
not ( n2474 , n2473 );
or ( n2475 , n2466 , n2474 );
not ( n2476 , n456 );
nand ( n2477 , n2476 , n486 );
nand ( n2478 , n456 , n470 );
nand ( n2479 , n2477 , n2478 , n489 );
nand ( n2480 , n2475 , n2479 );
nand ( n2481 , n1826 , n2480 );
nand ( n2482 , n2465 , n2481 );
xor ( n2483 , n2462 , n2482 );
and ( n2484 , n456 , n471 );
not ( n2485 , n456 );
and ( n2486 , n2485 , n487 );
nor ( n2487 , n2484 , n2486 );
not ( n2488 , n2487 );
and ( n2489 , n2488 , n489 );
and ( n2490 , n2483 , n2489 );
and ( n2491 , n2462 , n2482 );
or ( n2492 , n2490 , n2491 );
not ( n2493 , n1763 );
and ( n2494 , n495 , n1706 );
not ( n2495 , n495 );
and ( n2496 , n2495 , n1714 );
or ( n2497 , n2494 , n2496 );
not ( n2498 , n2497 );
or ( n2499 , n2493 , n2498 );
nand ( n2500 , n2380 , n1784 );
nand ( n2501 , n2499 , n2500 );
nand ( n2502 , n2149 , n2146 );
not ( n2503 , n2502 );
not ( n2504 , n2261 );
not ( n2505 , n1995 );
or ( n2506 , n2504 , n2505 );
and ( n2507 , n456 , n458 );
not ( n2508 , n456 );
and ( n2509 , n2508 , n474 );
nor ( n2510 , n2507 , n2509 );
nand ( n2511 , n501 , n2510 );
nand ( n2512 , n2506 , n2511 );
not ( n2513 , n2512 );
or ( n2514 , n2503 , n2513 );
nand ( n2515 , n2264 , n2272 );
nand ( n2516 , n2514 , n2515 );
xor ( n2517 , n2501 , n2516 );
not ( n2518 , n499 );
and ( n2519 , n456 , n460 );
not ( n2520 , n456 );
and ( n2521 , n2520 , n476 );
nor ( n2522 , n2519 , n2521 );
not ( n2523 , n2522 );
or ( n2524 , n2518 , n2523 );
not ( n2525 , n476 );
not ( n2526 , n456 );
nand ( n2527 , n2525 , n2526 );
not ( n2528 , n460 );
nand ( n2529 , n2528 , n456 );
nand ( n2530 , n2527 , n2529 , n70613 );
nand ( n2531 , n2524 , n2530 );
not ( n2532 , n2531 );
not ( n2533 , n2008 );
or ( n2534 , n2532 , n2533 );
nand ( n2535 , n2356 , n2018 );
nand ( n2536 , n2534 , n2535 );
and ( n2537 , n2517 , n2536 );
and ( n2538 , n2501 , n2516 );
or ( n2539 , n2537 , n2538 );
xor ( n2540 , n2492 , n2539 );
xor ( n2541 , n2306 , n2318 );
xor ( n2542 , n2541 , n2334 );
and ( n2543 , n2540 , n2542 );
and ( n2544 , n2492 , n2539 );
or ( n2545 , n2543 , n2544 );
xor ( n2546 , n2447 , n2545 );
xor ( n2547 , n2358 , n2365 );
xor ( n2548 , n2547 , n2382 );
not ( n2549 , n493 );
not ( n2550 , n1970 );
or ( n2551 , n2549 , n2550 );
not ( n2552 , n482 );
nand ( n2553 , n2351 , n2552 );
not ( n2554 , n466 );
nand ( n72505 , n2554 , n456 );
nand ( n2556 , n2553 , n72505 , n1976 );
nand ( n2557 , n2551 , n2556 );
nand ( n2558 , n2557 , n1908 );
not ( n2559 , n1976 );
not ( n2560 , n71767 );
or ( n2561 , n2559 , n2560 );
or ( n2562 , n71767 , n1976 );
nand ( n2563 , n2561 , n2562 );
nand ( n2564 , n1891 , n2563 );
nand ( n2565 , n2558 , n2564 );
not ( n2566 , n1739 );
not ( n2567 , n2325 );
or ( n2568 , n2566 , n2567 );
and ( n2569 , n456 , n468 );
not ( n2570 , n456 );
and ( n2571 , n2570 , n484 );
nor ( n2572 , n2569 , n2571 );
not ( n2573 , n2572 );
nand ( n2574 , n2573 , n1715 );
and ( n2575 , n456 , n468 );
not ( n2576 , n456 );
and ( n2577 , n2576 , n484 );
nor ( n2578 , n2575 , n2577 );
nand ( n2579 , n2578 , n491 );
nand ( n2580 , n2574 , n2579 );
nand ( n2581 , n2580 , n1700 );
nand ( n2582 , n2568 , n2581 );
xor ( n2583 , n2565 , n2582 );
and ( n2584 , n2583 , n2424 );
and ( n2585 , n2565 , n2582 );
or ( n2586 , n2584 , n2585 );
xor ( n2587 , n2548 , n2586 );
not ( n2588 , n1834 );
not ( n2589 , n2531 );
or ( n2590 , n2588 , n2589 );
and ( n2591 , n2164 , n499 );
and ( n2592 , n456 , n461 );
not ( n2593 , n456 );
and ( n2594 , n2593 , n477 );
or ( n2595 , n2592 , n2594 );
or ( n2596 , n2591 , n2595 );
and ( n2597 , n456 , n461 );
not ( n2598 , n456 );
and ( n2599 , n2598 , n477 );
nor ( n2600 , n2597 , n2599 );
not ( n2601 , n2600 );
not ( n2602 , n499 );
nand ( n2603 , n2602 , n501 , n500 );
nand ( n2604 , n2601 , n2603 );
nand ( n2605 , n2596 , n2604 );
nand ( n2606 , n2590 , n2605 );
not ( n2607 , n493 );
nor ( n2608 , n494 , n495 );
not ( n2609 , n2608 );
or ( n2610 , n2607 , n2609 );
nand ( n2611 , n2610 , n2297 );
not ( n2612 , n2611 );
not ( n2613 , n1976 );
not ( n2614 , n2102 );
or ( n2615 , n2613 , n2614 );
not ( n2616 , n456 );
nand ( n2617 , n2616 , n483 );
nand ( n2618 , n456 , n467 );
nand ( n2619 , n2617 , n2618 , n493 );
nand ( n2620 , n2615 , n2619 );
not ( n2621 , n2620 );
or ( n2622 , n2612 , n2621 );
nand ( n2623 , n2039 , n2557 );
nand ( n2624 , n2622 , n2623 );
xor ( n2625 , n2606 , n2624 );
not ( n2626 , n1928 );
not ( n2627 , n2580 );
or ( n2628 , n2626 , n2627 );
nand ( n2629 , n492 , n493 );
nor ( n2630 , n2629 , n491 );
or ( n2631 , n2192 , n2630 );
not ( n72582 , n491 );
nor ( n2636 , n492 , n493 );
not ( n2637 , n2636 );
or ( n2638 , n72582 , n2637 );
nand ( n2639 , n2638 , n2192 );
nand ( n2640 , n2631 , n2639 );
nand ( n2641 , n2628 , n2640 );
and ( n2642 , n2625 , n2641 );
and ( n2643 , n2606 , n2624 );
or ( n2644 , n2642 , n2643 );
not ( n2645 , n1826 );
not ( n2646 , n489 );
and ( n2647 , n456 , n471 );
not ( n2648 , n456 );
and ( n2649 , n2648 , n487 );
nor ( n2650 , n2647 , n2649 );
not ( n2651 , n2650 );
or ( n2652 , n2646 , n2651 );
or ( n2653 , n2650 , n489 );
nand ( n2654 , n2652 , n2653 );
not ( n2655 , n2654 );
or ( n2656 , n2645 , n2655 );
nand ( n2657 , n2480 , n1788 );
nand ( n2658 , n2656 , n2657 );
not ( n2659 , n2460 );
not ( n2660 , n498 );
not ( n2661 , n1077 );
or ( n2662 , n2660 , n2661 );
nand ( n2663 , n2662 , n1846 );
not ( n2664 , n2663 );
or ( n2665 , n2659 , n2664 );
not ( n2666 , n1760 );
and ( n2667 , n456 , n463 );
not ( n2668 , n456 );
and ( n2669 , n2668 , n479 );
nor ( n2670 , n2667 , n2669 );
not ( n2671 , n2670 );
not ( n2672 , n2671 );
or ( n2673 , n2666 , n2672 );
nand ( n2674 , n1735 , n497 );
nand ( n2675 , n2673 , n2674 );
nand ( n2676 , n2675 , n1869 );
nand ( n2677 , n2665 , n2676 );
xor ( n2678 , n2658 , n2677 );
not ( n2679 , n1763 );
not ( n2680 , n1801 );
not ( n2681 , n456 );
not ( n2682 , n481 );
and ( n2683 , n2681 , n2682 );
nor ( n2684 , n2683 , n495 );
not ( n2685 , n2684 );
or ( n2686 , n2680 , n2685 );
and ( n2687 , n456 , n465 );
not ( n2688 , n456 );
and ( n2689 , n2688 , n481 );
nor ( n2690 , n2687 , n2689 );
nand ( n2691 , n2690 , n495 );
nand ( n2692 , n2686 , n2691 );
not ( n2693 , n2692 );
or ( n2694 , n2679 , n2693 );
nand ( n2695 , n2497 , n1784 );
nand ( n2696 , n2694 , n2695 );
and ( n2697 , n2678 , n2696 );
and ( n2698 , n2658 , n2677 );
or ( n2699 , n2697 , n2698 );
xor ( n2700 , n2644 , n2699 );
and ( n2701 , n456 , n472 );
not ( n2702 , n456 );
and ( n2703 , n2702 , n488 );
or ( n2704 , n2701 , n2703 );
and ( n2705 , n2704 , n489 );
not ( n2706 , n2421 );
not ( n2707 , n2010 );
not ( n2708 , n2707 );
and ( n2709 , n2012 , n503 );
not ( n2710 , n2709 );
or ( n2711 , n2708 , n2710 );
not ( n2712 , n503 );
or ( n2713 , n456 , n473 );
not ( n2714 , n457 );
nand ( n2715 , n2714 , n456 );
nand ( n2716 , n2712 , n2713 , n2715 );
nand ( n2717 , n2711 , n2716 );
not ( n2718 , n2717 );
or ( n72666 , n2706 , n2718 );
nand ( n2720 , n72666 , n2423 );
xor ( n2721 , n2705 , n2720 );
buf ( n2722 , n2271 );
not ( n2723 , n2722 );
not ( n2724 , n2512 );
or ( n2725 , n2723 , n2724 );
and ( n2726 , n456 , n459 );
not ( n2727 , n456 );
and ( n2728 , n2727 , n475 );
nor ( n2729 , n2726 , n2728 );
not ( n2730 , n2729 );
and ( n2731 , n501 , n2730 );
not ( n2732 , n501 );
and ( n2733 , n2732 , n2729 );
nor ( n2734 , n2731 , n2733 );
buf ( n2735 , n2734 );
nand ( n2736 , n2735 , n2502 );
nand ( n2737 , n2725 , n2736 );
and ( n2738 , n2721 , n2737 );
and ( n2739 , n2705 , n2720 );
or ( n2740 , n2738 , n2739 );
and ( n2741 , n2700 , n2740 );
and ( n2742 , n2644 , n2699 );
or ( n2743 , n2741 , n2742 );
and ( n2744 , n2587 , n2743 );
and ( n2745 , n2548 , n2586 );
or ( n2746 , n2744 , n2745 );
and ( n2747 , n2546 , n2746 );
and ( n2748 , n2447 , n2545 );
or ( n2749 , n2747 , n2748 );
xor ( n2750 , n2445 , n2749 );
xor ( n2751 , n2394 , n2396 );
xor ( n2752 , n2751 , n2428 );
xor ( n2753 , n2416 , n2417 );
xor ( n2754 , n2753 , n2425 );
xor ( n2755 , n2492 , n2539 );
xor ( n2756 , n2755 , n2542 );
xor ( n2757 , n2754 , n2756 );
xor ( n2758 , n2462 , n2482 );
xor ( n2759 , n2758 , n2489 );
xor ( n2760 , n2501 , n2516 );
xor ( n2761 , n2760 , n2536 );
xor ( n2762 , n2759 , n2761 );
xor ( n2763 , n2565 , n2582 );
xor ( n2764 , n2763 , n2424 );
and ( n2765 , n2762 , n2764 );
and ( n2766 , n2759 , n2761 );
or ( n2767 , n2765 , n2766 );
and ( n2768 , n2757 , n2767 );
and ( n2769 , n2754 , n2756 );
or ( n2770 , n2768 , n2769 );
xor ( n2771 , n2752 , n2770 );
xor ( n2772 , n2447 , n2545 );
xor ( n2773 , n2772 , n2746 );
and ( n2774 , n2771 , n2773 );
and ( n2775 , n2752 , n2770 );
or ( n2776 , n2774 , n2775 );
nor ( n2777 , n2750 , n2776 );
xor ( n2778 , n2286 , n2288 );
xor ( n2779 , n2778 , n2434 );
xor ( n2780 , n2442 , n2444 );
and ( n2781 , n2780 , n2749 );
and ( n2782 , n2442 , n2444 );
or ( n2783 , n2781 , n2782 );
nor ( n2784 , n2779 , n2783 );
nor ( n2785 , n2777 , n2784 );
xor ( n2786 , n2752 , n2770 );
xor ( n2787 , n2786 , n2773 );
xor ( n2788 , n2548 , n2586 );
xor ( n2789 , n2788 , n2743 );
and ( n2790 , n456 , n472 );
not ( n2791 , n456 );
and ( n2792 , n2791 , n488 );
nor ( n2793 , n2790 , n2792 );
not ( n2794 , n2793 );
not ( n2795 , n1821 );
and ( n2796 , n2794 , n2795 );
nand ( n2797 , n490 , n491 );
nand ( n72745 , n2797 , n489 );
nor ( n2802 , n2796 , n72745 );
not ( n2803 , n504 );
not ( n2804 , n2717 );
or ( n2805 , n2803 , n2804 );
not ( n2806 , n503 );
and ( n2807 , n456 , n458 );
not ( n2808 , n456 );
and ( n2809 , n2808 , n474 );
nor ( n2810 , n2807 , n2809 );
and ( n2811 , n2806 , n2810 );
not ( n2812 , n2806 );
and ( n2813 , n2812 , n1881 );
nor ( n2814 , n2811 , n2813 );
nand ( n2815 , n2814 , n2421 );
nand ( n2816 , n2805 , n2815 );
and ( n2817 , n2802 , n2816 );
not ( n2818 , n2722 );
not ( n2819 , n2734 );
or ( n2820 , n2818 , n2819 );
not ( n2821 , n1746 );
nand ( n2822 , n2821 , n501 );
nand ( n2823 , n2149 , n2146 );
nand ( n2824 , n1981 , n2261 );
nand ( n2825 , n2822 , n2823 , n2824 );
nand ( n2826 , n2820 , n2825 );
not ( n2827 , n1788 );
not ( n2828 , n2654 );
or ( n2829 , n2827 , n2828 );
not ( n2830 , n489 );
and ( n2831 , n456 , n472 );
not ( n2832 , n456 );
and ( n2833 , n2832 , n488 );
nor ( n2834 , n2831 , n2833 );
not ( n2835 , n2834 );
or ( n2836 , n2830 , n2835 );
and ( n2837 , n456 , n472 );
not ( n2838 , n456 );
and ( n2839 , n2838 , n488 );
nor ( n2840 , n2837 , n2839 );
not ( n2841 , n2840 );
nand ( n2842 , n2841 , n1649 );
nand ( n2843 , n2836 , n2842 );
nand ( n2844 , n2843 , n1826 );
nand ( n2845 , n2829 , n2844 );
xor ( n2846 , n2826 , n2845 );
not ( n2847 , n497 );
not ( n2848 , n2847 );
not ( n2849 , n464 );
and ( n2850 , n456 , n2849 );
not ( n2851 , n456 );
not ( n2852 , n480 );
and ( n2853 , n2851 , n2852 );
nor ( n2854 , n2850 , n2853 );
not ( n2855 , n2854 );
or ( n2856 , n2848 , n2855 );
not ( n2857 , n464 );
and ( n2858 , n456 , n2857 );
not ( n2859 , n456 );
and ( n2860 , n2859 , n2852 );
nor ( n2861 , n2858 , n2860 );
or ( n2862 , n2861 , n2847 );
nand ( n2863 , n2856 , n2862 );
not ( n2864 , n2863 );
not ( n2865 , n1869 );
or ( n2866 , n2864 , n2865 );
nand ( n2867 , n2675 , n1848 );
nand ( n2868 , n2866 , n2867 );
and ( n2869 , n2846 , n2868 );
and ( n2870 , n2826 , n2845 );
or ( n2871 , n2869 , n2870 );
xor ( n2872 , n2817 , n2871 );
and ( n2873 , n496 , n497 );
not ( n2874 , n496 );
and ( n2875 , n2874 , n70541 );
nor ( n2876 , n2873 , n2875 );
not ( n2877 , n2876 );
not ( n2878 , n2692 );
or ( n2879 , n2877 , n2878 );
not ( n2880 , n495 );
and ( n2881 , n456 , n466 );
not ( n72826 , n456 );
and ( n2883 , n72826 , n482 );
nor ( n2884 , n2881 , n2883 );
not ( n2885 , n2884 );
or ( n2886 , n2880 , n2885 );
not ( n2887 , n2351 );
not ( n2888 , n2552 );
or ( n2889 , n2887 , n2888 );
and ( n2890 , n2554 , n456 );
nor ( n2891 , n2890 , n495 );
nand ( n2892 , n2889 , n2891 );
nand ( n2893 , n2886 , n2892 );
not ( n2894 , n70541 );
not ( n2895 , n495 );
nor ( n2896 , n2895 , n496 );
not ( n2897 , n2896 );
or ( n2898 , n2894 , n2897 );
nand ( n2899 , n2898 , n1759 );
nand ( n2900 , n2893 , n2899 );
nand ( n2901 , n2879 , n2900 );
not ( n2902 , n1840 );
and ( n2903 , n499 , n1917 );
not ( n2904 , n499 );
not ( n2905 , n478 );
not ( n2906 , n456 );
not ( n2907 , n2906 );
or ( n2908 , n2905 , n2907 );
nand ( n2909 , n456 , n462 );
nand ( n2910 , n2908 , n2909 );
and ( n2911 , n2904 , n2910 );
or ( n2912 , n2903 , n2911 );
not ( n2913 , n2912 );
or ( n2914 , n2902 , n2913 );
not ( n2915 , n499 );
nand ( n2916 , n2915 , n2088 );
not ( n2917 , n2916 );
nand ( n2918 , n2311 , n2312 , n499 );
not ( n2919 , n2918 );
or ( n2920 , n2917 , n2919 );
nand ( n2921 , n2920 , n1834 );
nand ( n2922 , n2914 , n2921 );
xor ( n2923 , n2901 , n2922 );
not ( n2924 , n1908 );
not ( n2925 , n493 );
nand ( n2926 , n2925 , n2573 );
and ( n2927 , n456 , n468 );
not ( n2928 , n456 );
and ( n2929 , n2928 , n484 );
nor ( n2930 , n2927 , n2929 );
nand ( n2931 , n2930 , n493 );
nand ( n2932 , n2926 , n2931 );
not ( n2933 , n2932 );
or ( n2934 , n2924 , n2933 );
nand ( n2935 , n2620 , n2039 );
nand ( n2936 , n2934 , n2935 );
and ( n2937 , n2923 , n2936 );
and ( n2938 , n2901 , n2922 );
or ( n2939 , n2937 , n2938 );
and ( n2940 , n2872 , n2939 );
and ( n2941 , n2817 , n2871 );
or ( n2942 , n2940 , n2941 );
xor ( n2943 , n2644 , n2699 );
xor ( n2944 , n2943 , n2740 );
xor ( n2945 , n2942 , n2944 );
xor ( n2946 , n2606 , n2624 );
xor ( n2947 , n2946 , n2641 );
xor ( n2948 , n2705 , n2720 );
xor ( n2949 , n2948 , n2737 );
xor ( n2950 , n2947 , n2949 );
xor ( n2951 , n2658 , n2677 );
xor ( n2952 , n2951 , n2696 );
and ( n2953 , n2950 , n2952 );
and ( n2954 , n2947 , n2949 );
or ( n2955 , n2953 , n2954 );
and ( n2956 , n2945 , n2955 );
and ( n72901 , n2942 , n2944 );
or ( n2961 , n2956 , n72901 );
xor ( n2962 , n2789 , n2961 );
xor ( n2963 , n2754 , n2756 );
xor ( n2964 , n2963 , n2767 );
and ( n2965 , n2962 , n2964 );
and ( n2966 , n2789 , n2961 );
or ( n2967 , n2965 , n2966 );
nor ( n2968 , n2787 , n2967 );
not ( n2969 , n2968 );
nand ( n2970 , n2785 , n2969 );
not ( n2971 , n2970 );
xor ( n2972 , n2947 , n2949 );
xor ( n2973 , n2972 , n2952 );
not ( n2974 , n1908 );
nand ( n2975 , n2526 , n485 );
nand ( n2976 , n456 , n469 );
nand ( n2977 , n2975 , n2976 );
xor ( n2978 , n493 , n2977 );
not ( n2979 , n2978 );
or ( n2980 , n2974 , n2979 );
nand ( n2981 , n2932 , n2039 );
nand ( n2982 , n2980 , n2981 );
not ( n2983 , n1928 );
not ( n2984 , n491 );
and ( n2985 , n456 , n470 );
not ( n2986 , n456 );
and ( n2987 , n2986 , n486 );
nor ( n2988 , n2985 , n2987 );
not ( n2989 , n2988 );
or ( n2990 , n2984 , n2989 );
and ( n2991 , n456 , n470 );
not ( n2992 , n456 );
and ( n2993 , n2992 , n486 );
nor ( n2994 , n2991 , n2993 );
not ( n2995 , n2994 );
nand ( n2996 , n2995 , n1715 );
nand ( n2997 , n2990 , n2996 );
not ( n2998 , n2997 );
or ( n2999 , n2983 , n2998 );
not ( n3000 , n491 );
and ( n3001 , n456 , n471 );
not ( n3002 , n456 );
and ( n3003 , n3002 , n487 );
nor ( n3004 , n3001 , n3003 );
not ( n3005 , n3004 );
or ( n3006 , n3000 , n3005 );
nand ( n3007 , n2488 , n1715 );
nand ( n3008 , n3006 , n3007 );
nand ( n3009 , n3008 , n1941 );
nand ( n3010 , n2999 , n3009 );
xor ( n3011 , n2982 , n3010 );
not ( n3012 , n488 );
or ( n3013 , n3012 , n456 );
nand ( n3014 , n456 , n472 );
nand ( n3015 , n3013 , n3014 );
or ( n3016 , n3015 , n492 );
nand ( n3017 , n3016 , n493 );
and ( n3018 , n3015 , n492 );
nor ( n3019 , n3018 , n1715 );
and ( n3020 , n3017 , n3019 );
not ( n3021 , n2421 );
and ( n3022 , n456 , n2528 );
not ( n3023 , n456 );
and ( n3024 , n3023 , n2525 );
nor ( n3025 , n3022 , n3024 );
not ( n3026 , n3025 );
not ( n3027 , n503 );
not ( n3028 , n3027 );
or ( n3029 , n3026 , n3028 );
nand ( n3030 , n1746 , n503 );
nand ( n3031 , n3029 , n3030 );
not ( n3032 , n3031 );
or ( n3033 , n3021 , n3032 );
and ( n3034 , n456 , n459 );
not ( n3035 , n456 );
and ( n3036 , n3035 , n475 );
nor ( n72978 , n3034 , n3036 );
and ( n3038 , n503 , n72978 );
not ( n3039 , n503 );
and ( n3040 , n3039 , n2345 );
or ( n3041 , n3038 , n3040 );
nand ( n3042 , n3041 , n504 );
nand ( n3043 , n3033 , n3042 );
and ( n3044 , n3020 , n3043 );
and ( n3045 , n3011 , n3044 );
and ( n3046 , n2982 , n3010 );
or ( n3047 , n3045 , n3046 );
not ( n3048 , n1928 );
and ( n3049 , n456 , n469 );
not ( n3050 , n456 );
and ( n3051 , n3050 , n485 );
or ( n3052 , n3049 , n3051 );
and ( n3053 , n491 , n3052 );
not ( n3054 , n491 );
and ( n3055 , n3054 , n2192 );
nor ( n3056 , n3053 , n3055 );
not ( n3057 , n3056 );
or ( n3058 , n3048 , n3057 );
nand ( n3059 , n2997 , n1941 );
nand ( n3060 , n3058 , n3059 );
xor ( n3061 , n2802 , n2816 );
xor ( n3062 , n3060 , n3061 );
not ( n3063 , n2840 );
and ( n3064 , n3063 , n1788 );
not ( n3065 , n503 );
nor ( n3066 , n3065 , n504 );
not ( n3067 , n3066 );
not ( n3068 , n3041 );
or ( n3069 , n3067 , n3068 );
nand ( n3070 , n2814 , n504 );
nand ( n3071 , n3069 , n3070 );
xor ( n3072 , n3064 , n3071 );
not ( n3073 , n2142 );
and ( n3074 , n2261 , n1981 );
not ( n3075 , n2261 );
not ( n3076 , n1746 );
and ( n3077 , n3075 , n3076 );
nor ( n3078 , n3074 , n3077 );
not ( n3079 , n3078 );
or ( n3080 , n3073 , n3079 );
not ( n3081 , n501 );
not ( n3082 , n2600 );
or ( n3083 , n3081 , n3082 );
not ( n3084 , n2616 );
not ( n3085 , n477 );
not ( n3086 , n3085 );
or ( n3087 , n3084 , n3086 );
not ( n3088 , n461 );
and ( n3089 , n3088 , n456 );
nor ( n3090 , n3089 , n501 );
nand ( n3091 , n3087 , n3090 );
nand ( n3092 , n3083 , n3091 );
nand ( n3093 , n2502 , n3092 );
nand ( n3094 , n3080 , n3093 );
and ( n3095 , n3072 , n3094 );
and ( n3096 , n3064 , n3071 );
or ( n3097 , n3095 , n3096 );
xor ( n3098 , n3062 , n3097 );
xor ( n3099 , n3047 , n3098 );
not ( n3100 , n2823 );
not ( n3101 , n501 );
and ( n3102 , n456 , n462 );
not ( n3103 , n456 );
and ( n3104 , n3103 , n478 );
nor ( n3105 , n3102 , n3104 );
not ( n3106 , n3105 );
or ( n3107 , n3101 , n3106 );
not ( n73049 , n462 );
and ( n3112 , n456 , n73049 );
not ( n3113 , n456 );
not ( n3114 , n478 );
and ( n3115 , n3113 , n3114 );
nor ( n3116 , n3112 , n3115 );
not ( n3117 , n501 );
nand ( n3118 , n3116 , n3117 );
nand ( n3119 , n3107 , n3118 );
not ( n3120 , n3119 );
or ( n3121 , n3100 , n3120 );
nand ( n3122 , n3092 , n2142 );
nand ( n3123 , n3121 , n3122 );
not ( n3124 , n1869 );
not ( n3125 , n497 );
not ( n3126 , n2884 );
or ( n3127 , n3125 , n3126 );
not ( n3128 , n2884 );
not ( n3129 , n497 );
nand ( n3130 , n3128 , n3129 );
nand ( n3131 , n3127 , n3130 );
not ( n3132 , n3131 );
or ( n3133 , n3124 , n3132 );
not ( n3134 , n2847 );
nand ( n3135 , n2906 , n481 );
nand ( n3136 , n456 , n465 );
nand ( n3137 , n3135 , n3136 );
not ( n3138 , n3137 );
or ( n3139 , n3134 , n3138 );
nand ( n3140 , n1795 , n497 );
nand ( n3141 , n3139 , n3140 );
xor ( n3142 , n498 , n499 );
nand ( n3143 , n3141 , n3142 );
nand ( n3144 , n3133 , n3143 );
xor ( n3145 , n3123 , n3144 );
not ( n3146 , n2876 );
not ( n3147 , n70594 );
not ( n3148 , n2102 );
or ( n3149 , n3147 , n3148 );
or ( n3150 , n70594 , n2102 );
nand ( n3151 , n3149 , n3150 );
not ( n3152 , n3151 );
or ( n3153 , n3146 , n3152 );
not ( n3154 , n495 );
and ( n3155 , n456 , n468 );
not ( n3156 , n456 );
and ( n3157 , n3156 , n484 );
nor ( n3158 , n3155 , n3157 );
not ( n3159 , n3158 );
or ( n3160 , n3154 , n3159 );
or ( n3161 , n495 , n2930 );
nand ( n3162 , n3160 , n3161 );
nand ( n3163 , n3162 , n1763 );
nand ( n3164 , n3153 , n3163 );
and ( n3165 , n3145 , n3164 );
and ( n3166 , n3123 , n3144 );
or ( n3167 , n3165 , n3166 );
not ( n3168 , n1258 );
not ( n3169 , n2861 );
or ( n3170 , n3168 , n3169 );
or ( n3171 , n1712 , n456 );
or ( n3172 , n1709 , n2086 );
nand ( n3173 , n3171 , n3172 , n499 );
nand ( n3174 , n3170 , n3173 );
not ( n3175 , n3174 );
not ( n3176 , n1840 );
or ( n3177 , n3175 , n3176 );
not ( n3178 , n499 );
not ( n3179 , n2670 );
or ( n3180 , n3178 , n3179 );
or ( n3181 , n2670 , n499 );
nand ( n73120 , n3180 , n3181 );
nand ( n3183 , n73120 , n1834 );
nand ( n3184 , n3177 , n3183 );
not ( n3185 , n2039 );
not ( n3186 , n2978 );
or ( n3187 , n3185 , n3186 );
not ( n3188 , n493 );
not ( n3189 , n3188 );
and ( n3190 , n456 , n2359 );
not ( n3191 , n456 );
and ( n3192 , n3191 , n2362 );
nor ( n3193 , n3190 , n3192 );
not ( n3194 , n3193 );
or ( n3195 , n3189 , n3194 );
or ( n3196 , n3193 , n3188 );
nand ( n3197 , n3195 , n3196 );
nand ( n3198 , n3197 , n2611 );
nand ( n3199 , n3187 , n3198 );
xor ( n3200 , n3184 , n3199 );
not ( n3201 , n1739 );
not ( n3202 , n3008 );
or ( n3203 , n3201 , n3202 );
not ( n3204 , n491 );
not ( n3205 , n2834 );
or ( n3206 , n3204 , n3205 );
or ( n3207 , n2834 , n491 );
nand ( n3208 , n3206 , n3207 );
nand ( n3209 , n1941 , n3208 );
nand ( n3210 , n3203 , n3209 );
and ( n3211 , n3200 , n3210 );
and ( n3212 , n3184 , n3199 );
or ( n3213 , n3211 , n3212 );
xor ( n3214 , n3167 , n3213 );
xor ( n3215 , n3064 , n3071 );
xor ( n3216 , n3215 , n3094 );
and ( n3217 , n3214 , n3216 );
and ( n3218 , n3167 , n3213 );
or ( n3219 , n3217 , n3218 );
and ( n3220 , n3099 , n3219 );
and ( n3221 , n3047 , n3098 );
or ( n3222 , n3220 , n3221 );
xor ( n3223 , n2973 , n3222 );
xor ( n3224 , n3060 , n3061 );
and ( n3225 , n3224 , n3097 );
and ( n3226 , n3060 , n3061 );
or ( n3227 , n3225 , n3226 );
xor ( n3228 , n2817 , n2871 );
xor ( n3229 , n3228 , n2939 );
xor ( n3230 , n3227 , n3229 );
nand ( n3231 , n1869 , n3141 );
nand ( n3232 , n2863 , n3142 );
nand ( n3233 , n3231 , n3232 );
not ( n3234 , n1763 );
not ( n3235 , n3151 );
or ( n3236 , n3234 , n3235 );
and ( n3237 , n496 , n497 );
not ( n3238 , n496 );
and ( n3239 , n3238 , n70541 );
nor ( n3240 , n3237 , n3239 );
nand ( n3241 , n2893 , n3240 );
nand ( n3242 , n3236 , n3241 );
xor ( n3243 , n3233 , n3242 );
not ( n3244 , n2167 );
not ( n3245 , n73120 );
or ( n3246 , n3244 , n3245 );
nand ( n73185 , n2912 , n1834 );
nand ( n3251 , n3246 , n73185 );
and ( n3252 , n3243 , n3251 );
and ( n3253 , n3233 , n3242 );
or ( n3254 , n3252 , n3253 );
xor ( n3255 , n2901 , n2922 );
xor ( n3256 , n3255 , n2936 );
xor ( n3257 , n3254 , n3256 );
xor ( n3258 , n2826 , n2845 );
xor ( n3259 , n3258 , n2868 );
and ( n3260 , n3257 , n3259 );
and ( n3261 , n3254 , n3256 );
or ( n3262 , n3260 , n3261 );
xor ( n3263 , n3230 , n3262 );
xor ( n3264 , n3223 , n3263 );
not ( n3265 , n3264 );
xor ( n3266 , n3254 , n3256 );
xor ( n3267 , n3266 , n3259 );
xor ( n3268 , n3233 , n3242 );
xor ( n3269 , n3268 , n3251 );
xor ( n3270 , n2982 , n3010 );
xor ( n3271 , n3270 , n3044 );
xor ( n3272 , n3269 , n3271 );
xor ( n3273 , n3020 , n3043 );
and ( n3274 , n456 , n472 );
not ( n3275 , n456 );
and ( n3276 , n3275 , n488 );
or ( n3277 , n3274 , n3276 );
and ( n3278 , n1928 , n3277 );
not ( n3279 , n501 );
not ( n3280 , n1735 );
or ( n3281 , n3279 , n3280 );
not ( n3282 , n479 );
nand ( n3283 , n3282 , n2351 );
not ( n3284 , n463 );
nand ( n3285 , n3284 , n456 );
nand ( n3286 , n3283 , n3285 , n2261 );
nand ( n3287 , n3281 , n3286 );
not ( n3288 , n3287 );
not ( n3289 , n2259 );
or ( n3290 , n3288 , n3289 );
not ( n3291 , n503 );
not ( n3292 , n2140 );
or ( n3293 , n3291 , n3292 );
nand ( n3294 , n2137 , n502 );
nand ( n3295 , n3293 , n3294 );
nand ( n3296 , n3119 , n3295 );
nand ( n3297 , n3290 , n3296 );
xor ( n3298 , n3278 , n3297 );
not ( n3299 , n1848 );
not ( n3300 , n3131 );
or ( n3301 , n3299 , n3300 );
not ( n3302 , n497 );
and ( n3303 , n456 , n467 );
not ( n3304 , n456 );
and ( n3305 , n3304 , n483 );
nor ( n3306 , n3303 , n3305 );
not ( n3307 , n3306 );
or ( n3308 , n3302 , n3307 );
or ( n3309 , n3306 , n497 );
nand ( n3310 , n3308 , n3309 );
nand ( n3311 , n3310 , n1869 );
nand ( n3312 , n3301 , n3311 );
and ( n3313 , n3298 , n3312 );
and ( n3314 , n3278 , n3297 );
or ( n3315 , n3313 , n3314 );
xor ( n3316 , n3273 , n3315 );
not ( n73252 , n3240 );
not ( n3318 , n3162 );
or ( n3319 , n73252 , n3318 );
not ( n3320 , n485 );
not ( n3321 , n71699 );
or ( n3322 , n3320 , n3321 );
nand ( n3323 , n456 , n469 );
nand ( n3324 , n3322 , n3323 );
not ( n3325 , n495 );
nand ( n3326 , n3324 , n3325 );
and ( n3327 , n456 , n469 );
not ( n3328 , n456 );
and ( n3329 , n3328 , n485 );
nor ( n3330 , n3327 , n3329 );
nand ( n3331 , n3330 , n495 );
nand ( n3332 , n3326 , n3331 );
nand ( n3333 , n2899 , n3332 );
nand ( n3334 , n3319 , n3333 );
not ( n3335 , n3066 );
not ( n3336 , n2269 );
not ( n3337 , n2088 );
or ( n3338 , n3336 , n3337 );
nand ( n3339 , n1896 , n503 );
nand ( n3340 , n3338 , n3339 );
not ( n3341 , n3340 );
or ( n3342 , n3335 , n3341 );
nand ( n3343 , n3031 , n504 );
nand ( n3344 , n3342 , n3343 );
xor ( n3345 , n3334 , n3344 );
not ( n3346 , n1891 );
not ( n3347 , n3197 );
or ( n3348 , n3346 , n3347 );
and ( n3349 , n493 , n3004 );
not ( n3350 , n493 );
and ( n3351 , n3350 , n2488 );
or ( n3352 , n3349 , n3351 );
nand ( n3353 , n3352 , n2611 );
nand ( n3354 , n3348 , n3353 );
and ( n3355 , n3345 , n3354 );
and ( n3356 , n3334 , n3344 );
or ( n3357 , n3355 , n3356 );
and ( n3358 , n3316 , n3357 );
and ( n3359 , n3273 , n3315 );
or ( n3360 , n3358 , n3359 );
and ( n3361 , n3272 , n3360 );
and ( n3362 , n3269 , n3271 );
or ( n3363 , n3361 , n3362 );
xor ( n3364 , n3267 , n3363 );
xor ( n3365 , n3047 , n3098 );
xor ( n3366 , n3365 , n3219 );
and ( n3367 , n3364 , n3366 );
and ( n3368 , n3267 , n3363 );
or ( n3369 , n3367 , n3368 );
not ( n3370 , n3369 );
nand ( n3371 , n3265 , n3370 );
buf ( n3372 , n3371 );
xor ( n3373 , n2789 , n2961 );
xor ( n3374 , n3373 , n2964 );
not ( n3375 , n3374 );
xor ( n3376 , n2759 , n2761 );
xor ( n3377 , n3376 , n2764 );
xor ( n73313 , n3227 , n3229 );
and ( n3382 , n73313 , n3262 );
and ( n3383 , n3227 , n3229 );
or ( n3384 , n3382 , n3383 );
xor ( n3385 , n3377 , n3384 );
xor ( n3386 , n2942 , n2944 );
xor ( n3387 , n3386 , n2955 );
and ( n3388 , n3385 , n3387 );
and ( n3389 , n3377 , n3384 );
or ( n3390 , n3388 , n3389 );
not ( n3391 , n3390 );
nand ( n3392 , n3375 , n3391 );
xor ( n3393 , n3377 , n3384 );
xor ( n3394 , n3393 , n3387 );
not ( n3395 , n3394 );
xor ( n3396 , n2973 , n3222 );
and ( n3397 , n3396 , n3263 );
and ( n3398 , n2973 , n3222 );
or ( n3399 , n3397 , n3398 );
not ( n3400 , n3399 );
nand ( n3401 , n3395 , n3400 );
and ( n3402 , n3372 , n3392 , n3401 );
xor ( n3403 , n3167 , n3213 );
xor ( n3404 , n3403 , n3216 );
xor ( n3405 , n3269 , n3271 );
xor ( n3406 , n3405 , n3360 );
xor ( n3407 , n3404 , n3406 );
xor ( n3408 , n3184 , n3199 );
xor ( n3409 , n3408 , n3210 );
xor ( n3410 , n3123 , n3144 );
xor ( n3411 , n3410 , n3164 );
xor ( n3412 , n3409 , n3411 );
not ( n3413 , n499 );
not ( n3414 , n2690 );
or ( n3415 , n3413 , n3414 );
nand ( n3416 , n3137 , n1864 );
nand ( n3417 , n3415 , n3416 );
not ( n3418 , n3417 );
not ( n3419 , n2008 );
or ( n3420 , n3418 , n3419 );
nand ( n3421 , n3174 , n2018 );
nand ( n3422 , n3420 , n3421 );
nand ( n3423 , n1888 , n70594 );
nand ( n3424 , n3423 , n3063 );
nand ( n3425 , n494 , n495 );
and ( n3426 , n3424 , n3425 , n493 );
not ( n3427 , n3295 );
not ( n3428 , n3287 );
or ( n3429 , n3427 , n3428 );
not ( n3430 , n2854 );
not ( n3431 , n2261 );
or ( n3432 , n3430 , n3431 );
nand ( n3433 , n1706 , n501 );
nand ( n3434 , n3432 , n3433 );
nand ( n3435 , n2259 , n3434 );
nand ( n3436 , n3429 , n3435 );
and ( n3437 , n3426 , n3436 );
xor ( n3438 , n3422 , n3437 );
not ( n3439 , n3142 );
not ( n3440 , n3310 );
or ( n3441 , n3439 , n3440 );
not ( n73374 , n2213 );
not ( n3443 , n3158 );
not ( n3444 , n3443 );
or ( n3445 , n73374 , n3444 );
nand ( n3446 , n2578 , n497 );
nand ( n3447 , n3445 , n3446 );
nand ( n3448 , n1869 , n3447 );
nand ( n3449 , n3441 , n3448 );
not ( n3450 , n1763 );
not ( n3451 , n495 );
not ( n3452 , n2988 );
or ( n3453 , n3451 , n3452 );
not ( n3454 , n495 );
and ( n3455 , n456 , n470 );
not ( n3456 , n456 );
and ( n3457 , n3456 , n486 );
or ( n3458 , n3455 , n3457 );
nand ( n3459 , n3454 , n3458 );
nand ( n3460 , n3453 , n3459 );
not ( n3461 , n3460 );
or ( n3462 , n3450 , n3461 );
nand ( n3463 , n3332 , n2876 );
nand ( n3464 , n3462 , n3463 );
xor ( n3465 , n3449 , n3464 );
not ( n3466 , n504 );
not ( n3467 , n3340 );
or ( n3468 , n3466 , n3467 );
not ( n3469 , n2909 );
nand ( n3470 , n3469 , n3027 );
nand ( n3471 , n3105 , n503 );
nand ( n3472 , n478 , n3027 , n2616 );
nand ( n3473 , n3470 , n3471 , n3472 );
nand ( n3474 , n3473 , n2421 );
nand ( n3475 , n3468 , n3474 );
and ( n3476 , n3465 , n3475 );
and ( n3477 , n3449 , n3464 );
or ( n3478 , n3476 , n3477 );
and ( n3479 , n3438 , n3478 );
and ( n3480 , n3422 , n3437 );
or ( n3481 , n3479 , n3480 );
and ( n3482 , n3412 , n3481 );
and ( n3483 , n3409 , n3411 );
or ( n3484 , n3482 , n3483 );
xor ( n3485 , n3407 , n3484 );
not ( n3486 , n3485 );
xor ( n3487 , n3273 , n3315 );
xor ( n3488 , n3487 , n3357 );
xor ( n3489 , n3334 , n3344 );
xor ( n3490 , n3489 , n3354 );
xor ( n3491 , n3278 , n3297 );
xor ( n3492 , n3491 , n3312 );
xor ( n3493 , n3490 , n3492 );
not ( n3494 , n2039 );
not ( n3495 , n3352 );
or ( n3496 , n3494 , n3495 );
and ( n3497 , n493 , n2834 );
not ( n3498 , n493 );
and ( n73431 , n3498 , n3277 );
or ( n3503 , n3497 , n73431 );
nand ( n3504 , n3503 , n2611 );
nand ( n3505 , n3496 , n3504 );
not ( n3506 , n2008 );
not ( n3507 , n1077 );
not ( n3508 , n1971 );
or ( n3509 , n3507 , n3508 );
nand ( n3510 , n1814 , n499 );
nand ( n3511 , n3509 , n3510 );
not ( n3512 , n3511 );
or ( n3513 , n3506 , n3512 );
nand ( n3514 , n3417 , n2018 );
nand ( n3515 , n3513 , n3514 );
xor ( n3516 , n3505 , n3515 );
xor ( n3517 , n3426 , n3436 );
and ( n3518 , n3516 , n3517 );
and ( n3519 , n3505 , n3515 );
or ( n3520 , n3518 , n3519 );
and ( n3521 , n3493 , n3520 );
and ( n3522 , n3490 , n3492 );
or ( n3523 , n3521 , n3522 );
xor ( n3524 , n3488 , n3523 );
xor ( n3525 , n3409 , n3411 );
xor ( n3526 , n3525 , n3481 );
and ( n3527 , n3524 , n3526 );
and ( n3528 , n3488 , n3523 );
or ( n3529 , n3527 , n3528 );
not ( n3530 , n3529 );
nor ( n3531 , n3486 , n3530 );
not ( n3532 , n3531 );
xor ( n3533 , n3267 , n3363 );
xor ( n3534 , n3533 , n3366 );
not ( n3535 , n3534 );
xor ( n3536 , n3404 , n3406 );
and ( n3537 , n3536 , n3484 );
and ( n3538 , n3404 , n3406 );
or ( n3539 , n3537 , n3538 );
not ( n3540 , n3539 );
nand ( n3541 , n3535 , n3540 );
not ( n3542 , n3541 );
or ( n3543 , n3532 , n3542 );
not ( n3544 , n3369 );
not ( n3545 , n3264 );
or ( n3546 , n3544 , n3545 );
nand ( n3547 , n3534 , n3539 );
nand ( n3548 , n3546 , n3547 );
not ( n3549 , n3548 );
nand ( n3550 , n3543 , n3549 );
not ( n3551 , n3550 );
not ( n3552 , n2876 );
not ( n3553 , n3460 );
or ( n3554 , n3552 , n3553 );
nor ( n3555 , n456 , n487 );
not ( n3556 , n3555 );
not ( n3557 , n471 );
nand ( n3558 , n3557 , n456 );
nand ( n73488 , n3556 , n3558 , n3325 );
not ( n3560 , n70594 );
nand ( n3561 , n3560 , n3004 );
nand ( n3562 , n73488 , n3561 );
nand ( n3563 , n3562 , n2899 );
nand ( n3564 , n3554 , n3563 );
not ( n3565 , n504 );
not ( n3566 , n3473 );
or ( n3567 , n3565 , n3566 );
xor ( n3568 , n503 , n2671 );
nand ( n3569 , n3568 , n3066 );
nand ( n3570 , n3567 , n3569 );
xor ( n3571 , n3564 , n3570 );
not ( n3572 , n2167 );
not ( n3573 , n499 );
not ( n3574 , n2005 );
or ( n3575 , n3573 , n3574 );
and ( n3576 , n456 , n467 );
not ( n3577 , n456 );
and ( n3578 , n3577 , n483 );
nor ( n3579 , n3576 , n3578 );
not ( n3580 , n3579 );
nand ( n3581 , n1077 , n3580 );
nand ( n3582 , n3575 , n3581 );
not ( n3583 , n3582 );
or ( n3584 , n3572 , n3583 );
nand ( n3585 , n3511 , n1834 );
nand ( n3586 , n3584 , n3585 );
xor ( n3587 , n3571 , n3586 );
not ( n3588 , n2018 );
not ( n3589 , n3582 );
or ( n3590 , n3588 , n3589 );
not ( n3591 , n499 );
not ( n3592 , n2118 );
or ( n3593 , n3591 , n3592 );
or ( n3594 , n499 , n2930 );
nand ( n3595 , n3593 , n3594 );
nand ( n3596 , n3595 , n1840 );
nand ( n3597 , n3590 , n3596 );
or ( n3598 , n496 , n497 );
and ( n3599 , n3598 , n3015 );
nand ( n3600 , n496 , n497 );
nand ( n3601 , n3600 , n495 );
nor ( n3602 , n3599 , n3601 );
not ( n3603 , n2259 );
not ( n3604 , n501 );
not ( n3605 , n1970 );
or ( n3606 , n3604 , n3605 );
not ( n3607 , n456 );
not ( n3608 , n482 );
and ( n3609 , n3607 , n3608 );
nor ( n3610 , n3609 , n501 );
nand ( n3611 , n2554 , n456 );
nand ( n73541 , n3610 , n3611 );
nand ( n3616 , n3606 , n73541 );
not ( n3617 , n3616 );
or ( n3618 , n3603 , n3617 );
not ( n3619 , n501 );
not ( n3620 , n2690 );
or ( n3621 , n3619 , n3620 );
not ( n3622 , n3136 );
not ( n3623 , n3135 );
or ( n3624 , n3622 , n3623 );
nand ( n3625 , n3624 , n2261 );
nand ( n3626 , n3621 , n3625 );
nand ( n3627 , n3626 , n2272 );
nand ( n3628 , n3618 , n3627 );
xor ( n3629 , n3602 , n3628 );
xor ( n3630 , n3597 , n3629 );
and ( n3631 , n3063 , n3240 );
not ( n3632 , n504 );
nand ( n3633 , n1706 , n503 );
nand ( n3634 , n2806 , n456 , n464 );
not ( n3635 , n503 );
nand ( n3636 , n3635 , n2202 , n480 );
nand ( n3637 , n3633 , n3634 , n3636 );
not ( n3638 , n3637 );
or ( n3639 , n3632 , n3638 );
not ( n3640 , n503 );
not ( n3641 , n2690 );
or ( n3642 , n3640 , n3641 );
and ( n3643 , n456 , n465 );
not ( n3644 , n456 );
and ( n3645 , n3644 , n481 );
or ( n3646 , n3643 , n3645 );
nand ( n3647 , n3646 , n3635 );
nand ( n3648 , n3642 , n3647 );
nand ( n3649 , n3648 , n3066 );
nand ( n3650 , n3639 , n3649 );
xor ( n3651 , n3631 , n3650 );
not ( n3652 , n1848 );
not ( n3653 , n2351 );
not ( n3654 , n486 );
or ( n3655 , n3653 , n3654 );
nand ( n3656 , n456 , n470 );
nand ( n3657 , n3655 , n3656 );
and ( n3658 , n497 , n3657 );
not ( n3659 , n497 );
and ( n3660 , n456 , n2359 );
not ( n3661 , n456 );
and ( n3662 , n3661 , n2362 );
nor ( n3663 , n3660 , n3662 );
not ( n3664 , n3663 );
and ( n3665 , n3659 , n3664 );
nor ( n73592 , n3658 , n3665 );
not ( n3667 , n73592 );
or ( n3668 , n3652 , n3667 );
not ( n3669 , n497 );
not ( n3670 , n3004 );
or ( n3671 , n3669 , n3670 );
and ( n3672 , n456 , n3557 );
not ( n3673 , n456 );
not ( n3674 , n487 );
and ( n3675 , n3673 , n3674 );
nor ( n3676 , n3672 , n3675 );
nand ( n3677 , n3676 , n3129 );
nand ( n3678 , n3671 , n3677 );
nand ( n3679 , n3678 , n1869 );
nand ( n3680 , n3668 , n3679 );
and ( n3681 , n3651 , n3680 );
and ( n3682 , n3631 , n3650 );
or ( n3683 , n3681 , n3682 );
and ( n3684 , n3630 , n3683 );
and ( n3685 , n3597 , n3629 );
or ( n3686 , n3684 , n3685 );
xor ( n3687 , n3587 , n3686 );
and ( n3688 , n3602 , n3628 );
not ( n3689 , n3142 );
and ( n3690 , n3330 , n497 );
not ( n3691 , n3330 );
and ( n3692 , n3691 , n1760 );
or ( n3693 , n3690 , n3692 );
not ( n3694 , n3693 );
or ( n3695 , n3689 , n3694 );
nand ( n3696 , n1869 , n73592 );
nand ( n3697 , n3695 , n3696 );
not ( n3698 , n1763 );
not ( n3699 , n495 );
not ( n3700 , n3699 );
not ( n3701 , n2841 );
or ( n3702 , n3700 , n3701 );
or ( n3703 , n3699 , n3063 );
nand ( n3704 , n3702 , n3703 );
not ( n3705 , n3704 );
or ( n3706 , n3698 , n3705 );
nand ( n3707 , n2876 , n3562 );
nand ( n3708 , n3706 , n3707 );
xor ( n3709 , n3697 , n3708 );
not ( n3710 , n2421 );
not ( n3711 , n3637 );
or ( n3712 , n3710 , n3711 );
nand ( n3713 , n3568 , n504 );
nand ( n73640 , n3712 , n3713 );
and ( n3718 , n3709 , n73640 );
and ( n3719 , n3697 , n3708 );
or ( n3720 , n3718 , n3719 );
xor ( n3721 , n3688 , n3720 );
not ( n3722 , n488 );
nor ( n3723 , n3722 , n456 );
not ( n3724 , n3723 );
and ( n3725 , n472 , n456 );
not ( n3726 , n3725 );
and ( n3727 , n3724 , n3726 );
nand ( n3728 , n70594 , n494 );
and ( n3729 , n3728 , n2037 );
nor ( n3730 , n3727 , n3729 );
not ( n3731 , n2722 );
not ( n3732 , n3434 );
or ( n3733 , n3731 , n3732 );
nand ( n3734 , n3626 , n2823 );
nand ( n3735 , n3733 , n3734 );
xor ( n3736 , n3730 , n3735 );
not ( n3737 , n1869 );
not ( n3738 , n3693 );
or ( n3739 , n3737 , n3738 );
nand ( n3740 , n3447 , n1848 );
nand ( n3741 , n3739 , n3740 );
xor ( n3742 , n3736 , n3741 );
xor ( n3743 , n3721 , n3742 );
xor ( n3744 , n3687 , n3743 );
not ( n3745 , n3744 );
xor ( n3746 , n3697 , n3708 );
xor ( n3747 , n3746 , n73640 );
not ( n3748 , n2259 );
and ( n3749 , n3579 , n3117 );
not ( n3750 , n3579 );
and ( n3751 , n3750 , n501 );
nor ( n3752 , n3749 , n3751 );
not ( n3753 , n3752 );
or ( n3754 , n3748 , n3753 );
nand ( n3755 , n3616 , n2272 );
nand ( n3756 , n3754 , n3755 );
not ( n3757 , n2167 );
nand ( n3758 , n499 , n2404 );
or ( n3759 , n456 , n485 );
not ( n3760 , n469 );
nand ( n3761 , n3760 , n456 );
nand ( n3762 , n3759 , n3761 , n1380 );
nand ( n3763 , n3758 , n3762 );
not ( n73687 , n3763 );
or ( n3765 , n3757 , n73687 );
nand ( n3766 , n3595 , n2018 );
nand ( n3767 , n3765 , n3766 );
xor ( n3768 , n3756 , n3767 );
nor ( n3769 , n498 , n499 );
not ( n3770 , n3769 );
and ( n3771 , n3770 , n3277 );
not ( n3772 , n498 );
not ( n3773 , n499 );
or ( n3774 , n3772 , n3773 );
nand ( n3775 , n3774 , n497 );
nor ( n3776 , n3771 , n3775 );
not ( n3777 , n504 );
not ( n3778 , n3648 );
or ( n3779 , n3777 , n3778 );
and ( n3780 , n3128 , n503 );
not ( n3781 , n3128 );
not ( n3782 , n503 );
and ( n3783 , n3781 , n3782 );
nor ( n3784 , n3780 , n3783 );
nand ( n3785 , n3784 , n2421 );
nand ( n3786 , n3779 , n3785 );
and ( n3787 , n3776 , n3786 );
and ( n3788 , n3768 , n3787 );
and ( n3789 , n3756 , n3767 );
or ( n3790 , n3788 , n3789 );
xor ( n3791 , n3747 , n3790 );
xor ( n3792 , n3597 , n3629 );
xor ( n3793 , n3792 , n3683 );
and ( n3794 , n3791 , n3793 );
and ( n3795 , n3747 , n3790 );
or ( n3796 , n3794 , n3795 );
not ( n3797 , n3796 );
nand ( n3798 , n3745 , n3797 );
not ( n3799 , n3798 );
xor ( n3800 , n3747 , n3790 );
xor ( n3801 , n3800 , n3793 );
nand ( n3802 , n3769 , n497 );
not ( n3803 , n3802 );
not ( n3804 , n2834 );
or ( n3805 , n3803 , n3804 );
not ( n3806 , n498 );
nor ( n3807 , n3806 , n1380 , n497 );
or ( n73731 , n2834 , n3807 );
nand ( n3812 , n3805 , n73731 );
and ( n3813 , n498 , n1077 );
not ( n3814 , n498 );
and ( n3815 , n3814 , n499 );
or ( n3816 , n3813 , n3815 );
nand ( n3817 , n3816 , n3678 );
nand ( n3818 , n3812 , n3817 );
not ( n3819 , n2259 );
not ( n3820 , n501 );
not ( n3821 , n2930 );
or ( n3822 , n3820 , n3821 );
nand ( n3823 , n2573 , n2261 );
nand ( n3824 , n3822 , n3823 );
not ( n3825 , n3824 );
or ( n3826 , n3819 , n3825 );
nand ( n3827 , n3752 , n3295 );
nand ( n3828 , n3826 , n3827 );
xor ( n3829 , n3818 , n3828 );
not ( n3830 , n1840 );
not ( n3831 , n499 );
and ( n3832 , n456 , n470 );
not ( n3833 , n456 );
and ( n3834 , n3833 , n486 );
nor ( n3835 , n3832 , n3834 );
not ( n3836 , n3835 );
or ( n3837 , n3831 , n3836 );
or ( n3838 , n3835 , n499 );
nand ( n3839 , n3837 , n3838 );
not ( n3840 , n3839 );
or ( n3841 , n3830 , n3840 );
nand ( n3842 , n3763 , n2018 );
nand ( n3843 , n3841 , n3842 );
and ( n3844 , n3829 , n3843 );
and ( n3845 , n3818 , n3828 );
or ( n3846 , n3844 , n3845 );
xor ( n3847 , n3631 , n3650 );
xor ( n3848 , n3847 , n3680 );
xor ( n3849 , n3846 , n3848 );
xor ( n3850 , n3756 , n3767 );
xor ( n3851 , n3850 , n3787 );
and ( n73772 , n3849 , n3851 );
and ( n3853 , n3846 , n3848 );
or ( n3854 , n73772 , n3853 );
nor ( n3855 , n3801 , n3854 );
xor ( n3856 , n3846 , n3848 );
xor ( n3857 , n3856 , n3851 );
xor ( n3858 , n3776 , n3786 );
and ( n3859 , n3063 , n3142 );
not ( n3860 , n504 );
not ( n3861 , n3784 );
or ( n3862 , n3860 , n3861 );
and ( n3863 , n456 , n467 );
not ( n3864 , n456 );
and ( n3865 , n3864 , n483 );
nor ( n3866 , n3863 , n3865 );
and ( n3867 , n3866 , n2269 );
not ( n3868 , n3866 );
and ( n3869 , n3868 , n503 );
nor ( n3870 , n3867 , n3869 );
nand ( n3871 , n3870 , n3066 );
nand ( n3872 , n3862 , n3871 );
xor ( n3873 , n3859 , n3872 );
not ( n3874 , n2259 );
not ( n3875 , n501 );
not ( n3876 , n2411 );
or ( n3877 , n3875 , n3876 );
not ( n3878 , n3323 );
not ( n3879 , n2975 );
or ( n3880 , n3878 , n3879 );
nand ( n3881 , n3880 , n2261 );
nand ( n3882 , n3877 , n3881 );
not ( n3883 , n3882 );
or ( n3884 , n3874 , n3883 );
nand ( n3885 , n3824 , n2272 );
nand ( n3886 , n3884 , n3885 );
and ( n3887 , n3873 , n3886 );
and ( n3888 , n3859 , n3872 );
or ( n3889 , n3887 , n3888 );
xor ( n73810 , n3858 , n3889 );
xor ( n3894 , n3818 , n3828 );
xor ( n3895 , n3894 , n3843 );
and ( n3896 , n73810 , n3895 );
and ( n3897 , n3858 , n3889 );
or ( n3898 , n3896 , n3897 );
nor ( n3899 , n3857 , n3898 );
nor ( n3900 , n3855 , n3899 );
not ( n3901 , n3900 );
xor ( n3902 , n3858 , n3889 );
xor ( n3903 , n3902 , n3895 );
not ( n3904 , n2008 );
xor ( n3905 , n499 , n2488 );
not ( n3906 , n3905 );
or ( n3907 , n3904 , n3906 );
nand ( n3908 , n3839 , n2018 );
nand ( n3909 , n3907 , n3908 );
not ( n3910 , n1836 );
nand ( n3911 , n3910 , n2704 );
nand ( n3912 , n500 , n501 );
and ( n3913 , n3911 , n3912 , n499 );
not ( n3914 , n3066 );
and ( n3915 , n503 , n2118 );
not ( n3916 , n503 );
and ( n3917 , n3916 , n2573 );
or ( n3918 , n3915 , n3917 );
not ( n3919 , n3918 );
or ( n3920 , n3914 , n3919 );
nand ( n3921 , n3870 , n504 );
nand ( n3922 , n3920 , n3921 );
and ( n3923 , n3913 , n3922 );
xor ( n3924 , n3909 , n3923 );
xor ( n3925 , n3859 , n3872 );
xor ( n3926 , n3925 , n3886 );
and ( n3927 , n3924 , n3926 );
and ( n3928 , n3909 , n3923 );
or ( n3929 , n3927 , n3928 );
nor ( n73847 , n3903 , n3929 );
xor ( n3931 , n3909 , n3923 );
xor ( n3932 , n3931 , n3926 );
not ( n3933 , n2259 );
not ( n3934 , n501 );
not ( n3935 , n2988 );
or ( n3936 , n3934 , n3935 );
nand ( n3937 , n2995 , n2261 );
nand ( n3938 , n3936 , n3937 );
not ( n3939 , n3938 );
or ( n3940 , n3933 , n3939 );
nand ( n3941 , n3882 , n3295 );
nand ( n3942 , n3940 , n3941 );
not ( n3943 , n499 );
not ( n3944 , n2793 );
or ( n3945 , n3943 , n3944 );
not ( n3946 , n499 );
nand ( n3947 , n3946 , n2704 );
nand ( n3948 , n3945 , n3947 );
not ( n3949 , n3948 );
not ( n3950 , n2167 );
or ( n3951 , n3949 , n3950 );
nand ( n3952 , n3905 , n2018 );
nand ( n3953 , n3951 , n3952 );
xor ( n3954 , n3942 , n3953 );
xor ( n3955 , n3913 , n3922 );
and ( n3956 , n3954 , n3955 );
and ( n3957 , n3942 , n3953 );
or ( n3958 , n3956 , n3957 );
nor ( n3959 , n3932 , n3958 );
nor ( n3960 , n73847 , n3959 );
and ( n3961 , n2988 , n503 );
and ( n3962 , n3961 , n1636 );
not ( n3963 , n2411 );
not ( n73881 , n2423 );
not ( n3968 , n73881 );
or ( n3969 , n3963 , n3968 );
not ( n3970 , n504 );
nor ( n3971 , n3970 , n503 );
nand ( n3972 , n2977 , n3971 );
nand ( n3973 , n3969 , n3972 );
nor ( n3974 , n3962 , n3973 );
not ( n3975 , n3974 );
not ( n3976 , n502 );
nand ( n3977 , n3976 , n2793 );
and ( n3978 , n3977 , n503 );
not ( n3979 , n502 );
not ( n3980 , n2841 );
or ( n3981 , n3979 , n3980 );
nand ( n3982 , n3981 , n501 );
nor ( n3983 , n3978 , n3982 );
not ( n3984 , n3983 );
and ( n3985 , n3975 , n3984 );
and ( n3986 , n3983 , n3974 );
nor ( n3987 , n3985 , n3986 );
not ( n3988 , n501 );
not ( n3989 , n2650 );
or ( n3990 , n3988 , n3989 );
nand ( n3991 , n2488 , n2261 );
nand ( n3992 , n3990 , n3991 );
not ( n3993 , n3992 );
not ( n3994 , n3993 );
not ( n3995 , n2143 );
and ( n3996 , n3994 , n3995 );
not ( n3997 , n501 );
not ( n73912 , n2834 );
or ( n3999 , n3997 , n73912 );
nand ( n4000 , n3063 , n2261 );
nand ( n4001 , n3999 , n4000 );
and ( n4002 , n4001 , n2502 );
nor ( n4003 , n3996 , n4002 );
nand ( n4004 , n3987 , n4003 );
not ( n4005 , n4004 );
nor ( n4006 , n2704 , n2423 );
not ( n4007 , n4006 );
buf ( n4008 , n3004 );
not ( n4009 , n4008 );
or ( n4010 , n4007 , n4009 );
nand ( n4011 , n2793 , n2421 );
nand ( n4012 , n4010 , n4011 );
and ( n4013 , n3015 , n3295 );
nor ( n4014 , n4012 , n4013 );
not ( n4015 , n2269 );
not ( n4016 , n2364 );
or ( n4017 , n4015 , n4016 );
not ( n4018 , n3961 );
nand ( n4019 , n4017 , n4018 );
and ( n4020 , n4019 , n504 );
not ( n4021 , n4008 );
nor ( n4022 , n4021 , n2420 );
nor ( n4023 , n4020 , n4022 );
or ( n4024 , n4014 , n4023 );
nand ( n4030 , n4024 , C1 );
not ( n4031 , n4030 );
or ( n4032 , n4005 , n4031 );
not ( n4033 , n3987 );
not ( n4034 , n4003 );
nand ( n4035 , n4033 , n4034 );
nand ( n4036 , n4032 , n4035 );
not ( n4037 , n4036 );
and ( n4038 , n1834 , n3277 );
not ( n4039 , n2722 );
not ( n4040 , n3938 );
or ( n4041 , n4039 , n4040 );
nand ( n4042 , n3992 , n2259 );
nand ( n4043 , n4041 , n4042 );
xor ( n4044 , n4038 , n4043 );
not ( n4045 , n2421 );
not ( n4046 , n503 );
not ( n4047 , n2411 );
or ( n4048 , n4046 , n4047 );
not ( n4049 , n503 );
nand ( n4050 , n4049 , n2977 );
nand ( n4051 , n4048 , n4050 );
not ( n4052 , n4051 );
or ( n4053 , n4045 , n4052 );
nand ( n4054 , n504 , n3918 );
nand ( n4055 , n4053 , n4054 );
xor ( n73965 , n4044 , n4055 );
not ( n4057 , n73965 );
and ( n4058 , n2988 , n503 , n1636 );
or ( n4059 , n4058 , n3973 );
nand ( n4060 , n4059 , n3983 );
nand ( n4061 , n4057 , n4060 );
not ( n4062 , n4061 );
or ( n4063 , n4037 , n4062 );
buf ( n4064 , n73965 );
not ( n4065 , n4060 );
nand ( n4066 , n4064 , n4065 );
nand ( n4067 , n4063 , n4066 );
xor ( n4068 , n3942 , n3953 );
xor ( n4069 , n4068 , n3955 );
not ( n4070 , n4069 );
xor ( n4071 , n4038 , n4043 );
and ( n4072 , n4071 , n4055 );
and ( n4073 , n4038 , n4043 );
or ( n4074 , n4072 , n4073 );
not ( n4075 , n4074 );
nand ( n4076 , n4070 , n4075 );
nand ( n4077 , n4067 , n4076 );
buf ( n4078 , n4069 );
nand ( n4079 , n4078 , n4074 );
nand ( n73989 , n3932 , n3958 );
nand ( n4084 , n4077 , n4079 , n73989 );
nand ( n4085 , n3960 , n4084 );
and ( n4086 , n3857 , n3898 );
and ( n4087 , n3903 , n3929 );
nor ( n4088 , n4086 , n4087 );
nand ( n4089 , n4085 , n4088 );
not ( n4090 , n4089 );
or ( n4091 , n3901 , n4090 );
buf ( n4092 , n3801 );
nand ( n4093 , n4092 , n3854 );
nand ( n4094 , n4091 , n4093 );
not ( n4095 , n4094 );
or ( n4096 , n3799 , n4095 );
buf ( n4097 , n3744 );
nand ( n4098 , n4097 , n3796 );
nand ( n4099 , n4096 , n4098 );
xor ( n4100 , n3505 , n3515 );
xor ( n4101 , n4100 , n3517 );
xor ( n4102 , n3730 , n3735 );
and ( n4103 , n4102 , n3741 );
and ( n74010 , n3730 , n3735 );
or ( n4105 , n4103 , n74010 );
xor ( n4106 , n3564 , n3570 );
and ( n4107 , n4106 , n3586 );
and ( n4108 , n3564 , n3570 );
or ( n4109 , n4107 , n4108 );
xor ( n4110 , n4105 , n4109 );
xor ( n4111 , n3449 , n3464 );
xor ( n4112 , n4111 , n3475 );
xor ( n4113 , n4110 , n4112 );
xor ( n4114 , n4101 , n4113 );
xor ( n4115 , n3688 , n3720 );
and ( n4116 , n4115 , n3742 );
and ( n4117 , n3688 , n3720 );
or ( n4118 , n4116 , n4117 );
xor ( n4119 , n4114 , n4118 );
not ( n4120 , n4119 );
xor ( n4121 , n3587 , n3686 );
and ( n74028 , n4121 , n3743 );
and ( n4126 , n3587 , n3686 );
or ( n74030 , n74028 , n4126 );
not ( n74031 , n74030 );
and ( n4129 , n4120 , n74031 );
xor ( n74033 , n3422 , n3437 );
xor ( n74034 , n74033 , n3478 );
xor ( n4132 , n4105 , n4109 );
and ( n74036 , n4132 , n4112 );
and ( n4134 , n4105 , n4109 );
or ( n4135 , n74036 , n4134 );
xor ( n4136 , n74034 , n4135 );
xor ( n74040 , n3490 , n3492 );
xor ( n74041 , n74040 , n3520 );
xor ( n4139 , n4136 , n74041 );
xor ( n74043 , n4101 , n4113 );
and ( n74044 , n74043 , n4118 );
and ( n4142 , n4101 , n4113 );
or ( n74046 , n74044 , n4142 );
nor ( n74047 , n4139 , n74046 );
nor ( n4145 , n4129 , n74047 );
xor ( n4146 , n3488 , n3523 );
xor ( n4147 , n4146 , n3526 );
not ( n74051 , n4147 );
xor ( n74052 , n74034 , n4135 );
and ( n4150 , n74052 , n74041 );
and ( n74054 , n74034 , n4135 );
or ( n4152 , n4150 , n74054 );
not ( n74056 , n4152 );
nand ( n4154 , n74051 , n74056 );
nand ( n4155 , n4099 , n4145 , n4154 );
nand ( n4156 , n4147 , n4152 );
not ( n4157 , n4156 );
nand ( n4158 , n4119 , n74030 );
not ( n74062 , n4158 );
nand ( n4160 , n74046 , n4139 );
not ( n4161 , n4160 );
or ( n4162 , n74062 , n4161 );
not ( n4163 , n4139 );
not ( n74067 , n74046 );
nand ( n4165 , n4163 , n74067 );
nand ( n74069 , n4162 , n4165 );
not ( n4167 , n74069 );
or ( n74071 , n4157 , n4167 );
not ( n4169 , n4147 );
nand ( n4170 , n4169 , n74056 );
nand ( n4171 , n74071 , n4170 );
nand ( n4172 , n4155 , n4171 );
not ( n4173 , n3534 );
nand ( n4174 , n4173 , n3540 );
nand ( n74078 , n3486 , n3530 );
nand ( n4176 , n4172 , n4174 , n74078 );
nand ( n4177 , n3551 , n4176 );
nand ( n4178 , n2971 , n3402 , n4177 );
not ( n4179 , n2783 );
not ( n4180 , n2779 );
and ( n4181 , n4179 , n4180 );
nand ( n4182 , n2750 , n2776 );
or ( n4183 , n4181 , n4182 );
not ( n74087 , n4179 );
not ( n4185 , n4180 );
nand ( n74089 , n74087 , n4185 );
nand ( n4187 , n4183 , n74089 );
not ( n4188 , n4187 );
not ( n4189 , n2750 );
not ( n4190 , n2776 );
and ( n4191 , n4189 , n4190 );
nor ( n4192 , n4191 , n2784 );
and ( n4193 , n2787 , n2967 );
nand ( n4194 , n4192 , n4193 );
nor ( n4195 , n2787 , n2967 );
not ( n4196 , n4195 );
nor ( n4197 , n3390 , n3374 );
nand ( n4198 , n3394 , n3399 );
or ( n4199 , n4197 , n4198 );
nand ( n4200 , n3374 , n3390 );
nand ( n4201 , n4199 , n4200 );
nand ( n4202 , n4196 , n2785 , n4201 );
nand ( n4203 , n4178 , n4188 , n4194 , n4202 );
xor ( n4204 , n2440 , n4203 );
nand ( n4205 , n4204 , n455 );
buf ( n4206 , n3857 );
nor ( n4207 , n4206 , n3898 );
not ( n4208 , n4207 );
buf ( n4209 , n4089 );
nand ( n4210 , n4208 , n4209 );
or ( n4211 , n4092 , n3854 );
nand ( n4212 , n4211 , n4093 );
xor ( n4213 , n4210 , n4212 );
nand ( n4214 , n4213 , n455 );
not ( n4215 , n454 );
and ( n4216 , n539 , n540 );
and ( n4217 , n540 , n541 );
not ( n4218 , n540 );
not ( n4219 , n541 );
and ( n4220 , n4218 , n4219 );
nor ( n4221 , n4217 , n4220 );
nor ( n4222 , n539 , n540 );
nor ( n4223 , n4216 , n4221 , n4222 );
buf ( n4224 , n4223 );
not ( n4225 , n4224 );
not ( n74129 , n539 );
buf ( n74130 , n74078 );
not ( n4228 , n74130 );
nand ( n74132 , n4155 , n4171 );
buf ( n4230 , n74132 );
not ( n74134 , n4230 );
or ( n4232 , n4228 , n74134 );
nand ( n4233 , n3485 , n3529 );
nand ( n4234 , n4232 , n4233 );
not ( n4235 , n4174 );
nand ( n4236 , n3534 , n3539 );
not ( n4237 , n4236 );
nor ( n4238 , n4235 , n4237 );
not ( n4239 , n455 );
nor ( n4240 , n4238 , n4239 );
and ( n4241 , n4234 , n4240 );
not ( n74145 , n4234 );
and ( n4243 , n455 , n4174 , n4236 );
and ( n4244 , n74145 , n4243 );
nor ( n4245 , n4241 , n4244 );
nand ( n4246 , n4245 , n1685 );
buf ( n4247 , n4246 );
not ( n74151 , n4247 );
not ( n4249 , n74151 );
or ( n4250 , n74129 , n4249 );
not ( n4251 , n539 );
nand ( n4252 , n4247 , n4251 );
nand ( n4253 , n4250 , n4252 );
not ( n4254 , n4253 );
or ( n4255 , n4225 , n4254 );
nand ( n4256 , n4236 , n4233 );
not ( n4257 , n4256 );
not ( n4258 , n4174 );
or ( n4259 , n4257 , n4258 );
nand ( n4260 , n4259 , n4176 );
nand ( n4261 , n3369 , n3264 );
buf ( n4262 , n4261 );
nor ( n4263 , n3264 , n3369 );
not ( n4264 , n4263 );
and ( n4265 , n4262 , n4264 );
and ( n4266 , n4260 , n4265 );
not ( n4267 , n455 );
nor ( n4268 , n4266 , n4267 );
not ( n4269 , n4268 );
not ( n4270 , n4260 );
nand ( n4271 , n3372 , n4262 );
nand ( n4272 , n4270 , n4271 );
not ( n74176 , n4272 );
or ( n74177 , n4269 , n74176 );
not ( n4275 , n1682 );
not ( n4276 , n1522 );
or ( n4277 , n4275 , n4276 );
nand ( n4278 , n4277 , n1679 );
not ( n4279 , n1633 );
nand ( n74183 , n4279 , n1655 );
not ( n74184 , n74183 );
not ( n4282 , n1624 );
or ( n74186 , n74184 , n4282 );
not ( n4284 , n1655 );
nand ( n74188 , n4284 , n1633 );
nand ( n4286 , n74186 , n74188 );
not ( n4287 , n1654 );
not ( n4288 , n1557 );
not ( n4289 , n1543 );
or ( n74193 , n4288 , n4289 );
or ( n4291 , n1543 , n1557 );
nand ( n4292 , n4291 , n1532 );
nand ( n4293 , n74193 , n4292 );
xor ( n4294 , n4287 , n4293 );
xor ( n4295 , n1575 , n1585 );
and ( n4296 , n4295 , n1595 );
and ( n4297 , n1575 , n1585 );
or ( n4298 , n4296 , n4297 );
xor ( n4299 , n4294 , n4298 );
xor ( n4300 , n4286 , n4299 );
or ( n74204 , n1596 , n1563 );
nand ( n74205 , n74204 , n1526 );
nand ( n4303 , n1596 , n1563 );
nand ( n4304 , n74205 , n4303 );
xor ( n4305 , n4300 , n4304 );
not ( n4306 , n4305 );
not ( n4307 , n1618 );
not ( n74211 , n4307 );
not ( n4309 , n1659 );
not ( n4310 , n4309 );
or ( n4311 , n74211 , n4310 );
not ( n4312 , n1618 );
not ( n4313 , n1659 );
or ( n4314 , n4312 , n4313 );
nand ( n4315 , n4314 , n1664 );
nand ( n4316 , n4311 , n4315 );
not ( n4317 , n4316 );
not ( n4318 , n4317 );
not ( n4319 , n1573 );
not ( n4320 , n1268 );
or ( n4321 , n4319 , n4320 );
xor ( n4322 , n514 , n493 );
nand ( n4323 , n70491 , n4322 );
nand ( n4324 , n4321 , n4323 );
not ( n4325 , n1593 );
not ( n4326 , n70652 );
or ( n74230 , n4325 , n4326 );
and ( n74231 , n508 , n499 );
not ( n4329 , n508 );
not ( n4330 , n499 );
and ( n4331 , n4329 , n4330 );
nor ( n4332 , n74231 , n4331 );
nand ( n4333 , n70426 , n4332 );
nand ( n4334 , n74230 , n4333 );
xor ( n4335 , n4324 , n4334 );
not ( n4336 , n1631 );
nor ( n4337 , n1626 , n1247 );
not ( n4338 , n4337 );
or ( n4339 , n4336 , n4338 );
xor ( n74243 , n516 , n491 );
nand ( n74244 , n1630 , n74243 );
nand ( n4342 , n4339 , n74244 );
xor ( n4343 , n4335 , n4342 );
not ( n4344 , n1541 );
not ( n4345 , n70413 );
or ( n4346 , n4344 , n4345 );
xor ( n4347 , n506 , n501 );
nand ( n4348 , n4347 , n70371 );
nand ( n4349 , n4346 , n4348 );
nand ( n4350 , n520 , n489 );
not ( n4351 , n70360 );
not ( n4352 , n1640 );
or ( n4353 , n4351 , n4352 );
nand ( n4354 , n4353 , n70376 );
xnor ( n4355 , n4350 , n4354 );
xor ( n4356 , n4349 , n4355 );
not ( n4357 , n4356 );
and ( n4358 , n4343 , n4357 );
not ( n4359 , n4343 );
and ( n4360 , n4359 , n4356 );
nor ( n4361 , n4358 , n4360 );
not ( n4362 , n1555 );
not ( n4363 , n1550 );
nor ( n4364 , n4363 , n1448 );
not ( n4365 , n4364 );
or ( n4366 , n4362 , n4365 );
xor ( n4367 , n518 , n489 );
nand ( n4368 , n1553 , n4367 );
nand ( n4369 , n4366 , n4368 );
not ( n4370 , n1579 );
not ( n4371 , n70536 );
or ( n4372 , n4370 , n4371 );
xor ( n4373 , n512 , n495 );
nand ( n4374 , n70544 , n4373 );
nand ( n4375 , n4372 , n4374 );
xor ( n4376 , n4369 , n4375 );
not ( n4377 , n1530 );
not ( n4378 , n70640 );
or ( n4379 , n4377 , n4378 );
xor ( n4380 , n510 , n497 );
nand ( n4381 , n70513 , n4380 );
nand ( n4382 , n4379 , n4381 );
xor ( n4383 , n4376 , n4382 );
buf ( n74287 , n4383 );
and ( n74288 , n4361 , n74287 );
not ( n4386 , n4361 );
not ( n74290 , n74287 );
and ( n4388 , n4386 , n74290 );
nor ( n74292 , n74288 , n4388 );
not ( n4390 , n74292 );
not ( n4391 , n4390 );
or ( n4392 , n4318 , n4391 );
nand ( n4393 , n4316 , n74292 );
nand ( n74297 , n4392 , n4393 );
not ( n4395 , n74297 );
not ( n4396 , n4395 );
or ( n4397 , n4306 , n4396 );
not ( n4398 , n4305 );
nand ( n4399 , n74297 , n4398 );
nand ( n4400 , n4397 , n4399 );
not ( n4401 , n4400 );
not ( n4402 , n1597 );
not ( n4403 , n1668 );
or ( n74307 , n4402 , n4403 );
not ( n4405 , n1665 );
not ( n4406 , n1597 );
not ( n4407 , n4406 );
or ( n4408 , n4405 , n4407 );
nand ( n4409 , n4408 , n1606 );
nand ( n74313 , n74307 , n4409 );
not ( n4411 , n74313 );
not ( n74315 , n4411 );
and ( n4413 , n4401 , n74315 );
not ( n74317 , n4401 );
and ( n4415 , n74317 , n4411 );
nor ( n4416 , n4413 , n4415 );
not ( n4417 , n4416 );
and ( n4418 , n4278 , n4417 );
not ( n4419 , n4278 );
and ( n74323 , n4419 , n4416 );
nor ( n4421 , n4418 , n74323 );
nand ( n4422 , n4421 , n70470 );
nand ( n4423 , n74177 , n4422 );
not ( n4424 , n4423 );
not ( n4425 , n4424 );
not ( n74329 , n4425 );
not ( n4427 , n4251 );
and ( n74331 , n74329 , n4427 );
buf ( n4429 , n4423 );
and ( n4430 , n4429 , n4251 );
nor ( n4431 , n74331 , n4430 );
not ( n4432 , n4431 );
buf ( n4433 , n4221 );
buf ( n4434 , n4433 );
nand ( n74338 , n4432 , n4434 );
nand ( n4436 , n4255 , n74338 );
xnor ( n4437 , n543 , n544 );
not ( n4438 , n544 );
or ( n4439 , n4438 , n545 );
not ( n4440 , n545 );
or ( n4441 , n4440 , n544 );
nand ( n4442 , n4439 , n4441 );
buf ( n4443 , n4442 );
nor ( n4444 , n4437 , n4443 );
buf ( n4445 , n4444 );
not ( n4446 , n4445 );
not ( n4447 , n543 );
xor ( n4448 , n507 , n499 );
not ( n4449 , n4448 );
not ( n4450 , n70652 );
or ( n4451 , n4449 , n4450 );
and ( n4452 , n506 , n499 );
not ( n4453 , n506 );
and ( n4454 , n4453 , n1864 );
nor ( n4455 , n4452 , n4454 );
nand ( n4456 , n70704 , n4455 );
nand ( n4457 , n4451 , n4456 );
nand ( n4458 , n518 , n489 );
not ( n4459 , n4458 );
and ( n4460 , n4457 , n4459 );
not ( n4461 , n4457 );
and ( n4462 , n4461 , n4458 );
nor ( n4463 , n4460 , n4462 );
xor ( n4464 , n511 , n495 );
not ( n4465 , n4464 );
not ( n4466 , n1028 );
not ( n4467 , n4466 );
or ( n4468 , n4465 , n4467 );
xor ( n4469 , n510 , n495 );
nand ( n4470 , n70544 , n4469 );
nand ( n4471 , n4468 , n4470 );
xor ( n4472 , n4463 , n4471 );
xor ( n4473 , n505 , n501 );
not ( n4474 , n4473 );
not ( n4475 , n70413 );
or ( n4476 , n4474 , n4475 );
nand ( n4477 , n70371 , n501 );
nand ( n4478 , n4476 , n4477 );
xor ( n4479 , n517 , n489 );
not ( n4480 , n4479 );
not ( n4481 , n4364 );
or ( n4482 , n4480 , n4481 );
xor ( n4483 , n516 , n489 );
nand ( n4484 , n1553 , n4483 );
nand ( n4485 , n4482 , n4484 );
and ( n4486 , n4478 , n4485 );
not ( n4487 , n4478 );
not ( n4488 , n4485 );
and ( n4489 , n4487 , n4488 );
or ( n4490 , n4486 , n4489 );
not ( n4491 , n4380 );
not ( n4492 , n70640 );
or ( n4493 , n4491 , n4492 );
xor ( n4494 , n509 , n497 );
nand ( n4495 , n70513 , n4494 );
nand ( n4496 , n4493 , n4495 );
not ( n74400 , n4496 );
and ( n4501 , n4490 , n74400 );
not ( n74402 , n4490 );
and ( n4503 , n74402 , n4496 );
nor ( n74404 , n4501 , n4503 );
not ( n4505 , n74404 );
xor ( n4506 , n4472 , n4505 );
not ( n74407 , n4354 );
nand ( n4508 , n74407 , n4350 );
not ( n4509 , n4508 );
not ( n4513 , n4349 );
or ( n74411 , n4509 , n4513 );
not ( n74412 , n4350 );
nand ( n4516 , n74412 , n4354 );
nand ( n4517 , n74411 , n4516 );
xor ( n4518 , n4324 , n4334 );
and ( n74416 , n4518 , n4342 );
and ( n74417 , n4324 , n4334 );
or ( n4521 , n74416 , n74417 );
xor ( n4522 , n4517 , n4521 );
xor ( n4523 , n4369 , n4375 );
and ( n4524 , n4523 , n4382 );
and ( n4525 , n4369 , n4375 );
or ( n74423 , n4524 , n4525 );
and ( n4527 , n4522 , n74423 );
and ( n4528 , n4517 , n4521 );
or ( n4529 , n4527 , n4528 );
xnor ( n4530 , n4506 , n4529 );
not ( n4531 , n4496 );
not ( n74429 , n1268 );
not ( n74430 , n4322 );
or ( n4534 , n74429 , n74430 );
xor ( n4535 , n513 , n493 );
nand ( n4536 , n70491 , n4535 );
nand ( n74434 , n4534 , n4536 );
not ( n74435 , n74434 );
not ( n4539 , n74243 );
not ( n4540 , n1627 );
or ( n4541 , n4539 , n4540 );
and ( n4542 , n515 , n1693 );
not ( n4543 , n515 );
and ( n4544 , n4543 , n491 );
or ( n4545 , n4542 , n4544 );
nand ( n74443 , n1630 , n4545 );
nand ( n74444 , n4541 , n74443 );
not ( n4548 , n74444 );
not ( n4549 , n4548 );
or ( n4550 , n74435 , n4549 );
or ( n4551 , n4548 , n74434 );
nand ( n4552 , n4550 , n4551 );
not ( n4553 , n4552 );
or ( n4554 , n4531 , n4553 );
or ( n74452 , n4552 , n4496 );
nand ( n74453 , n4554 , n74452 );
not ( n4557 , n74453 );
xor ( n4558 , n4517 , n4521 );
xor ( n4559 , n4558 , n74423 );
not ( n4560 , n4559 );
or ( n4561 , n4557 , n4560 );
or ( n4562 , n74453 , n4559 );
not ( n4563 , n4356 );
not ( n4564 , n4343 );
or ( n4565 , n4563 , n4564 );
or ( n4566 , n4356 , n4343 );
nand ( n74464 , n4566 , n4383 );
nand ( n4568 , n4565 , n74464 );
nand ( n4569 , n4562 , n4568 );
nand ( n4570 , n4561 , n4569 );
not ( n4571 , n4570 );
xor ( n4572 , n4530 , n4571 );
not ( n4573 , n74444 );
not ( n4574 , n74434 );
or ( n4575 , n4573 , n4574 );
not ( n4576 , n4548 );
not ( n74474 , n74434 );
not ( n4578 , n74474 );
or ( n4579 , n4576 , n4578 );
nand ( n4580 , n4579 , n74400 );
nand ( n4581 , n4575 , n4580 );
not ( n4582 , n4581 );
not ( n4583 , n1630 );
xor ( n4584 , n514 , n491 );
not ( n4585 , n4584 );
or ( n4586 , n4583 , n4585 );
xnor ( n4587 , n491 , n492 );
not ( n4588 , n4587 );
not ( n4589 , n1247 );
nand ( n4590 , n4588 , n4545 , n4589 );
nand ( n4591 , n4586 , n4590 );
not ( n74489 , n4591 );
not ( n74490 , n4535 );
not ( n4594 , n1157 );
or ( n4595 , n74490 , n4594 );
xor ( n4596 , n512 , n493 );
nand ( n4597 , n70491 , n4596 );
nand ( n4598 , n4595 , n4597 );
not ( n4599 , n4598 );
and ( n4600 , n74489 , n4599 );
not ( n4601 , n74489 );
and ( n4602 , n4601 , n4598 );
nor ( n4603 , n4600 , n4602 );
not ( n4604 , n4494 );
not ( n4605 , n70640 );
or ( n4606 , n4604 , n4605 );
xor ( n4607 , n508 , n497 );
nand ( n4608 , n70513 , n4607 );
nand ( n74506 , n4606 , n4608 );
xor ( n4610 , n4603 , n74506 );
not ( n4611 , n4610 );
or ( n4612 , n4582 , n4611 );
not ( n4613 , n4610 );
not ( n4614 , n4581 );
nand ( n4615 , n4613 , n4614 );
nand ( n4616 , n4612 , n4615 );
nand ( n4617 , n519 , n489 );
not ( n4618 , n4617 );
not ( n4619 , n503 );
not ( n4620 , n70360 );
or ( n4621 , n4619 , n4620 );
nand ( n4622 , n4621 , n70376 );
not ( n4623 , n4622 );
or ( n74521 , n4618 , n4623 );
not ( n4625 , n4367 );
not ( n4626 , n4364 );
or ( n4627 , n4625 , n4626 );
nand ( n4628 , n1553 , n4479 );
nand ( n4629 , n4627 , n4628 );
nand ( n74527 , n74521 , n4629 );
not ( n4631 , n4622 );
not ( n4632 , n4617 );
nand ( n4633 , n4631 , n4632 );
nand ( n4634 , n74527 , n4633 );
not ( n4635 , n4634 );
not ( n4636 , n4373 );
not ( n4637 , n70536 );
or ( n4638 , n4636 , n4637 );
nand ( n4639 , n70544 , n4464 );
nand ( n4640 , n4638 , n4639 );
not ( n4641 , n4640 );
not ( n4642 , n4448 );
not ( n4643 , n70426 );
or ( n4644 , n4642 , n4643 );
nand ( n4645 , n70611 , n70615 , n4332 , n70614 );
nand ( n74543 , n4644 , n4645 );
not ( n4647 , n74543 );
or ( n4648 , n4641 , n4647 );
not ( n4649 , n4640 );
not ( n4650 , n4649 );
not ( n4651 , n74543 );
not ( n4652 , n4651 );
or ( n4653 , n4650 , n4652 );
not ( n4654 , n4347 );
not ( n4655 , n70413 );
or ( n4656 , n4654 , n4655 );
nand ( n74554 , n70371 , n4473 );
nand ( n4661 , n4656 , n74554 );
nand ( n74556 , n4653 , n4661 );
nand ( n4663 , n4648 , n74556 );
not ( n4664 , n4663 );
not ( n4665 , n4664 );
or ( n74560 , n4635 , n4665 );
not ( n4670 , n4634 );
nand ( n4671 , n4670 , n4663 );
nand ( n4672 , n74560 , n4671 );
and ( n74564 , n4616 , n4672 );
not ( n74565 , n4616 );
not ( n4675 , n4672 );
and ( n4676 , n74565 , n4675 );
nor ( n4677 , n74564 , n4676 );
xor ( n4678 , n4632 , n4622 );
xnor ( n4679 , n4678 , n4629 );
not ( n4680 , n4651 );
not ( n74572 , n4649 );
nand ( n74573 , n4680 , n74572 , n4661 );
not ( n4683 , n4661 );
nand ( n4684 , n74572 , n4683 , n4651 );
not ( n4685 , n4651 );
not ( n4686 , n4640 );
nand ( n74578 , n4685 , n4686 , n4683 );
nand ( n4688 , n4686 , n4651 , n4661 );
nand ( n4689 , n74573 , n4684 , n74578 , n4688 );
or ( n4690 , n4679 , n4689 );
not ( n4691 , n4690 );
xor ( n4692 , n4287 , n4293 );
and ( n4693 , n4692 , n4298 );
and ( n74585 , n4287 , n4293 );
or ( n74586 , n4693 , n74585 );
not ( n4696 , n74586 );
or ( n4697 , n4691 , n4696 );
nand ( n4698 , n4679 , n4689 );
nand ( n4699 , n4697 , n4698 );
and ( n74591 , n4677 , n4699 );
not ( n74592 , n4677 );
not ( n4702 , n4699 );
and ( n4703 , n74592 , n4702 );
nor ( n4704 , n74591 , n4703 );
xor ( n4705 , n4572 , n4704 );
or ( n4706 , n4679 , n4689 );
nand ( n4707 , n4706 , n4698 );
not ( n74599 , n4707 );
not ( n74600 , n74586 );
and ( n4710 , n74599 , n74600 );
and ( n4711 , n74586 , n4707 );
nor ( n4712 , n4710 , n4711 );
not ( n4713 , n4712 );
not ( n4714 , n4713 );
xor ( n4715 , n74453 , n4568 );
xnor ( n74607 , n4715 , n4559 );
not ( n4717 , n74607 );
not ( n4718 , n4717 );
or ( n4719 , n4714 , n4718 );
not ( n4720 , n4712 );
not ( n4721 , n74607 );
or ( n4722 , n4720 , n4721 );
xor ( n74614 , n4286 , n4299 );
and ( n4724 , n74614 , n4304 );
and ( n4725 , n4286 , n4299 );
or ( n4726 , n4724 , n4725 );
buf ( n4727 , n4726 );
nand ( n4728 , n4722 , n4727 );
nand ( n74620 , n4719 , n4728 );
not ( n4730 , n74620 );
nand ( n4731 , n4705 , n4730 );
not ( n4732 , n4731 );
not ( n4733 , n4712 );
not ( n4734 , n4726 );
or ( n4735 , n4733 , n4734 );
not ( n4736 , n4726 );
nand ( n4737 , n4736 , n4713 );
nand ( n4738 , n4735 , n4737 );
or ( n4739 , n4717 , n4738 );
nand ( n4740 , n4738 , n4717 );
nand ( n4741 , n4739 , n4740 );
not ( n4742 , n4398 );
buf ( n4743 , n74292 );
not ( n4744 , n4743 );
and ( n4745 , n4742 , n4744 );
nand ( n4746 , n4398 , n4743 );
buf ( n4747 , n4316 );
and ( n4748 , n4746 , n4747 );
nor ( n4749 , n4745 , n4748 );
nand ( n4750 , n4741 , n4749 );
not ( n4751 , n4750 );
not ( n4752 , n1680 );
not ( n4753 , n1681 );
or ( n4754 , n4752 , n4753 );
or ( n4755 , n74297 , n4398 );
nand ( n4756 , n4755 , n4399 );
not ( n4757 , n4756 );
not ( n4758 , n74313 );
nand ( n4759 , n4757 , n4758 );
nand ( n4760 , n4754 , n4759 );
nor ( n4761 , n4751 , n4760 );
not ( n4762 , n4761 );
not ( n4763 , n1522 );
or ( n4764 , n4762 , n4763 );
or ( n4765 , n4741 , n4749 );
nand ( n4766 , n4401 , n4758 );
not ( n4767 , n74313 );
not ( n74659 , n4756 );
or ( n74660 , n4767 , n74659 );
nand ( n4770 , n74660 , n1678 );
nand ( n4771 , n4750 , n4766 , n4770 );
nand ( n4772 , n4765 , n4771 );
not ( n4773 , n4772 );
nand ( n4774 , n4764 , n4773 );
not ( n4775 , n4774 );
or ( n4776 , n4732 , n4775 );
not ( n4777 , n4705 );
nand ( n4778 , n4777 , n74620 );
nand ( n4779 , n4776 , n4778 );
not ( n74671 , n455 );
not ( n4781 , n74671 );
not ( n4782 , n4485 );
nand ( n4783 , n4782 , n4478 );
not ( n4784 , n4783 );
not ( n4785 , n4496 );
or ( n4786 , n4784 , n4785 );
not ( n4787 , n4478 );
nand ( n4788 , n4787 , n4485 );
nand ( n4789 , n4786 , n4788 );
not ( n4790 , n4596 );
not ( n4791 , n1268 );
or ( n4792 , n4790 , n4791 );
and ( n4793 , n493 , n1261 );
not ( n4794 , n493 );
and ( n4795 , n4794 , n511 );
or ( n4796 , n4793 , n4795 );
nand ( n4797 , n70491 , n4796 );
nand ( n4798 , n4792 , n4797 );
nand ( n4799 , n517 , n489 );
xor ( n4800 , n4798 , n4799 );
not ( n4801 , n70513 );
xor ( n4802 , n497 , n507 );
not ( n4803 , n4802 );
or ( n4804 , n4801 , n4803 );
nand ( n4805 , n4607 , n70640 );
nand ( n4806 , n4804 , n4805 );
xnor ( n4807 , n4800 , n4806 );
xor ( n4808 , n4789 , n4807 );
not ( n4809 , n4584 );
not ( n74701 , n1627 );
or ( n4811 , n4809 , n74701 );
xor ( n4812 , n491 , n513 );
nand ( n4813 , n1630 , n4812 );
nand ( n4814 , n4811 , n4813 );
not ( n4815 , n4483 );
not ( n74707 , n4364 );
or ( n4817 , n4815 , n74707 );
xor ( n4818 , n515 , n489 );
nand ( n4819 , n1553 , n4818 );
nand ( n4820 , n4817 , n4819 );
xnor ( n4821 , n4814 , n4820 );
and ( n4822 , n4821 , n4787 );
not ( n4823 , n4821 );
and ( n4824 , n4823 , n4478 );
nor ( n4825 , n4822 , n4824 );
xor ( n4826 , n4808 , n4825 );
xnor ( n74718 , n4672 , n4610 );
nand ( n4828 , n74718 , n4614 );
not ( n4829 , n4828 );
not ( n4830 , n4699 );
or ( n4831 , n4829 , n4830 );
not ( n4832 , n74718 );
nand ( n4833 , n4832 , n4581 );
nand ( n4834 , n4831 , n4833 );
xor ( n4835 , n4826 , n4834 );
not ( n4836 , n4670 );
not ( n4837 , n4664 );
or ( n4838 , n4836 , n4837 );
nand ( n4839 , n4838 , n4610 );
nand ( n4840 , n4663 , n4634 );
nand ( n4841 , n4839 , n4840 );
not ( n4842 , n74506 );
nand ( n4843 , n4599 , n74489 );
not ( n4844 , n4843 );
or ( n4845 , n4842 , n4844 );
nand ( n4846 , n4591 , n4598 );
nand ( n4847 , n4845 , n4846 );
or ( n4848 , n4457 , n4459 );
nand ( n4849 , n4848 , n4471 );
nand ( n4850 , n4457 , n4459 );
nand ( n4851 , n4849 , n4850 );
not ( n4852 , n4851 );
and ( n4853 , n4847 , n4852 );
not ( n4854 , n4847 );
and ( n4855 , n4854 , n4851 );
or ( n4856 , n4853 , n4855 );
not ( n74748 , n70704 );
and ( n4861 , n499 , n505 );
not ( n74750 , n499 );
not ( n4863 , n505 );
and ( n4864 , n74750 , n4863 );
nor ( n74753 , n4861 , n4864 );
not ( n4866 , n74753 );
or ( n4867 , n74748 , n4866 );
nand ( n4868 , n4455 , n70650 , n1376 );
nand ( n4869 , n4867 , n4868 );
not ( n4870 , n4869 );
not ( n4871 , n70411 );
nand ( n4872 , n4871 , n70478 , n70479 );
nand ( n74761 , n4872 , n501 );
and ( n4877 , n4870 , n74761 );
not ( n4878 , n4870 );
not ( n4879 , n74761 );
and ( n74765 , n4878 , n4879 );
nor ( n74766 , n4877 , n74765 );
not ( n4882 , n4469 );
not ( n4883 , n70536 );
or ( n4884 , n4882 , n4883 );
xor ( n4885 , n509 , n495 );
nand ( n4886 , n70544 , n4885 );
nand ( n4887 , n4884 , n4886 );
xor ( n74773 , n74766 , n4887 );
not ( n74774 , n74773 );
and ( n4890 , n4856 , n74774 );
not ( n4891 , n4856 );
and ( n4892 , n4891 , n74773 );
nor ( n4893 , n4890 , n4892 );
xor ( n74779 , n4841 , n4893 );
not ( n4895 , n4472 );
nand ( n4896 , n74404 , n4895 );
not ( n4897 , n4896 );
not ( n4898 , n4529 );
or ( n4899 , n4897 , n4898 );
not ( n4900 , n4895 );
nand ( n4901 , n4900 , n4505 );
nand ( n4902 , n4899 , n4901 );
xor ( n4903 , n74779 , n4902 );
xnor ( n4904 , n4835 , n4903 );
not ( n4905 , n4904 );
xor ( n4906 , n4530 , n4571 );
and ( n4907 , n4906 , n4704 );
and ( n4908 , n4530 , n4571 );
or ( n4909 , n4907 , n4908 );
not ( n4910 , n4909 );
xnor ( n4911 , n4905 , n4910 );
nor ( n4912 , n4781 , n4911 );
and ( n4913 , n4779 , n4912 );
not ( n74799 , n4779 );
and ( n74800 , n4911 , n4267 );
and ( n4916 , n74799 , n74800 );
nor ( n4917 , n4913 , n4916 );
not ( n4918 , n4177 );
not ( n4919 , n3402 );
or ( n4920 , n4918 , n4919 );
not ( n74806 , n4201 );
nand ( n74807 , n4920 , n74806 );
not ( n4923 , n4193 );
and ( n4924 , n2969 , n4923 , n455 );
and ( n4925 , n74807 , n4924 );
not ( n4926 , n74807 );
not ( n4927 , n4193 );
nand ( n4928 , n4927 , n2969 );
not ( n74814 , n4928 );
nor ( n74815 , n74814 , n4267 );
and ( n4931 , n4926 , n74815 );
nor ( n4932 , n4925 , n4931 );
nand ( n4933 , n4917 , n4932 );
not ( n4934 , n4933 );
or ( n4935 , n4447 , n4934 );
nand ( n4936 , n4917 , n4932 );
not ( n4937 , n4936 );
not ( n4938 , n543 );
nand ( n4939 , n4937 , n4938 );
nand ( n4940 , n4935 , n4939 );
not ( n4941 , n4940 );
or ( n4942 , n4446 , n4941 );
not ( n4943 , n543 );
nand ( n4944 , n4904 , n4909 );
nand ( n4945 , n4944 , n4731 );
not ( n4946 , n4945 );
not ( n4947 , n4946 );
and ( n4948 , n1522 , n4761 );
not ( n74834 , n4948 );
or ( n4950 , n4947 , n74834 );
buf ( n4951 , n4772 );
and ( n4952 , n4951 , n4946 );
not ( n4953 , n4910 );
not ( n4954 , n4905 );
or ( n4955 , n4953 , n4954 );
not ( n4956 , n4909 );
not ( n4957 , n4904 );
or ( n4958 , n4956 , n4957 );
nor ( n4959 , n4705 , n4730 );
nand ( n4960 , n4958 , n4959 );
nand ( n4961 , n4955 , n4960 );
nor ( n4962 , n4952 , n4961 );
nand ( n4963 , n4950 , n4962 );
not ( n74849 , n4963 );
xor ( n4965 , n4789 , n4807 );
and ( n4966 , n4965 , n4825 );
and ( n4967 , n4789 , n4807 );
or ( n4968 , n4966 , n4967 );
not ( n4969 , n74753 );
not ( n4970 , n699 );
or ( n4971 , n4969 , n4970 );
nand ( n4972 , n70655 , n499 );
nand ( n4973 , n4971 , n4972 );
not ( n74859 , n4973 );
not ( n4975 , n4879 );
not ( n4976 , n4870 );
or ( n4977 , n4975 , n4976 );
nand ( n4978 , n4977 , n4887 );
nand ( n4979 , n74761 , n4869 );
nand ( n4980 , n4978 , n4979 );
xor ( n4981 , n74859 , n4980 );
not ( n4982 , n4798 );
nand ( n4983 , n4982 , n4799 );
not ( n4984 , n4983 );
not ( n4985 , n4806 );
or ( n4986 , n4984 , n4985 );
not ( n4987 , n4799 );
nand ( n4988 , n4798 , n4987 );
nand ( n4989 , n4986 , n4988 );
xor ( n4990 , n4981 , n4989 );
not ( n4991 , n4851 );
not ( n4992 , n74774 );
or ( n4993 , n4991 , n4992 );
not ( n4994 , n74773 );
not ( n4995 , n4852 );
or ( n4996 , n4994 , n4995 );
nand ( n74882 , n4996 , n4847 );
nand ( n74883 , n4993 , n74882 );
xor ( n4999 , n4990 , n74883 );
and ( n5000 , n516 , n489 );
not ( n5001 , n4818 );
not ( n5002 , n1550 );
nor ( n5003 , n5002 , n1448 );
not ( n5004 , n5003 );
or ( n5005 , n5001 , n5004 );
xor ( n5006 , n514 , n489 );
nand ( n5007 , n1448 , n5006 );
nand ( n5008 , n5005 , n5007 );
xor ( n5009 , n5000 , n5008 );
not ( n5010 , n4885 );
not ( n5011 , n4466 );
or ( n5012 , n5010 , n5011 );
xor ( n5013 , n508 , n495 );
nand ( n5014 , n70544 , n5013 );
nand ( n5015 , n5012 , n5014 );
xor ( n5016 , n5009 , n5015 );
not ( n5017 , n4812 );
not ( n5018 , n1627 );
or ( n74904 , n5017 , n5018 );
xor ( n5020 , n512 , n491 );
nand ( n5021 , n1630 , n5020 );
nand ( n5022 , n74904 , n5021 );
buf ( n5023 , n5022 );
not ( n5024 , n4802 );
not ( n5025 , n70509 );
or ( n5026 , n5024 , n5025 );
and ( n5027 , n506 , n497 );
not ( n5028 , n506 );
and ( n5029 , n5028 , n1760 );
nor ( n5030 , n5027 , n5029 );
nand ( n5031 , n70513 , n5030 );
nand ( n5032 , n5026 , n5031 );
not ( n5033 , n5032 );
not ( n5034 , n4796 );
not ( n74920 , n71126 );
or ( n5036 , n5034 , n74920 );
not ( n5037 , n991 );
xor ( n5038 , n510 , n493 );
nand ( n5039 , n5037 , n5038 );
nand ( n5040 , n5036 , n5039 );
not ( n74926 , n5040 );
or ( n5042 , n5033 , n74926 );
or ( n5043 , n5040 , n5032 );
nand ( n5044 , n5042 , n5043 );
and ( n5045 , n5023 , n5044 );
not ( n5046 , n5023 );
not ( n5047 , n5040 );
not ( n5048 , n5032 );
not ( n5049 , n5048 );
or ( n5050 , n5047 , n5049 );
not ( n5051 , n4796 );
not ( n5052 , n71126 );
or ( n5053 , n5051 , n5052 );
nand ( n5054 , n5053 , n5039 );
not ( n5055 , n5032 );
or ( n5056 , n5054 , n5055 );
nand ( n5057 , n5050 , n5056 );
and ( n5058 , n5046 , n5057 );
nor ( n5059 , n5045 , n5058 );
xor ( n5060 , n5016 , n5059 );
not ( n5061 , n4814 );
not ( n74947 , n4820 );
or ( n5063 , n5061 , n74947 );
or ( n5064 , n4820 , n4814 );
nand ( n5065 , n5064 , n4478 );
nand ( n5066 , n5063 , n5065 );
xnor ( n5067 , n5060 , n5066 );
xor ( n5068 , n4999 , n5067 );
xor ( n5069 , n4968 , n5068 );
xor ( n5070 , n4841 , n4893 );
and ( n5071 , n5070 , n4902 );
and ( n5072 , n4841 , n4893 );
or ( n5073 , n5071 , n5072 );
xor ( n5074 , n5069 , n5073 );
not ( n5075 , n4826 );
not ( n5076 , n4903 );
or ( n5077 , n5075 , n5076 );
or ( n74963 , n4903 , n4826 );
not ( n5082 , n4828 );
not ( n74965 , n4699 );
or ( n5084 , n5082 , n74965 );
nand ( n5085 , n5084 , n4833 );
nand ( n5086 , n74963 , n5085 );
nand ( n5087 , n5077 , n5086 );
nand ( n74970 , n5074 , n5087 );
not ( n5089 , n5074 );
not ( n5090 , n5087 );
nand ( n5091 , n5089 , n5090 );
nand ( n5092 , n74970 , n5091 );
not ( n5093 , n5092 );
nand ( n5094 , n74849 , n5093 );
nand ( n5095 , n4963 , n5092 );
not ( n5096 , n455 );
nand ( n5097 , n5094 , n5095 , n5096 );
not ( n5098 , n3394 );
nand ( n5099 , n5098 , n3400 );
nand ( n74982 , n5099 , n3371 );
not ( n5104 , n74982 );
and ( n5105 , n2969 , n5104 , n3392 );
nand ( n5106 , n5105 , n4177 );
and ( n5107 , n4201 , n2969 );
nor ( n5108 , n5107 , n4193 );
nand ( n5109 , n5106 , n5108 );
not ( n5110 , n5109 );
nand ( n74990 , n2776 , n2750 );
or ( n74991 , n2750 , n2776 );
nand ( n5113 , n74990 , n74991 );
and ( n5114 , n5113 , n455 );
nand ( n5115 , n5110 , n5114 );
not ( n5116 , n5113 );
nand ( n5117 , n5116 , n5109 , n455 );
nand ( n5118 , n5097 , n5115 , n5117 );
not ( n74998 , n5118 );
not ( n74999 , n74998 );
not ( n5121 , n74999 );
or ( n5122 , n4943 , n5121 );
nand ( n5123 , n5097 , n5115 , n5117 );
not ( n5124 , n5123 );
nand ( n5125 , n5124 , n4938 );
nand ( n5126 , n5122 , n5125 );
buf ( n5127 , n4443 );
buf ( n5128 , n5127 );
nand ( n5129 , n5126 , n5128 );
nand ( n75009 , n4942 , n5129 );
xor ( n5131 , n4436 , n75009 );
xor ( n5132 , n546 , n547 );
not ( n5133 , n5132 );
and ( n5134 , n545 , n546 );
nor ( n5135 , n545 , n546 );
nor ( n5136 , n5134 , n5135 );
and ( n5137 , n5133 , n5136 );
not ( n75017 , n5137 );
not ( n75018 , n75017 );
not ( n5140 , n75018 );
not ( n5141 , n545 );
not ( n5142 , n455 );
not ( n5143 , n74990 );
not ( n5144 , n74991 );
not ( n5145 , n5144 );
or ( n5146 , n5143 , n5145 );
not ( n5147 , n4181 );
nand ( n5148 , n74087 , n4185 );
nand ( n5149 , n5147 , n5148 );
nand ( n75029 , n5146 , n5149 );
not ( n75030 , n75029 );
not ( n5152 , n75030 );
nand ( n5153 , n5108 , n5106 , n74990 );
not ( n5154 , n5153 );
or ( n5155 , n5152 , n5154 );
not ( n5156 , n74991 );
not ( n5157 , n5109 );
or ( n75037 , n5156 , n5157 );
not ( n75038 , n74990 );
nor ( n5160 , n75038 , n5149 );
nand ( n5161 , n75037 , n5160 );
nand ( n5162 , n5155 , n5161 );
not ( n5163 , n5162 );
or ( n5164 , n5142 , n5163 );
not ( n5165 , n5091 );
not ( n5166 , n4946 );
not ( n5167 , n4948 );
or ( n5168 , n5166 , n5167 );
nand ( n75048 , n5168 , n4962 );
not ( n5170 , n75048 );
or ( n5171 , n5165 , n5170 );
nand ( n5172 , n5171 , n74970 );
xor ( n5173 , n4968 , n5068 );
and ( n5174 , n5173 , n5073 );
and ( n5175 , n4968 , n5068 );
or ( n5176 , n5174 , n5175 );
xor ( n5177 , n5000 , n5008 );
and ( n5178 , n5177 , n5015 );
and ( n5179 , n5000 , n5008 );
or ( n5180 , n5178 , n5179 );
not ( n5181 , n5180 );
not ( n5182 , n5006 );
not ( n5183 , n4364 );
or ( n5184 , n5182 , n5183 );
xor ( n5185 , n513 , n489 );
nand ( n5186 , n1553 , n5185 );
nand ( n5187 , n5184 , n5186 );
not ( n5188 , n5013 );
not ( n5189 , n4466 );
or ( n5190 , n5188 , n5189 );
xor ( n5191 , n507 , n495 );
nand ( n5192 , n70544 , n5191 );
nand ( n5193 , n5190 , n5192 );
xor ( n75073 , n5187 , n5193 );
not ( n5195 , n5020 );
not ( n5196 , n1627 );
or ( n5197 , n5195 , n5196 );
xor ( n5198 , n511 , n491 );
nand ( n5199 , n1630 , n5198 );
nand ( n5200 , n5197 , n5199 );
xor ( n5201 , n75073 , n5200 );
xor ( n5202 , n5181 , n5201 );
or ( n5203 , n70655 , n699 );
nand ( n75083 , n5203 , n499 );
not ( n5205 , n5038 );
not ( n5206 , n1157 );
or ( n5207 , n5205 , n5206 );
xor ( n5208 , n509 , n493 );
nand ( n5209 , n992 , n5208 );
nand ( n5210 , n5207 , n5209 );
xor ( n5211 , n75083 , n5210 );
not ( n5212 , n5030 );
not ( n5213 , n70640 );
or ( n5214 , n5212 , n5213 );
xor ( n5215 , n497 , n505 );
nand ( n5216 , n70513 , n5215 );
nand ( n5217 , n5214 , n5216 );
xor ( n5218 , n5211 , n5217 );
xnor ( n5219 , n5202 , n5218 );
not ( n5220 , n5040 );
not ( n5221 , n5022 );
or ( n5222 , n5220 , n5221 );
or ( n5223 , n5022 , n5040 );
nand ( n5224 , n5223 , n5032 );
nand ( n5225 , n5222 , n5224 );
nand ( n5226 , n515 , n489 );
and ( n5227 , n5226 , n74859 );
not ( n5228 , n5226 );
and ( n5229 , n5228 , n4973 );
nor ( n5230 , n5227 , n5229 );
xor ( n5231 , n5225 , n5230 );
xor ( n5232 , n74859 , n4980 );
and ( n5233 , n5232 , n4989 );
and ( n5234 , n74859 , n4980 );
or ( n5235 , n5233 , n5234 );
xor ( n5236 , n5231 , n5235 );
not ( n5237 , n5016 );
not ( n5238 , n5237 );
not ( n5239 , n5066 );
not ( n5240 , n5239 );
or ( n5241 , n5238 , n5240 );
not ( n5242 , n5059 );
nand ( n5243 , n5241 , n5242 );
not ( n5244 , n5237 );
nand ( n75124 , n5244 , n5066 );
nand ( n75125 , n5243 , n75124 );
xor ( n5247 , n5236 , n75125 );
xor ( n5248 , n5219 , n5247 );
xor ( n5249 , n4990 , n74883 );
and ( n5250 , n5249 , n5067 );
and ( n5251 , n4990 , n74883 );
or ( n5252 , n5250 , n5251 );
xor ( n5253 , n5248 , n5252 );
or ( n5254 , n5176 , n5253 );
nand ( n5255 , n5176 , n5253 );
nand ( n5256 , n5254 , n5255 );
not ( n5257 , n5256 );
and ( n5258 , n5172 , n5257 );
not ( n5259 , n5172 );
and ( n5260 , n5259 , n5256 );
nor ( n5261 , n5258 , n5260 );
nand ( n75141 , n5261 , n70470 );
nand ( n5263 , n5164 , n75141 );
buf ( n5264 , n5263 );
not ( n5265 , n5264 );
not ( n5266 , n5265 );
or ( n5267 , n5141 , n5266 );
not ( n5268 , n545 );
nand ( n5269 , n5268 , n5264 );
nand ( n5270 , n5267 , n5269 );
not ( n5271 , n5270 );
or ( n5272 , n5140 , n5271 );
not ( n5273 , n545 );
not ( n5274 , n70470 );
xor ( n5275 , n5187 , n5193 );
and ( n5276 , n5275 , n5200 );
and ( n5277 , n5187 , n5193 );
or ( n5278 , n5276 , n5277 );
not ( n5279 , n5185 );
not ( n5280 , n5003 );
or ( n5281 , n5279 , n5280 );
xor ( n5282 , n512 , n489 );
nand ( n5283 , n1448 , n5282 );
nand ( n5284 , n5281 , n5283 );
not ( n5285 , n5198 );
nor ( n5286 , n4587 , n1247 );
not ( n5287 , n5286 );
or ( n5288 , n5285 , n5287 );
xor ( n5289 , n510 , n491 );
nand ( n5290 , n1129 , n5289 );
nand ( n5291 , n5288 , n5290 );
xor ( n5292 , n5284 , n5291 );
not ( n75172 , n70509 );
not ( n5294 , n75172 );
and ( n5295 , n5294 , n5215 );
and ( n5296 , n70513 , n497 );
nor ( n5297 , n5295 , n5296 );
xnor ( n5298 , n5292 , n5297 );
xor ( n75178 , n5278 , n5298 );
xor ( n5300 , n75083 , n5210 );
and ( n5301 , n5300 , n5217 );
and ( n5302 , n75083 , n5210 );
or ( n5303 , n5301 , n5302 );
xor ( n5304 , n75178 , n5303 );
xor ( n5305 , n5231 , n5235 );
and ( n5306 , n5305 , n75125 );
and ( n5307 , n5231 , n5235 );
or ( n5308 , n5306 , n5307 );
xor ( n5309 , n5304 , n5308 );
not ( n5310 , n5180 );
not ( n5311 , n5201 );
or ( n5312 , n5310 , n5311 );
not ( n5313 , n5181 );
not ( n5314 , n5201 );
not ( n75194 , n5314 );
or ( n5316 , n5313 , n75194 );
nand ( n5317 , n5316 , n5218 );
nand ( n5318 , n5312 , n5317 );
nand ( n5319 , n514 , n489 );
not ( n5320 , n5191 );
not ( n5321 , n70536 );
or ( n5322 , n5320 , n5321 );
xor ( n5323 , n506 , n495 );
nand ( n5324 , n70544 , n5323 );
nand ( n5325 , n5322 , n5324 );
xor ( n5326 , n5319 , n5325 );
xor ( n5327 , n508 , n493 );
and ( n5328 , n5327 , n992 );
not ( n5329 , n5208 );
not ( n5330 , n1157 );
nor ( n5331 , n5329 , n5330 );
nor ( n5332 , n5328 , n5331 );
xor ( n5333 , n5326 , n5332 );
not ( n5334 , n5333 );
nand ( n5335 , n74859 , n5226 );
not ( n5336 , n5335 );
not ( n5337 , n5225 );
or ( n5338 , n5336 , n5337 );
or ( n5339 , n74859 , n5226 );
nand ( n5340 , n5338 , n5339 );
not ( n5341 , n5340 );
not ( n5342 , n5341 );
or ( n5343 , n5334 , n5342 );
not ( n5344 , n5333 );
nand ( n5345 , n5344 , n5340 );
nand ( n5346 , n5343 , n5345 );
not ( n5347 , n5346 );
and ( n5348 , n5318 , n5347 );
not ( n5349 , n5318 );
and ( n75229 , n5349 , n5346 );
nor ( n5354 , n5348 , n75229 );
xor ( n75231 , n5309 , n5354 );
not ( n5356 , n75231 );
xor ( n5357 , n5219 , n5247 );
and ( n5358 , n5357 , n5252 );
and ( n5359 , n5219 , n5247 );
or ( n5360 , n5358 , n5359 );
not ( n5361 , n5360 );
nand ( n5362 , n5356 , n5361 );
and ( n5363 , n5360 , n75231 );
not ( n5364 , n5363 );
nand ( n5365 , n5362 , n5364 );
not ( n75242 , n4761 );
not ( n5370 , n1522 );
or ( n5371 , n75242 , n5370 );
nand ( n5372 , n5371 , n4773 );
not ( n5373 , n5372 );
and ( n5374 , n4944 , n5254 , n5091 , n4731 );
not ( n5375 , n5374 );
or ( n5376 , n5373 , n5375 );
not ( n75250 , n5087 );
not ( n75251 , n5074 );
and ( n5379 , n75250 , n75251 );
nor ( n5380 , n5176 , n5253 );
nor ( n5381 , n5379 , n5380 );
and ( n5382 , n4961 , n5381 );
or ( n5383 , n74970 , n5380 );
nand ( n5384 , n5383 , n5255 );
buf ( n75258 , n5384 );
nor ( n75259 , n5382 , n75258 );
nand ( n5387 , n5376 , n75259 );
xnor ( n5388 , n5365 , n5387 );
not ( n5389 , n5388 );
or ( n5390 , n5274 , n5389 );
nand ( n5391 , n5390 , n4205 );
buf ( n5392 , n5391 );
not ( n5393 , n5392 );
not ( n5394 , n5393 );
or ( n5395 , n5273 , n5394 );
nand ( n5396 , n5392 , n4440 );
nand ( n75270 , n5395 , n5396 );
buf ( n5398 , n5132 );
buf ( n5399 , n5398 );
nand ( n5400 , n75270 , n5399 );
nand ( n5401 , n5272 , n5400 );
xor ( n5402 , n5131 , n5401 );
not ( n5403 , n538 );
not ( n5404 , n5403 );
not ( n5405 , n539 );
and ( n5406 , n5404 , n5405 );
nor ( n5407 , n4251 , n538 );
nor ( n5408 , n5406 , n5407 );
not ( n5409 , n537 );
and ( n5410 , n5403 , n5409 );
and ( n5411 , n537 , n538 );
nor ( n5412 , n5410 , n5411 );
and ( n5413 , n5408 , n5412 );
not ( n5414 , n5413 );
not ( n5415 , n537 );
not ( n5416 , n70470 );
not ( n75290 , n1507 );
nand ( n75291 , n75290 , n1222 );
not ( n5419 , n695 );
not ( n5420 , n979 );
or ( n5421 , n5419 , n5420 );
nand ( n5422 , n5421 , n989 );
not ( n5423 , n5422 );
not ( n75297 , n5423 );
and ( n75298 , n75291 , n75297 );
not ( n5426 , n75291 );
and ( n5427 , n5426 , n5423 );
nor ( n5428 , n75298 , n5427 );
not ( n5429 , n5428 );
or ( n5430 , n5416 , n5429 );
buf ( n5431 , n4099 );
not ( n75305 , n5431 );
buf ( n75306 , n4119 );
not ( n5434 , n75306 );
not ( n5435 , n74030 );
nand ( n5436 , n5434 , n5435 );
nand ( n5437 , n75306 , n74030 );
nand ( n5438 , n5436 , n5437 );
or ( n5439 , n5438 , n70470 );
not ( n5440 , n5439 );
or ( n5441 , n75305 , n5440 );
not ( n5442 , n455 );
not ( n5443 , n5438 );
or ( n5444 , n5442 , n5443 );
not ( n5445 , n5431 );
nand ( n5446 , n5444 , n5445 );
nand ( n5447 , n5441 , n5446 );
nand ( n5448 , n5430 , n5447 );
not ( n5449 , n5448 );
or ( n5450 , n5415 , n5449 );
not ( n5451 , n5448 );
nand ( n5452 , n5451 , n5409 );
nand ( n5453 , n5450 , n5452 );
not ( n5454 , n5453 );
or ( n5455 , n5414 , n5454 );
not ( n5456 , n537 );
not ( n5457 , n455 );
not ( n5458 , n4163 );
not ( n5459 , n5458 );
not ( n5460 , n74067 );
not ( n5461 , n5460 );
or ( n75335 , n5459 , n5461 );
buf ( n5463 , n4165 );
nand ( n5464 , n75335 , n5463 );
not ( n5465 , n5464 );
not ( n5466 , n5465 );
not ( n5467 , n5436 );
not ( n5468 , n4099 );
or ( n5469 , n5467 , n5468 );
nand ( n5470 , n5469 , n5437 );
not ( n5471 , n5470 );
not ( n5472 , n5471 );
or ( n5473 , n5466 , n5472 );
not ( n5474 , n74047 );
not ( n5475 , n5474 );
nand ( n5476 , n5458 , n5460 );
not ( n5477 , n5476 );
or ( n5478 , n5475 , n5477 );
nand ( n5479 , n5478 , n5470 );
nand ( n5480 , n5473 , n5479 );
not ( n5481 , n5480 );
or ( n5482 , n5457 , n5481 );
not ( n5483 , n5422 );
not ( n5484 , n1222 );
or ( n5485 , n5483 , n5484 );
nand ( n75359 , n5485 , n75290 );
nand ( n5487 , n1511 , n1204 );
not ( n5488 , n5487 );
and ( n5489 , n75359 , n5488 );
not ( n5490 , n75359 );
buf ( n5491 , n5487 );
and ( n5492 , n5490 , n5491 );
nor ( n5493 , n5489 , n5492 );
nand ( n5494 , n5493 , n70470 );
nand ( n5495 , n5482 , n5494 );
not ( n5496 , n5495 );
not ( n5497 , n5496 );
or ( n5498 , n5456 , n5497 );
or ( n5499 , n537 , n5496 );
nand ( n5500 , n5498 , n5499 );
not ( n5501 , n5408 );
nand ( n5502 , n5500 , n5501 );
nand ( n5503 , n5455 , n5502 );
not ( n5504 , n3744 );
nand ( n5505 , n5504 , n3797 );
nand ( n5506 , n4098 , n5505 );
not ( n5507 , n5506 );
buf ( n5508 , n4094 );
not ( n5509 , n455 );
nor ( n5510 , n5508 , n5509 );
not ( n5511 , n5510 );
or ( n5512 , n5507 , n5511 );
nand ( n5513 , n4098 , n5505 , n455 );
not ( n5514 , n5508 );
or ( n5515 , n5513 , n5514 );
nand ( n5516 , n5512 , n5515 );
not ( n75390 , n979 );
and ( n5518 , n988 , n982 );
not ( n5519 , n988 );
not ( n5520 , n982 );
and ( n5521 , n5519 , n5520 );
nor ( n5522 , n5518 , n5521 );
not ( n5523 , n5522 );
and ( n5524 , n75390 , n5523 );
not ( n5525 , n75390 );
and ( n5526 , n5525 , n5522 );
nor ( n5527 , n5524 , n5526 );
nor ( n5528 , n5527 , n455 );
nor ( n5529 , n5516 , n5528 );
not ( n5530 , n5529 );
not ( n5531 , n5530 );
and ( n5532 , n5531 , n537 );
and ( n75406 , n5503 , n5532 );
not ( n75407 , n541 );
not ( n5535 , n4429 );
not ( n5536 , n5535 );
or ( n5537 , n75407 , n5536 );
not ( n5538 , n541 );
nand ( n5539 , n4425 , n5538 );
nand ( n5540 , n5537 , n5539 );
not ( n5541 , n5540 );
and ( n5542 , n542 , n543 );
not ( n5543 , n542 );
and ( n5544 , n5543 , n4938 );
nor ( n5545 , n5542 , n5544 );
not ( n5546 , n5545 );
and ( n5547 , n541 , n542 );
nor ( n5548 , n541 , n542 );
nor ( n5549 , n5547 , n5548 );
and ( n5550 , n5546 , n5549 );
buf ( n5551 , n5550 );
not ( n5552 , n5551 );
or ( n5553 , n5541 , n5552 );
and ( n5554 , n4401 , n4758 );
and ( n5555 , n1680 , n1681 );
nor ( n5556 , n5554 , n5555 );
not ( n5557 , n5556 );
not ( n5558 , n1522 );
or ( n5559 , n5557 , n5558 );
nand ( n5560 , n4766 , n4770 );
nand ( n5561 , n5559 , n5560 );
not ( n5562 , n5561 );
nand ( n5563 , n4765 , n4750 );
and ( n75437 , n5563 , n4239 );
nand ( n5565 , n5562 , n75437 );
nand ( n5566 , n4172 , n3371 , n4174 , n74078 );
nand ( n5567 , n3550 , n3371 );
nand ( n5568 , n5566 , n5567 );
not ( n5569 , n5568 );
nand ( n5570 , n3401 , n4198 );
and ( n5571 , n5570 , n455 );
nand ( n5572 , n5569 , n5571 );
nor ( n5573 , n5563 , n455 );
nand ( n5574 , n5561 , n5573 );
not ( n5575 , n5567 );
not ( n5576 , n5566 );
or ( n75450 , n5575 , n5576 );
and ( n5578 , n3401 , n4198 , n455 );
nand ( n5579 , n75450 , n5578 );
nand ( n5580 , n5565 , n5572 , n5574 , n5579 );
not ( n5581 , n5580 );
not ( n5582 , n5581 );
nand ( n5583 , n5582 , n541 );
not ( n5584 , n5583 );
nand ( n5585 , n5581 , n4219 );
not ( n5586 , n5585 );
or ( n75460 , n5584 , n5586 );
buf ( n5588 , n5545 );
buf ( n5589 , n5588 );
buf ( n5590 , n5589 );
nand ( n5591 , n75460 , n5590 );
nand ( n5592 , n5553 , n5591 );
xor ( n5593 , n75406 , n5592 );
not ( n5594 , n5501 );
not ( n5595 , n455 );
not ( n5596 , n5595 );
buf ( n5597 , n1367 );
or ( n5598 , n1517 , n1366 );
nand ( n5599 , n5597 , n5598 );
not ( n5600 , n1223 );
not ( n5601 , n5422 );
or ( n5602 , n5600 , n5601 );
not ( n5603 , n1512 );
nand ( n5604 , n5602 , n5603 );
and ( n5605 , n5599 , n5604 );
not ( n5606 , n5599 );
not ( n5607 , n5604 );
and ( n5608 , n5606 , n5607 );
nor ( n5609 , n5605 , n5608 );
not ( n5610 , n5609 );
or ( n5611 , n5596 , n5610 );
not ( n5612 , n5463 );
not ( n5613 , n5470 );
or ( n75487 , n5612 , n5613 );
nand ( n5615 , n5458 , n74046 );
buf ( n5616 , n5615 );
nand ( n5617 , n75487 , n5616 );
nand ( n5618 , n4170 , n4156 );
not ( n5619 , n5618 );
and ( n5620 , n5619 , n455 );
and ( n5621 , n5617 , n5620 );
and ( n5622 , n5615 , n5618 , n455 );
nand ( n5623 , n5463 , n5470 );
and ( n5624 , n5622 , n5623 );
nor ( n5625 , n5621 , n5624 );
nand ( n5626 , n5611 , n5625 );
not ( n5627 , n5626 );
not ( n5628 , n5627 );
not ( n5629 , n5628 );
not ( n75503 , n537 );
nand ( n5634 , n5629 , n75503 );
nand ( n75505 , n5628 , n537 );
nand ( n5636 , n5634 , n75505 );
not ( n5637 , n5636 );
or ( n5638 , n5594 , n5637 );
nand ( n5639 , n5413 , n5500 );
nand ( n5640 , n5638 , n5639 );
not ( n5641 , n455 );
nand ( n5642 , n5641 , n5428 );
nand ( n5643 , n5642 , n5447 );
not ( n5644 , n5643 );
nand ( n5645 , n5644 , n537 );
xnor ( n5646 , n5640 , n5645 );
and ( n5647 , n5593 , n5646 );
and ( n5648 , n75406 , n5592 );
or ( n5649 , n5647 , n5648 );
not ( n5650 , n541 );
not ( n75521 , n5595 );
nand ( n5655 , n4778 , n4731 );
xor ( n5656 , n5372 , n5655 );
not ( n5657 , n5656 );
or ( n5658 , n75521 , n5657 );
not ( n5659 , n74132 );
nor ( n5660 , n3485 , n3529 );
nor ( n5661 , n4263 , n5660 );
nand ( n75529 , n4174 , n5099 , n5661 );
nor ( n75530 , n5659 , n75529 );
not ( n5664 , n75530 );
not ( n5665 , n5664 );
not ( n5666 , n3541 );
nor ( n5667 , n5666 , n4233 );
nor ( n5668 , n5667 , n4237 );
or ( n5669 , n5668 , n74982 );
not ( n75537 , n4261 );
nand ( n75538 , n3399 , n3394 );
not ( n5672 , n75538 );
or ( n5673 , n75537 , n5672 );
nand ( n5674 , n5673 , n3401 );
nand ( n5675 , n5669 , n5674 );
not ( n5676 , n5675 );
not ( n5677 , n5676 );
or ( n5678 , n5665 , n5677 );
nand ( n5679 , n3374 , n3390 );
nand ( n5680 , n3392 , n5679 );
not ( n5681 , n5680 );
not ( n5682 , n5681 );
nand ( n5683 , n5678 , n5682 );
nand ( n5684 , n5681 , n5664 , n5676 );
nand ( n5685 , n5683 , n5684 , n455 );
nand ( n5686 , n5658 , n5685 );
not ( n75554 , n5686 );
or ( n5688 , n5650 , n75554 );
not ( n5689 , n5372 );
nand ( n5690 , n5689 , n5655 , n5096 );
not ( n5691 , n5664 );
not ( n5692 , n5676 );
or ( n5693 , n5691 , n5692 );
not ( n5694 , n455 );
nor ( n5695 , n5694 , n5680 );
nand ( n5696 , n5693 , n5695 );
nand ( n5697 , n5676 , n5664 , n5680 , n455 );
nor ( n75565 , n5655 , n455 );
nand ( n75566 , n75565 , n5372 );
nand ( n5700 , n5690 , n5696 , n5697 , n75566 );
not ( n5701 , n5700 );
nand ( n5702 , n5701 , n5538 );
nand ( n5703 , n5688 , n5702 );
nand ( n5704 , n5703 , n5589 );
not ( n5705 , n5585 );
nand ( n5706 , n5582 , n541 );
not ( n5707 , n5706 );
or ( n5708 , n5705 , n5707 );
nand ( n5709 , n5708 , n5551 );
nand ( n5710 , n5704 , n5709 );
not ( n5711 , n5500 );
not ( n5712 , n5711 );
not ( n5713 , n5413 );
not ( n5714 , n5713 );
and ( n5715 , n5712 , n5714 );
and ( n5716 , n5636 , n5501 );
nor ( n5717 , n5715 , n5716 );
nor ( n5718 , n5717 , n5645 );
xor ( n75586 , n5710 , n5718 );
not ( n75587 , n455 );
not ( n5721 , n5480 );
or ( n5722 , n75587 , n5721 );
nand ( n5723 , n5722 , n5494 );
buf ( n5724 , n5723 );
and ( n5725 , n5724 , n537 );
not ( n5726 , n5501 );
not ( n75594 , n537 );
not ( n75595 , n455 );
nand ( n5729 , n74078 , n4233 );
not ( n5730 , n5729 );
and ( n5731 , n4230 , n5730 );
not ( n5732 , n4230 );
and ( n5733 , n5732 , n5729 );
nor ( n5734 , n5731 , n5733 );
not ( n5735 , n5734 );
or ( n5736 , n75595 , n5735 );
not ( n5737 , n5597 );
not ( n5738 , n5604 );
or ( n75606 , n5737 , n5738 );
buf ( n5740 , n5598 );
nand ( n5741 , n75606 , n5740 );
and ( n5742 , n1502 , n1491 );
not ( n5743 , n1502 );
and ( n5744 , n5743 , n1520 );
nor ( n5745 , n5742 , n5744 );
not ( n5746 , n5745 );
and ( n5747 , n5741 , n5746 );
not ( n5748 , n5741 );
and ( n5749 , n5748 , n5745 );
nor ( n5750 , n5747 , n5749 );
nand ( n5751 , n5750 , n70470 );
nand ( n5752 , n5736 , n5751 );
buf ( n5753 , n5752 );
not ( n5754 , n5753 );
not ( n5755 , n5754 );
or ( n5756 , n75594 , n5755 );
nand ( n5757 , n5753 , n5409 );
nand ( n5758 , n5756 , n5757 );
not ( n75626 , n5758 );
or ( n5760 , n5726 , n75626 );
nand ( n5761 , n5413 , n5636 );
nand ( n5762 , n5760 , n5761 );
xor ( n5763 , n5725 , n5762 );
xor ( n5764 , n75586 , n5763 );
xor ( n5765 , n5649 , n5764 );
not ( n5766 , n4434 );
not ( n5767 , n4253 );
or ( n5768 , n5766 , n5767 );
not ( n5769 , n5753 );
not ( n5770 , n5769 );
not ( n5771 , n4224 );
nor ( n5772 , n5771 , n539 );
and ( n5773 , n5770 , n5772 );
nand ( n5774 , n4224 , n539 );
not ( n5775 , n5774 );
and ( n5776 , n5769 , n5775 );
nor ( n5777 , n5773 , n5776 );
nand ( n5778 , n5768 , n5777 );
not ( n5779 , n5753 );
not ( n5780 , n4434 );
nor ( n5781 , n5780 , n4251 );
nand ( n5782 , n5779 , n5781 );
not ( n5783 , n455 );
not ( n5784 , n5734 );
or ( n5785 , n5783 , n5784 );
nand ( n5786 , n5785 , n5751 );
nor ( n5787 , n5780 , n539 );
nand ( n5788 , n5786 , n5787 );
and ( n5789 , n5627 , n539 );
not ( n75657 , n5627 );
and ( n5791 , n75657 , n4251 );
nor ( n5792 , n5789 , n5791 );
nand ( n5793 , n5792 , n4224 );
nand ( n5794 , n5782 , n5788 , n5793 );
not ( n5795 , n537 );
not ( n5796 , n5530 );
or ( n5797 , n5795 , n5796 );
nand ( n5798 , n5409 , n5529 );
nand ( n5799 , n5797 , n5798 );
not ( n5800 , n5799 );
not ( n5801 , n5800 );
not ( n5802 , n5713 );
and ( n5803 , n5801 , n5802 );
and ( n5804 , n5453 , n5501 );
nor ( n5805 , n5803 , n5804 );
not ( n5806 , n70470 );
not ( n5807 , n965 );
buf ( n5808 , n905 );
not ( n5809 , n5808 );
or ( n5810 , n5807 , n5809 );
nand ( n5811 , n972 , n973 );
nand ( n5812 , n5810 , n5811 );
nand ( n5813 , n970 , n977 );
not ( n5814 , n5813 );
and ( n5815 , n5812 , n5814 );
not ( n75683 , n5812 );
and ( n75684 , n75683 , n5813 );
nor ( n5818 , n5815 , n75684 );
not ( n5819 , n5818 );
or ( n5820 , n5806 , n5819 );
nand ( n5821 , n5820 , n4214 );
buf ( n5822 , n5821 );
not ( n5823 , n5822 );
not ( n5824 , n5823 );
nand ( n5825 , n5824 , n537 );
nor ( n5826 , n5805 , n5825 );
xor ( n5827 , n5794 , n5826 );
and ( n5828 , n5413 , n5453 );
and ( n5829 , n5500 , n5501 );
nor ( n5830 , n5828 , n5829 );
and ( n5831 , n5532 , n5830 );
not ( n5832 , n5532 );
and ( n5833 , n5832 , n5503 );
or ( n5834 , n5831 , n5833 );
and ( n5835 , n5827 , n5834 );
and ( n5836 , n5794 , n5826 );
or ( n5837 , n5835 , n5836 );
xor ( n5838 , n5778 , n5837 );
not ( n5839 , n5128 );
not ( n5840 , n4940 );
or ( n5841 , n5839 , n5840 );
not ( n75709 , n4938 );
not ( n5843 , n5701 );
not ( n5844 , n5843 );
not ( n5845 , n5844 );
or ( n5846 , n75709 , n5845 );
nand ( n5847 , n5843 , n543 );
nand ( n5848 , n5846 , n5847 );
nand ( n5849 , n5848 , n4445 );
nand ( n5850 , n5841 , n5849 );
and ( n5851 , n5838 , n5850 );
and ( n5852 , n5778 , n5837 );
or ( n5853 , n5851 , n5852 );
xor ( n5854 , n5765 , n5853 );
xor ( n5855 , n5402 , n5854 );
not ( n5856 , n5399 );
not ( n5857 , n5270 );
or ( n5858 , n5856 , n5857 );
xor ( n5859 , n545 , n74998 );
nand ( n5860 , n5859 , n75018 );
nand ( n5861 , n5858 , n5860 );
xor ( n5862 , n75406 , n5592 );
xor ( n5863 , n5862 , n5646 );
xor ( n5864 , n5861 , n5863 );
not ( n5865 , n4445 );
buf ( n5866 , n5580 );
and ( n5867 , n4938 , n5866 );
not ( n5868 , n4938 );
not ( n5869 , n5866 );
and ( n5870 , n5868 , n5869 );
nor ( n5871 , n5867 , n5870 );
not ( n5872 , n5871 );
or ( n5873 , n5865 , n5872 );
nand ( n5874 , n5848 , n5128 );
nand ( n5875 , n5873 , n5874 );
not ( n5876 , n5551 );
and ( n5877 , n4247 , n5538 );
not ( n75745 , n4247 );
and ( n5879 , n75745 , n541 );
or ( n5880 , n5877 , n5879 );
not ( n5881 , n5880 );
or ( n5882 , n5876 , n5881 );
nand ( n5883 , n5540 , n5590 );
nand ( n5884 , n5882 , n5883 );
xor ( n5885 , n5875 , n5884 );
not ( n5886 , n5137 );
not ( n5887 , n545 );
not ( n5888 , n4933 );
or ( n5889 , n5887 , n5888 );
nand ( n5890 , n4937 , n4440 );
nand ( n5891 , n5889 , n5890 );
not ( n75759 , n5891 );
or ( n5893 , n5886 , n75759 );
nand ( n5894 , n5859 , n5399 );
nand ( n5895 , n5893 , n5894 );
and ( n5896 , n5885 , n5895 );
and ( n5897 , n5875 , n5884 );
or ( n5898 , n5896 , n5897 );
and ( n5899 , n5864 , n5898 );
and ( n5900 , n5861 , n5863 );
or ( n5901 , n5899 , n5900 );
xor ( n5902 , n5855 , n5901 );
xor ( n5903 , n5861 , n5863 );
xor ( n5904 , n5903 , n5898 );
xor ( n5905 , n550 , n551 );
not ( n5906 , n5905 );
not ( n5907 , n2437 );
not ( n5908 , n2284 );
and ( n5909 , n5907 , n5908 );
xor ( n5910 , n1966 , n2132 );
and ( n5911 , n5910 , n2283 );
and ( n5912 , n1966 , n2132 );
or ( n5913 , n5911 , n5912 );
xor ( n75781 , n1833 , n1926 );
and ( n5915 , n75781 , n1965 );
and ( n5916 , n1833 , n1926 );
or ( n5917 , n5915 , n5916 );
or ( n5918 , n1848 , n1870 );
nand ( n5919 , n5918 , n497 );
not ( n5920 , n1784 );
and ( n5921 , n495 , n1855 );
not ( n5922 , n495 );
and ( n5923 , n5922 , n1858 );
or ( n5924 , n5921 , n5923 );
not ( n5925 , n5924 );
or ( n5926 , n5920 , n5925 );
nand ( n5927 , n1997 , n1763 );
nand ( n5928 , n5926 , n5927 );
xor ( n5929 , n5919 , n5928 );
not ( n5930 , n1700 );
not ( n5931 , n1938 );
or ( n5932 , n5930 , n5931 );
not ( n5933 , n491 );
not ( n5934 , n1896 );
or ( n5935 , n5933 , n5934 );
nand ( n5936 , n1899 , n1715 );
nand ( n5937 , n5935 , n5936 );
nand ( n5938 , n5937 , n1739 );
nand ( n5939 , n5932 , n5938 );
xor ( n5940 , n5929 , n5939 );
xor ( n5941 , n1972 , n1988 );
and ( n5942 , n5941 , n2000 );
and ( n5943 , n1972 , n1988 );
or ( n5944 , n5942 , n5943 );
xor ( n75812 , n5940 , n5944 );
xor ( n5949 , n1943 , n1957 );
and ( n75814 , n5949 , n1964 );
and ( n5951 , n1943 , n1957 );
or ( n5952 , n75814 , n5951 );
xor ( n5953 , n1999 , n5952 );
not ( n5954 , n1826 );
not ( n5955 , n1954 );
or ( n5956 , n5954 , n5955 );
xor ( n5957 , n489 , n1726 );
nand ( n5958 , n5957 , n1955 );
nand ( n5959 , n5956 , n5958 );
not ( n5960 , n1986 );
not ( n5961 , n1908 );
or ( n5962 , n5960 , n5961 );
not ( n5963 , n72978 );
not ( n5964 , n5963 );
nand ( n5965 , n1891 , n1976 );
not ( n5966 , n5965 );
or ( n5967 , n5964 , n5966 );
not ( n5968 , n493 );
not ( n5969 , n1891 );
or ( n5970 , n5968 , n5969 );
nand ( n5971 , n5970 , n1770 );
nand ( n5972 , n5967 , n5971 );
nand ( n5973 , n5962 , n5972 );
xor ( n75838 , n5959 , n5973 );
and ( n5978 , n71767 , n489 );
xor ( n5979 , n75838 , n5978 );
xor ( n5980 , n5953 , n5979 );
xor ( n5981 , n75812 , n5980 );
xor ( n5982 , n5917 , n5981 );
xor ( n5983 , n2001 , n2075 );
and ( n5984 , n5983 , n2131 );
and ( n75846 , n2001 , n2075 );
or ( n75847 , n5984 , n75846 );
xor ( n5987 , n5982 , n75847 );
nor ( n5988 , n5913 , n5987 );
nor ( n5989 , n5909 , n5988 );
buf ( n5990 , n5989 );
xor ( n5991 , n1999 , n5952 );
and ( n5992 , n5991 , n5979 );
and ( n75854 , n1999 , n5952 );
or ( n75855 , n5992 , n75854 );
xor ( n5995 , n5919 , n5928 );
and ( n5996 , n5995 , n5939 );
and ( n5997 , n5919 , n5928 );
or ( n5998 , n5996 , n5997 );
not ( n5999 , n71761 );
not ( n75861 , n489 );
not ( n6001 , n1917 );
or ( n6002 , n75861 , n6001 );
nand ( n6003 , n1936 , n1649 );
nand ( n6004 , n6002 , n6003 );
not ( n6005 , n6004 );
or ( n6006 , n5999 , n6005 );
nand ( n6007 , n5957 , n1828 );
nand ( n6008 , n6006 , n6007 );
and ( n6009 , n2199 , n489 );
xor ( n6010 , n6008 , n6009 );
not ( n6011 , n1763 );
not ( n6012 , n5924 );
or ( n6013 , n6011 , n6012 );
nand ( n6014 , n1784 , n495 );
nand ( n6015 , n6013 , n6014 );
xor ( n6016 , n6010 , n6015 );
xor ( n6017 , n5998 , n6016 );
not ( n6018 , n1700 );
not ( n6019 , n5937 );
or ( n6020 , n6018 , n6019 );
not ( n6021 , n491 );
not ( n6022 , n1982 );
not ( n6023 , n6022 );
or ( n6024 , n6021 , n6023 );
nand ( n6025 , n1982 , n1715 );
nand ( n6026 , n6024 , n6025 );
nand ( n6027 , n6026 , n1739 );
nand ( n6028 , n6020 , n6027 );
and ( n6029 , n1976 , n72978 );
not ( n6030 , n1976 );
and ( n6031 , n6030 , n5963 );
nor ( n6032 , n6029 , n6031 );
not ( n6033 , n6032 );
not ( n6034 , n1909 );
or ( n75896 , n6033 , n6034 );
and ( n75897 , n456 , n458 );
not ( n6037 , n456 );
and ( n6038 , n6037 , n474 );
nor ( n6039 , n75897 , n6038 );
and ( n6040 , n493 , n6039 );
not ( n6041 , n493 );
and ( n6042 , n6041 , n1995 );
or ( n6043 , n6040 , n6042 );
nand ( n6044 , n6043 , n1891 );
nand ( n6045 , n75896 , n6044 );
not ( n6046 , n6045 );
xor ( n6047 , n6028 , n6046 );
xor ( n6048 , n5959 , n5973 );
and ( n6049 , n6048 , n5978 );
and ( n6050 , n5959 , n5973 );
or ( n75912 , n6049 , n6050 );
xor ( n75913 , n6047 , n75912 );
xor ( n6053 , n6017 , n75913 );
xor ( n6054 , n75855 , n6053 );
xor ( n6055 , n5940 , n5944 );
and ( n6056 , n6055 , n5980 );
and ( n6057 , n5940 , n5944 );
or ( n6058 , n6056 , n6057 );
xor ( n75920 , n6054 , n6058 );
xor ( n75921 , n5917 , n5981 );
and ( n6061 , n75921 , n75847 );
and ( n6062 , n5917 , n5981 );
or ( n6063 , n6061 , n6062 );
nor ( n6064 , n75920 , n6063 );
not ( n6065 , n6064 );
and ( n6066 , n5990 , n6065 );
not ( n6067 , n6066 );
not ( n6068 , n4203 );
or ( n6069 , n6067 , n6068 );
not ( n6070 , n5913 );
not ( n6071 , n5987 );
or ( n6072 , n6070 , n6071 );
nor ( n6073 , n5987 , n5913 );
nand ( n6074 , n2284 , n2437 );
or ( n6075 , n6073 , n6074 );
nand ( n6076 , n6072 , n6075 );
buf ( n6077 , n6076 );
not ( n6078 , n6063 );
not ( n6079 , n75920 );
nand ( n6080 , n6078 , n6079 );
and ( n6081 , n6077 , n6080 );
nand ( n6082 , n6063 , n75920 );
not ( n6083 , n6082 );
nor ( n6084 , n6081 , n6083 );
nand ( n6085 , n6069 , n6084 );
xor ( n6086 , n6028 , n6046 );
and ( n6087 , n6086 , n75912 );
and ( n6088 , n6028 , n6046 );
or ( n6089 , n6087 , n6088 );
xor ( n75951 , n6008 , n6009 );
and ( n6091 , n75951 , n6015 );
and ( n6092 , n6008 , n6009 );
or ( n6093 , n6091 , n6092 );
or ( n6094 , n1784 , n1763 );
nand ( n6095 , n6094 , n495 );
not ( n6096 , n1891 );
and ( n6097 , n493 , n1855 );
not ( n6098 , n493 );
and ( n6099 , n6098 , n1858 );
or ( n6100 , n6097 , n6099 );
not ( n6101 , n6100 );
or ( n6102 , n6096 , n6101 );
nand ( n6103 , n6043 , n1909 );
nand ( n6104 , n6102 , n6103 );
xor ( n6105 , n6095 , n6104 );
not ( n6106 , n71761 );
xor ( n6107 , n489 , n1899 );
not ( n6108 , n6107 );
or ( n6109 , n6106 , n6108 );
nand ( n6110 , n6004 , n1828 );
nand ( n6111 , n6109 , n6110 );
xor ( n6112 , n6105 , n6111 );
xor ( n75974 , n6093 , n6112 );
and ( n6114 , n489 , n1726 );
not ( n6115 , n1739 );
not ( n6116 , n491 );
not ( n6117 , n1770 );
or ( n6118 , n6116 , n6117 );
not ( n75980 , n1778 );
not ( n6120 , n75980 );
nand ( n6121 , n6120 , n1715 );
nand ( n6122 , n6118 , n6121 );
not ( n6123 , n6122 );
or ( n6124 , n6115 , n6123 );
nand ( n6125 , n6026 , n1700 );
nand ( n6126 , n6124 , n6125 );
xor ( n6127 , n6114 , n6126 );
xor ( n6128 , n6127 , n6045 );
xor ( n6129 , n75974 , n6128 );
xor ( n6130 , n6089 , n6129 );
xor ( n6131 , n5998 , n6016 );
and ( n6132 , n6131 , n75913 );
and ( n6133 , n5998 , n6016 );
or ( n6134 , n6132 , n6133 );
xor ( n6135 , n6130 , n6134 );
not ( n6136 , n6135 );
xor ( n6137 , n75855 , n6053 );
and ( n6138 , n6137 , n6058 );
and ( n6139 , n75855 , n6053 );
or ( n6140 , n6138 , n6139 );
not ( n6141 , n6140 );
nand ( n6142 , n6136 , n6141 );
not ( n6143 , n6141 );
nand ( n6144 , n6143 , n6135 );
nand ( n6145 , n6142 , n6144 );
not ( n6146 , n6145 );
and ( n6147 , n6146 , n455 );
and ( n6148 , n6085 , n6147 );
not ( n6149 , n6085 );
and ( n6150 , n6145 , n455 );
and ( n6151 , n6149 , n6150 );
nor ( n6152 , n6148 , n6151 );
not ( n6153 , n5361 );
not ( n6154 , n5356 );
or ( n6155 , n6153 , n6154 );
xor ( n6156 , n5304 , n5308 );
and ( n6157 , n6156 , n5354 );
and ( n6158 , n5304 , n5308 );
or ( n6159 , n6157 , n6158 );
not ( n6160 , n6159 );
xor ( n6161 , n5278 , n5298 );
and ( n6162 , n6161 , n5303 );
and ( n6163 , n5278 , n5298 );
or ( n6164 , n6162 , n6163 );
not ( n6165 , n6164 );
not ( n76027 , n6165 );
xor ( n76028 , n5319 , n5325 );
and ( n6168 , n76028 , n5332 );
and ( n6169 , n5319 , n5325 );
or ( n6170 , n6168 , n6169 );
not ( n6171 , n6170 );
not ( n6172 , n6171 );
not ( n6173 , n5323 );
not ( n6174 , n70536 );
or ( n6175 , n6173 , n6174 );
xor ( n6176 , n505 , n495 );
nand ( n6177 , n70544 , n6176 );
nand ( n6178 , n6175 , n6177 );
not ( n6179 , n70513 );
not ( n6180 , n6179 );
not ( n6181 , n75172 );
or ( n6182 , n6180 , n6181 );
nand ( n6183 , n6182 , n497 );
xor ( n6184 , n6178 , n6183 );
not ( n6185 , n5289 );
not ( n6186 , n1627 );
or ( n6187 , n6185 , n6186 );
xor ( n6188 , n509 , n491 );
nand ( n6189 , n1630 , n6188 );
nand ( n6190 , n6187 , n6189 );
not ( n6191 , n6190 );
and ( n6192 , n6184 , n6191 );
not ( n6193 , n6184 );
and ( n6194 , n6193 , n6190 );
nor ( n6195 , n6192 , n6194 );
not ( n6196 , n6195 );
not ( n6197 , n6196 );
or ( n6198 , n6172 , n6197 );
nand ( n6199 , n6195 , n6170 );
nand ( n6200 , n6198 , n6199 );
not ( n6201 , n5325 );
not ( n6202 , n6201 );
not ( n76064 , n5291 );
not ( n6204 , n5284 );
or ( n6205 , n76064 , n6204 );
nor ( n6206 , n5291 , n5284 );
or ( n6207 , n5297 , n6206 );
nand ( n6208 , n6205 , n6207 );
not ( n6209 , n6208 );
not ( n6210 , n6209 );
or ( n6211 , n6202 , n6210 );
not ( n6212 , n6201 );
nand ( n6213 , n6212 , n6208 );
nand ( n6214 , n6211 , n6213 );
nand ( n6215 , n513 , n489 );
xor ( n6216 , n489 , n511 );
nand ( n6217 , n1553 , n6216 );
nand ( n6218 , n5003 , n5282 );
and ( n6219 , n6217 , n6218 );
xor ( n76081 , n6215 , n6219 );
not ( n6221 , n5330 );
xnor ( n6222 , n508 , n493 );
not ( n6223 , n6222 );
and ( n6224 , n6221 , n6223 );
xor ( n6225 , n493 , n507 );
and ( n6226 , n70491 , n6225 );
nor ( n6227 , n6224 , n6226 );
xor ( n6228 , n76081 , n6227 );
not ( n6229 , n6228 );
not ( n6230 , n6229 );
and ( n6231 , n6214 , n6230 );
not ( n6232 , n6214 );
and ( n6233 , n6232 , n6229 );
nor ( n76095 , n6231 , n6233 );
and ( n6235 , n6200 , n76095 );
not ( n6236 , n6200 );
not ( n6237 , n76095 );
and ( n6238 , n6236 , n6237 );
nor ( n6239 , n6235 , n6238 );
not ( n6240 , n6239 );
or ( n6241 , n76027 , n6240 );
or ( n6242 , n6239 , n6165 );
nand ( n6243 , n6241 , n6242 );
not ( n6244 , n5340 );
nand ( n6245 , n6244 , n5333 );
not ( n6246 , n6245 );
not ( n6247 , n5318 );
or ( n6248 , n6246 , n6247 );
nand ( n6249 , n6248 , n5345 );
xor ( n6250 , n6243 , n6249 );
nand ( n6251 , n6160 , n6250 );
nand ( n6252 , n6155 , n6251 );
buf ( n6253 , n6252 );
nand ( n6254 , n6239 , n6165 );
not ( n6255 , n6254 );
not ( n6256 , n6249 );
or ( n6257 , n6255 , n6256 );
or ( n6258 , n6165 , n6239 );
nand ( n6259 , n6257 , n6258 );
not ( n6260 , n6201 );
not ( n6261 , n6228 );
or ( n6262 , n6260 , n6261 );
nand ( n6263 , n6262 , n6208 );
nand ( n6264 , n6229 , n5325 );
nand ( n6265 , n6263 , n6264 );
not ( n6266 , n6265 );
nand ( n6267 , n512 , n489 );
not ( n6268 , n6267 );
not ( n6269 , n6216 );
not ( n76131 , n4364 );
or ( n6271 , n6269 , n76131 );
xor ( n6272 , n489 , n510 );
nand ( n6273 , n1553 , n6272 );
nand ( n6274 , n6271 , n6273 );
not ( n6275 , n6274 );
xor ( n6276 , n6268 , n6275 );
not ( n6277 , n6176 );
not ( n6278 , n4466 );
or ( n6279 , n6277 , n6278 );
nand ( n6280 , n70544 , n495 );
nand ( n6281 , n6279 , n6280 );
xor ( n6282 , n6276 , n6281 );
not ( n76144 , n6190 );
not ( n6287 , n6178 );
or ( n76146 , n76144 , n6287 );
not ( n6289 , n6191 );
not ( n6290 , n6178 );
not ( n6291 , n6290 );
or ( n6292 , n6289 , n6291 );
nand ( n6293 , n6292 , n6183 );
nand ( n6294 , n76146 , n6293 );
not ( n6295 , n6294 );
xor ( n6296 , n6282 , n6295 );
not ( n6297 , n6225 );
not ( n6298 , n1157 );
or ( n6299 , n6297 , n6298 );
xor ( n6300 , n506 , n493 );
nand ( n6301 , n70491 , n6300 );
nand ( n6302 , n6299 , n6301 );
not ( n6303 , n6188 );
not ( n6304 , n1627 );
or ( n6305 , n6303 , n6304 );
xor ( n6306 , n508 , n491 );
nand ( n6307 , n1630 , n6306 );
nand ( n6308 , n6305 , n6307 );
xor ( n6309 , n6302 , n6308 );
xor ( n6310 , n6215 , n6219 );
and ( n6311 , n6310 , n6227 );
and ( n76170 , n6215 , n6219 );
or ( n6316 , n6311 , n76170 );
not ( n6317 , n6316 );
and ( n6318 , n6309 , n6317 );
not ( n6319 , n6309 );
and ( n6320 , n6319 , n6316 );
nor ( n76176 , n6318 , n6320 );
xor ( n76177 , n6296 , n76176 );
xor ( n6323 , n6266 , n76177 );
not ( n6324 , n6199 );
not ( n6325 , n76095 );
or ( n6326 , n6324 , n6325 );
or ( n6327 , n6195 , n6170 );
nand ( n6328 , n6326 , n6327 );
xnor ( n76184 , n6323 , n6328 );
not ( n76185 , n76184 );
nor ( n6331 , n6259 , n76185 );
nor ( n6332 , n6253 , n6331 );
and ( n6333 , n6332 , n5091 , n5254 );
not ( n6334 , n6333 );
not ( n6335 , n75048 );
or ( n6336 , n6334 , n6335 );
nor ( n6337 , n6252 , n6331 );
not ( n6338 , n6337 );
not ( n6339 , n5384 );
or ( n6340 , n6338 , n6339 );
not ( n6341 , n6251 );
not ( n6342 , n5363 );
or ( n76198 , n6341 , n6342 );
not ( n76199 , n6250 );
nand ( n6345 , n76199 , n6159 );
nand ( n6346 , n76198 , n6345 );
not ( n6347 , n6259 );
buf ( n6348 , n76184 );
nand ( n6349 , n6347 , n6348 );
and ( n6350 , n6346 , n6349 );
nand ( n76206 , n6259 , n76185 );
not ( n76207 , n76206 );
nor ( n6353 , n6350 , n76207 );
nand ( n6354 , n6340 , n6353 );
not ( n6355 , n6354 );
nand ( n6356 , n6336 , n6355 );
and ( n6357 , n489 , n511 );
xor ( n6358 , n6357 , n6302 );
xor ( n6359 , n507 , n491 );
nand ( n6360 , n1630 , n6359 );
nand ( n6361 , n6306 , n1627 );
nand ( n6362 , n6360 , n6361 );
xor ( n6363 , n6358 , n6362 );
not ( n6364 , n6363 );
not ( n6365 , n6364 );
not ( n6366 , n6267 );
not ( n6367 , n6275 );
or ( n6368 , n6366 , n6367 );
nand ( n6369 , n6368 , n6281 );
nand ( n6370 , n6268 , n6274 );
nand ( n6371 , n6369 , n6370 );
not ( n6372 , n6371 );
or ( n6373 , n6365 , n6372 );
not ( n6374 , n6371 );
nand ( n6375 , n6363 , n6374 );
nand ( n6376 , n6373 , n6375 );
not ( n76232 , n6300 );
not ( n6378 , n1268 );
or ( n6379 , n76232 , n6378 );
xor ( n6380 , n505 , n493 );
nand ( n6381 , n992 , n6380 );
nand ( n6382 , n6379 , n6381 );
not ( n6383 , n6272 );
buf ( n6384 , n4364 );
not ( n6385 , n6384 );
or ( n6386 , n6383 , n6385 );
xor ( n6387 , n489 , n509 );
nand ( n6388 , n1553 , n6387 );
nand ( n76244 , n6386 , n6388 );
not ( n76245 , n76244 );
xor ( n6391 , n6382 , n76245 );
or ( n6392 , n4466 , n70544 );
nand ( n6393 , n6392 , n495 );
xnor ( n6394 , n6391 , n6393 );
xor ( n6395 , n6376 , n6394 );
not ( n6396 , n6395 );
not ( n6397 , n6308 );
nand ( n6398 , n6397 , n6302 );
not ( n6399 , n6398 );
not ( n6400 , n6317 );
or ( n6401 , n6399 , n6400 );
not ( n6402 , n6302 );
nand ( n6403 , n6402 , n6308 );
nand ( n6404 , n6401 , n6403 );
not ( n6405 , n6404 );
not ( n6406 , n6405 );
and ( n6407 , n6396 , n6406 );
and ( n6408 , n6395 , n6405 );
nor ( n6409 , n6407 , n6408 );
not ( n6410 , n76176 );
not ( n6411 , n6282 );
or ( n6412 , n6410 , n6411 );
nand ( n6413 , n6412 , n6294 );
not ( n6414 , n76176 );
nand ( n6415 , n6414 , n6411 );
nand ( n6416 , n6413 , n6415 );
xor ( n6417 , n6409 , n6416 );
not ( n6418 , n6266 );
not ( n6419 , n76177 );
or ( n76275 , n6418 , n6419 );
nand ( n6421 , n76275 , n6328 );
not ( n6422 , n76177 );
nand ( n6423 , n6422 , n6265 );
and ( n6424 , n6421 , n6423 );
nor ( n6425 , n6417 , n6424 );
not ( n6426 , n6425 );
not ( n6427 , n6424 );
not ( n6428 , n6427 );
nand ( n6429 , n6428 , n6417 );
nand ( n6430 , n6426 , n6429 );
not ( n6431 , n6430 );
and ( n6432 , n6431 , n74671 );
and ( n6433 , n6356 , n6432 );
not ( n6434 , n6356 );
not ( n6435 , n6430 );
nor ( n6436 , n6435 , n455 );
and ( n6437 , n6434 , n6436 );
nor ( n6438 , n6433 , n6437 );
nand ( n6439 , n6152 , n6438 );
not ( n6440 , n6439 );
xor ( n6441 , n549 , n6440 );
not ( n6442 , n6441 );
or ( n76298 , n5906 , n6442 );
not ( n6444 , n549 );
not ( n6445 , n5990 );
not ( n6446 , n3401 );
nor ( n6447 , n6446 , n4197 );
nand ( n6448 , n5568 , n6447 , n4192 , n2969 );
nand ( n76304 , n6448 , n4202 , n4194 );
not ( n6450 , n76304 );
or ( n6451 , n6445 , n6450 );
not ( n6452 , n4188 );
and ( n6453 , n6452 , n5990 );
nor ( n6454 , n6453 , n6077 );
nand ( n6455 , n6451 , n6454 );
not ( n6456 , n6455 );
nand ( n6457 , n6082 , n6080 );
nand ( n6458 , n6456 , n6457 );
not ( n6459 , n6458 );
not ( n6460 , n6457 );
and ( n6461 , n6455 , n6460 );
nor ( n6462 , n6461 , n5509 );
not ( n6463 , n6462 );
or ( n6464 , n6459 , n6463 );
not ( n6465 , n6252 );
not ( n6466 , n6465 );
not ( n6467 , n5387 );
or ( n6468 , n6466 , n6467 );
not ( n6469 , n6346 );
nand ( n6470 , n6468 , n6469 );
nand ( n6471 , n6349 , n76206 );
not ( n6472 , n6471 );
and ( n6473 , n6470 , n6472 );
not ( n6474 , n6470 );
and ( n6475 , n6474 , n6471 );
nor ( n6476 , n6473 , n6475 );
nand ( n6477 , n6476 , n70470 );
nand ( n6478 , n6464 , n6477 );
not ( n6479 , n6478 );
not ( n6480 , n6479 );
or ( n6481 , n6444 , n6480 );
not ( n6482 , n549 );
nand ( n6483 , n6482 , n6478 );
nand ( n6484 , n6481 , n6483 );
and ( n6485 , n549 , n550 );
nor ( n6486 , n549 , n550 );
nor ( n6487 , n6485 , n5905 , n6486 );
not ( n6488 , n6487 );
not ( n6489 , n6488 );
nand ( n6490 , n6484 , n6489 );
nand ( n6491 , n76298 , n6490 );
not ( n6492 , n552 );
not ( n6493 , n4946 );
not ( n6494 , n4774 );
or ( n6495 , n6493 , n6494 );
not ( n6496 , n4961 );
nand ( n6497 , n6495 , n6496 );
nor ( n6498 , n6252 , n6331 );
nand ( n6499 , n5381 , n6429 , n6498 );
not ( n6500 , n6499 );
and ( n6501 , n6497 , n6500 );
not ( n6502 , n6429 );
not ( n6503 , n6354 );
or ( n6504 , n6502 , n6503 );
buf ( n6505 , n6426 );
nand ( n6506 , n6504 , n6505 );
or ( n6507 , n6501 , n6506 );
not ( n6508 , n6404 );
not ( n6509 , n6395 );
or ( n6510 , n6508 , n6509 );
not ( n6511 , n6405 );
not ( n6512 , n6395 );
not ( n6513 , n6512 );
or ( n76369 , n6511 , n6513 );
nand ( n76370 , n76369 , n6416 );
nand ( n6516 , n6510 , n76370 );
xor ( n6517 , n6357 , n6302 );
and ( n6518 , n6517 , n6362 );
and ( n6519 , n6357 , n6302 );
or ( n6520 , n6518 , n6519 );
not ( n6521 , n6520 );
not ( n6522 , n6363 );
not ( n6523 , n6371 );
or ( n6524 , n6522 , n6523 );
not ( n6525 , n6374 );
not ( n6526 , n6364 );
or ( n6527 , n6525 , n6526 );
nand ( n6528 , n6527 , n6394 );
nand ( n6529 , n6524 , n6528 );
xor ( n6530 , n6521 , n6529 );
not ( n6531 , n6380 );
not ( n6532 , n1157 );
or ( n6533 , n6531 , n6532 );
nand ( n6534 , n992 , n493 );
nand ( n6535 , n6533 , n6534 );
not ( n6536 , n6535 );
and ( n6537 , n489 , n510 );
not ( n6538 , n6387 );
not ( n6539 , n6384 );
or ( n6540 , n6538 , n6539 );
xnor ( n6541 , n489 , n508 );
not ( n6542 , n6541 );
nand ( n6543 , n6542 , n1553 );
nand ( n6544 , n6540 , n6543 );
xor ( n6545 , n6537 , n6544 );
not ( n76401 , n6359 );
not ( n6547 , n4337 );
or ( n6548 , n76401 , n6547 );
xnor ( n6549 , n491 , n506 );
not ( n6550 , n6549 );
nand ( n6551 , n6550 , n1630 );
nand ( n6552 , n6548 , n6551 );
xor ( n6553 , n6545 , n6552 );
xor ( n6554 , n6536 , n6553 );
not ( n6555 , n76245 );
not ( n6556 , n6393 );
not ( n6557 , n6556 );
or ( n6558 , n6555 , n6557 );
nand ( n6559 , n6558 , n6382 );
nand ( n6560 , n6393 , n76244 );
nand ( n6561 , n6559 , n6560 );
xor ( n6562 , n6554 , n6561 );
not ( n6563 , n6562 );
not ( n6564 , n6563 );
xnor ( n6565 , n6530 , n6564 );
nor ( n6566 , n6516 , n6565 );
not ( n6567 , n6566 );
nand ( n6568 , n6507 , n6567 );
nand ( n6569 , n6565 , n6516 );
buf ( n6570 , n6569 );
not ( n6571 , n6564 );
not ( n6572 , n6520 );
or ( n6573 , n6571 , n6572 );
not ( n6574 , n6563 );
not ( n6575 , n6521 );
or ( n6576 , n6574 , n6575 );
nand ( n6577 , n6576 , n6529 );
nand ( n76433 , n6573 , n6577 );
and ( n6579 , n489 , n509 );
not ( n6580 , n4337 );
or ( n6581 , n6580 , n6549 );
not ( n6582 , n1630 );
and ( n6583 , n491 , n4863 );
not ( n6584 , n491 );
and ( n6585 , n6584 , n505 );
nor ( n6586 , n6583 , n6585 );
or ( n6587 , n6582 , n6586 );
nand ( n6588 , n6581 , n6587 );
xor ( n6589 , n6579 , n6588 );
not ( n6590 , n991 );
not ( n6591 , n5330 );
or ( n6592 , n6590 , n6591 );
nand ( n6593 , n6592 , n493 );
xor ( n6594 , n6589 , n6593 );
not ( n6595 , n6384 );
or ( n6596 , n6595 , n6541 );
not ( n6597 , n1553 );
xnor ( n6598 , n507 , n489 );
or ( n6599 , n6597 , n6598 );
nand ( n6600 , n6596 , n6599 );
and ( n6601 , n6600 , n6535 );
not ( n6602 , n6600 );
and ( n76458 , n6602 , n6536 );
nor ( n6604 , n6601 , n76458 );
xor ( n6605 , n6537 , n6544 );
and ( n6606 , n6605 , n6552 );
and ( n6607 , n6537 , n6544 );
or ( n6608 , n6606 , n6607 );
and ( n6609 , n6604 , n6608 );
not ( n6610 , n6604 );
not ( n6611 , n6608 );
and ( n6612 , n6610 , n6611 );
or ( n6613 , n6609 , n6612 );
xor ( n6614 , n6594 , n6613 );
xor ( n6615 , n6536 , n6553 );
and ( n6616 , n6615 , n6561 );
and ( n6617 , n6536 , n6553 );
or ( n6618 , n6616 , n6617 );
xnor ( n76474 , n6614 , n6618 );
nor ( n6620 , n76433 , n76474 );
not ( n6621 , n6620 );
nand ( n6622 , n76433 , n76474 );
and ( n6623 , n6570 , n6621 , n6622 , n70470 );
and ( n6624 , n6568 , n6623 );
and ( n6625 , n6570 , n6568 );
not ( n6626 , n6621 );
not ( n6627 , n6622 );
or ( n6628 , n6626 , n6627 );
nand ( n6629 , n6628 , n70470 );
nor ( n6630 , n6625 , n6629 );
nor ( n6631 , n6624 , n6630 );
nor ( n6632 , n6140 , n6135 );
nor ( n6633 , n6064 , n6632 );
nand ( n6634 , n5989 , n6633 );
xor ( n6635 , n6089 , n6129 );
and ( n6636 , n6635 , n6134 );
and ( n6637 , n6089 , n6129 );
or ( n6638 , n6636 , n6637 );
xor ( n6639 , n6114 , n6126 );
and ( n6640 , n6639 , n6045 );
and ( n6641 , n6114 , n6126 );
or ( n6642 , n6640 , n6641 );
and ( n6643 , n6100 , n1909 );
and ( n6644 , n1891 , n493 );
nor ( n6645 , n6643 , n6644 );
xor ( n6646 , n6095 , n6104 );
and ( n6647 , n6646 , n6111 );
and ( n6648 , n6095 , n6104 );
or ( n6649 , n6647 , n6648 );
xor ( n6650 , n6645 , n6649 );
and ( n6651 , n1936 , n489 );
not ( n6652 , n1739 );
not ( n6653 , n491 );
not ( n6654 , n1874 );
or ( n76510 , n6653 , n6654 );
nand ( n6659 , n1995 , n1715 );
nand ( n76512 , n76510 , n6659 );
not ( n6661 , n76512 );
or ( n6662 , n6652 , n6661 );
nand ( n6663 , n6122 , n1700 );
nand ( n6664 , n6662 , n6663 );
xor ( n6665 , n6651 , n6664 );
not ( n6666 , n1828 );
not ( n6667 , n6107 );
or ( n6668 , n6666 , n6667 );
xor ( n6669 , n489 , n1982 );
nand ( n6670 , n6669 , n71761 );
nand ( n6671 , n6668 , n6670 );
xor ( n6672 , n6665 , n6671 );
xor ( n6673 , n6650 , n6672 );
xor ( n6674 , n6642 , n6673 );
xor ( n6675 , n6093 , n6112 );
and ( n6676 , n6675 , n6128 );
and ( n6677 , n6093 , n6112 );
or ( n6678 , n6676 , n6677 );
xor ( n6679 , n6674 , n6678 );
nor ( n6680 , n6638 , n6679 );
nor ( n6681 , n6634 , n6680 );
not ( n6682 , n6681 );
not ( n6683 , n4203 );
or ( n76536 , n6682 , n6683 );
not ( n6688 , n6680 );
not ( n6689 , n6633 );
not ( n6690 , n6076 );
or ( n6691 , n6689 , n6690 );
or ( n6692 , n6082 , n6632 );
nand ( n6693 , n6140 , n6135 );
nand ( n76543 , n6692 , n6693 );
not ( n76544 , n76543 );
nand ( n6696 , n6691 , n76544 );
and ( n6697 , n6688 , n6696 );
nand ( n6698 , n6679 , n6638 );
not ( n6699 , n6698 );
nor ( n6700 , n6697 , n6699 );
nand ( n6701 , n76536 , n6700 );
or ( n76551 , n1891 , n1909 );
nand ( n76552 , n76551 , n493 );
not ( n6704 , n1700 );
not ( n6705 , n76512 );
or ( n6706 , n6704 , n6705 );
not ( n6707 , n491 );
not ( n6708 , n1855 );
or ( n6709 , n6707 , n6708 );
nand ( n6710 , n1858 , n1715 );
nand ( n6711 , n6709 , n6710 );
nand ( n6712 , n6711 , n1739 );
nand ( n6713 , n6706 , n6712 );
xor ( n6714 , n76552 , n6713 );
and ( n6715 , n489 , n1899 );
xor ( n6716 , n6714 , n6715 );
not ( n6717 , n71761 );
xor ( n6718 , n489 , n6120 );
not ( n6719 , n6718 );
or ( n6720 , n6717 , n6719 );
nand ( n6721 , n6669 , n1828 );
nand ( n6722 , n6720 , n6721 );
not ( n6723 , n6645 );
xor ( n6724 , n6722 , n6723 );
xor ( n6725 , n6651 , n6664 );
and ( n6726 , n6725 , n6671 );
and ( n6727 , n6651 , n6664 );
or ( n6728 , n6726 , n6727 );
xor ( n6729 , n6724 , n6728 );
xor ( n6730 , n6716 , n6729 );
xor ( n6731 , n6645 , n6649 );
and ( n6732 , n6731 , n6672 );
and ( n6733 , n6645 , n6649 );
or ( n6734 , n6732 , n6733 );
xor ( n6735 , n6730 , n6734 );
xor ( n6736 , n6642 , n6673 );
and ( n6737 , n6736 , n6678 );
and ( n76587 , n6642 , n6673 );
or ( n76588 , n6737 , n76587 );
nor ( n6740 , n6735 , n76588 );
not ( n6741 , n6740 );
nand ( n6742 , n6735 , n76588 );
nand ( n6743 , n6741 , n6742 );
and ( n6744 , n6743 , n455 );
and ( n6745 , n6701 , n6744 );
not ( n76595 , n6701 );
not ( n76596 , n455 );
nor ( n6748 , n76596 , n6743 );
and ( n6749 , n76595 , n6748 );
nor ( n6750 , n6745 , n6749 );
nand ( n6751 , n6631 , n6750 );
not ( n6752 , n551 );
and ( n76602 , n6751 , n6752 );
not ( n6754 , n6751 );
and ( n6755 , n6754 , n551 );
or ( n6756 , n76602 , n6755 );
not ( n6757 , n6756 );
or ( n6758 , n6492 , n6757 );
not ( n6759 , n551 );
not ( n6760 , n70470 );
not ( n6761 , n6496 );
nand ( n6762 , n6500 , n6761 );
not ( n6763 , n6499 );
buf ( n6764 , n4774 );
nand ( n6765 , n6763 , n6764 , n4946 );
not ( n6766 , n6417 );
not ( n6767 , n6424 );
and ( n6768 , n6766 , n6767 );
and ( n6769 , n6354 , n6429 );
nor ( n6770 , n6768 , n6769 );
nand ( n6771 , n6762 , n6765 , n6770 );
nand ( n6772 , n6567 , n6569 );
not ( n6773 , n6772 );
and ( n6774 , n6771 , n6773 );
not ( n6775 , n6771 );
and ( n6776 , n6775 , n6772 );
nor ( n6777 , n6774 , n6776 );
not ( n6778 , n6777 );
or ( n6779 , n6760 , n6778 );
not ( n6780 , n6634 );
not ( n6781 , n6780 );
not ( n6782 , n4203 );
or ( n6783 , n6781 , n6782 );
not ( n6784 , n6696 );
nand ( n6785 , n6783 , n6784 );
nand ( n6786 , n6688 , n6698 );
and ( n6787 , n455 , n6786 );
and ( n6788 , n6785 , n6787 );
not ( n6789 , n6785 );
not ( n6790 , n455 );
nor ( n6791 , n6790 , n6786 );
and ( n6792 , n6789 , n6791 );
nor ( n6793 , n6788 , n6792 );
nand ( n76643 , n6779 , n6793 );
buf ( n76644 , n76643 );
not ( n6796 , n76644 );
not ( n6797 , n6796 );
or ( n6798 , n6759 , n6797 );
nand ( n6799 , n76644 , n6752 );
nand ( n6800 , n6798 , n6799 );
not ( n6801 , n552 );
and ( n6802 , n6801 , n551 );
nand ( n6803 , n6800 , n6802 );
nand ( n6804 , n6758 , n6803 );
xor ( n6805 , n6491 , n6804 );
not ( n6806 , n549 );
not ( n6807 , n548 );
or ( n6808 , n6806 , n6807 );
or ( n6809 , n548 , n549 );
nand ( n6810 , n6808 , n6809 );
not ( n6811 , n6810 );
not ( n6812 , n6811 );
not ( n6813 , n6448 );
nand ( n6814 , n4202 , n4194 );
nor ( n6815 , n6813 , n6814 );
not ( n6816 , n2438 );
or ( n6817 , n6815 , n6816 );
not ( n6818 , n2439 );
nor ( n76668 , n4188 , n6816 );
nor ( n6820 , n6818 , n76668 );
nand ( n6821 , n6817 , n6820 );
not ( n6822 , n5988 );
nand ( n6823 , n5913 , n5987 );
nand ( n6824 , n6822 , n6823 );
nand ( n6825 , n6824 , n455 );
nor ( n6826 , n6821 , n6825 );
not ( n6827 , n6826 );
not ( n6828 , n5362 );
not ( n6829 , n5387 );
or ( n6830 , n6828 , n6829 );
nand ( n6831 , n6830 , n5364 );
not ( n6832 , n6831 );
nand ( n6833 , n6251 , n6345 );
not ( n6834 , n6833 );
nor ( n6835 , n6834 , n455 );
nand ( n6836 , n6832 , n6835 );
nor ( n6837 , n6833 , n455 );
nand ( n6838 , n6831 , n6837 );
not ( n6839 , n455 );
nor ( n6840 , n6839 , n6824 );
nand ( n6841 , n6840 , n6821 );
nand ( n6842 , n6827 , n6836 , n6838 , n6841 );
not ( n6843 , n6842 );
not ( n6844 , n6843 );
and ( n6845 , n547 , n6844 );
not ( n6846 , n547 );
not ( n6847 , n6843 );
not ( n6848 , n6847 );
and ( n6849 , n6846 , n6848 );
or ( n6850 , n6845 , n6849 );
not ( n6851 , n6850 );
or ( n76701 , n6812 , n6851 );
xor ( n6853 , n548 , n547 );
and ( n6854 , n6853 , n6810 );
and ( n6855 , n5392 , n547 );
not ( n6856 , n5392 );
not ( n6857 , n547 );
and ( n6858 , n6856 , n6857 );
nor ( n6859 , n6855 , n6858 );
nand ( n6860 , n6854 , n6859 );
nand ( n6861 , n76701 , n6860 );
xor ( n76711 , n6805 , n6861 );
xor ( n6863 , n5904 , n76711 );
not ( n6864 , n6800 );
not ( n6865 , n552 );
or ( n6866 , n6864 , n6865 );
not ( n6867 , n6440 );
buf ( n6868 , n6802 );
nand ( n6869 , n6867 , n6868 );
nand ( n6870 , n6866 , n6869 );
not ( n6871 , n5399 );
not ( n6872 , n5891 );
or ( n6873 , n6871 , n6872 );
not ( n6874 , n545 );
not ( n6875 , n5701 );
not ( n6876 , n6875 );
or ( n6877 , n6874 , n6876 );
nand ( n6878 , n5701 , n4440 );
nand ( n6879 , n6877 , n6878 );
nand ( n6880 , n6879 , n5137 );
nand ( n6881 , n6873 , n6880 );
not ( n6882 , n5501 );
not ( n6883 , n5799 );
or ( n6884 , n6882 , n6883 );
not ( n6885 , n537 );
or ( n6886 , n6885 , n5822 );
nand ( n6887 , n5822 , n5409 );
nand ( n6888 , n6886 , n6887 );
nand ( n6889 , n6888 , n5413 );
nand ( n6890 , n6884 , n6889 );
not ( n6891 , n6890 );
not ( n6892 , n70470 );
nand ( n6893 , n5811 , n965 );
xor ( n6894 , n6893 , n5808 );
not ( n6895 , n6894 );
or ( n6896 , n6892 , n6895 );
and ( n6897 , n4206 , n3898 );
nor ( n6898 , n6897 , n4207 );
not ( n6899 , n6898 );
buf ( n6900 , n4085 );
nand ( n6901 , n3903 , n3929 );
buf ( n6902 , n6901 );
nand ( n6903 , n6900 , n6902 );
or ( n6904 , n6899 , n6903 );
not ( n76754 , n6898 );
nand ( n76755 , n76754 , n6903 );
nand ( n6907 , n6904 , n76755 , n455 );
nand ( n6908 , n6896 , n6907 );
buf ( n6909 , n6908 );
not ( n6910 , n6909 );
nand ( n6911 , n6910 , n537 );
nor ( n6912 , n6891 , n6911 );
not ( n6913 , n4433 );
not ( n6914 , n5792 );
or ( n6915 , n6913 , n6914 );
not ( n6916 , n5723 );
and ( n6917 , n539 , n6916 );
not ( n6918 , n539 );
and ( n6919 , n6918 , n5723 );
nor ( n6920 , n6917 , n6919 );
not ( n6921 , n6920 );
nand ( n6922 , n6921 , n4224 );
nand ( n6923 , n6915 , n6922 );
xor ( n6924 , n6912 , n6923 );
xor ( n6925 , n5805 , n5825 );
xor ( n6926 , n6924 , n6925 );
xor ( n6927 , n6881 , n6926 );
not ( n6928 , n6811 );
and ( n6929 , n5264 , n547 );
not ( n6930 , n5264 );
and ( n6931 , n6930 , n6857 );
nor ( n6932 , n6929 , n6931 );
not ( n6933 , n6932 );
or ( n6934 , n6928 , n6933 );
and ( n6935 , n547 , n5123 );
not ( n6936 , n547 );
buf ( n6937 , n74998 );
and ( n6938 , n6936 , n6937 );
nor ( n6939 , n6935 , n6938 );
not ( n6940 , n6939 );
nand ( n6941 , n6940 , n6854 );
nand ( n6942 , n6934 , n6941 );
and ( n6943 , n6927 , n6942 );
and ( n6944 , n6881 , n6926 );
or ( n6945 , n6943 , n6944 );
xor ( n6946 , n6870 , n6945 );
xor ( n6947 , n6912 , n6923 );
and ( n6948 , n6947 , n6925 );
and ( n6949 , n6912 , n6923 );
or ( n6950 , n6948 , n6949 );
not ( n76800 , n6811 );
not ( n6952 , n6859 );
or ( n6953 , n76800 , n6952 );
not ( n6954 , n6854 );
not ( n6955 , n6954 );
nand ( n6956 , n6932 , n6955 );
nand ( n6957 , n6953 , n6956 );
xor ( n6958 , n6950 , n6957 );
not ( n6959 , n6911 );
not ( n6960 , n6890 );
not ( n6961 , n6960 );
or ( n6962 , n6959 , n6961 );
not ( n6963 , n6911 );
nand ( n6964 , n6963 , n6890 );
nand ( n6965 , n6962 , n6964 );
not ( n6966 , n6920 );
not ( n6967 , n5780 );
and ( n6968 , n6966 , n6967 );
not ( n76818 , n539 );
not ( n6970 , n5448 );
or ( n6971 , n76818 , n6970 );
not ( n6972 , n70470 );
not ( n6973 , n5428 );
or ( n6974 , n6972 , n6973 );
nand ( n6975 , n6974 , n5447 );
not ( n6976 , n6975 );
nand ( n6977 , n6976 , n4251 );
nand ( n6978 , n6971 , n6977 );
and ( n6979 , n6978 , n4224 );
nor ( n6980 , n6968 , n6979 );
nor ( n6981 , n6965 , n6980 );
not ( n6982 , n5128 );
not ( n6983 , n5871 );
or ( n6984 , n6982 , n6983 );
not ( n6985 , n4938 );
not ( n6986 , n4429 );
or ( n6987 , n6985 , n6986 );
nand ( n6988 , n4424 , n543 );
nand ( n6989 , n6987 , n6988 );
nand ( n6990 , n6989 , n4445 );
nand ( n6991 , n6984 , n6990 );
xor ( n6992 , n6981 , n6991 );
not ( n6993 , n5590 );
not ( n76843 , n5880 );
or ( n6995 , n6993 , n76843 );
and ( n6996 , n5538 , n5779 );
not ( n6997 , n5538 );
and ( n6998 , n6997 , n5753 );
nor ( n6999 , n6996 , n6998 );
nand ( n7000 , n6999 , n5551 );
nand ( n7001 , n6995 , n7000 );
and ( n7002 , n6992 , n7001 );
and ( n7003 , n6981 , n6991 );
or ( n7004 , n7002 , n7003 );
xor ( n7005 , n6958 , n7004 );
and ( n7006 , n6946 , n7005 );
and ( n7007 , n6870 , n6945 );
or ( n7008 , n7006 , n7007 );
and ( n7009 , n6863 , n7008 );
and ( n7010 , n5904 , n76711 );
or ( n7011 , n7009 , n7010 );
xor ( n7012 , n5902 , n7011 );
xor ( n7013 , n6491 , n6804 );
and ( n7014 , n7013 , n6861 );
and ( n7015 , n6491 , n6804 );
or ( n7016 , n7014 , n7015 );
not ( n7017 , n5905 );
not ( n7018 , n549 );
nor ( n7019 , n7017 , n7018 );
not ( n7020 , n7019 );
not ( n7021 , n7020 );
not ( n7022 , n76644 );
not ( n7023 , n7022 );
or ( n76873 , n7021 , n7023 );
nor ( n7025 , n7017 , n549 );
or ( n7026 , n7022 , n7025 );
nand ( n7027 , n76873 , n7026 );
nand ( n7028 , n6441 , n6489 );
nand ( n7029 , n7027 , n7028 );
not ( n7030 , n6802 );
not ( n7031 , n6756 );
or ( n7032 , n7030 , n7031 );
not ( n7033 , n6752 );
not ( n7034 , n6638 );
not ( n7035 , n6679 );
and ( n7036 , n7034 , n7035 );
nor ( n7037 , n7036 , n6740 );
not ( n7038 , n7037 );
nor ( n7039 , n7038 , n6634 );
not ( n7040 , n7039 );
not ( n7041 , n4203 );
or ( n76891 , n7040 , n7041 );
and ( n7046 , n6696 , n7037 );
nor ( n76893 , n76588 , n6735 );
or ( n7048 , n76893 , n6698 );
nand ( n7049 , n7048 , n6742 );
nor ( n7050 , n7046 , n7049 );
nand ( n7051 , n76891 , n7050 );
not ( n7052 , n7051 );
xor ( n7053 , n6716 , n6729 );
and ( n7054 , n7053 , n6734 );
and ( n7055 , n6716 , n6729 );
or ( n7056 , n7054 , n7055 );
xor ( n7057 , n76552 , n6713 );
and ( n7058 , n7057 , n6715 );
and ( n7059 , n76552 , n6713 );
or ( n7060 , n7058 , n7059 );
not ( n7061 , n1828 );
not ( n7062 , n6718 );
or ( n7063 , n7061 , n7062 );
not ( n7064 , n489 );
not ( n7065 , n1874 );
or ( n7066 , n7064 , n7065 );
nand ( n7067 , n1995 , n1649 );
nand ( n7068 , n7066 , n7067 );
nand ( n7069 , n7068 , n71761 );
nand ( n7070 , n7063 , n7069 );
and ( n76917 , n489 , n1982 );
xor ( n7075 , n7070 , n76917 );
not ( n7076 , n6711 );
not ( n7077 , n7076 );
not ( n7078 , n1699 );
and ( n7079 , n7077 , n7078 );
and ( n7080 , n1739 , n491 );
nor ( n7081 , n7079 , n7080 );
xor ( n76925 , n7075 , n7081 );
xor ( n76926 , n7060 , n76925 );
xor ( n7084 , n6722 , n6723 );
and ( n7085 , n7084 , n6728 );
and ( n7086 , n6722 , n6723 );
or ( n7087 , n7085 , n7086 );
xor ( n7088 , n76926 , n7087 );
or ( n7089 , n7056 , n7088 );
nand ( n76933 , n7056 , n7088 );
nand ( n76934 , n7089 , n76933 );
and ( n7092 , n76934 , n455 );
nand ( n7093 , n7052 , n7092 );
nor ( n7094 , n6566 , n6620 );
not ( n7095 , n7094 );
not ( n7096 , n6771 );
or ( n7097 , n7095 , n7096 );
or ( n7098 , n6569 , n6620 );
nand ( n7099 , n7098 , n6622 );
not ( n7100 , n7099 );
nand ( n7101 , n7097 , n7100 );
not ( n7102 , n7101 );
not ( n7103 , n6600 );
nand ( n7104 , n7103 , n6536 );
not ( n76948 , n7104 );
not ( n7106 , n6608 );
or ( n7107 , n76948 , n7106 );
nand ( n7108 , n6535 , n6600 );
nand ( n7109 , n7107 , n7108 );
and ( n7110 , n508 , n489 );
xor ( n7111 , n489 , n506 );
not ( n7112 , n7111 );
not ( n7113 , n1553 );
or ( n7114 , n7112 , n7113 );
not ( n7115 , n6598 );
nand ( n7116 , n7115 , n6384 );
nand ( n7117 , n7114 , n7116 );
xor ( n7118 , n7110 , n7117 );
not ( n7119 , n6580 );
not ( n7120 , n6586 );
and ( n7121 , n7119 , n7120 );
and ( n7122 , n1630 , n491 );
nor ( n7123 , n7121 , n7122 );
xor ( n7124 , n7118 , n7123 );
xor ( n7125 , n6579 , n6588 );
and ( n7126 , n7125 , n6593 );
and ( n7127 , n6579 , n6588 );
or ( n7128 , n7126 , n7127 );
and ( n7129 , n7124 , n7128 );
not ( n7130 , n7124 );
not ( n7131 , n7128 );
and ( n7132 , n7130 , n7131 );
nor ( n7133 , n7129 , n7132 );
xor ( n7134 , n7109 , n7133 );
not ( n7135 , n7134 );
not ( n7136 , n6618 );
not ( n7137 , n7136 );
not ( n7138 , n6594 );
not ( n7139 , n7138 );
and ( n7140 , n7137 , n7139 );
nand ( n7141 , n7136 , n7138 );
not ( n7142 , n6613 );
and ( n7143 , n7141 , n7142 );
nor ( n76987 , n7140 , n7143 );
nand ( n76988 , n7135 , n76987 );
not ( n7146 , n7134 );
nor ( n7147 , n7146 , n76987 );
not ( n7148 , n7147 );
nand ( n7149 , n76988 , n7148 );
not ( n7150 , n7149 );
nor ( n7151 , n7150 , n455 );
nand ( n7152 , n7102 , n7151 );
not ( n7153 , n76934 );
and ( n7154 , n7153 , n455 );
nand ( n7155 , n7051 , n7154 );
not ( n7156 , n74671 );
nor ( n7157 , n7156 , n7149 );
nand ( n7158 , n7157 , n7101 );
nand ( n7159 , n7093 , n7152 , n7155 , n7158 );
not ( n7160 , n7159 );
not ( n7161 , n7160 );
or ( n7162 , n7033 , n7161 );
or ( n7163 , n7160 , n6752 );
nand ( n7164 , n7162 , n7163 );
nand ( n7165 , n7164 , n552 );
nand ( n7166 , n7032 , n7165 );
xor ( n7167 , n7029 , n7166 );
not ( n7168 , n6955 );
not ( n7169 , n6850 );
or ( n7170 , n7168 , n7169 );
not ( n7171 , n6462 );
not ( n7172 , n6458 );
or ( n7173 , n7171 , n7172 );
nand ( n7174 , n7173 , n6477 );
not ( n7175 , n7174 );
and ( n7176 , n547 , n7175 );
not ( n77020 , n547 );
and ( n77021 , n77020 , n6478 );
or ( n7179 , n7176 , n77021 );
nand ( n7180 , n7179 , n6811 );
nand ( n7181 , n7170 , n7180 );
xor ( n7182 , n7167 , n7181 );
xor ( n7183 , n7016 , n7182 );
xor ( n7184 , n5778 , n5837 );
xor ( n77028 , n7184 , n5850 );
xor ( n77029 , n6950 , n6957 );
and ( n7187 , n77029 , n7004 );
and ( n7188 , n6950 , n6957 );
or ( n7189 , n7187 , n7188 );
xor ( n7190 , n77028 , n7189 );
xor ( n7191 , n5794 , n5826 );
xor ( n7192 , n7191 , n5834 );
xor ( n7193 , n5875 , n5884 );
xor ( n7194 , n7193 , n5895 );
xor ( n7195 , n7192 , n7194 );
not ( n7196 , n6489 );
and ( n7197 , n549 , n6843 );
not ( n7198 , n549 );
and ( n7199 , n7198 , n6847 );
nor ( n7200 , n7197 , n7199 );
not ( n7201 , n7200 );
or ( n7202 , n7196 , n7201 );
nand ( n77046 , n6484 , n5905 );
nand ( n7204 , n7202 , n77046 );
and ( n7205 , n7195 , n7204 );
and ( n7206 , n7192 , n7194 );
or ( n7207 , n7205 , n7206 );
and ( n7208 , n7190 , n7207 );
and ( n7209 , n77028 , n7189 );
or ( n7210 , n7208 , n7209 );
xor ( n7211 , n7183 , n7210 );
xor ( n7212 , n7012 , n7211 );
not ( n7213 , n7212 );
xor ( n7214 , n77028 , n7189 );
xor ( n7215 , n7214 , n7207 );
not ( n7216 , n5589 );
not ( n7217 , n6999 );
or ( n7218 , n7216 , n7217 );
not ( n7219 , n5626 );
not ( n7220 , n7219 );
not ( n7221 , n5538 );
or ( n7222 , n7220 , n7221 );
nand ( n7223 , n5628 , n541 );
nand ( n7224 , n7222 , n7223 );
nand ( n7225 , n7224 , n5551 );
nand ( n7226 , n7218 , n7225 );
not ( n7227 , n5128 );
not ( n7228 , n6989 );
or ( n7229 , n7227 , n7228 );
nand ( n7230 , n4444 , n543 );
not ( n7231 , n7230 );
not ( n7232 , n4247 );
and ( n7233 , n7231 , n7232 );
buf ( n7234 , n4247 );
not ( n7235 , n4444 );
nor ( n7236 , n7235 , n543 );
and ( n7237 , n7234 , n7236 );
nor ( n7238 , n7233 , n7237 );
nand ( n7239 , n7229 , n7238 );
xor ( n7240 , n7226 , n7239 );
not ( n7241 , n5413 );
not ( n7242 , n5409 );
not ( n7243 , n6909 );
not ( n7244 , n7243 );
or ( n7245 , n7242 , n7244 );
nand ( n7246 , n537 , n6909 );
nand ( n7247 , n7245 , n7246 );
not ( n7248 , n7247 );
or ( n7249 , n7241 , n7248 );
nand ( n7250 , n6888 , n5501 );
nand ( n7251 , n7249 , n7250 );
not ( n7252 , n824 );
nand ( n7253 , n7252 , n901 );
not ( n7254 , n455 );
nand ( n7255 , n7253 , n889 , n897 , n7254 );
nand ( n7256 , n3932 , n3958 );
not ( n7257 , n7256 );
not ( n7258 , n3959 );
not ( n7259 , n4074 );
not ( n7260 , n4078 );
or ( n7261 , n7259 , n7260 );
nand ( n7262 , n7261 , n4077 );
nand ( n7263 , n7258 , n7262 );
not ( n7264 , n7263 );
or ( n7265 , n7257 , n7264 );
nor ( n7266 , n7254 , n73847 );
and ( n7267 , n6901 , n7266 );
nand ( n7268 , n7265 , n7267 );
not ( n7269 , n73847 );
nand ( n7270 , n7269 , n6901 );
nand ( n7271 , n7270 , n7256 , n455 , n7263 );
not ( n7272 , n7253 );
nand ( n77116 , n889 , n897 );
nand ( n7274 , n7272 , n77116 , n7254 );
nand ( n7275 , n7255 , n7268 , n7271 , n7274 );
not ( n7276 , n7275 );
not ( n7277 , n7276 );
not ( n7278 , n7277 );
and ( n7279 , n7278 , n537 );
xor ( n7280 , n7251 , n7279 );
not ( n7281 , n4433 );
not ( n7282 , n6978 );
or ( n7283 , n7281 , n7282 );
not ( n7284 , n539 );
not ( n7285 , n5530 );
or ( n7286 , n7284 , n7285 );
nand ( n7287 , n5531 , n4251 );
nand ( n7288 , n7286 , n7287 );
nand ( n7289 , n7288 , n4224 );
nand ( n7290 , n7283 , n7289 );
and ( n7291 , n7280 , n7290 );
and ( n7292 , n7251 , n7279 );
or ( n7293 , n7291 , n7292 );
and ( n7294 , n7240 , n7293 );
and ( n7295 , n7226 , n7239 );
or ( n7296 , n7294 , n7295 );
xor ( n7297 , n6981 , n6991 );
xor ( n77141 , n7297 , n7001 );
xor ( n7299 , n7296 , n77141 );
not ( n7300 , n5905 );
not ( n7301 , n7200 );
or ( n7302 , n7300 , n7301 );
not ( n7303 , n5392 );
not ( n7304 , n7303 );
nor ( n7305 , n6488 , n549 );
and ( n7306 , n7304 , n7305 );
nor ( n7307 , n6488 , n7018 );
and ( n7308 , n7303 , n7307 );
nor ( n7309 , n7306 , n7308 );
nand ( n7310 , n7302 , n7309 );
and ( n7311 , n7299 , n7310 );
and ( n7312 , n7296 , n77141 );
or ( n7313 , n7311 , n7312 );
xor ( n7314 , n7192 , n7194 );
xor ( n7315 , n7314 , n7204 );
xor ( n7316 , n7313 , n7315 );
not ( n7317 , n551 );
not ( n7318 , n7174 );
not ( n7319 , n7318 );
or ( n7320 , n7317 , n7319 );
nand ( n7321 , n6478 , n6752 );
nand ( n77165 , n7320 , n7321 );
nand ( n77166 , n77165 , n6802 );
not ( n7324 , n6440 );
nor ( n7325 , n6752 , n6801 );
nand ( n7326 , n7324 , n7325 );
not ( n7327 , n7324 );
nor ( n7328 , n6801 , n551 );
nand ( n7329 , n7327 , n7328 );
nand ( n7330 , n77166 , n7326 , n7329 );
not ( n7331 , n5137 );
not ( n7332 , n545 );
not ( n7333 , n5869 );
not ( n7334 , n7333 );
or ( n7335 , n7332 , n7334 );
not ( n7336 , n5866 );
nand ( n7337 , n7336 , n4440 );
nand ( n7338 , n7335 , n7337 );
not ( n7339 , n7338 );
or ( n7340 , n7331 , n7339 );
nand ( n7341 , n5399 , n6879 );
nand ( n7342 , n7340 , n7341 );
xor ( n7343 , n6965 , n6980 );
xor ( n7344 , n7342 , n7343 );
and ( n7345 , n547 , n4933 );
not ( n7346 , n547 );
and ( n7347 , n7346 , n4937 );
or ( n77191 , n7345 , n7347 );
not ( n7349 , n77191 );
or ( n7350 , n7349 , n6954 );
or ( n7351 , n6939 , n6810 );
nand ( n7352 , n7350 , n7351 );
and ( n7353 , n7344 , n7352 );
and ( n7354 , n7342 , n7343 );
or ( n7355 , n7353 , n7354 );
xor ( n7356 , n7330 , n7355 );
xor ( n7357 , n6881 , n6926 );
xor ( n7358 , n7357 , n6942 );
and ( n7359 , n7356 , n7358 );
and ( n7360 , n7330 , n7355 );
or ( n7361 , n7359 , n7360 );
and ( n7362 , n7316 , n7361 );
and ( n7363 , n7313 , n7315 );
or ( n7364 , n7362 , n7363 );
xor ( n7365 , n7215 , n7364 );
xor ( n7366 , n5904 , n76711 );
xor ( n7367 , n7366 , n7008 );
and ( n7368 , n7365 , n7367 );
and ( n7369 , n7215 , n7364 );
or ( n7370 , n7368 , n7369 );
not ( n7371 , n7370 );
and ( n7372 , n7213 , n7371 );
xor ( n7373 , n7215 , n7364 );
xor ( n7374 , n7373 , n7367 );
not ( n7375 , n7374 );
xor ( n7376 , n6870 , n6945 );
xor ( n7377 , n7376 , n7005 );
not ( n7378 , n5264 );
nand ( n7379 , n7378 , n7307 );
nand ( n7380 , n5393 , n7019 );
nand ( n77224 , n5392 , n7025 );
nand ( n7382 , n5264 , n7305 );
nand ( n7383 , n7379 , n7380 , n77224 , n7382 );
not ( n7384 , n5501 );
not ( n7385 , n7247 );
or ( n7386 , n7384 , n7385 );
not ( n7387 , n537 );
not ( n7388 , n7275 );
or ( n7389 , n7387 , n7388 );
nand ( n7390 , n7276 , n5409 );
nand ( n7391 , n7389 , n7390 );
nand ( n7392 , n7391 , n5413 );
nand ( n7393 , n7386 , n7392 );
buf ( n7394 , n7262 );
nand ( n7395 , n7258 , n7256 );
not ( n7396 , n7395 );
and ( n7397 , n7394 , n7396 );
not ( n7398 , n7394 );
and ( n7399 , n7398 , n7395 );
nor ( n7400 , n7397 , n7399 );
and ( n7401 , n455 , n7400 );
not ( n7402 , n455 );
not ( n7403 , n762 );
buf ( n7404 , n751 );
not ( n7405 , n7404 );
or ( n7406 , n7403 , n7405 );
nand ( n7407 , n7406 , n745 );
nand ( n7408 , n822 , n901 );
or ( n7409 , n7407 , n7408 );
nand ( n7410 , n7407 , n7408 );
nand ( n7411 , n7409 , n7410 );
and ( n7412 , n7402 , n7411 );
nor ( n7413 , n7401 , n7412 );
not ( n7414 , n7413 );
and ( n7415 , n7414 , n537 );
xor ( n77259 , n7393 , n7415 );
not ( n7417 , n4434 );
not ( n7418 , n7288 );
or ( n7419 , n7417 , n7418 );
not ( n7420 , n539 );
not ( n7421 , n5822 );
not ( n7422 , n7421 );
or ( n7423 , n7420 , n7422 );
nand ( n7424 , n5822 , n4251 );
nand ( n7425 , n7423 , n7424 );
nand ( n7426 , n7425 , n4224 );
nand ( n7427 , n7419 , n7426 );
and ( n7428 , n77259 , n7427 );
and ( n7429 , n7393 , n7415 );
or ( n7430 , n7428 , n7429 );
not ( n7431 , n541 );
not ( n7432 , n6916 );
or ( n7433 , n7431 , n7432 );
nand ( n7434 , n5538 , n5495 );
nand ( n7435 , n7433 , n7434 );
not ( n77279 , n7435 );
not ( n7437 , n5551 );
or ( n7438 , n77279 , n7437 );
not ( n7439 , n7224 );
not ( n7440 , n5590 );
or ( n7441 , n7439 , n7440 );
nand ( n7442 , n7438 , n7441 );
xor ( n7443 , n7430 , n7442 );
nand ( n7444 , n4443 , n543 );
or ( n7445 , n7444 , n7234 );
not ( n7446 , n74151 );
not ( n7447 , n4443 );
nor ( n7448 , n7447 , n543 );
nand ( n7449 , n7446 , n7448 );
not ( n7450 , n543 );
not ( n7451 , n5753 );
not ( n7452 , n7451 );
or ( n7453 , n7450 , n7452 );
nand ( n7454 , n5753 , n4938 );
nand ( n7455 , n7453 , n7454 );
nand ( n7456 , n7455 , n4445 );
nand ( n7457 , n7445 , n7449 , n7456 );
and ( n7458 , n7443 , n7457 );
and ( n7459 , n7430 , n7442 );
or ( n7460 , n7458 , n7459 );
xor ( n7461 , n7383 , n7460 );
xor ( n7462 , n7251 , n7279 );
xor ( n7463 , n7462 , n7290 );
not ( n7464 , n5399 );
not ( n7465 , n7338 );
or ( n7466 , n7464 , n7465 );
not ( n7467 , n545 );
not ( n77311 , n5535 );
or ( n7472 , n7467 , n77311 );
nand ( n77313 , n4429 , n4440 );
nand ( n7474 , n7472 , n77313 );
nand ( n7475 , n7474 , n5137 );
nand ( n7476 , n7466 , n7475 );
xor ( n7477 , n7463 , n7476 );
not ( n7478 , n7435 );
not ( n7479 , n5588 );
or ( n7480 , n7478 , n7479 );
not ( n7481 , n541 );
not ( n7482 , n6975 );
or ( n7483 , n7481 , n7482 );
nand ( n7484 , n5538 , n5642 , n5447 );
nand ( n7485 , n7483 , n7484 );
nand ( n7486 , n7485 , n5551 );
nand ( n7487 , n7480 , n7486 );
not ( n7488 , n5501 );
not ( n7489 , n7391 );
or ( n7490 , n7488 , n7489 );
and ( n7491 , n7414 , n537 );
not ( n7492 , n7414 );
and ( n7493 , n7492 , n6885 );
nor ( n7494 , n7491 , n7493 );
nand ( n7495 , n7494 , n5413 );
nand ( n7496 , n7490 , n7495 );
not ( n77337 , n455 );
not ( n7501 , n4074 );
not ( n7502 , n4078 );
or ( n7503 , n7501 , n7502 );
nand ( n7504 , n7503 , n4076 );
not ( n7505 , n4036 );
not ( n7506 , n4061 );
or ( n7507 , n7505 , n7506 );
nand ( n7508 , n7507 , n4066 );
not ( n7509 , n7508 );
and ( n7510 , n7504 , n7509 );
not ( n7511 , n7504 );
and ( n7512 , n7511 , n7508 );
nor ( n7513 , n7510 , n7512 );
not ( n7514 , n7513 );
or ( n7515 , n77337 , n7514 );
not ( n7516 , n724 );
not ( n7517 , n7516 );
not ( n7518 , n760 );
not ( n7519 , n730 );
and ( n7520 , n7518 , n7519 );
and ( n77358 , n760 , n730 );
nor ( n77359 , n7520 , n77358 );
not ( n7523 , n77359 );
not ( n7524 , n7523 );
or ( n7525 , n7517 , n7524 );
not ( n7526 , n7516 );
nand ( n7527 , n7526 , n77359 );
nand ( n7528 , n7525 , n7527 );
and ( n77366 , n7528 , n7404 );
not ( n77367 , n7528 );
not ( n7531 , n7404 );
and ( n7532 , n77367 , n7531 );
nor ( n7533 , n77366 , n7532 );
nand ( n7534 , n7533 , n70470 );
nand ( n7535 , n7515 , n7534 );
buf ( n7536 , n7535 );
buf ( n7537 , n7536 );
and ( n7538 , n7537 , n537 );
xor ( n7539 , n7496 , n7538 );
not ( n7540 , n4434 );
not ( n7541 , n7425 );
or ( n7542 , n7540 , n7541 );
or ( n7543 , n539 , n6909 );
nand ( n7544 , n6909 , n539 );
nand ( n7545 , n7543 , n7544 );
nand ( n7546 , n7545 , n4224 );
nand ( n7547 , n7542 , n7546 );
and ( n7548 , n7539 , n7547 );
and ( n7549 , n7496 , n7538 );
or ( n7550 , n7548 , n7549 );
xor ( n77388 , n7487 , n7550 );
not ( n7552 , n4445 );
not ( n7553 , n543 );
not ( n7554 , n7219 );
not ( n7555 , n7554 );
or ( n7556 , n7553 , n7555 );
nand ( n7557 , n7219 , n4938 );
nand ( n7558 , n7556 , n7557 );
not ( n7559 , n7558 );
or ( n7560 , n7552 , n7559 );
nand ( n7561 , n7455 , n5128 );
nand ( n7562 , n7560 , n7561 );
and ( n7563 , n77388 , n7562 );
and ( n7564 , n7487 , n7550 );
or ( n7565 , n7563 , n7564 );
and ( n7566 , n7477 , n7565 );
and ( n7567 , n7463 , n7476 );
or ( n7568 , n7566 , n7567 );
and ( n7569 , n7461 , n7568 );
and ( n7570 , n7383 , n7460 );
or ( n7571 , n7569 , n7570 );
xor ( n7572 , n7296 , n77141 );
xor ( n7573 , n7572 , n7310 );
xor ( n7574 , n7571 , n7573 );
xor ( n7575 , n7226 , n7239 );
xor ( n7576 , n7575 , n7293 );
not ( n7577 , n6802 );
and ( n7578 , n6844 , n551 );
not ( n7579 , n6844 );
and ( n7580 , n7579 , n6752 );
or ( n7581 , n7578 , n7580 );
not ( n7582 , n7581 );
or ( n7583 , n7577 , n7582 );
nand ( n7584 , n77165 , n552 );
nand ( n77422 , n7583 , n7584 );
xor ( n77423 , n7576 , n77422 );
xor ( n7587 , n7342 , n7343 );
xor ( n7588 , n7587 , n7352 );
and ( n7589 , n77423 , n7588 );
and ( n7590 , n7576 , n77422 );
or ( n7591 , n7589 , n7590 );
and ( n7592 , n7574 , n7591 );
and ( n7593 , n7571 , n7573 );
or ( n7594 , n7592 , n7593 );
xor ( n7595 , n7377 , n7594 );
xor ( n7596 , n7313 , n7315 );
xor ( n7597 , n7596 , n7361 );
and ( n7598 , n7595 , n7597 );
and ( n7599 , n7377 , n7594 );
or ( n7600 , n7598 , n7599 );
not ( n7601 , n7600 );
and ( n7602 , n7375 , n7601 );
nor ( n7603 , n7372 , n7602 );
not ( n7604 , n7603 );
xor ( n7605 , n7576 , n77422 );
xor ( n7606 , n7605 , n7588 );
not ( n7607 , n552 );
not ( n7608 , n7581 );
or ( n7609 , n7607 , n7608 );
not ( n7610 , n551 );
not ( n7611 , n7303 );
or ( n7612 , n7610 , n7611 );
nand ( n77450 , n5392 , n6752 );
nand ( n77451 , n7612 , n77450 );
nand ( n7615 , n77451 , n6802 );
nand ( n7616 , n7609 , n7615 );
not ( n7617 , n6811 );
not ( n7618 , n77191 );
or ( n7619 , n7617 , n7618 );
not ( n7620 , n5843 );
buf ( n77458 , n7620 );
nor ( n77459 , n6954 , n547 );
and ( n7623 , n77458 , n77459 );
not ( n7624 , n7620 );
not ( n7625 , n547 );
nor ( n7626 , n7625 , n6954 );
and ( n7627 , n7624 , n7626 );
nor ( n7628 , n7623 , n7627 );
nand ( n7629 , n7619 , n7628 );
xor ( n7630 , n7393 , n7415 );
xor ( n7631 , n7630 , n7427 );
nand ( n7632 , n7333 , n7626 );
not ( n7633 , n5843 );
nor ( n7634 , n6810 , n547 );
nand ( n7635 , n7633 , n7634 );
nand ( n7636 , n5869 , n77459 );
nand ( n7637 , n6811 , n547 );
not ( n7638 , n7637 );
nand ( n7639 , n7638 , n6875 );
nand ( n7640 , n7632 , n7635 , n7636 , n7639 );
xor ( n7641 , n7631 , n7640 );
and ( n7642 , n4247 , n4440 );
not ( n7643 , n4247 );
and ( n7644 , n7643 , n545 );
or ( n7645 , n7642 , n7644 );
not ( n7646 , n7645 );
or ( n7647 , n7646 , n75017 );
not ( n7648 , n7474 );
not ( n7649 , n5399 );
or ( n7650 , n7648 , n7649 );
nand ( n7651 , n7647 , n7650 );
and ( n7652 , n7641 , n7651 );
and ( n7653 , n7631 , n7640 );
or ( n7654 , n7652 , n7653 );
xor ( n7655 , n7629 , n7654 );
xor ( n7656 , n7430 , n7442 );
xor ( n7657 , n7656 , n7457 );
xor ( n77495 , n7655 , n7657 );
xor ( n7659 , n7616 , n77495 );
not ( n7660 , n6802 );
not ( n7661 , n551 );
not ( n7662 , n5265 );
or ( n7663 , n7661 , n7662 );
nand ( n7664 , n6752 , n5264 );
nand ( n7665 , n7663 , n7664 );
not ( n7666 , n7665 );
or ( n7667 , n7660 , n7666 );
nand ( n7668 , n77451 , n552 );
nand ( n7669 , n7667 , n7668 );
not ( n7670 , n5128 );
not ( n7671 , n7558 );
or ( n7672 , n7670 , n7671 );
not ( n7673 , n543 );
not ( n7674 , n6916 );
or ( n7675 , n7673 , n7674 );
nand ( n7676 , n4938 , n5495 );
nand ( n7677 , n7675 , n7676 );
nand ( n7678 , n7677 , n4445 );
nand ( n7679 , n7672 , n7678 );
not ( n7680 , n70419 );
nand ( n7681 , n7680 , n70423 );
not ( n7682 , n70386 );
and ( n7683 , n7681 , n7682 );
not ( n7684 , n7681 );
and ( n7685 , n7684 , n70386 );
nor ( n7686 , n7683 , n7685 );
nand ( n7687 , n7686 , n70470 );
nand ( n7688 , n4035 , n4004 );
not ( n7689 , n7688 );
nor ( n7690 , n4030 , n5595 );
and ( n7691 , n7689 , n7690 );
and ( n7692 , n4030 , n455 );
and ( n7693 , n7692 , n7688 );
nor ( n7694 , n7691 , n7693 );
nand ( n7695 , n7687 , n7694 );
buf ( n7696 , n7695 );
and ( n7697 , n537 , n7696 );
not ( n7698 , n5501 );
not ( n7699 , n537 );
not ( n7700 , n7536 );
not ( n7701 , n7700 );
or ( n7702 , n7699 , n7701 );
nand ( n7703 , n7536 , n5409 );
nand ( n7704 , n7702 , n7703 );
not ( n7705 , n7704 );
or ( n7706 , n7698 , n7705 );
not ( n7707 , n4065 );
not ( n7708 , n4064 );
or ( n7709 , n7707 , n7708 );
nand ( n7710 , n7709 , n4061 );
not ( n7711 , n7710 );
buf ( n7712 , n4036 );
nand ( n7713 , n7711 , n7712 );
not ( n7714 , n7712 );
nand ( n7715 , n7710 , n7714 );
nand ( n7716 , n7713 , n7715 , n455 );
nand ( n7717 , n7716 , n70471 );
buf ( n7718 , n7717 );
xor ( n7719 , n537 , n7718 );
nand ( n7720 , n7719 , n5413 );
nand ( n7721 , n7706 , n7720 );
xor ( n7722 , n7697 , n7721 );
not ( n7723 , n5501 );
not ( n7724 , n7719 );
or ( n7725 , n7723 , n7724 );
xor ( n7726 , n537 , n7696 );
nand ( n7727 , n7726 , n5413 );
nand ( n7728 , n7725 , n7727 );
not ( n7729 , n7728 );
not ( n7730 , n5403 );
not ( n7731 , n7696 );
not ( n7732 , n7731 );
or ( n7733 , n7730 , n7732 );
nand ( n7734 , n7733 , n539 );
not ( n7735 , n7696 );
not ( n7736 , n7735 );
and ( n7737 , n7736 , n538 );
nor ( n7738 , n7737 , n5409 );
nand ( n7739 , n7734 , n7738 );
nor ( n7740 , n7729 , n7739 );
and ( n7741 , n7722 , n7740 );
and ( n7742 , n7697 , n7721 );
or ( n7743 , n7741 , n7742 );
not ( n7744 , n5550 );
not ( n7745 , n541 );
not ( n7746 , n7421 );
or ( n7747 , n7745 , n7746 );
nand ( n7748 , n5822 , n5538 );
nand ( n7749 , n7747 , n7748 );
not ( n77587 , n7749 );
or ( n77588 , n7744 , n77587 );
not ( n7752 , n541 );
not ( n7753 , n5530 );
or ( n7754 , n7752 , n7753 );
not ( n7755 , n5516 );
nor ( n7756 , n5527 , n455 );
not ( n7757 , n7756 );
nand ( n7758 , n7755 , n7757 , n5538 );
nand ( n7759 , n7754 , n7758 );
nand ( n7760 , n7759 , n5545 );
nand ( n7761 , n77588 , n7760 );
xor ( n7762 , n7743 , n7761 );
and ( n7763 , n537 , n7718 );
not ( n7764 , n5501 );
not ( n7765 , n7494 );
or ( n7766 , n7764 , n7765 );
nand ( n7767 , n7704 , n5413 );
nand ( n7768 , n7766 , n7767 );
xor ( n7769 , n7763 , n7768 );
not ( n7770 , n4434 );
not ( n7771 , n7545 );
or ( n7772 , n7770 , n7771 );
not ( n7773 , n539 );
not ( n7774 , n7275 );
or ( n7775 , n7773 , n7774 );
nand ( n7776 , n7276 , n4251 );
nand ( n7777 , n7775 , n7776 );
nand ( n7778 , n7777 , n4224 );
nand ( n7779 , n7772 , n7778 );
xor ( n7780 , n7769 , n7779 );
and ( n7781 , n7762 , n7780 );
and ( n7782 , n7743 , n7761 );
or ( n7783 , n7781 , n7782 );
xor ( n7784 , n7679 , n7783 );
not ( n7785 , n6811 );
not ( n7786 , n5866 );
and ( n7787 , n547 , n7786 );
not ( n7788 , n547 );
buf ( n7789 , n5866 );
and ( n7790 , n7788 , n7789 );
nor ( n7791 , n7787 , n7790 );
not ( n7792 , n7791 );
or ( n7793 , n7785 , n7792 );
not ( n7794 , n547 );
not ( n7795 , n5535 );
or ( n7796 , n7794 , n7795 );
not ( n7797 , n547 );
not ( n7798 , n4424 );
nand ( n7799 , n7797 , n7798 );
nand ( n7800 , n7796 , n7799 );
nand ( n7801 , n7800 , n6955 );
nand ( n7802 , n7793 , n7801 );
and ( n7803 , n7784 , n7802 );
and ( n7804 , n7679 , n7783 );
or ( n7805 , n7803 , n7804 );
xor ( n7806 , n7669 , n7805 );
not ( n7807 , n5399 );
not ( n7808 , n7645 );
or ( n7809 , n7807 , n7808 );
and ( n7810 , n5786 , n4440 );
not ( n7811 , n5786 );
and ( n7812 , n7811 , n545 );
or ( n7813 , n7810 , n7812 );
nand ( n7814 , n7813 , n5137 );
nand ( n7815 , n7809 , n7814 );
xor ( n7816 , n7763 , n7768 );
and ( n7817 , n7816 , n7779 );
and ( n7818 , n7763 , n7768 );
or ( n7819 , n7817 , n7818 );
not ( n7820 , n5589 );
not ( n77658 , n7485 );
or ( n7822 , n7820 , n77658 );
nand ( n7823 , n5551 , n7759 );
nand ( n7824 , n7822 , n7823 );
xor ( n7825 , n7819 , n7824 );
xor ( n7826 , n7496 , n7538 );
xor ( n7827 , n7826 , n7547 );
xor ( n7828 , n7825 , n7827 );
xor ( n7829 , n7815 , n7828 );
not ( n7830 , n4444 );
not ( n7831 , n543 );
not ( n7832 , n5643 );
or ( n7833 , n7831 , n7832 );
nand ( n7834 , n5644 , n4938 );
nand ( n7835 , n7833 , n7834 );
not ( n7836 , n7835 );
or ( n7837 , n7830 , n7836 );
nand ( n7838 , n7677 , n5127 );
nand ( n7839 , n7837 , n7838 );
not ( n7840 , n5399 );
not ( n7841 , n7813 );
or ( n7842 , n7840 , n7841 );
not ( n7843 , n545 );
not ( n7844 , n7554 );
or ( n7845 , n7843 , n7844 );
nand ( n7846 , n7219 , n4440 );
nand ( n7847 , n7845 , n7846 );
nand ( n7848 , n7847 , n5137 );
nand ( n7849 , n7842 , n7848 );
xor ( n7850 , n7839 , n7849 );
not ( n7851 , n4434 );
not ( n7852 , n7777 );
or ( n7853 , n7851 , n7852 );
and ( n7854 , n4239 , n7411 );
not ( n7855 , n4239 );
and ( n77693 , n7855 , n7400 );
nor ( n7857 , n7854 , n77693 );
and ( n7858 , n7857 , n539 );
not ( n7859 , n7857 );
and ( n7860 , n7859 , n4251 );
or ( n7861 , n7858 , n7860 );
nand ( n7862 , n7861 , n4224 );
nand ( n7863 , n7853 , n7862 );
xor ( n7864 , n7697 , n7721 );
xor ( n7865 , n7864 , n7740 );
xor ( n7866 , n7863 , n7865 );
not ( n7867 , n5545 );
not ( n7868 , n7749 );
or ( n7869 , n7867 , n7868 );
not ( n7870 , n541 );
not ( n7871 , n6909 );
or ( n7872 , n7870 , n7871 );
nand ( n7873 , n7243 , n5538 );
nand ( n7874 , n7872 , n7873 );
nand ( n7875 , n7874 , n5551 );
nand ( n7876 , n7869 , n7875 );
and ( n7877 , n7866 , n7876 );
and ( n7878 , n7863 , n7865 );
or ( n7879 , n7877 , n7878 );
and ( n7880 , n7850 , n7879 );
and ( n7881 , n7839 , n7849 );
or ( n7882 , n7880 , n7881 );
and ( n7883 , n7829 , n7882 );
and ( n7884 , n7815 , n7828 );
or ( n7885 , n7883 , n7884 );
and ( n7886 , n7806 , n7885 );
and ( n7887 , n7669 , n7805 );
or ( n7888 , n7886 , n7887 );
and ( n7889 , n7659 , n7888 );
and ( n7890 , n7616 , n77495 );
or ( n7891 , n7889 , n7890 );
xor ( n7892 , n7606 , n7891 );
xor ( n7893 , n7629 , n7654 );
and ( n7894 , n7893 , n7657 );
and ( n7895 , n7629 , n7654 );
or ( n7896 , n7894 , n7895 );
xor ( n7897 , n7383 , n7460 );
xor ( n7898 , n7897 , n7568 );
xor ( n7899 , n7896 , n7898 );
not ( n7900 , n5905 );
and ( n77738 , n549 , n5264 );
not ( n7905 , n549 );
and ( n77740 , n7905 , n7378 );
nor ( n7907 , n77738 , n77740 );
not ( n7908 , n7907 );
or ( n7909 , n7900 , n7908 );
not ( n7910 , n549 );
not ( n7911 , n6937 );
not ( n7912 , n7911 );
or ( n7913 , n7910 , n7912 );
not ( n7914 , n549 );
nand ( n7915 , n7914 , n6937 );
nand ( n7916 , n7913 , n7915 );
nand ( n7917 , n7916 , n6489 );
nand ( n7918 , n7909 , n7917 );
xor ( n7919 , n7463 , n7476 );
xor ( n7920 , n7919 , n7565 );
xor ( n7921 , n7918 , n7920 );
xor ( n7922 , n7819 , n7824 );
and ( n7923 , n7922 , n7827 );
and ( n7924 , n7819 , n7824 );
or ( n7925 , n7923 , n7924 );
xor ( n7926 , n7487 , n7550 );
xor ( n7927 , n7926 , n7562 );
xor ( n7928 , n7925 , n7927 );
not ( n7929 , n6489 );
not ( n77764 , n4937 );
and ( n7934 , n549 , n77764 );
not ( n7935 , n549 );
not ( n7936 , n4933 );
and ( n7937 , n7935 , n7936 );
or ( n7938 , n7934 , n7937 );
not ( n7939 , n7938 );
or ( n7940 , n7929 , n7939 );
nand ( n7941 , n7916 , n5905 );
nand ( n7942 , n7940 , n7941 );
and ( n7943 , n7928 , n7942 );
and ( n7944 , n7925 , n7927 );
or ( n7945 , n7943 , n7944 );
and ( n7946 , n7921 , n7945 );
and ( n7947 , n7918 , n7920 );
or ( n7948 , n7946 , n7947 );
xor ( n7949 , n7899 , n7948 );
xor ( n7950 , n7892 , n7949 );
xor ( n7951 , n7918 , n7920 );
xor ( n7952 , n7951 , n7945 );
xor ( n7953 , n7631 , n7640 );
xor ( n7954 , n7953 , n7651 );
not ( n7955 , n5905 );
not ( n7956 , n7938 );
or ( n7957 , n7955 , n7956 );
and ( n7958 , n549 , n6875 );
not ( n77790 , n549 );
and ( n77791 , n77790 , n7633 );
or ( n7961 , n7958 , n77791 );
nand ( n7962 , n7961 , n6489 );
nand ( n7963 , n7957 , n7962 );
xor ( n7964 , n7743 , n7761 );
xor ( n7965 , n7964 , n7780 );
not ( n7966 , n6854 );
xor ( n77798 , n4247 , n547 );
not ( n77799 , n77798 );
or ( n7969 , n7966 , n77799 );
nand ( n7970 , n7800 , n6811 );
nand ( n7971 , n7969 , n7970 );
xor ( n7972 , n7965 , n7971 );
not ( n7973 , n6489 );
not ( n7974 , n549 );
not ( n7975 , n7333 );
or ( n7976 , n7974 , n7975 );
not ( n7977 , n549 );
nand ( n7978 , n7977 , n7786 );
nand ( n7979 , n7976 , n7978 );
not ( n7980 , n7979 );
or ( n7981 , n7973 , n7980 );
nand ( n7982 , n7961 , n5905 );
nand ( n7983 , n7981 , n7982 );
and ( n7984 , n7972 , n7983 );
and ( n7985 , n7965 , n7971 );
or ( n7986 , n7984 , n7985 );
xor ( n7987 , n7963 , n7986 );
not ( n7988 , n551 );
not ( n7989 , n7911 );
or ( n7990 , n7988 , n7989 );
nand ( n77822 , n6937 , n6752 );
nand ( n77823 , n7990 , n77822 );
not ( n7993 , n77823 );
not ( n7994 , n6802 );
or ( n7995 , n7993 , n7994 );
not ( n7996 , n7665 );
or ( n7997 , n7996 , n6801 );
nand ( n7998 , n7995 , n7997 );
and ( n77830 , n7987 , n7998 );
and ( n77831 , n7963 , n7986 );
or ( n8001 , n77830 , n77831 );
xor ( n8002 , n7954 , n8001 );
xor ( n8003 , n7925 , n7927 );
xor ( n8004 , n8003 , n7942 );
and ( n8005 , n8002 , n8004 );
and ( n8006 , n7954 , n8001 );
or ( n8007 , n8005 , n8006 );
xor ( n8008 , n7952 , n8007 );
xor ( n8009 , n7616 , n77495 );
xor ( n8010 , n8009 , n7888 );
and ( n8011 , n8008 , n8010 );
and ( n8012 , n7952 , n8007 );
or ( n8013 , n8011 , n8012 );
nor ( n8014 , n7950 , n8013 );
xor ( n8015 , n7952 , n8007 );
xor ( n8016 , n8015 , n8010 );
xor ( n8017 , n7669 , n7805 );
xor ( n8018 , n8017 , n7885 );
xor ( n8019 , n7679 , n7783 );
xor ( n8020 , n8019 , n7802 );
xor ( n8021 , n7815 , n7828 );
xor ( n8022 , n8021 , n7882 );
xor ( n8023 , n8020 , n8022 );
xnor ( n8024 , n7728 , n7739 );
not ( n8025 , n4434 );
not ( n8026 , n7861 );
or ( n8027 , n8025 , n8026 );
not ( n8028 , n539 );
not ( n8029 , n7700 );
or ( n8030 , n8028 , n8029 );
nand ( n8031 , n7536 , n4251 );
nand ( n8032 , n8030 , n8031 );
nand ( n8033 , n4224 , n8032 );
nand ( n8034 , n8027 , n8033 );
xor ( n8035 , n8024 , n8034 );
buf ( n8036 , n7696 );
and ( n8037 , n8036 , n5501 );
not ( n8038 , n4433 );
not ( n8039 , n8032 );
or ( n77871 , n8038 , n8039 );
not ( n8041 , n539 );
not ( n8042 , n7718 );
not ( n8043 , n8042 );
or ( n8044 , n8041 , n8043 );
nand ( n8045 , n7718 , n4251 );
nand ( n8046 , n8044 , n8045 );
nand ( n8047 , n8046 , n4224 );
nand ( n8048 , n77871 , n8047 );
xor ( n8049 , n8037 , n8048 );
not ( n8050 , n540 );
nand ( n8051 , n8050 , n7731 );
and ( n8052 , n8051 , n541 );
not ( n8053 , n540 );
not ( n8054 , n7696 );
or ( n77886 , n8053 , n8054 );
nand ( n77887 , n77886 , n539 );
nor ( n8057 , n8052 , n77887 );
not ( n8058 , n4434 );
not ( n8059 , n8046 );
or ( n8060 , n8058 , n8059 );
and ( n8061 , n7736 , n5772 );
nor ( n8062 , n7695 , n5774 );
nor ( n8063 , n8061 , n8062 );
nand ( n8064 , n8060 , n8063 );
and ( n8065 , n8057 , n8064 );
and ( n8066 , n8049 , n8065 );
and ( n8067 , n8037 , n8048 );
or ( n8068 , n8066 , n8067 );
and ( n8069 , n8035 , n8068 );
and ( n8070 , n8024 , n8034 );
or ( n8071 , n8069 , n8070 );
not ( n8072 , n4443 );
not ( n8073 , n7835 );
or ( n8074 , n8072 , n8073 );
not ( n8075 , n543 );
nor ( n8076 , n7756 , n5516 );
not ( n8077 , n8076 );
not ( n8078 , n8077 );
or ( n8079 , n8075 , n8078 );
nand ( n8080 , n8076 , n4938 );
nand ( n8081 , n8079 , n8080 );
nand ( n8082 , n8081 , n4444 );
nand ( n77914 , n8074 , n8082 );
xor ( n8084 , n8071 , n77914 );
not ( n8085 , n5399 );
not ( n8086 , n7847 );
or ( n8087 , n8085 , n8086 );
not ( n8088 , n545 );
not ( n8089 , n6916 );
or ( n8090 , n8088 , n8089 );
nand ( n8091 , n5724 , n4440 );
nand ( n8092 , n8090 , n8091 );
nand ( n8093 , n8092 , n5137 );
nand ( n8094 , n8087 , n8093 );
and ( n8095 , n8084 , n8094 );
and ( n8096 , n8071 , n77914 );
or ( n8097 , n8095 , n8096 );
not ( n8098 , n6802 );
not ( n8099 , n551 );
not ( n8100 , n77764 );
or ( n8101 , n8099 , n8100 );
nand ( n8102 , n7936 , n6752 );
nand ( n8103 , n8101 , n8102 );
not ( n8104 , n8103 );
or ( n8105 , n8098 , n8104 );
nand ( n8106 , n77823 , n552 );
nand ( n8107 , n8105 , n8106 );
xor ( n8108 , n8097 , n8107 );
xor ( n8109 , n7839 , n7849 );
xor ( n8110 , n8109 , n7879 );
and ( n8111 , n8108 , n8110 );
and ( n8112 , n8097 , n8107 );
or ( n8113 , n8111 , n8112 );
and ( n8114 , n8023 , n8113 );
and ( n8115 , n8020 , n8022 );
or ( n8116 , n8114 , n8115 );
xor ( n8117 , n8018 , n8116 );
xor ( n8118 , n7954 , n8001 );
xor ( n8119 , n8118 , n8004 );
and ( n8120 , n8117 , n8119 );
and ( n8121 , n8018 , n8116 );
or ( n8122 , n8120 , n8121 );
nand ( n8123 , n8016 , n8122 );
or ( n8124 , n8014 , n8123 );
nand ( n8125 , n7950 , n8013 );
nand ( n8126 , n8124 , n8125 );
not ( n8127 , n8126 );
xor ( n8128 , n7377 , n7594 );
xor ( n8129 , n8128 , n7597 );
xor ( n8130 , n7330 , n7355 );
xor ( n8131 , n8130 , n7358 );
xor ( n8132 , n7896 , n7898 );
and ( n8133 , n8132 , n7948 );
and ( n8134 , n7896 , n7898 );
or ( n8135 , n8133 , n8134 );
xor ( n8136 , n8131 , n8135 );
xor ( n8137 , n7571 , n7573 );
xor ( n8138 , n8137 , n7591 );
and ( n8139 , n8136 , n8138 );
and ( n8140 , n8131 , n8135 );
or ( n8141 , n8139 , n8140 );
nor ( n8142 , n8129 , n8141 );
xor ( n8143 , n8131 , n8135 );
xor ( n8144 , n8143 , n8138 );
xor ( n8145 , n7606 , n7891 );
and ( n8146 , n8145 , n7949 );
and ( n8147 , n7606 , n7891 );
or ( n8148 , n8146 , n8147 );
nor ( n8149 , n8144 , n8148 );
nor ( n8150 , n8142 , n8149 );
not ( n8151 , n8150 );
or ( n8152 , n8127 , n8151 );
not ( n8153 , n8142 );
nand ( n8154 , n8144 , n8148 );
not ( n8155 , n8154 );
and ( n8156 , n8153 , n8155 );
not ( n8157 , n8129 );
not ( n8158 , n8141 );
nor ( n8159 , n8157 , n8158 );
nor ( n8160 , n8156 , n8159 );
nand ( n8161 , n8152 , n8160 );
not ( n8162 , n8161 );
or ( n8163 , n7604 , n8162 );
nor ( n8164 , n7212 , n7370 );
not ( n8165 , n8164 );
nand ( n8166 , n7374 , n7600 );
not ( n8167 , n8166 );
and ( n8168 , n8165 , n8167 );
and ( n8169 , n7212 , n7370 );
nor ( n8170 , n8168 , n8169 );
nand ( n8171 , n8163 , n8170 );
not ( n8172 , n8129 );
nand ( n8173 , n8172 , n8158 );
not ( n8174 , n8144 );
not ( n8175 , n8148 );
nand ( n8176 , n8174 , n8175 );
nand ( n78008 , n8173 , n8176 );
not ( n78009 , n78008 );
not ( n8179 , n7950 );
not ( n8180 , n8013 );
nand ( n8181 , n8179 , n8180 );
not ( n8182 , n8016 );
not ( n8183 , n8122 );
nand ( n8184 , n8182 , n8183 );
nand ( n8185 , n8181 , n8184 );
not ( n8186 , n8185 );
not ( n8187 , n552 );
not ( n8188 , n551 );
not ( n8189 , n7789 );
or ( n8190 , n8188 , n8189 );
nand ( n8191 , n7786 , n6752 );
nand ( n8192 , n8190 , n8191 );
not ( n8193 , n8192 );
or ( n8194 , n8187 , n8193 );
buf ( n8195 , n4425 );
nand ( n8196 , n8195 , n6752 );
nand ( n8197 , n551 , n5535 );
nand ( n8198 , n8196 , n8197 );
nand ( n8199 , n8198 , n6802 );
nand ( n8200 , n8194 , n8199 );
not ( n8201 , n6854 );
and ( n8202 , n547 , n6975 );
not ( n8203 , n547 );
and ( n8204 , n8203 , n5644 );
or ( n8205 , n8202 , n8204 );
not ( n8206 , n8205 );
or ( n8207 , n8201 , n8206 );
and ( n8208 , n5724 , n6857 );
not ( n8209 , n5724 );
and ( n8210 , n8209 , n547 );
or ( n8211 , n8208 , n8210 );
nand ( n8212 , n8211 , n6811 );
nand ( n8213 , n8207 , n8212 );
not ( n8214 , n543 );
not ( n8215 , n7277 );
or ( n8216 , n8214 , n8215 );
nand ( n8217 , n7276 , n4938 );
nand ( n8218 , n8216 , n8217 );
nand ( n8219 , n8218 , n4443 );
not ( n8220 , n543 );
not ( n8221 , n7857 );
or ( n8222 , n8220 , n8221 );
not ( n8223 , n7857 );
nand ( n8224 , n8223 , n4938 );
nand ( n8225 , n8222 , n8224 );
nand ( n8226 , n8225 , n4444 );
nand ( n8227 , n8219 , n8226 );
and ( n8228 , n8036 , n4433 );
not ( n8229 , n5545 );
not ( n8230 , n5538 );
not ( n8231 , n7536 );
or ( n8232 , n8230 , n8231 );
or ( n8233 , n7536 , n4219 );
nand ( n8234 , n8232 , n8233 );
not ( n8235 , n8234 );
or ( n8236 , n8229 , n8235 );
not ( n8237 , n541 );
not ( n8238 , n8042 );
or ( n8239 , n8237 , n8238 );
nand ( n8240 , n7718 , n5538 );
nand ( n8241 , n8239 , n8240 );
nand ( n8242 , n8241 , n5550 );
nand ( n8243 , n8236 , n8242 );
xor ( n8244 , n8228 , n8243 );
not ( n8245 , n5545 );
not ( n8246 , n8241 );
or ( n8247 , n8245 , n8246 );
not ( n8248 , n7696 );
not ( n8249 , n4219 );
or ( n8250 , n8248 , n8249 );
or ( n78082 , n7696 , n4219 );
nand ( n8252 , n8250 , n78082 );
nand ( n8253 , n8252 , n5550 );
nand ( n8254 , n8247 , n8253 );
not ( n8255 , n8254 );
not ( n8256 , n542 );
not ( n8257 , n8256 );
not ( n8258 , n7731 );
or ( n8259 , n8257 , n8258 );
nand ( n8260 , n8259 , n543 );
and ( n8261 , n7736 , n542 );
nor ( n8262 , n8261 , n5538 );
nand ( n8263 , n8260 , n8262 );
nor ( n8264 , n8255 , n8263 );
xor ( n8265 , n8244 , n8264 );
xor ( n8266 , n8227 , n8265 );
not ( n8267 , n5399 );
not ( n8268 , n545 );
not ( n8269 , n5822 );
not ( n8270 , n8269 );
or ( n8271 , n8268 , n8270 );
nand ( n8272 , n5822 , n4440 );
nand ( n8273 , n8271 , n8272 );
not ( n8274 , n8273 );
or ( n8275 , n8267 , n8274 );
not ( n8276 , n545 );
not ( n8277 , n6909 );
or ( n8278 , n8276 , n8277 );
nand ( n8279 , n7243 , n4440 );
nand ( n8280 , n8278 , n8279 );
nand ( n8281 , n8280 , n5137 );
nand ( n8282 , n8275 , n8281 );
and ( n8283 , n8266 , n8282 );
and ( n8284 , n8227 , n8265 );
or ( n8285 , n8283 , n8284 );
xor ( n8286 , n8213 , n8285 );
not ( n8287 , n5905 );
and ( n8288 , n549 , n5769 );
not ( n8289 , n549 );
not ( n8290 , n7451 );
and ( n8291 , n8289 , n8290 );
or ( n8292 , n8288 , n8291 );
not ( n8293 , n8292 );
or ( n8294 , n8287 , n8293 );
not ( n8295 , n549 );
not ( n8296 , n7554 );
or ( n8297 , n8295 , n8296 );
not ( n8298 , n549 );
not ( n8299 , n7554 );
nand ( n8300 , n8298 , n8299 );
nand ( n8301 , n8297 , n8300 );
nand ( n78133 , n8301 , n6489 );
nand ( n8303 , n8294 , n78133 );
and ( n8304 , n8286 , n8303 );
and ( n8305 , n8213 , n8285 );
or ( n8306 , n8304 , n8305 );
xor ( n8307 , n8200 , n8306 );
xor ( n8308 , n8057 , n8064 );
xor ( n8309 , n7414 , n541 );
not ( n8310 , n8309 );
not ( n8311 , n5545 );
or ( n8312 , n8310 , n8311 );
nand ( n8313 , n8234 , n5550 );
nand ( n8314 , n8312 , n8313 );
xor ( n8315 , n8308 , n8314 );
xor ( n8316 , n8228 , n8243 );
and ( n8317 , n8316 , n8264 );
and ( n8318 , n8228 , n8243 );
or ( n8319 , n8317 , n8318 );
and ( n8320 , n8315 , n8319 );
and ( n8321 , n8308 , n8314 );
or ( n8322 , n8320 , n8321 );
not ( n8323 , n5399 );
not ( n8324 , n545 );
not ( n8325 , n5643 );
or ( n8326 , n8324 , n8325 );
nand ( n8327 , n5644 , n4440 );
nand ( n8328 , n8326 , n8327 );
not ( n8329 , n8328 );
or ( n8330 , n8323 , n8329 );
not ( n8331 , n545 );
not ( n8332 , n8077 );
or ( n8333 , n8331 , n8332 );
nand ( n78165 , n8076 , n4440 );
nand ( n8338 , n8333 , n78165 );
nand ( n78167 , n8338 , n5137 );
nand ( n8340 , n8330 , n78167 );
xor ( n8341 , n8322 , n8340 );
not ( n8342 , n5588 );
not ( n8343 , n541 );
not ( n8344 , n7277 );
or ( n8345 , n8343 , n8344 );
nand ( n8346 , n7276 , n5538 );
nand ( n8347 , n8345 , n8346 );
not ( n8348 , n8347 );
or ( n8349 , n8342 , n8348 );
nand ( n8350 , n8309 , n5551 );
nand ( n8351 , n8349 , n8350 );
xor ( n8352 , n8037 , n8048 );
xor ( n8353 , n8352 , n8065 );
xor ( n8354 , n8351 , n8353 );
not ( n8355 , n543 );
not ( n8356 , n6909 );
or ( n8357 , n8355 , n8356 );
nand ( n8358 , n7243 , n4938 );
nand ( n8359 , n8357 , n8358 );
nand ( n8360 , n8359 , n4444 );
not ( n8361 , n543 );
not ( n8362 , n8269 );
or ( n78191 , n8361 , n8362 );
nand ( n8367 , n5822 , n4938 );
nand ( n8368 , n78191 , n8367 );
nand ( n8369 , n8368 , n4443 );
nand ( n8370 , n8360 , n8369 );
xor ( n8371 , n8354 , n8370 );
xor ( n8372 , n8341 , n8371 );
and ( n8373 , n8307 , n8372 );
and ( n78199 , n8200 , n8306 );
or ( n8375 , n8373 , n78199 );
not ( n8376 , n5545 );
not ( n8377 , n7874 );
or ( n8378 , n8376 , n8377 );
nand ( n8379 , n8347 , n5550 );
nand ( n8380 , n8378 , n8379 );
not ( n8381 , n4444 );
not ( n8382 , n8368 );
or ( n8383 , n8381 , n8382 );
nand ( n8384 , n8081 , n4443 );
nand ( n8385 , n8383 , n8384 );
xor ( n8386 , n8380 , n8385 );
xor ( n8387 , n8024 , n8034 );
xor ( n8388 , n8387 , n8068 );
xor ( n8389 , n8386 , n8388 );
not ( n8390 , n6489 );
not ( n8391 , n549 );
not ( n8392 , n74151 );
or ( n8393 , n8391 , n8392 );
not ( n8394 , n549 );
nand ( n8395 , n8394 , n7446 );
nand ( n8396 , n8393 , n8395 );
not ( n8397 , n8396 );
or ( n8398 , n8390 , n8397 );
and ( n78224 , n549 , n5535 );
not ( n78225 , n549 );
and ( n8401 , n78225 , n4425 );
or ( n8402 , n78224 , n8401 );
nand ( n8403 , n8402 , n5905 );
nand ( n8404 , n8398 , n8403 );
xor ( n8405 , n8389 , n8404 );
not ( n8406 , n552 );
not ( n78232 , n6752 );
not ( n78233 , n77458 );
or ( n8409 , n78232 , n78233 );
nand ( n8410 , n7624 , n551 );
nand ( n8411 , n8409 , n8410 );
not ( n8412 , n8411 );
or ( n8413 , n8406 , n8412 );
nand ( n8414 , n8192 , n6802 );
nand ( n8415 , n8413 , n8414 );
xor ( n8416 , n8405 , n8415 );
xor ( n8417 , n8375 , n8416 );
xor ( n8418 , n8322 , n8340 );
and ( n8419 , n8418 , n8371 );
and ( n8420 , n8322 , n8340 );
or ( n8421 , n8419 , n8420 );
not ( n8422 , n5137 );
not ( n8423 , n8328 );
or ( n8424 , n8422 , n8423 );
nand ( n8425 , n8092 , n5399 );
nand ( n8426 , n8424 , n8425 );
not ( n8427 , n6854 );
not ( n8428 , n547 );
not ( n8429 , n8428 );
not ( n8430 , n8299 );
or ( n8431 , n8429 , n8430 );
nand ( n8432 , n7554 , n547 );
nand ( n8433 , n8431 , n8432 );
not ( n8434 , n8433 );
or ( n8435 , n8427 , n8434 );
and ( n8436 , n547 , n5754 );
not ( n8437 , n547 );
and ( n8438 , n8437 , n5786 );
or ( n8439 , n8436 , n8438 );
nand ( n8440 , n8439 , n6811 );
nand ( n8441 , n8435 , n8440 );
xor ( n8442 , n8426 , n8441 );
xor ( n8443 , n8351 , n8353 );
and ( n8444 , n8443 , n8370 );
and ( n8445 , n8351 , n8353 );
or ( n8446 , n8444 , n8445 );
xor ( n8447 , n8442 , n8446 );
xor ( n8448 , n8421 , n8447 );
not ( n8449 , n6811 );
not ( n8450 , n8433 );
or ( n8451 , n8449 , n8450 );
nand ( n8452 , n8211 , n6955 );
nand ( n8453 , n8451 , n8452 );
not ( n8454 , n5127 );
not ( n8455 , n8359 );
or ( n8456 , n8454 , n8455 );
nand ( n8457 , n8218 , n4444 );
nand ( n8458 , n8456 , n8457 );
not ( n8459 , n5137 );
not ( n78285 , n8273 );
or ( n78286 , n8459 , n78285 );
nand ( n8462 , n8338 , n5399 );
nand ( n8463 , n78286 , n8462 );
xor ( n8464 , n8458 , n8463 );
xor ( n8465 , n8308 , n8314 );
xor ( n8466 , n8465 , n8319 );
and ( n8467 , n8464 , n8466 );
and ( n8468 , n8458 , n8463 );
or ( n8469 , n8467 , n8468 );
xor ( n8470 , n8453 , n8469 );
not ( n8471 , n5905 );
not ( n8472 , n8396 );
or ( n8473 , n8471 , n8472 );
nand ( n8474 , n6489 , n8292 );
nand ( n8475 , n8473 , n8474 );
and ( n8476 , n8470 , n8475 );
and ( n8477 , n8453 , n8469 );
or ( n8478 , n8476 , n8477 );
xor ( n8479 , n8448 , n8478 );
and ( n8480 , n8417 , n8479 );
and ( n8481 , n8375 , n8416 );
or ( n8482 , n8480 , n8481 );
not ( n8483 , n5905 );
not ( n8484 , n7979 );
or ( n78310 , n8483 , n8484 );
nand ( n78311 , n8402 , n6489 );
nand ( n8487 , n78310 , n78311 );
xor ( n8488 , n8071 , n77914 );
xor ( n8489 , n8488 , n8094 );
xor ( n8490 , n8487 , n8489 );
xor ( n8491 , n8426 , n8441 );
and ( n8492 , n8491 , n8446 );
and ( n78318 , n8426 , n8441 );
or ( n78319 , n8492 , n78318 );
xor ( n8495 , n8490 , n78319 );
xor ( n8496 , n8421 , n8447 );
and ( n8497 , n8496 , n8478 );
and ( n8498 , n8421 , n8447 );
or ( n8499 , n8497 , n8498 );
xor ( n8500 , n8495 , n8499 );
not ( n8501 , n552 );
not ( n8502 , n8103 );
or ( n8503 , n8501 , n8502 );
nand ( n8504 , n8411 , n6802 );
nand ( n8505 , n8503 , n8504 );
xor ( n8506 , n7863 , n7865 );
xor ( n8507 , n8506 , n7876 );
xor ( n8508 , n8380 , n8385 );
and ( n8509 , n8508 , n8388 );
and ( n8510 , n8380 , n8385 );
or ( n8511 , n8509 , n8510 );
xor ( n8512 , n8507 , n8511 );
not ( n8513 , n6811 );
not ( n8514 , n77798 );
or ( n8515 , n8513 , n8514 );
nand ( n8516 , n8439 , n6955 );
nand ( n8517 , n8515 , n8516 );
xor ( n8518 , n8512 , n8517 );
xor ( n8519 , n8505 , n8518 );
xor ( n8520 , n8389 , n8404 );
and ( n8521 , n8520 , n8415 );
and ( n8522 , n8389 , n8404 );
or ( n8523 , n8521 , n8522 );
xor ( n8524 , n8519 , n8523 );
xor ( n8525 , n8500 , n8524 );
nor ( n8526 , n8482 , n8525 );
xor ( n8527 , n8375 , n8416 );
xor ( n8528 , n8527 , n8479 );
xor ( n8529 , n8453 , n8469 );
xor ( n8530 , n8529 , n8475 );
xor ( n8531 , n8458 , n8463 );
xor ( n8532 , n8531 , n8466 );
not ( n8533 , n6802 );
not ( n8534 , n551 );
not ( n8535 , n74151 );
or ( n8536 , n8534 , n8535 );
nand ( n8537 , n7446 , n6752 );
nand ( n8538 , n8536 , n8537 );
not ( n8539 , n8538 );
or ( n8540 , n8533 , n8539 );
not ( n8541 , n8197 );
not ( n8542 , n8196 );
or ( n8543 , n8541 , n8542 );
nand ( n78369 , n8543 , n552 );
nand ( n8545 , n8540 , n78369 );
xor ( n8546 , n8532 , n8545 );
xnor ( n8547 , n8254 , n8263 );
not ( n8548 , n4443 );
not ( n8549 , n8225 );
or ( n8550 , n8548 , n8549 );
not ( n8551 , n543 );
not ( n8552 , n7700 );
or ( n8553 , n8551 , n8552 );
nand ( n8554 , n7536 , n4938 );
nand ( n8555 , n8553 , n8554 );
nand ( n8556 , n8555 , n4444 );
nand ( n8557 , n8550 , n8556 );
xor ( n8558 , n8547 , n8557 );
and ( n8559 , n8036 , n5545 );
not ( n8560 , n4443 );
not ( n8561 , n8555 );
or ( n8562 , n8560 , n8561 );
not ( n8563 , n543 );
not ( n8564 , n8042 );
or ( n8565 , n8563 , n8564 );
nand ( n8566 , n7718 , n4938 );
nand ( n8567 , n8565 , n8566 );
nand ( n8568 , n8567 , n4444 );
nand ( n8569 , n8562 , n8568 );
xor ( n8570 , n8559 , n8569 );
not ( n8571 , n4438 );
not ( n8572 , n7731 );
or ( n8573 , n8571 , n8572 );
nand ( n8574 , n8573 , n545 );
and ( n8575 , n7736 , n544 );
nor ( n8576 , n8575 , n4938 );
and ( n8577 , n8574 , n8576 );
not ( n8578 , n4443 );
not ( n8579 , n8567 );
or ( n8580 , n8578 , n8579 );
not ( n8581 , n7731 );
not ( n8582 , n7236 );
not ( n8583 , n8582 );
and ( n8584 , n8581 , n8583 );
nor ( n8585 , n7736 , n7230 );
nor ( n8586 , n8584 , n8585 );
nand ( n8587 , n8580 , n8586 );
and ( n8588 , n8577 , n8587 );
and ( n8589 , n8570 , n8588 );
and ( n8590 , n8559 , n8569 );
or ( n8591 , n8589 , n8590 );
and ( n8592 , n8558 , n8591 );
and ( n8593 , n8547 , n8557 );
or ( n8594 , n8592 , n8593 );
not ( n8595 , n6811 );
not ( n8596 , n8205 );
or ( n8597 , n8595 , n8596 );
and ( n8598 , n547 , n5530 );
not ( n8599 , n547 );
and ( n8600 , n8599 , n8076 );
or ( n8601 , n8598 , n8600 );
nand ( n8602 , n8601 , n6955 );
nand ( n8603 , n8597 , n8602 );
xor ( n8604 , n8594 , n8603 );
xor ( n8605 , n8227 , n8265 );
xor ( n8606 , n8605 , n8282 );
and ( n8607 , n8604 , n8606 );
and ( n8608 , n8594 , n8603 );
or ( n8609 , n8607 , n8608 );
and ( n8610 , n8546 , n8609 );
and ( n8611 , n8532 , n8545 );
or ( n8612 , n8610 , n8611 );
xor ( n8613 , n8530 , n8612 );
xor ( n8614 , n8200 , n8306 );
xor ( n8615 , n8614 , n8372 );
and ( n8616 , n8613 , n8615 );
and ( n8617 , n8530 , n8612 );
or ( n8618 , n8616 , n8617 );
nor ( n8619 , n8528 , n8618 );
nor ( n8620 , n8526 , n8619 );
not ( n8621 , n8620 );
xor ( n8622 , n8530 , n8612 );
xor ( n8623 , n8622 , n8615 );
not ( n8624 , n8623 );
xor ( n8625 , n8213 , n8285 );
xor ( n8626 , n8625 , n8303 );
not ( n8627 , n5905 );
not ( n8628 , n8301 );
or ( n8629 , n8627 , n8628 );
not ( n8630 , n549 );
not ( n8631 , n6916 );
or ( n8632 , n8630 , n8631 );
nand ( n8633 , n5724 , n7018 );
nand ( n8634 , n8632 , n8633 );
nand ( n8635 , n8634 , n6489 );
nand ( n8636 , n8629 , n8635 );
not ( n8637 , n5399 );
not ( n78463 , n8280 );
or ( n78464 , n8637 , n78463 );
not ( n8640 , n545 );
not ( n8641 , n7277 );
or ( n8642 , n8640 , n8641 );
nand ( n8643 , n4440 , n7278 );
nand ( n8644 , n8642 , n8643 );
nand ( n8645 , n5137 , n8644 );
nand ( n8646 , n78464 , n8645 );
not ( n8647 , n6811 );
not ( n8648 , n8601 );
or ( n8649 , n8647 , n8648 );
not ( n8650 , n5822 );
not ( n8651 , n8428 );
or ( n8652 , n8650 , n8651 );
or ( n8653 , n8428 , n5822 );
nand ( n8654 , n8652 , n8653 );
nand ( n8655 , n8654 , n6854 );
nand ( n8656 , n8649 , n8655 );
xor ( n8657 , n8646 , n8656 );
xor ( n8658 , n8547 , n8557 );
xor ( n8659 , n8658 , n8591 );
and ( n8660 , n8657 , n8659 );
and ( n8661 , n8646 , n8656 );
or ( n8662 , n8660 , n8661 );
xor ( n8663 , n8636 , n8662 );
not ( n8664 , n552 );
not ( n8665 , n8538 );
or ( n8666 , n8664 , n8665 );
not ( n8667 , n551 );
not ( n8668 , n5754 );
or ( n8669 , n8667 , n8668 );
nand ( n8670 , n5753 , n6752 );
nand ( n8671 , n8669 , n8670 );
nand ( n8672 , n8671 , n6802 );
nand ( n8673 , n8666 , n8672 );
and ( n8674 , n8663 , n8673 );
and ( n8675 , n8636 , n8662 );
or ( n8676 , n8674 , n8675 );
xor ( n8677 , n8626 , n8676 );
xor ( n8678 , n8532 , n8545 );
xor ( n8679 , n8678 , n8609 );
and ( n8680 , n8677 , n8679 );
and ( n8681 , n8626 , n8676 );
or ( n8682 , n8680 , n8681 );
not ( n8683 , n8682 );
nand ( n8684 , n8624 , n8683 );
not ( n8685 , n8684 );
xor ( n8686 , n8626 , n8676 );
xor ( n8687 , n8686 , n8679 );
not ( n8688 , n8687 );
not ( n8689 , n5905 );
not ( n8690 , n8634 );
or ( n8691 , n8689 , n8690 );
not ( n8692 , n5448 );
not ( n8693 , n549 );
or ( n8694 , n8692 , n8693 );
or ( n8695 , n6975 , n549 );
nand ( n8696 , n8694 , n8695 );
nand ( n8697 , n8696 , n6489 );
nand ( n8698 , n8691 , n8697 );
not ( n8699 , n552 );
not ( n8700 , n8671 );
or ( n8701 , n8699 , n8700 );
and ( n8702 , n7554 , n6868 );
nor ( n8703 , C0 , n8702 );
nand ( n8704 , n8701 , n8703 );
xor ( n8705 , n8698 , n8704 );
not ( n8706 , n5399 );
not ( n8707 , n8644 );
or ( n8708 , n8706 , n8707 );
not ( n8709 , n545 );
not ( n8710 , n7857 );
or ( n8711 , n8709 , n8710 );
nand ( n8712 , n8223 , n4440 );
nand ( n8713 , n8711 , n8712 );
nand ( n8714 , n8713 , n5137 );
nand ( n8715 , n8708 , n8714 );
xor ( n78541 , n8559 , n8569 );
xor ( n8717 , n78541 , n8588 );
xor ( n8718 , n8715 , n8717 );
not ( n8719 , n6811 );
not ( n8720 , n8654 );
or ( n8721 , n8719 , n8720 );
and ( n8722 , n547 , n6909 );
not ( n8723 , n547 );
and ( n8724 , n8723 , n7243 );
or ( n8725 , n8722 , n8724 );
nand ( n8726 , n8725 , n6854 );
nand ( n78552 , n8721 , n8726 );
and ( n8728 , n8718 , n78552 );
and ( n8729 , n8715 , n8717 );
or ( n8730 , n8728 , n8729 );
and ( n8731 , n8705 , n8730 );
and ( n8732 , n8698 , n8704 );
or ( n8733 , n8731 , n8732 );
xor ( n8734 , n8594 , n8603 );
xor ( n8735 , n8734 , n8606 );
xor ( n8736 , n8733 , n8735 );
xor ( n8737 , n8636 , n8662 );
xor ( n8738 , n8737 , n8673 );
and ( n8739 , n8736 , n8738 );
and ( n8740 , n8733 , n8735 );
or ( n8741 , n8739 , n8740 );
not ( n8742 , n8741 );
and ( n8743 , n8688 , n8742 );
xor ( n8744 , n8733 , n8735 );
xor ( n8745 , n8744 , n8738 );
xor ( n8746 , n8646 , n8656 );
xor ( n8747 , n8746 , n8659 );
xor ( n8748 , n8577 , n8587 );
not ( n8749 , n5398 );
not ( n8750 , n8713 );
or ( n8751 , n8749 , n8750 );
not ( n8752 , n545 );
not ( n8753 , n7700 );
or ( n8754 , n8752 , n8753 );
nand ( n8755 , n7536 , n4440 );
nand ( n8756 , n8754 , n8755 );
nand ( n8757 , n8756 , n5137 );
nand ( n8758 , n8751 , n8757 );
xor ( n8759 , n8748 , n8758 );
not ( n8760 , n6811 );
not ( n8761 , n8725 );
or ( n8762 , n8760 , n8761 );
not ( n8763 , n547 );
not ( n8764 , n7277 );
or ( n8765 , n8763 , n8764 );
not ( n8766 , n547 );
nand ( n8767 , n8766 , n7276 );
nand ( n8768 , n8765 , n8767 );
nand ( n8769 , n8768 , n6955 );
nand ( n8770 , n8762 , n8769 );
and ( n8771 , n8759 , n8770 );
and ( n8772 , n8748 , n8758 );
or ( n8773 , n8771 , n8772 );
not ( n8774 , n5905 );
not ( n8775 , n8696 );
or ( n8776 , n8774 , n8775 );
and ( n8777 , n549 , n8076 );
not ( n8778 , n549 );
and ( n8779 , n8778 , n5530 );
nor ( n8780 , n8777 , n8779 );
nand ( n8781 , n8780 , n6489 );
nand ( n8782 , n8776 , n8781 );
xor ( n8783 , n8773 , n8782 );
nand ( n8784 , n8299 , n7328 );
nand ( n8785 , n7554 , n7325 );
and ( n8786 , n6752 , n6916 );
not ( n8787 , n6752 );
and ( n8788 , n8787 , n5724 );
nor ( n8789 , n8786 , n8788 );
nand ( n8790 , n8789 , n6802 );
nand ( n8791 , n8784 , n8785 , n8790 );
and ( n8792 , n8783 , n8791 );
and ( n8793 , n8773 , n8782 );
or ( n8794 , n8792 , n8793 );
xor ( n8795 , n8747 , n8794 );
xor ( n8796 , n8698 , n8704 );
xor ( n8797 , n8796 , n8730 );
and ( n8798 , n8795 , n8797 );
and ( n78624 , n8747 , n8794 );
or ( n8803 , n8798 , n78624 );
nor ( n78626 , n8745 , n8803 );
nor ( n8805 , n8743 , n78626 );
not ( n8806 , n8805 );
xor ( n8807 , n8747 , n8794 );
xor ( n8808 , n8807 , n8797 );
not ( n8809 , n8808 );
xor ( n8810 , n8715 , n8717 );
xor ( n8811 , n8810 , n78552 );
and ( n8812 , n8036 , n4443 );
not ( n8813 , n5398 );
not ( n8814 , n8756 );
or ( n8815 , n8813 , n8814 );
not ( n8816 , n545 );
not ( n8817 , n8042 );
or ( n8818 , n8816 , n8817 );
nand ( n8819 , n7718 , n4440 );
nand ( n8820 , n8818 , n8819 );
nand ( n8821 , n5137 , n8820 );
nand ( n8822 , n8815 , n8821 );
xor ( n78645 , n8812 , n8822 );
and ( n8827 , n7736 , n546 );
nor ( n8828 , n8827 , n4440 );
not ( n8829 , n546 );
not ( n8830 , n8829 );
not ( n8831 , n7731 );
or ( n8832 , n8830 , n8831 );
nand ( n8833 , n8832 , n547 );
and ( n8834 , n8828 , n8833 );
not ( n8835 , n5398 );
not ( n8836 , n8820 );
or ( n8837 , n8835 , n8836 );
and ( n8838 , n545 , n7696 );
not ( n8839 , n545 );
and ( n8840 , n8839 , n7731 );
nor ( n8841 , n8838 , n8840 );
nand ( n8842 , n8841 , n5137 );
nand ( n8843 , n8837 , n8842 );
and ( n8844 , n8834 , n8843 );
and ( n8845 , n78645 , n8844 );
and ( n8846 , n8812 , n8822 );
or ( n8847 , n8845 , n8846 );
not ( n8848 , n5822 );
and ( n8849 , n549 , n8848 );
not ( n8850 , n549 );
and ( n8851 , n8850 , n5822 );
or ( n8852 , n8849 , n8851 );
not ( n8853 , n8852 );
not ( n8854 , n6489 );
or ( n8855 , n8853 , n8854 );
nand ( n8856 , n8780 , n5905 );
nand ( n8857 , n8855 , n8856 );
xor ( n8858 , n8847 , n8857 );
xor ( n8859 , n8748 , n8758 );
xor ( n8860 , n8859 , n8770 );
and ( n78680 , n8858 , n8860 );
and ( n78681 , n8847 , n8857 );
or ( n8863 , n78680 , n78681 );
xor ( n8864 , n8811 , n8863 );
xor ( n8865 , n8773 , n8782 );
xor ( n8866 , n8865 , n8791 );
and ( n8867 , n8864 , n8866 );
and ( n8868 , n8811 , n8863 );
or ( n78688 , n8867 , n8868 );
not ( n78689 , n78688 );
nand ( n8871 , n8809 , n78689 );
not ( n8872 , n8871 );
xor ( n8873 , n8811 , n8863 );
xor ( n8874 , n8873 , n8866 );
not ( n8875 , n8789 );
not ( n8876 , n552 );
or ( n8877 , n8875 , n8876 );
not ( n8878 , n6868 );
or ( n8879 , n5644 , n8878 );
nand ( n8880 , n8877 , n8879 );
not ( n8881 , n6811 );
not ( n8882 , n8768 );
or ( n8883 , n8881 , n8882 );
and ( n8884 , n547 , n7857 );
not ( n8885 , n547 );
and ( n8886 , n8885 , n7414 );
or ( n8887 , n8884 , n8886 );
nand ( n8888 , n8887 , n6955 );
nand ( n8889 , n8883 , n8888 );
xor ( n78709 , n8812 , n8822 );
xor ( n78710 , n78709 , n8844 );
xor ( n8892 , n8889 , n78710 );
not ( n8893 , n5905 );
not ( n8894 , n8852 );
or ( n8895 , n8893 , n8894 );
and ( n8896 , n549 , n6909 );
not ( n8897 , n549 );
and ( n78717 , n8897 , n6910 );
or ( n78718 , n8896 , n78717 );
nand ( n8900 , n78718 , n6489 );
nand ( n8901 , n8895 , n8900 );
and ( n8902 , n8892 , n8901 );
and ( n8903 , n8889 , n78710 );
or ( n8904 , n8902 , n8903 );
xor ( n8905 , n8880 , n8904 );
xor ( n8906 , n8847 , n8857 );
xor ( n8907 , n8906 , n8860 );
and ( n8908 , n8905 , n8907 );
and ( n8909 , n8880 , n8904 );
or ( n8910 , n8908 , n8909 );
nor ( n8911 , n8874 , n8910 );
xor ( n8912 , n8880 , n8904 );
xor ( n8913 , n8912 , n8907 );
not ( n8914 , n8913 );
xor ( n8915 , n8834 , n8843 );
not ( n8916 , n6811 );
not ( n8917 , n8887 );
or ( n8918 , n8916 , n8917 );
xor ( n8919 , n547 , n7536 );
nand ( n8920 , n8919 , n6854 );
nand ( n8921 , n8918 , n8920 );
xor ( n8922 , n8915 , n8921 );
and ( n8923 , n8036 , n5398 );
not ( n8924 , n6811 );
not ( n8925 , n8919 );
or ( n8926 , n8924 , n8925 );
xor ( n8927 , n7718 , n547 );
nand ( n8928 , n8927 , n6854 );
nand ( n8929 , n8926 , n8928 );
xor ( n8930 , n8923 , n8929 );
and ( n8931 , n8927 , n6811 );
not ( n8932 , n7626 );
not ( n8933 , n7731 );
or ( n8934 , n8932 , n8933 );
nand ( n8935 , n7696 , n77459 );
nand ( n8936 , n8934 , n8935 );
nor ( n8937 , n8931 , n8936 );
and ( n8938 , n7696 , n548 );
nor ( n8939 , n8938 , n8428 );
not ( n8940 , n548 );
not ( n8941 , n8940 );
not ( n8942 , n7731 );
or ( n8943 , n8941 , n8942 );
nand ( n8944 , n8943 , n549 );
nand ( n8945 , n8939 , n8944 );
nor ( n8946 , n8937 , n8945 );
and ( n8947 , n8930 , n8946 );
and ( n8948 , n8923 , n8929 );
or ( n8949 , n8947 , n8948 );
and ( n8950 , n8922 , n8949 );
and ( n8951 , n8915 , n8921 );
or ( n8952 , n8950 , n8951 );
not ( n8953 , n552 );
and ( n8954 , n551 , n5644 );
not ( n8955 , n551 );
and ( n8956 , n8955 , n5643 );
nor ( n8957 , n8954 , n8956 );
not ( n8958 , n8957 );
or ( n8959 , n8953 , n8958 );
not ( n8960 , n551 );
not ( n8961 , n5530 );
or ( n8962 , n8960 , n8961 );
nand ( n8963 , n8076 , n6752 );
nand ( n8964 , n8962 , n8963 );
nand ( n8965 , n8964 , n6802 );
nand ( n78785 , n8959 , n8965 );
xor ( n78786 , n8952 , n78785 );
xor ( n8968 , n8889 , n78710 );
xor ( n8969 , n8968 , n8901 );
and ( n8970 , n78786 , n8969 );
and ( n8971 , n8952 , n78785 );
or ( n8972 , n8970 , n8971 );
not ( n8973 , n8972 );
nand ( n8974 , n8914 , n8973 );
xor ( n8975 , n8952 , n78785 );
xor ( n8976 , n8975 , n8969 );
not ( n8977 , n5905 );
not ( n8978 , n78718 );
or ( n8979 , n8977 , n8978 );
and ( n8980 , n549 , n7277 );
not ( n8981 , n549 );
and ( n8982 , n8981 , n7276 );
or ( n8983 , n8980 , n8982 );
nand ( n8984 , n8983 , n6489 );
nand ( n8985 , n8979 , n8984 );
not ( n8986 , n6802 );
not ( n8987 , n5823 );
or ( n8988 , n8986 , n8987 );
nand ( n8989 , n8964 , n552 );
nand ( n8990 , n8988 , n8989 );
xor ( n8991 , n8985 , n8990 );
xor ( n8992 , n8915 , n8921 );
xor ( n78812 , n8992 , n8949 );
and ( n8994 , n8991 , n78812 );
and ( n8995 , n8985 , n8990 );
or ( n8996 , n8994 , n8995 );
nor ( n8997 , n8976 , n8996 );
not ( n8998 , n5905 );
not ( n8999 , n8983 );
or ( n9000 , n8998 , n8999 );
and ( n9001 , n549 , n7857 );
not ( n9002 , n549 );
and ( n9003 , n9002 , n7414 );
or ( n9004 , n9001 , n9003 );
nand ( n9005 , n9004 , n6489 );
nand ( n9006 , n9000 , n9005 );
xor ( n9007 , n8923 , n8929 );
xor ( n9008 , n9007 , n8946 );
xor ( n9009 , n9006 , n9008 );
not ( n9010 , n7328 );
not ( n9011 , n9010 );
nand ( n9012 , n9011 , n5822 );
nand ( n9013 , n6909 , n6802 );
nand ( n9014 , n8848 , n7325 );
nand ( n9015 , n9012 , n9013 , n9014 );
and ( n9016 , n9009 , n9015 );
and ( n9017 , n9006 , n9008 );
or ( n9018 , n9016 , n9017 );
not ( n9019 , n9018 );
xor ( n9020 , n8985 , n8990 );
xor ( n9021 , n9020 , n78812 );
not ( n9022 , n9021 );
nand ( n9023 , n9019 , n9022 );
nor ( n9024 , n7735 , n6810 );
not ( n9025 , n5905 );
and ( n9026 , n549 , n7700 );
not ( n9027 , n549 );
and ( n9028 , n9027 , n7536 );
or ( n9029 , n9026 , n9028 );
not ( n9030 , n9029 );
or ( n9031 , n9025 , n9030 );
not ( n9032 , n549 );
not ( n9033 , n8042 );
or ( n9034 , n9032 , n9033 );
not ( n9035 , n549 );
nand ( n9036 , n9035 , n7718 );
nand ( n9037 , n9034 , n9036 );
nand ( n9038 , n9037 , n6489 );
nand ( n9039 , n9031 , n9038 );
xor ( n9040 , n9024 , n9039 );
and ( n9041 , n7736 , n550 );
nor ( n9042 , n9041 , n7018 );
not ( n9043 , n550 );
not ( n9044 , n9043 );
not ( n9045 , n7731 );
or ( n9046 , n9044 , n9045 );
nand ( n9047 , n9046 , n551 );
and ( n9048 , n9042 , n9047 );
not ( n9049 , n5905 );
not ( n9050 , n9037 );
or ( n9051 , n9049 , n9050 );
and ( n9052 , n7736 , n7305 );
and ( n9053 , n7731 , n7307 );
nor ( n9054 , n9052 , n9053 );
nand ( n9055 , n9051 , n9054 );
and ( n9056 , n9048 , n9055 );
xor ( n9057 , n9040 , n9056 );
not ( n9058 , n552 );
and ( n9059 , n7275 , n551 );
not ( n9060 , n7275 );
and ( n9061 , n9060 , n6752 );
or ( n9062 , n9059 , n9061 );
not ( n9063 , n9062 );
or ( n9064 , n9058 , n9063 );
and ( n9065 , n7414 , n6752 );
not ( n9066 , n7414 );
and ( n9067 , n9066 , n551 );
or ( n9068 , n9065 , n9067 );
nand ( n9069 , n9068 , n6802 );
nand ( n9070 , n9064 , n9069 );
or ( n9071 , n9057 , n9070 );
xor ( n9072 , n9048 , n9055 );
not ( n9073 , n9072 );
not ( n9074 , n7537 );
not ( n9075 , n6802 );
not ( n9076 , n9075 );
and ( n9077 , n9074 , n9076 );
and ( n9078 , n9068 , n552 );
nor ( n9079 , n9077 , n9078 );
nand ( n9080 , n9073 , n9079 );
not ( n9081 , n9080 );
and ( n9082 , n8036 , n5905 );
not ( n9083 , n551 );
not ( n9084 , n8042 );
or ( n9085 , n9083 , n9084 );
nand ( n9086 , n7718 , n6752 );
nand ( n9087 , n9085 , n9086 );
and ( n9088 , n552 , n9087 );
and ( n9089 , n7731 , n6868 );
nor ( n9090 , n9088 , n9089 );
nand ( n9091 , n7695 , n552 );
nand ( n9092 , n551 , n9091 );
nor ( n9093 , n9090 , n9092 );
xor ( n9094 , n9082 , n9093 );
not ( n9095 , n7537 );
nand ( n9096 , n9095 , n7325 );
nand ( n9097 , n9087 , n6802 );
nand ( n9098 , n7537 , n7328 );
nand ( n9099 , n9096 , n9097 , n9098 );
and ( n9100 , n9094 , n9099 );
or ( n9102 , n9100 , C0 );
not ( n9103 , n9102 );
or ( n9104 , n9081 , n9103 );
not ( n9105 , n9079 );
nand ( n9106 , n9105 , n9072 );
nand ( n9107 , n9104 , n9106 );
and ( n78926 , n9071 , n9107 );
and ( n78927 , n9057 , n9070 );
nor ( n9110 , n78926 , n78927 );
xor ( n9111 , n8937 , n8945 );
not ( n9112 , n5905 );
not ( n9113 , n9004 );
or ( n9114 , n9112 , n9113 );
nand ( n9115 , n9029 , n6489 );
nand ( n9116 , n9114 , n9115 );
xor ( n9117 , n9111 , n9116 );
nand ( n9118 , n7328 , n7243 );
nand ( n9119 , n6909 , n7325 );
nand ( n9120 , n9062 , n6802 );
nand ( n9121 , n9118 , n9119 , n9120 );
xor ( n9122 , n9117 , n9121 );
xor ( n9123 , n9024 , n9039 );
and ( n9124 , n9123 , n9056 );
and ( n9125 , n9024 , n9039 );
or ( n9126 , n9124 , n9125 );
nor ( n9127 , n9122 , n9126 );
or ( n9128 , n9110 , n9127 );
nand ( n9129 , n9122 , n9126 );
nand ( n9130 , n9128 , n9129 );
not ( n9131 , n9130 );
xor ( n9132 , n9006 , n9008 );
xor ( n9133 , n9132 , n9015 );
not ( n9134 , n9133 );
xor ( n9135 , n9111 , n9116 );
and ( n9136 , n9135 , n9121 );
and ( n9137 , n9111 , n9116 );
or ( n9138 , n9136 , n9137 );
not ( n9139 , n9138 );
nand ( n9140 , n9134 , n9139 );
not ( n9141 , n9140 );
or ( n9142 , n9131 , n9141 );
nand ( n9143 , n9133 , n9138 );
nand ( n9144 , n9142 , n9143 );
and ( n9145 , n9023 , n9144 );
nand ( n9146 , n9021 , n9018 );
not ( n9147 , n9146 );
nor ( n9148 , n9145 , n9147 );
or ( n9149 , n8997 , n9148 );
nand ( n9150 , n8976 , n8996 );
nand ( n9151 , n9149 , n9150 );
and ( n9152 , n8974 , n9151 );
nand ( n9153 , n8913 , n8972 );
not ( n9154 , n9153 );
nor ( n9155 , n9152 , n9154 );
or ( n9156 , n8911 , n9155 );
nand ( n78975 , n8874 , n8910 );
nand ( n9158 , n9156 , n78975 );
not ( n9159 , n9158 );
or ( n9160 , n8872 , n9159 );
nand ( n9161 , n8808 , n78688 );
nand ( n9162 , n9160 , n9161 );
not ( n78981 , n9162 );
or ( n9164 , n8806 , n78981 );
not ( n9165 , n8687 );
not ( n9166 , n8741 );
nand ( n9167 , n9165 , n9166 );
and ( n9168 , n8745 , n8803 );
and ( n9169 , n9167 , n9168 );
not ( n9170 , n8687 );
nor ( n9171 , n9170 , n9166 );
nor ( n9172 , n9169 , n9171 );
nand ( n9173 , n9164 , n9172 );
not ( n9174 , n9173 );
or ( n9175 , n8685 , n9174 );
buf ( n9176 , n8623 );
nand ( n9177 , n9176 , n8682 );
nand ( n9178 , n9175 , n9177 );
not ( n9179 , n9178 );
or ( n9180 , n8621 , n9179 );
nand ( n9181 , n8528 , n8618 );
not ( n9182 , n9181 );
nor ( n9183 , n8525 , n8482 );
not ( n9184 , n9183 );
and ( n9185 , n9182 , n9184 );
nand ( n9186 , n8525 , n8482 );
not ( n9187 , n9186 );
nor ( n9188 , n9185 , n9187 );
nand ( n9189 , n9180 , n9188 );
not ( n9190 , n9189 );
xor ( n9191 , n8505 , n8518 );
and ( n9192 , n9191 , n8523 );
and ( n9193 , n8505 , n8518 );
or ( n9194 , n9192 , n9193 );
xor ( n9195 , n8097 , n8107 );
xor ( n9196 , n9195 , n8110 );
xor ( n9197 , n9194 , n9196 );
xor ( n9198 , n8507 , n8511 );
and ( n9199 , n9198 , n8517 );
and ( n9200 , n8507 , n8511 );
or ( n9201 , n9199 , n9200 );
xor ( n9202 , n7965 , n7971 );
xor ( n9203 , n9202 , n7983 );
xor ( n9204 , n9201 , n9203 );
xor ( n9205 , n8487 , n8489 );
and ( n9206 , n9205 , n78319 );
and ( n9207 , n8487 , n8489 );
or ( n9208 , n9206 , n9207 );
xor ( n9209 , n9204 , n9208 );
and ( n9210 , n9197 , n9209 );
and ( n9211 , n9194 , n9196 );
or ( n9212 , n9210 , n9211 );
not ( n9213 , n9212 );
not ( n9214 , n9213 );
xor ( n9215 , n9201 , n9203 );
and ( n9216 , n9215 , n9208 );
and ( n9217 , n9201 , n9203 );
or ( n9218 , n9216 , n9217 );
xor ( n9219 , n7963 , n7986 );
xor ( n9220 , n9219 , n7998 );
xor ( n9221 , n9218 , n9220 );
xor ( n9222 , n8020 , n8022 );
xor ( n9223 , n9222 , n8113 );
xor ( n9224 , n9221 , n9223 );
not ( n9225 , n9224 );
not ( n9226 , n9225 );
or ( n9227 , n9214 , n9226 );
xor ( n9228 , n9194 , n9196 );
xor ( n9229 , n9228 , n9209 );
xor ( n9230 , n8495 , n8499 );
and ( n9231 , n9230 , n8524 );
and ( n9232 , n8495 , n8499 );
or ( n9233 , n9231 , n9232 );
or ( n9234 , n9229 , n9233 );
nand ( n9235 , n9227 , n9234 );
xor ( n9236 , n8018 , n8116 );
xor ( n9237 , n9236 , n8119 );
xor ( n9238 , n9218 , n9220 );
and ( n9239 , n9238 , n9223 );
and ( n9240 , n9218 , n9220 );
or ( n9241 , n9239 , n9240 );
nor ( n9242 , n9237 , n9241 );
nor ( n79061 , n9235 , n9242 );
not ( n9247 , n79061 );
or ( n79063 , n9190 , n9247 );
not ( n9249 , n9237 );
not ( n9250 , n9241 );
nand ( n9251 , n9249 , n9250 );
nor ( n9252 , n9212 , n9224 );
nand ( n9253 , n9229 , n9233 );
or ( n9254 , n9252 , n9253 );
nand ( n9255 , n9224 , n9212 );
nand ( n9256 , n9254 , n9255 );
and ( n9257 , n9251 , n9256 );
nand ( n9258 , n9237 , n9241 );
not ( n9259 , n9258 );
nor ( n9260 , n9257 , n9259 );
nand ( n9261 , n79063 , n9260 );
and ( n9262 , n7603 , n78009 , n8186 , n9261 );
nor ( n9263 , n8171 , n9262 );
not ( n9264 , n545 );
not ( n9265 , n6826 );
nand ( n9266 , n9265 , n6836 , n6838 , n6841 );
not ( n9267 , n9266 );
or ( n9268 , n9264 , n9267 );
nand ( n9269 , n6843 , n4440 );
nand ( n9270 , n9268 , n9269 );
nand ( n9271 , n9270 , n5399 );
nand ( n79087 , n75270 , n75018 );
nand ( n9276 , n9271 , n79087 );
not ( n9277 , n552 );
and ( n9278 , n7094 , n76988 );
not ( n9279 , n9278 );
not ( n9280 , n6771 );
or ( n9281 , n9279 , n9280 );
not ( n9282 , n76988 );
not ( n9283 , n7099 );
or ( n9284 , n9282 , n9283 );
nand ( n9285 , n9284 , n7148 );
not ( n9286 , n9285 );
nand ( n79099 , n9281 , n9286 );
not ( n79100 , n79099 );
xor ( n9289 , n7110 , n7117 );
and ( n9290 , n9289 , n7123 );
and ( n9291 , n7110 , n7117 );
or ( n9292 , n9290 , n9291 );
and ( n9293 , n507 , n489 );
not ( n9294 , n7111 );
not ( n79107 , n6384 );
or ( n79108 , n9294 , n79107 );
xnor ( n9297 , n489 , n505 );
not ( n9298 , n9297 );
nand ( n9299 , n9298 , n1553 );
nand ( n9300 , n79108 , n9299 );
xor ( n9301 , n9293 , n9300 );
not ( n9302 , n6582 );
not ( n9303 , n6580 );
or ( n9304 , n9302 , n9303 );
nand ( n9305 , n9304 , n491 );
xor ( n9306 , n9301 , n9305 );
xor ( n9307 , n9292 , n9306 );
not ( n9308 , n7123 );
xor ( n9309 , n9307 , n9308 );
not ( n9310 , n9309 );
not ( n9311 , n7124 );
nand ( n9312 , n9311 , n7131 );
and ( n9313 , n7109 , n9312 );
and ( n9314 , n7128 , n7124 );
nor ( n9315 , n9313 , n9314 );
nand ( n9316 , n9310 , n9315 );
or ( n9317 , n9310 , n9315 );
nand ( n9318 , n9316 , n9317 );
nor ( n9319 , n9318 , n455 );
nand ( n9320 , n79100 , n9319 );
nand ( n9321 , n7037 , n7089 );
nor ( n9322 , n6634 , n9321 );
not ( n9323 , n9322 );
not ( n9324 , n76304 );
or ( n9325 , n9323 , n9324 );
not ( n9326 , n5989 );
not ( n9327 , n4187 );
or ( n9328 , n9326 , n9327 );
nor ( n9329 , n6076 , n76543 );
nand ( n9330 , n9328 , n9329 );
nand ( n9331 , n6080 , n6142 );
and ( n9332 , n76544 , n9331 );
nor ( n9333 , n9332 , n9321 );
and ( n9334 , n9330 , n9333 );
not ( n9335 , n7089 );
not ( n9336 , n7049 );
or ( n9337 , n9335 , n9336 );
nand ( n9338 , n9337 , n76933 );
nor ( n9339 , n9334 , n9338 );
nand ( n9340 , n9325 , n9339 );
not ( n9341 , n9340 );
xor ( n9342 , n7060 , n76925 );
and ( n9343 , n9342 , n7087 );
and ( n9344 , n7060 , n76925 );
or ( n9345 , n9343 , n9344 );
not ( n9346 , n9345 );
not ( n9347 , n7081 );
not ( n9348 , n1738 );
not ( n9349 , n1699 );
or ( n9350 , n9348 , n9349 );
nand ( n9351 , n9350 , n491 );
not ( n9352 , n1828 );
not ( n9353 , n7068 );
or ( n9354 , n9352 , n9353 );
xor ( n9355 , n489 , n1858 );
nand ( n9356 , n9355 , n71761 );
nand ( n9357 , n9354 , n9356 );
xor ( n9358 , n9351 , n9357 );
and ( n9359 , n489 , n6120 );
xor ( n9360 , n9358 , n9359 );
xor ( n9361 , n9347 , n9360 );
xor ( n9362 , n7070 , n76917 );
and ( n9363 , n9362 , n7081 );
and ( n9364 , n7070 , n76917 );
or ( n79177 , n9363 , n9364 );
xor ( n79178 , n9361 , n79177 );
not ( n9367 , n79178 );
xnor ( n9368 , n9346 , n9367 );
nor ( n9369 , n9368 , n5595 );
nand ( n9370 , n9341 , n9369 );
not ( n9371 , n9318 );
nor ( n9372 , n9371 , n455 );
nand ( n9373 , n9372 , n79099 );
nand ( n9374 , n9340 , n9368 , n455 );
nand ( n9375 , n9320 , n9370 , n9373 , n9374 );
and ( n9376 , n9375 , n6752 );
not ( n9377 , n9375 );
and ( n9378 , n9377 , n551 );
or ( n9379 , n9376 , n9378 );
not ( n9380 , n9379 );
or ( n9381 , n9277 , n9380 );
nand ( n9382 , n7093 , n7152 , n7155 , n7158 );
nand ( n9383 , n9382 , n6868 );
nand ( n9384 , n9381 , n9383 );
xor ( n9385 , n9276 , n9384 );
and ( n9386 , n76644 , n7305 );
not ( n9387 , n76644 );
and ( n9388 , n9387 , n7307 );
nor ( n9389 , n9386 , n9388 );
xor ( n79202 , n549 , n6751 );
nand ( n79203 , n79202 , n5905 );
nand ( n9392 , n9389 , n79203 );
and ( n9393 , n9385 , n9392 );
and ( n9394 , n9276 , n9384 );
or ( n9395 , n9393 , n9394 );
not ( n9396 , n541 );
not ( n9397 , n74999 );
or ( n79210 , n9396 , n9397 );
nand ( n79211 , n6937 , n5538 );
nand ( n9400 , n79210 , n79211 );
not ( n9401 , n9400 );
not ( n9402 , n5590 );
or ( n9403 , n9401 , n9402 );
not ( n9404 , n4937 );
not ( n9405 , n5538 );
or ( n9406 , n9404 , n9405 );
nand ( n9407 , n541 , n4933 );
nand ( n9408 , n9406 , n9407 );
nand ( n9409 , n9408 , n5551 );
nand ( n9410 , n9403 , n9409 );
not ( n9411 , n4445 );
not ( n9412 , n543 );
not ( n9413 , n7378 );
or ( n9414 , n9412 , n9413 );
nand ( n9415 , n4938 , n5264 );
nand ( n9416 , n9414 , n9415 );
not ( n9417 , n9416 );
or ( n9418 , n9411 , n9417 );
not ( n9419 , n543 );
not ( n9420 , n5393 );
or ( n9421 , n9419 , n9420 );
nand ( n9422 , n5392 , n4938 );
nand ( n9423 , n9421 , n9422 );
nand ( n9424 , n9423 , n5128 );
nand ( n9425 , n9418 , n9424 );
xor ( n9426 , n9410 , n9425 );
not ( n9427 , n545 );
not ( n9428 , n6479 );
or ( n9429 , n9427 , n9428 );
nand ( n9430 , n6478 , n4440 );
nand ( n9431 , n9429 , n9430 );
nand ( n9432 , n9431 , n5399 );
nand ( n9433 , n9270 , n75018 );
nand ( n9434 , n9432 , n9433 );
xor ( n9435 , n9426 , n9434 );
xor ( n9436 , n9395 , n9435 );
not ( n9437 , n6811 );
and ( n9438 , n547 , n6867 );
not ( n9439 , n547 );
and ( n9440 , n9439 , n7327 );
or ( n9441 , n9438 , n9440 );
not ( n9442 , n9441 );
or ( n9443 , n9437 , n9442 );
nand ( n9444 , n7179 , n6955 );
nand ( n9445 , n9443 , n9444 );
not ( n9446 , n5501 );
not ( n9447 , n537 );
not ( n9448 , n74151 );
or ( n9449 , n9447 , n9448 );
nand ( n9450 , n4247 , n5409 );
nand ( n9451 , n9449 , n9450 );
not ( n9452 , n9451 );
or ( n9453 , n9446 , n9452 );
nand ( n9454 , n5413 , n5758 );
nand ( n9455 , n9453 , n9454 );
and ( n9456 , n5725 , n5762 );
xor ( n9457 , n9455 , n9456 );
not ( n9458 , n539 );
not ( n9459 , n5866 );
or ( n9460 , n9458 , n9459 );
nand ( n79273 , n5581 , n4251 );
nand ( n9462 , n9460 , n79273 );
and ( n9463 , n9462 , n4433 );
not ( n9464 , n4224 );
nor ( n9465 , n9464 , n4431 );
nor ( n9466 , n9463 , n9465 );
nand ( n9467 , n8299 , n537 );
and ( n9468 , n9466 , n9467 );
not ( n9469 , n9466 );
not ( n9470 , n9467 );
and ( n9471 , n9469 , n9470 );
nor ( n9472 , n9468 , n9471 );
xor ( n9473 , n9457 , n9472 );
xor ( n9474 , n9445 , n9473 );
xor ( n9475 , n4436 , n75009 );
and ( n9476 , n9475 , n5401 );
and ( n9477 , n4436 , n75009 );
or ( n9478 , n9476 , n9477 );
and ( n9479 , n9474 , n9478 );
and ( n9480 , n9445 , n9473 );
or ( n9481 , n9479 , n9480 );
xor ( n9482 , n9436 , n9481 );
and ( n9483 , n76988 , n9316 );
and ( n9484 , n7094 , n9483 );
not ( n9485 , n9484 );
not ( n9486 , n6771 );
or ( n9487 , n9485 , n9486 );
and ( n9488 , n9285 , n9316 );
not ( n9489 , n9317 );
nor ( n9490 , n9488 , n9489 );
nand ( n9491 , n9487 , n9490 );
xor ( n9492 , n9292 , n9306 );
not ( n9493 , n7123 );
and ( n9494 , n9492 , n9493 );
and ( n9495 , n9292 , n9306 );
or ( n9496 , n9494 , n9495 );
or ( n9497 , n6595 , n9297 );
or ( n9498 , n6597 , n1824 );
nand ( n9499 , n9497 , n9498 );
nand ( n9500 , n506 , n489 );
xor ( n9501 , n9499 , n9500 );
xor ( n9502 , n9293 , n9300 );
and ( n9503 , n9502 , n9305 );
and ( n9504 , n9293 , n9300 );
or ( n9505 , n9503 , n9504 );
xor ( n9506 , n9501 , n9505 );
or ( n9507 , n9496 , n9506 );
nand ( n9508 , n9496 , n9506 );
nand ( n9509 , n9507 , n9508 );
and ( n9510 , n9491 , n9509 );
nor ( n9511 , n9510 , n455 );
not ( n9512 , n9511 );
not ( n9513 , n9491 );
not ( n9514 , n9509 );
nand ( n9515 , n9513 , n9514 );
not ( n9516 , n9515 );
or ( n9517 , n9512 , n9516 );
nor ( n9518 , n9367 , n9346 );
nor ( n9519 , n9340 , n9518 );
xor ( n9520 , n9347 , n9360 );
and ( n9521 , n9520 , n79177 );
and ( n9522 , n9347 , n9360 );
or ( n9523 , n9521 , n9522 );
not ( n9524 , n9523 );
not ( n9525 , n1828 );
not ( n9526 , n9355 );
or ( n9527 , n9525 , n9526 );
or ( n9528 , n1789 , n1649 );
nand ( n9529 , n9527 , n9528 );
nand ( n9530 , n1995 , n489 );
xor ( n9531 , n9529 , n9530 );
xor ( n9532 , n9351 , n9357 );
and ( n9533 , n9532 , n9359 );
and ( n9534 , n9351 , n9357 );
or ( n9535 , n9533 , n9534 );
xor ( n9536 , n9531 , n9535 );
not ( n9537 , n9536 );
or ( n9538 , n9524 , n9537 );
not ( n9539 , n9538 );
nand ( n9540 , n9524 , n9537 );
not ( n9541 , n9540 );
or ( n9542 , n9539 , n9541 );
nand ( n9543 , n9542 , n455 );
nand ( n9544 , n9519 , n9543 );
nand ( n9545 , n9540 , n9538 , n455 );
nand ( n9546 , n9346 , n9367 );
nand ( n9547 , n9340 , n9545 , n9546 );
nor ( n9548 , n9518 , n9546 );
nand ( n9549 , n9543 , n9548 );
nand ( n9550 , n9545 , n9518 );
nand ( n9551 , n9544 , n9547 , n9549 , n9550 );
nand ( n9552 , n9517 , n9551 );
not ( n9553 , n9552 );
not ( n9554 , n9553 );
nand ( n9555 , n9554 , n7325 );
nand ( n9556 , n9553 , n7328 );
not ( n9557 , n9375 );
nand ( n9558 , n9557 , n6868 );
nand ( n9559 , n9555 , n9556 , n9558 );
not ( n9560 , n5905 );
not ( n9561 , n549 );
not ( n9562 , n9561 );
not ( n9563 , n7160 );
or ( n9564 , n9562 , n9563 );
not ( n9565 , n7159 );
or ( n9566 , n9561 , n9565 );
nand ( n9567 , n9564 , n9566 );
not ( n9568 , n9567 );
or ( n9569 , n9560 , n9568 );
nand ( n9570 , n79202 , n6489 );
nand ( n9571 , n9569 , n9570 );
xor ( n9572 , n9559 , n9571 );
xor ( n9573 , n9455 , n9456 );
and ( n9574 , n9573 , n9472 );
and ( n9575 , n9455 , n9456 );
or ( n9576 , n9574 , n9575 );
xor ( n9577 , n9572 , n9576 );
not ( n9578 , n6955 );
not ( n9579 , n9441 );
or ( n9580 , n9578 , n9579 );
xor ( n79393 , n547 , n76644 );
nand ( n79394 , n79393 , n6811 );
nand ( n9583 , n9580 , n79394 );
not ( n9584 , n5590 );
not ( n9585 , n9408 );
or ( n9586 , n9584 , n9585 );
buf ( n9587 , n5703 );
nand ( n9588 , n5551 , n9587 );
nand ( n9589 , n9586 , n9588 );
xor ( n9590 , n5710 , n5718 );
and ( n9591 , n9590 , n5763 );
and ( n9592 , n5710 , n5718 );
or ( n9593 , n9591 , n9592 );
xor ( n9594 , n9589 , n9593 );
buf ( n9595 , n5128 );
not ( n9596 , n9595 );
not ( n9597 , n9416 );
or ( n9598 , n9596 , n9597 );
nand ( n9599 , n5126 , n4445 );
nand ( n9600 , n9598 , n9599 );
and ( n9601 , n9594 , n9600 );
and ( n9602 , n9589 , n9593 );
or ( n9603 , n9601 , n9602 );
xor ( n9604 , n9583 , n9603 );
not ( n9605 , n5413 );
not ( n9606 , n9451 );
or ( n9607 , n9605 , n9606 );
not ( n9608 , n4425 );
not ( n9609 , n5409 );
and ( n9610 , n9608 , n9609 );
and ( n9611 , n7798 , n5409 );
nor ( n9612 , n9610 , n9611 );
not ( n9613 , n9612 );
nand ( n9614 , n9613 , n5501 );
nand ( n9615 , n9607 , n9614 );
nor ( n9616 , n9466 , n9467 );
xor ( n9617 , n9615 , n9616 );
and ( n9618 , n8290 , n537 );
not ( n9619 , n9618 );
not ( n9620 , n9619 );
not ( n9621 , n4433 );
not ( n9622 , n539 );
not ( n9623 , n5843 );
or ( n9624 , n9622 , n9623 );
nand ( n9625 , n5701 , n4251 );
nand ( n79438 , n9624 , n9625 );
not ( n9627 , n79438 );
or ( n79440 , n9621 , n9627 );
nand ( n9629 , n9462 , n4224 );
nand ( n9630 , n79440 , n9629 );
not ( n9631 , n9630 );
or ( n9632 , n9620 , n9631 );
buf ( n9633 , n9619 );
or ( n9634 , n9633 , n9630 );
nand ( n9635 , n9632 , n9634 );
xor ( n9636 , n9617 , n9635 );
xor ( n9637 , n9604 , n9636 );
xor ( n9638 , n9577 , n9637 );
xor ( n9639 , n9589 , n9593 );
xor ( n9640 , n9639 , n9600 );
xor ( n9641 , n5649 , n5764 );
and ( n9642 , n9641 , n5853 );
and ( n9643 , n5649 , n5764 );
or ( n9644 , n9642 , n9643 );
xor ( n9645 , n9640 , n9644 );
xor ( n9646 , n7029 , n7166 );
and ( n9647 , n9646 , n7181 );
and ( n9648 , n7029 , n7166 );
or ( n9649 , n9647 , n9648 );
and ( n9650 , n9645 , n9649 );
and ( n9651 , n9640 , n9644 );
or ( n9652 , n9650 , n9651 );
xor ( n9653 , n9638 , n9652 );
xor ( n9654 , n9482 , n9653 );
xor ( n9655 , n9445 , n9473 );
xor ( n9656 , n9655 , n9478 );
xor ( n9657 , n9276 , n9384 );
xor ( n9658 , n9657 , n9392 );
xor ( n9659 , n9656 , n9658 );
xor ( n9660 , n5402 , n5854 );
and ( n9661 , n9660 , n5901 );
and ( n9662 , n5402 , n5854 );
or ( n9663 , n9661 , n9662 );
and ( n9664 , n9659 , n9663 );
and ( n9665 , n9656 , n9658 );
or ( n9666 , n9664 , n9665 );
xor ( n9667 , n9654 , n9666 );
xor ( n9668 , n9640 , n9644 );
xor ( n9669 , n9668 , n9649 );
xor ( n9670 , n9656 , n9658 );
xor ( n9671 , n9670 , n9663 );
xor ( n9672 , n9669 , n9671 );
xor ( n9673 , n7016 , n7182 );
and ( n9674 , n9673 , n7210 );
and ( n9675 , n7016 , n7182 );
or ( n9676 , n9674 , n9675 );
and ( n9677 , n9672 , n9676 );
and ( n9678 , n9669 , n9671 );
or ( n9679 , n9677 , n9678 );
nor ( n9680 , n9667 , n9679 );
not ( n9681 , n9680 );
xor ( n9682 , n9410 , n9425 );
and ( n9683 , n9682 , n9434 );
and ( n9684 , n9410 , n9425 );
or ( n9685 , n9683 , n9684 );
not ( n9686 , n5590 );
not ( n9687 , n541 );
not ( n9688 , n5265 );
or ( n9689 , n9687 , n9688 );
nand ( n9690 , n5264 , n5538 );
nand ( n9691 , n9689 , n9690 );
not ( n9692 , n9691 );
or ( n9693 , n9686 , n9692 );
nand ( n9694 , n9400 , n5551 );
nand ( n9695 , n9693 , n9694 );
not ( n9696 , n5399 );
not ( n9697 , n545 );
not ( n9698 , n7324 );
or ( n9699 , n9697 , n9698 );
nand ( n9700 , n6440 , n4440 );
nand ( n9701 , n9699 , n9700 );
not ( n9702 , n9701 );
or ( n9703 , n9696 , n9702 );
nand ( n9704 , n9431 , n75018 );
nand ( n9705 , n9703 , n9704 );
xor ( n9706 , n9695 , n9705 );
not ( n9707 , n5905 );
and ( n9708 , n549 , n9557 );
not ( n9709 , n549 );
and ( n9710 , n9709 , n9375 );
or ( n9711 , n9708 , n9710 );
not ( n79524 , n9711 );
or ( n9716 , n9707 , n79524 );
nand ( n79526 , n9567 , n6489 );
nand ( n9718 , n9716 , n79526 );
xor ( n9719 , n9706 , n9718 );
xor ( n9720 , n9685 , n9719 );
nand ( n9721 , n6848 , n7448 );
nand ( n9722 , n9423 , n4445 );
not ( n9723 , n7444 );
nand ( n9724 , n9723 , n6847 );
nand ( n9725 , n9721 , n9722 , n9724 );
xor ( n9726 , n9615 , n9616 );
and ( n9727 , n9726 , n9635 );
and ( n9728 , n9615 , n9616 );
or ( n9729 , n9727 , n9728 );
xor ( n9730 , n9725 , n9729 );
not ( n9731 , n6955 );
not ( n9732 , n79393 );
or ( n9733 , n9731 , n9732 );
nand ( n9734 , n6750 , n6631 );
not ( n9735 , n9734 );
and ( n79545 , n547 , n9735 );
not ( n9740 , n547 );
and ( n9741 , n9740 , n6751 );
or ( n9742 , n79545 , n9741 );
nand ( n9743 , n9742 , n6811 );
nand ( n9744 , n9733 , n9743 );
xor ( n9745 , n9730 , n9744 );
xor ( n9746 , n9720 , n9745 );
xor ( n9747 , n9577 , n9637 );
and ( n9748 , n9747 , n9652 );
and ( n9749 , n9577 , n9637 );
or ( n9750 , n9748 , n9749 );
xor ( n9751 , n9746 , n9750 );
xor ( n9752 , n9583 , n9603 );
and ( n9753 , n9752 , n9636 );
and ( n9754 , n9583 , n9603 );
or ( n9755 , n9753 , n9754 );
not ( n9756 , n6868 );
not ( n9757 , n9554 );
not ( n9758 , n9757 );
not ( n9759 , n9758 );
or ( n9760 , n9756 , n9759 );
not ( n9761 , n551 );
not ( n9762 , n455 );
not ( n9763 , n9340 );
not ( n9764 , n9540 );
not ( n9765 , n9518 );
or ( n9766 , n9764 , n9765 );
nand ( n9767 , n9766 , n9538 );
or ( n9768 , n1828 , n71761 );
nand ( n9769 , n9768 , n489 );
and ( n9770 , n489 , n1858 );
xor ( n9771 , n9769 , n9770 );
not ( n9772 , n9530 );
xor ( n9773 , n9771 , n9772 );
not ( n9774 , n9773 );
xor ( n9775 , n9529 , n9530 );
and ( n9776 , n9775 , n9535 );
and ( n9777 , n9529 , n9530 );
or ( n9778 , n9776 , n9777 );
not ( n9779 , n9778 );
or ( n9780 , n9774 , n9779 );
or ( n9781 , n9778 , n9773 );
nand ( n9782 , n9780 , n9781 );
nor ( n9783 , n9767 , n9782 );
nand ( n9784 , n9763 , n9783 );
nand ( n9785 , n9546 , n9540 );
not ( n9786 , n9782 );
nor ( n9787 , n9785 , n9786 );
nand ( n79594 , n9787 , n9340 );
not ( n79595 , n9782 );
not ( n9790 , n9767 );
nand ( n9791 , n79595 , n9790 , n9785 );
not ( n9792 , n9786 );
nand ( n9793 , n9792 , n9767 );
nand ( n9794 , n9784 , n79594 , n9791 , n9793 );
not ( n9795 , n9794 );
or ( n9796 , n9762 , n9795 );
xor ( n9797 , n9499 , n9500 );
and ( n9798 , n9797 , n9505 );
and ( n9799 , n9499 , n9500 );
or ( n9800 , n9798 , n9799 );
not ( n9801 , n9800 );
not ( n9802 , n9500 );
nand ( n9803 , n505 , n489 );
not ( n9804 , n9803 );
or ( n9805 , n6384 , n1553 );
nand ( n9806 , n9805 , n489 );
not ( n9807 , n9806 );
or ( n9808 , n9804 , n9807 );
or ( n9809 , n9806 , n9803 );
nand ( n9810 , n9808 , n9809 );
not ( n9811 , n9810 );
or ( n9812 , n9802 , n9811 );
or ( n9813 , n9810 , n9500 );
nand ( n9814 , n9812 , n9813 );
not ( n9815 , n9814 );
and ( n9816 , n9801 , n9815 );
and ( n9817 , n9800 , n9814 );
nor ( n9818 , n9816 , n9817 );
not ( n9819 , n9818 );
not ( n9820 , n9819 );
not ( n9821 , n6762 );
not ( n9822 , n6765 );
or ( n9823 , n9821 , n9822 );
and ( n9824 , n9483 , n9507 );
and ( n9825 , n9824 , n7094 );
nand ( n9826 , n9823 , n9825 );
not ( n9827 , n7094 );
not ( n9828 , n6506 );
or ( n9829 , n9827 , n9828 );
nand ( n9830 , n9829 , n7100 );
nand ( n9831 , n9830 , n9824 );
not ( n9832 , n9316 );
not ( n9833 , n7147 );
or ( n9834 , n9832 , n9833 );
nand ( n9835 , n9834 , n9317 );
and ( n9836 , n9835 , n9507 );
not ( n9837 , n9508 );
nor ( n9838 , n9836 , n9837 );
nand ( n9839 , n9826 , n9831 , n9838 );
not ( n9840 , n9839 );
or ( n9841 , n9820 , n9840 );
not ( n9842 , n9838 );
nor ( n9843 , n9842 , n9819 );
nand ( n9844 , n9826 , n9831 , n9843 );
nand ( n9845 , n9841 , n9844 );
nand ( n79652 , n9845 , n70470 );
nand ( n79653 , n9796 , n79652 );
not ( n9848 , n79653 );
not ( n9849 , n9848 );
or ( n9850 , n9761 , n9849 );
or ( n9851 , n551 , n9848 );
nand ( n9852 , n9850 , n9851 );
nand ( n9853 , n9852 , n552 );
nand ( n9854 , n9760 , n9853 );
buf ( n9855 , n4224 );
nand ( n9856 , n79438 , n9855 );
nand ( n9857 , n4933 , n5781 );
nand ( n9858 , n4937 , n5787 );
nand ( n9859 , n9856 , n9857 , n9858 );
not ( n9860 , n4224 );
not ( n9861 , n9462 );
or ( n9862 , n9860 , n9861 );
nand ( n9863 , n79438 , n4433 );
nand ( n9864 , n9862 , n9863 );
nand ( n9865 , n9864 , n9618 );
not ( n9866 , n9865 );
xor ( n9867 , n9859 , n9866 );
and ( n9868 , n7234 , n537 );
not ( n9869 , n9868 );
not ( n9870 , n9869 );
or ( n9871 , n9612 , n5713 );
not ( n9872 , n537 );
not ( n9873 , n5866 );
or ( n9874 , n9872 , n9873 );
nand ( n9875 , n5869 , n5409 );
nand ( n9876 , n9874 , n9875 );
nand ( n9877 , n9876 , n5501 );
nand ( n9878 , n9871 , n9877 );
not ( n9879 , n9878 );
or ( n9880 , n9870 , n9879 );
nand ( n9881 , n9877 , n9868 , n9871 );
nand ( n9882 , n9880 , n9881 );
xor ( n79689 , n9867 , n9882 );
xor ( n79690 , n9854 , n79689 );
xor ( n9885 , n9559 , n9571 );
and ( n9886 , n9885 , n9576 );
and ( n9887 , n9559 , n9571 );
or ( n9888 , n9886 , n9887 );
xor ( n9889 , n79690 , n9888 );
xor ( n9890 , n9755 , n9889 );
xor ( n9891 , n9395 , n9435 );
and ( n9892 , n9891 , n9481 );
and ( n9893 , n9395 , n9435 );
or ( n9894 , n9892 , n9893 );
xor ( n9895 , n9890 , n9894 );
xor ( n9896 , n9751 , n9895 );
xor ( n9897 , n9482 , n9653 );
and ( n9898 , n9897 , n9666 );
and ( n9899 , n9482 , n9653 );
or ( n9900 , n9898 , n9899 );
nor ( n9901 , n9896 , n9900 );
not ( n9902 , n9901 );
xor ( n9903 , n9669 , n9671 );
xor ( n9904 , n9903 , n9676 );
not ( n9905 , n9904 );
xor ( n9906 , n5902 , n7011 );
and ( n9907 , n9906 , n7211 );
and ( n9908 , n5902 , n7011 );
or ( n9909 , n9907 , n9908 );
not ( n79716 , n9909 );
nand ( n9911 , n9905 , n79716 );
nand ( n9912 , n9681 , n9902 , n9911 );
or ( n9913 , n9263 , n9912 );
nor ( n9914 , n9901 , n9680 );
nand ( n9915 , n9904 , n9909 );
nand ( n9916 , n9667 , n9679 );
nand ( n9917 , n9915 , n9916 );
and ( n9918 , n9914 , n9917 );
nand ( n9919 , n9896 , n9900 );
not ( n9920 , n9919 );
nor ( n9921 , n9918 , n9920 );
nand ( n9922 , n9913 , n9921 );
buf ( n9923 , n9922 );
buf ( n9924 , n9923 );
xor ( n9925 , n9695 , n9705 );
and ( n9926 , n9925 , n9718 );
and ( n9927 , n9695 , n9705 );
or ( n9928 , n9926 , n9927 );
not ( n9929 , n5590 );
not ( n9930 , n541 );
not ( n9931 , n5392 );
not ( n9932 , n9931 );
or ( n9933 , n9930 , n9932 );
nand ( n9934 , n5392 , n5538 );
nand ( n9935 , n9933 , n9934 );
not ( n9936 , n9935 );
or ( n9937 , n9929 , n9936 );
buf ( n9938 , n5551 );
nand ( n9939 , n9691 , n9938 );
nand ( n9940 , n9937 , n9939 );
not ( n9941 , n75018 );
not ( n9942 , n9701 );
or ( n9943 , n9941 , n9942 );
not ( n9944 , n545 );
not ( n9945 , n76644 );
not ( n9946 , n9945 );
or ( n9947 , n9944 , n9946 );
nand ( n9948 , n76644 , n4440 );
nand ( n9949 , n9947 , n9948 );
nand ( n9950 , n9949 , n5399 );
nand ( n9951 , n9943 , n9950 );
xor ( n9952 , n9940 , n9951 );
not ( n9953 , n5905 );
xor ( n9954 , n549 , n9553 );
not ( n9955 , n9954 );
or ( n9956 , n9953 , n9955 );
nand ( n9957 , n9711 , n6489 );
nand ( n9958 , n9956 , n9957 );
xor ( n9959 , n9952 , n9958 );
xor ( n9960 , n9928 , n9959 );
not ( n9961 , n543 );
not ( n9962 , n7318 );
or ( n9963 , n9961 , n9962 );
nand ( n9964 , n7174 , n4938 );
nand ( n9965 , n9963 , n9964 );
nand ( n9966 , n9965 , n5128 );
not ( n9967 , n7230 );
nand ( n9968 , n9967 , n6844 );
nand ( n9969 , n6843 , n7236 );
nand ( n9970 , n9966 , n9968 , n9969 );
xor ( n9971 , n9859 , n9866 );
and ( n9972 , n9971 , n9882 );
and ( n9973 , n9859 , n9866 );
or ( n9974 , n9972 , n9973 );
xor ( n9975 , n9970 , n9974 );
not ( n9976 , n6854 );
not ( n9977 , n9742 );
or ( n9978 , n9976 , n9977 );
not ( n9979 , n8428 );
not ( n9980 , n7160 );
or ( n9981 , n9979 , n9980 );
or ( n9982 , n7160 , n8428 );
nand ( n9983 , n9981 , n9982 );
nand ( n9984 , n9983 , n6811 );
nand ( n9985 , n9978 , n9984 );
xor ( n9986 , n9975 , n9985 );
xor ( n79793 , n9960 , n9986 );
not ( n79794 , n6802 );
not ( n9989 , n9852 );
or ( n9990 , n79794 , n9989 );
not ( n9991 , n7325 );
nand ( n9992 , n9990 , n9991 );
not ( n9993 , n4434 );
not ( n9994 , n539 );
not ( n9995 , n74999 );
or ( n9996 , n9994 , n9995 );
nand ( n9997 , n74998 , n4251 );
nand ( n9998 , n9996 , n9997 );
not ( n9999 , n9998 );
or ( n10000 , n9993 , n9999 );
not ( n10001 , n4937 );
not ( n10002 , n5774 );
and ( n10003 , n10001 , n10002 );
and ( n10004 , n7936 , n5772 );
nor ( n10005 , n10003 , n10004 );
nand ( n10006 , n10000 , n10005 );
and ( n10007 , n9877 , n9871 );
nor ( n10008 , n10007 , n9869 );
xor ( n10009 , n10006 , n10008 );
and ( n10010 , n4429 , n537 );
not ( n10011 , n5501 );
not ( n10012 , n537 );
not ( n10013 , n7624 );
or ( n10014 , n10012 , n10013 );
nand ( n10015 , n7620 , n5409 );
nand ( n10016 , n10014 , n10015 );
not ( n10017 , n10016 );
or ( n10018 , n10011 , n10017 );
nand ( n10019 , n9876 , n5413 );
nand ( n10020 , n10018 , n10019 );
xor ( n10021 , n10010 , n10020 );
xor ( n10022 , n10009 , n10021 );
xor ( n10023 , n9992 , n10022 );
xor ( n10024 , n9725 , n9729 );
and ( n10025 , n10024 , n9744 );
and ( n10026 , n9725 , n9729 );
or ( n10027 , n10025 , n10026 );
xor ( n10028 , n10023 , n10027 );
xor ( n10029 , n9854 , n79689 );
and ( n10030 , n10029 , n9888 );
and ( n10031 , n9854 , n79689 );
or ( n10032 , n10030 , n10031 );
xor ( n10033 , n10028 , n10032 );
xor ( n10034 , n9685 , n9719 );
and ( n10035 , n10034 , n9745 );
and ( n10036 , n9685 , n9719 );
or ( n10037 , n10035 , n10036 );
xor ( n10038 , n10033 , n10037 );
xor ( n10039 , n79793 , n10038 );
xor ( n10040 , n9755 , n9889 );
and ( n10041 , n10040 , n9894 );
and ( n10042 , n9755 , n9889 );
or ( n10043 , n10041 , n10042 );
xor ( n10044 , n10039 , n10043 );
xor ( n10045 , n9746 , n9750 );
and ( n10046 , n10045 , n9895 );
and ( n10047 , n9746 , n9750 );
or ( n10048 , n10046 , n10047 );
nor ( n10049 , n10044 , n10048 );
not ( n10050 , n10049 );
nand ( n10051 , n10044 , n10048 );
buf ( n10052 , n10051 );
nand ( n10053 , n10050 , n10052 );
not ( n10054 , n10053 );
and ( n10055 , n9924 , n10054 );
not ( n10056 , n9924 );
and ( n10057 , n10056 , n10053 );
nor ( n10058 , n10055 , n10057 );
not ( n10059 , n10058 );
or ( n10060 , n4215 , n10059 );
not ( n10061 , n454 );
not ( n10062 , n504 );
not ( n10063 , n503 );
xor ( n10064 , n529 , n457 );
not ( n79871 , n10064 );
xor ( n10066 , n458 , n459 );
not ( n10067 , n10066 );
not ( n10068 , n10067 );
not ( n10069 , n10068 );
or ( n10070 , n79871 , n10069 );
xnor ( n79877 , n458 , n457 );
xor ( n10072 , n458 , n459 );
nor ( n10073 , n79877 , n10072 );
and ( n10074 , n530 , n457 );
not ( n10075 , n530 );
and ( n10076 , n10075 , n2714 );
nor ( n10077 , n10074 , n10076 );
nand ( n10078 , n10073 , n10077 );
nand ( n10079 , n10070 , n10078 );
xor ( n10080 , n528 , n459 );
not ( n10081 , n10080 );
not ( n10082 , n460 );
nand ( n10083 , n3088 , n10082 , n459 );
nand ( n10084 , n2348 , n460 , n461 );
nand ( n10085 , n10083 , n10084 );
not ( n10086 , n10085 );
not ( n10087 , n10086 );
not ( n10088 , n10087 );
or ( n10089 , n10081 , n10088 );
and ( n10090 , n461 , n460 );
not ( n10091 , n461 );
and ( n10092 , n10091 , n2528 );
nor ( n10093 , n10090 , n10092 );
buf ( n10094 , n10093 );
xor ( n10095 , n527 , n459 );
nand ( n10096 , n10094 , n10095 );
nand ( n10097 , n10089 , n10096 );
xor ( n10098 , n10079 , n10097 );
xor ( n10099 , n524 , n463 );
not ( n10100 , n10099 );
not ( n10101 , n465 );
and ( n10102 , n464 , n10101 );
not ( n10103 , n464 );
and ( n10104 , n10103 , n465 );
nor ( n10105 , n10102 , n10104 );
xor ( n10106 , n464 , n463 );
nand ( n10107 , n10105 , n10106 );
not ( n10108 , n10107 );
not ( n10109 , n10108 );
or ( n10110 , n10100 , n10109 );
xor ( n10111 , n464 , n465 );
buf ( n10112 , n10111 );
xor ( n10113 , n463 , n523 );
nand ( n10114 , n10112 , n10113 );
nand ( n10115 , n10110 , n10114 );
and ( n10116 , n10098 , n10115 );
and ( n10117 , n10079 , n10097 );
or ( n10118 , n10116 , n10117 );
not ( n10119 , n10095 );
not ( n10120 , n10085 );
or ( n10121 , n10119 , n10120 );
xor ( n10122 , n526 , n459 );
nand ( n10123 , n10094 , n10122 );
nand ( n10124 , n10121 , n10123 );
not ( n10125 , n10064 );
nor ( n10126 , n79877 , n10072 );
buf ( n10127 , n10126 );
not ( n10128 , n10127 );
or ( n10129 , n10125 , n10128 );
xor ( n10130 , n457 , n528 );
nand ( n10131 , n10068 , n10130 );
nand ( n10132 , n10129 , n10131 );
xor ( n10133 , n10124 , n10132 );
xor ( n10134 , n521 , n465 );
not ( n10135 , n10134 );
nand ( n10136 , n2554 , n467 );
not ( n10137 , n467 );
nand ( n10138 , n10137 , n466 );
nand ( n10139 , n10136 , n10138 );
not ( n10140 , n10139 );
xor ( n10141 , n466 , n465 );
and ( n10142 , n10140 , n10141 );
not ( n10143 , n10142 );
or ( n10144 , n10135 , n10143 );
xor ( n10145 , n466 , n467 );
nand ( n10146 , n10145 , n465 );
nand ( n10147 , n10144 , n10146 );
xor ( n10148 , n10133 , n10147 );
xor ( n10149 , n10118 , n10148 );
not ( n79956 , n468 );
and ( n10154 , n79956 , n469 );
not ( n79958 , n469 );
and ( n10156 , n79958 , n468 );
nor ( n10157 , n10154 , n10156 );
not ( n10158 , n10157 );
xnor ( n10159 , n468 , n469 );
xor ( n10160 , n468 , n467 );
nand ( n10161 , n10159 , n10160 );
not ( n10162 , n10161 );
buf ( n10163 , n10162 );
not ( n10164 , n10163 );
not ( n10165 , n10164 );
or ( n10166 , n10158 , n10165 );
nand ( n10167 , n10166 , n467 );
not ( n10168 , n10167 );
xor ( n10169 , n522 , n465 );
not ( n10170 , n10169 );
not ( n10171 , n10142 );
or ( n10172 , n10170 , n10171 );
nand ( n10173 , n10145 , n10134 );
nand ( n10174 , n10172 , n10173 );
not ( n10175 , n10174 );
or ( n10176 , n10168 , n10175 );
nor ( n10177 , n10167 , n10174 );
xor ( n10178 , n526 , n461 );
not ( n79982 , n10178 );
xor ( n10183 , n461 , n462 );
not ( n10184 , n10183 );
and ( n10185 , n462 , n463 );
not ( n10186 , n462 );
not ( n10187 , n463 );
and ( n10188 , n10186 , n10187 );
nor ( n10189 , n10185 , n10188 );
or ( n10190 , n10184 , n10189 );
not ( n10191 , n10190 );
not ( n10192 , n10191 );
or ( n10193 , n79982 , n10192 );
xor ( n10194 , n462 , n463 );
xor ( n10195 , n525 , n461 );
nand ( n10196 , n10194 , n10195 );
nand ( n10197 , n10193 , n10196 );
not ( n10198 , n10197 );
or ( n10199 , n10177 , n10198 );
nand ( n10200 , n10176 , n10199 );
and ( n10201 , n10149 , n10200 );
and ( n10202 , n10118 , n10148 );
or ( n10203 , n10201 , n10202 );
not ( n10204 , n10122 );
not ( n10205 , n10085 );
or ( n10206 , n10204 , n10205 );
xor ( n10207 , n525 , n459 );
nand ( n10208 , n10094 , n10207 );
nand ( n10209 , n10206 , n10208 );
xor ( n10210 , n522 , n463 );
not ( n10211 , n10210 );
not ( n10212 , n10108 );
or ( n10213 , n10211 , n10212 );
xor ( n10214 , n521 , n463 );
nand ( n10215 , n10112 , n10214 );
nand ( n10216 , n10213 , n10215 );
xor ( n10217 , n10209 , n10216 );
not ( n10218 , n10145 );
not ( n10219 , n10218 );
xnor ( n10220 , n466 , n467 );
nand ( n10221 , n10220 , n10141 );
not ( n10222 , n10221 );
or ( n10223 , n10219 , n10222 );
nand ( n10224 , n10223 , n465 );
xor ( n10225 , n10217 , n10224 );
not ( n10226 , n10225 );
nand ( n10227 , n530 , n457 );
not ( n10228 , n10227 );
not ( n10229 , n10228 );
not ( n10230 , n10113 );
not ( n10231 , n10108 );
or ( n10232 , n10230 , n10231 );
nand ( n10233 , n10112 , n10210 );
nand ( n10234 , n10232 , n10233 );
not ( n10235 , n10234 );
not ( n10236 , n10235 );
or ( n10237 , n10229 , n10236 );
not ( n10238 , n10227 );
not ( n10239 , n10234 );
or ( n10240 , n10238 , n10239 );
not ( n10241 , n463 );
nand ( n10242 , n10241 , n462 );
nand ( n10243 , n1933 , n463 );
nand ( n10244 , n10242 , n10243 );
xor ( n10245 , n524 , n461 );
nand ( n10246 , n10244 , n10245 );
and ( n10247 , n462 , n463 );
not ( n10248 , n462 );
and ( n10249 , n10248 , n10187 );
nor ( n10250 , n10247 , n10249 );
not ( n10251 , n10250 );
nand ( n10252 , n10251 , n10183 );
not ( n10253 , n10252 );
nand ( n10254 , n10195 , n10253 );
nand ( n10255 , n10246 , n10254 );
nand ( n10256 , n10240 , n10255 );
nand ( n10257 , n10237 , n10256 );
not ( n10258 , n10257 );
not ( n10259 , n10258 );
and ( n10260 , n10226 , n10259 );
and ( n10261 , n10225 , n10258 );
nor ( n10262 , n10260 , n10261 );
nand ( n10263 , n529 , n457 );
not ( n10264 , n10130 );
not ( n10265 , n10127 );
or ( n10266 , n10264 , n10265 );
xor ( n10267 , n457 , n527 );
nand ( n10268 , n10068 , n10267 );
nand ( n10269 , n10266 , n10268 );
xor ( n10270 , n10263 , n10269 );
not ( n10271 , n10245 );
not ( n10272 , n10191 );
or ( n10273 , n10271 , n10272 );
xor ( n10274 , n523 , n461 );
nand ( n10275 , n10194 , n10274 );
nand ( n10276 , n10273 , n10275 );
xnor ( n10277 , n10270 , n10276 );
xor ( n10278 , n10234 , n10277 );
or ( n10279 , n10124 , n10132 );
nand ( n10280 , n10279 , n10147 );
nand ( n10281 , n10124 , n10132 );
nand ( n10282 , n10280 , n10281 );
xor ( n10283 , n10278 , n10282 );
or ( n10284 , n10262 , n10283 );
nand ( n80085 , n10283 , n10262 );
nand ( n80086 , n10284 , n80085 );
xor ( n10287 , n10203 , n80086 );
xor ( n10288 , n10079 , n10097 );
xor ( n10289 , n10288 , n10115 );
not ( n10290 , n10289 );
and ( n10291 , n532 , n457 );
xnor ( n10292 , n458 , n457 );
nor ( n10293 , n10292 , n10072 );
not ( n10294 , n10293 );
xor ( n10295 , n531 , n457 );
not ( n10296 , n10295 );
or ( n10297 , n10294 , n10296 );
nand ( n10298 , n10066 , n10077 );
nand ( n10299 , n10297 , n10298 );
xor ( n10300 , n10291 , n10299 );
xor ( n10301 , n525 , n463 );
not ( n10302 , n10301 );
not ( n10303 , n10108 );
or ( n10304 , n10302 , n10303 );
nand ( n10305 , n10112 , n10099 );
nand ( n10306 , n10304 , n10305 );
and ( n10307 , n10300 , n10306 );
and ( n10308 , n10291 , n10299 );
or ( n10309 , n10307 , n10308 );
not ( n10310 , n10309 );
or ( n10311 , n10290 , n10310 );
nor ( n10312 , n10289 , n10309 );
xor ( n10313 , n10174 , n10167 );
and ( n10314 , n10313 , n10198 );
not ( n10315 , n10313 );
and ( n10316 , n10315 , n10197 );
nor ( n10317 , n10314 , n10316 );
or ( n10318 , n10312 , n10317 );
nand ( n10319 , n10311 , n10318 );
not ( n10320 , n10319 );
xor ( n10321 , n521 , n467 );
not ( n10322 , n10321 );
not ( n10323 , n10162 );
or ( n10324 , n10322 , n10323 );
not ( n10325 , n468 );
not ( n10326 , n79958 );
or ( n10327 , n10325 , n10326 );
nand ( n10328 , n79956 , n469 );
nand ( n10329 , n10327 , n10328 );
nand ( n10330 , n10329 , n467 );
nand ( n10331 , n10324 , n10330 );
not ( n10332 , n10331 );
nand ( n10333 , n531 , n457 );
nand ( n10334 , n10332 , n10333 );
not ( n10335 , n10334 );
not ( n10336 , n3088 );
not ( n10337 , n463 );
and ( n10338 , n10336 , n10337 );
nor ( n10339 , n10338 , n462 );
not ( n10340 , n10339 );
xor ( n10341 , n527 , n461 );
not ( n10342 , n462 );
not ( n10343 , n463 );
nor ( n10344 , n10343 , n461 );
nor ( n10345 , n10342 , n10344 );
not ( n10346 , n10345 );
nand ( n10347 , n10340 , n10341 , n10346 );
nand ( n80148 , n10242 , n10243 );
nand ( n10349 , n80148 , n10178 );
nand ( n10350 , n10347 , n10349 );
xor ( n10351 , n465 , n523 );
not ( n10352 , n10351 );
not ( n10353 , n10221 );
not ( n10354 , n10353 );
or ( n10355 , n10352 , n10354 );
xor ( n10356 , n467 , n466 );
buf ( n10357 , n10356 );
nand ( n10358 , n10357 , n10169 );
nand ( n10359 , n10355 , n10358 );
xor ( n10360 , n10350 , n10359 );
xor ( n10361 , n529 , n459 );
not ( n10362 , n10361 );
not ( n10363 , n10085 );
or ( n10364 , n10362 , n10363 );
nand ( n10365 , n10094 , n10080 );
nand ( n10366 , n10364 , n10365 );
and ( n10367 , n10360 , n10366 );
and ( n10368 , n10350 , n10359 );
or ( n10369 , n10367 , n10368 );
not ( n10370 , n10369 );
or ( n10371 , n10335 , n10370 );
not ( n10372 , n10333 );
nand ( n10373 , n10331 , n10372 );
nand ( n10374 , n10371 , n10373 );
not ( n10375 , n10374 );
xor ( n10376 , n10228 , n10235 );
xor ( n10377 , n10376 , n10255 );
not ( n10378 , n10377 );
nand ( n10379 , n10375 , n10378 );
not ( n10380 , n10379 );
or ( n10381 , n10320 , n10380 );
not ( n10382 , n10378 );
nand ( n10383 , n10382 , n10374 );
nand ( n10384 , n10381 , n10383 );
and ( n10385 , n10287 , n10384 );
and ( n10386 , n10203 , n80086 );
or ( n10387 , n10385 , n10386 );
not ( n10388 , n10387 );
not ( n10389 , n10225 );
nand ( n10390 , n10389 , n10258 );
not ( n10391 , n10390 );
not ( n10392 , n10283 );
or ( n10393 , n10391 , n10392 );
nand ( n10394 , n10225 , n10257 );
nand ( n10395 , n10393 , n10394 );
not ( n10396 , n10395 );
not ( n10397 , n10396 );
xor ( n10398 , n10234 , n10277 );
and ( n10399 , n10398 , n10282 );
and ( n10400 , n10234 , n10277 );
or ( n10401 , n10399 , n10400 );
not ( n10402 , n10401 );
not ( n10403 , n10402 );
xor ( n10404 , n10209 , n10216 );
and ( n10405 , n10404 , n10224 );
and ( n10406 , n10209 , n10216 );
or ( n10407 , n10405 , n10406 );
and ( n10408 , n457 , n528 );
not ( n10409 , n10267 );
not ( n10410 , n10127 );
or ( n10411 , n10409 , n10410 );
xor ( n10412 , n457 , n526 );
nand ( n10413 , n10068 , n10412 );
nand ( n10414 , n10411 , n10413 );
xor ( n10415 , n10408 , n10414 );
not ( n10416 , n10214 );
not ( n10417 , n10108 );
or ( n10418 , n10416 , n10417 );
nand ( n10419 , n463 , n10112 );
nand ( n10420 , n10418 , n10419 );
xor ( n10421 , n10415 , n10420 );
xor ( n10422 , n10407 , n10421 );
not ( n10423 , n10207 );
not ( n10424 , n10087 );
or ( n10425 , n10423 , n10424 );
xor ( n10426 , n459 , n524 );
nand ( n10427 , n10094 , n10426 );
nand ( n10428 , n10425 , n10427 );
not ( n10429 , n10428 );
not ( n10430 , n10274 );
not ( n10431 , n10253 );
or ( n10432 , n10430 , n10431 );
xor ( n10433 , n522 , n461 );
nand ( n10434 , n10433 , n80148 );
nand ( n80235 , n10432 , n10434 );
not ( n80236 , n80235 );
and ( n10437 , n10429 , n80236 );
and ( n10438 , n10428 , n80235 );
nor ( n10439 , n10437 , n10438 );
not ( n10440 , n10439 );
not ( n10441 , n10263 );
not ( n10442 , n10441 );
not ( n10443 , n10276 );
or ( n10444 , n10442 , n10443 );
or ( n10445 , n10276 , n10441 );
not ( n10446 , n10130 );
not ( n10447 , n10127 );
or ( n10448 , n10446 , n10447 );
nand ( n10449 , n10448 , n10268 );
nand ( n10450 , n10445 , n10449 );
nand ( n10451 , n10444 , n10450 );
not ( n10452 , n10451 );
or ( n10453 , n10440 , n10452 );
or ( n10454 , n10451 , n10439 );
nand ( n10455 , n10453 , n10454 );
xor ( n10456 , n10422 , n10455 );
not ( n10457 , n10456 );
or ( n10458 , n10403 , n10457 );
not ( n10459 , n10456 );
nand ( n10460 , n10459 , n10401 );
nand ( n10461 , n10458 , n10460 );
not ( n10462 , n10461 );
not ( n10463 , n10462 );
or ( n10464 , n10397 , n10463 );
nand ( n10465 , n10395 , n10461 );
nand ( n10466 , n10464 , n10465 );
nand ( n10467 , n10388 , n10466 );
not ( n10468 , n10467 );
xor ( n10469 , n468 , n469 );
not ( n10470 , n10469 );
not ( n10471 , n10321 );
or ( n10472 , n10470 , n10471 );
xor ( n10473 , n468 , n469 );
not ( n10474 , n10473 );
xor ( n10475 , n522 , n467 );
nand ( n10476 , n10474 , n10475 , n10160 );
nand ( n10477 , n10472 , n10476 );
xor ( n10478 , n526 , n463 );
not ( n10479 , n10478 );
and ( n10480 , n10105 , n10106 );
not ( n10481 , n10480 );
or ( n10482 , n10479 , n10481 );
nand ( n10483 , n10112 , n10301 );
nand ( n10484 , n10482 , n10483 );
xor ( n10485 , n10477 , n10484 );
xor ( n10486 , n470 , n471 );
not ( n10487 , n10486 );
not ( n10488 , n10487 );
xor ( n10489 , n470 , n469 );
not ( n10490 , n10489 );
xor ( n10491 , n470 , n471 );
nor ( n10492 , n10490 , n10491 );
not ( n10493 , n10492 );
not ( n10494 , n10493 );
or ( n10495 , n10488 , n10494 );
nand ( n10496 , n10495 , n469 );
and ( n10497 , n10485 , n10496 );
and ( n10498 , n10477 , n10484 );
or ( n10499 , n10497 , n10498 );
xor ( n10500 , n10332 , n10499 );
and ( n10501 , n524 , n465 );
not ( n10502 , n524 );
not ( n10503 , n465 );
and ( n80304 , n10502 , n10503 );
nor ( n10505 , n10501 , n80304 );
not ( n10506 , n10505 );
not ( n10507 , n10142 );
or ( n10508 , n10506 , n10507 );
nand ( n10509 , n10357 , n10351 );
nand ( n10510 , n10508 , n10509 );
and ( n10511 , n533 , n457 );
or ( n10512 , n10510 , n10511 );
xor ( n10513 , n528 , n461 );
not ( n10514 , n10513 );
not ( n10515 , n10253 );
or ( n10516 , n10514 , n10515 );
nand ( n10517 , n10244 , n10341 );
nand ( n10518 , n10516 , n10517 );
nand ( n10519 , n10512 , n10518 );
nand ( n10520 , n10510 , n10511 );
nand ( n10521 , n10519 , n10520 );
and ( n10522 , n10500 , n10521 );
and ( n10523 , n10332 , n10499 );
or ( n10524 , n10522 , n10523 );
not ( n10525 , n10369 );
not ( n10526 , n10332 );
not ( n10527 , n10372 );
and ( n10528 , n10526 , n10527 );
and ( n10529 , n10332 , n10372 );
nor ( n10530 , n10528 , n10529 );
not ( n10531 , n10530 );
or ( n10532 , n10525 , n10531 );
or ( n80333 , n10369 , n10530 );
nand ( n10534 , n10532 , n80333 );
xor ( n10535 , n10524 , n10534 );
xor ( n10536 , n10291 , n10299 );
xor ( n10537 , n10536 , n10306 );
xor ( n10538 , n532 , n457 );
not ( n10539 , n10538 );
not ( n10540 , n10127 );
or ( n10541 , n10539 , n10540 );
nand ( n10542 , n10068 , n10295 );
nand ( n10543 , n10541 , n10542 );
not ( n10544 , n10543 );
not ( n10545 , n10085 );
xor ( n10546 , n530 , n459 );
not ( n10547 , n10546 );
or ( n10548 , n10545 , n10547 );
nand ( n10549 , n10094 , n10361 );
nand ( n10550 , n10548 , n10549 );
not ( n10551 , n10550 );
or ( n10552 , n10544 , n10551 );
or ( n10553 , n10550 , n10543 );
xor ( n10554 , n521 , n469 );
not ( n10555 , n10554 );
not ( n10556 , n470 );
nand ( n10557 , n10556 , n471 );
not ( n10558 , n471 );
nand ( n10559 , n10558 , n470 );
and ( n10560 , n10557 , n10559 , n10489 );
not ( n10561 , n10560 );
or ( n10562 , n10555 , n10561 );
buf ( n10563 , n10486 );
nand ( n10564 , n469 , n10563 );
nand ( n10565 , n10562 , n10564 );
nand ( n10566 , n10553 , n10565 );
nand ( n10567 , n10552 , n10566 );
xor ( n10568 , n10537 , n10567 );
xor ( n10569 , n10350 , n10359 );
xor ( n10570 , n10569 , n10366 );
and ( n10571 , n10568 , n10570 );
and ( n10572 , n10537 , n10567 );
or ( n10573 , n10571 , n10572 );
xnor ( n10574 , n10535 , n10573 );
not ( n10575 , n10574 );
not ( n10576 , n10575 );
not ( n10577 , n10317 );
not ( n10578 , n10577 );
not ( n10579 , n10578 );
xor ( n10580 , n10289 , n10309 );
not ( n10581 , n10580 );
not ( n10582 , n10581 );
or ( n10583 , n10579 , n10582 );
nand ( n10584 , n10580 , n10577 );
nand ( n10585 , n10583 , n10584 );
not ( n10586 , n10585 );
not ( n10587 , n10586 );
or ( n10588 , n10576 , n10587 );
not ( n10589 , n10585 );
not ( n10590 , n10574 );
or ( n80391 , n10589 , n10590 );
xor ( n10595 , n527 , n463 );
not ( n80393 , n10595 );
not ( n10597 , n10480 );
or ( n10598 , n80393 , n10597 );
nand ( n10599 , n10112 , n10478 );
nand ( n10600 , n10598 , n10599 );
not ( n10601 , n10600 );
not ( n10602 , n10469 );
and ( n10603 , n467 , n523 );
not ( n10604 , n467 );
not ( n10605 , n523 );
and ( n10606 , n10604 , n10605 );
nor ( n10607 , n10603 , n10606 );
nand ( n10608 , n10607 , n10160 );
and ( n10609 , n10602 , n10608 );
not ( n10610 , n10602 );
not ( n10611 , n10475 );
and ( n10612 , n10610 , n10611 );
nor ( n10613 , n10609 , n10612 );
nand ( n10614 , n534 , n457 );
not ( n80412 , n10614 );
nor ( n10619 , n10613 , n80412 );
not ( n10620 , n10619 );
not ( n10621 , n10620 );
or ( n10622 , n10601 , n10621 );
not ( n10623 , n10614 );
nand ( n10624 , n10623 , n10613 );
nand ( n10625 , n10622 , n10624 );
not ( n10626 , n10139 );
not ( n10627 , n10505 );
or ( n10628 , n10626 , n10627 );
xor ( n10629 , n525 , n465 );
nand ( n10630 , n10629 , n10141 );
or ( n10631 , n10630 , n10356 );
nand ( n10632 , n10628 , n10631 );
xor ( n10633 , n529 , n461 );
not ( n10634 , n10633 );
not ( n10635 , n10253 );
or ( n10636 , n10634 , n10635 );
nand ( n10637 , n80148 , n10513 );
nand ( n10638 , n10636 , n10637 );
xor ( n10639 , n10632 , n10638 );
xor ( n10640 , n531 , n459 );
not ( n10641 , n10640 );
not ( n10642 , n10085 );
or ( n10643 , n10641 , n10642 );
nand ( n10644 , n10093 , n10546 );
nand ( n10645 , n10643 , n10644 );
and ( n10646 , n10639 , n10645 );
and ( n10647 , n10632 , n10638 );
or ( n10648 , n10646 , n10647 );
xor ( n10649 , n10625 , n10648 );
xor ( n10650 , n10477 , n10484 );
xor ( n10651 , n10650 , n10496 );
and ( n10652 , n10649 , n10651 );
and ( n10653 , n10625 , n10648 );
or ( n10654 , n10652 , n10653 );
xor ( n10655 , n10332 , n10499 );
xor ( n10656 , n10655 , n10521 );
xor ( n10657 , n10654 , n10656 );
xor ( n10658 , n10537 , n10567 );
xor ( n10659 , n10658 , n10570 );
and ( n10660 , n10657 , n10659 );
and ( n10661 , n10654 , n10656 );
or ( n10662 , n10660 , n10661 );
nand ( n10663 , n80391 , n10662 );
nand ( n10664 , n10588 , n10663 );
not ( n10665 , n10664 );
xor ( n10666 , n10118 , n10148 );
xor ( n10667 , n10666 , n10200 );
not ( n10668 , n10378 );
not ( n10669 , n10374 );
or ( n10670 , n10668 , n10669 );
or ( n10671 , n10374 , n10378 );
nand ( n10672 , n10670 , n10671 );
xor ( n10673 , n10672 , n10319 );
xor ( n10674 , n10667 , n10673 );
buf ( n10675 , n10524 );
not ( n10676 , n10675 );
not ( n10677 , n10534 );
or ( n10678 , n10676 , n10677 );
or ( n10679 , n10534 , n10675 );
nand ( n10680 , n10679 , n10573 );
nand ( n10681 , n10678 , n10680 );
xor ( n10682 , n10674 , n10681 );
not ( n10683 , n10682 );
and ( n10684 , n10665 , n10683 );
xor ( n10685 , n10667 , n10673 );
and ( n10686 , n10685 , n10681 );
and ( n10687 , n10667 , n10673 );
or ( n10688 , n10686 , n10687 );
xor ( n10689 , n10203 , n80086 );
xor ( n10690 , n10689 , n10384 );
nor ( n10691 , n10688 , n10690 );
nor ( n10692 , n10684 , n10691 );
buf ( n10693 , n10692 );
not ( n10694 , n10693 );
nor ( n10695 , n10468 , n10694 );
not ( n10696 , n10695 );
xor ( n10697 , n524 , n467 );
not ( n10698 , n10697 );
not ( n10699 , n10160 );
nor ( n10700 , n10699 , n10469 );
not ( n10701 , n10700 );
or ( n10702 , n10698 , n10701 );
nand ( n10703 , n10473 , n10607 );
nand ( n80498 , n10702 , n10703 );
xor ( n80499 , n528 , n463 );
not ( n10706 , n80499 );
not ( n10707 , n10108 );
or ( n10708 , n10706 , n10707 );
nand ( n10709 , n10112 , n10595 );
nand ( n10710 , n10708 , n10709 );
xor ( n10711 , n80498 , n10710 );
xor ( n10712 , n522 , n469 );
not ( n10713 , n10712 );
buf ( n10714 , n10560 );
not ( n10715 , n10714 );
or ( n10716 , n10713 , n10715 );
nand ( n10717 , n10563 , n10554 );
nand ( n10718 , n10716 , n10717 );
xor ( n10719 , n10711 , n10718 );
not ( n10720 , n10719 );
and ( n10721 , n534 , n2714 );
not ( n10722 , n534 );
and ( n10723 , n10722 , n457 );
nor ( n10724 , n10721 , n10723 );
not ( n10725 , n10724 );
not ( n10726 , n10725 );
not ( n10727 , n10073 );
or ( n10728 , n10726 , n10727 );
xor ( n10729 , n533 , n457 );
nand ( n10730 , n10066 , n10729 );
nand ( n10731 , n10728 , n10730 );
nand ( n10732 , n535 , n457 );
not ( n10733 , n10732 );
not ( n10734 , n471 );
and ( n10735 , n10733 , n10734 );
not ( n10736 , n10733 );
not ( n10737 , n10558 );
and ( n10738 , n10736 , n10737 );
or ( n10739 , n10735 , n10738 );
and ( n10740 , n10731 , n10739 );
not ( n10741 , n10731 );
not ( n10742 , n471 );
and ( n10743 , n10732 , n10742 );
not ( n10744 , n10732 );
not ( n10745 , n10558 );
and ( n10746 , n10744 , n10745 );
or ( n10747 , n10743 , n10746 );
and ( n10748 , n10741 , n10747 );
or ( n10749 , n10740 , n10748 );
not ( n10750 , n10749 );
nand ( n10751 , n10720 , n10750 );
nand ( n10752 , n10719 , n10749 );
nand ( n10753 , n10751 , n10752 );
xor ( n10754 , n461 , n532 );
not ( n10755 , n10754 );
not ( n10756 , n10253 );
or ( n10757 , n10755 , n10756 );
and ( n10758 , n461 , n531 );
not ( n10759 , n461 );
not ( n10760 , n531 );
and ( n10761 , n10759 , n10760 );
nor ( n10762 , n10758 , n10761 );
nand ( n10763 , n10194 , n10762 );
nand ( n10764 , n10757 , n10763 );
not ( n10765 , n10764 );
not ( n10766 , n10473 );
xor ( n10767 , n525 , n467 );
not ( n10768 , n10767 );
or ( n10769 , n10766 , n10768 );
xor ( n10770 , n526 , n467 );
nand ( n10771 , n10157 , n10160 , n10770 );
nand ( n10772 , n10769 , n10771 );
xor ( n10773 , n529 , n463 );
not ( n10774 , n10773 );
not ( n10775 , n10105 );
not ( n10776 , n10775 );
or ( n10777 , n10774 , n10776 );
and ( n10778 , n530 , n463 );
not ( n10779 , n530 );
and ( n10780 , n10779 , n2374 );
nor ( n10781 , n10778 , n10780 );
and ( n10782 , n10106 , n10781 );
not ( n10783 , n10111 );
nand ( n80578 , n10782 , n10783 );
nand ( n10785 , n10777 , n80578 );
or ( n10786 , n10772 , n10785 );
not ( n10787 , n10786 );
or ( n10788 , n10765 , n10787 );
nand ( n10789 , n10772 , n10785 );
nand ( n10790 , n10788 , n10789 );
not ( n10791 , n10790 );
or ( n10792 , n536 , n458 );
nand ( n10793 , n10792 , n459 );
nand ( n10794 , n536 , n458 );
and ( n10795 , n10793 , n10794 , n457 );
and ( n10796 , n522 , n471 );
not ( n10797 , n522 );
not ( n10798 , n471 );
and ( n10799 , n10797 , n10798 );
nor ( n10800 , n10796 , n10799 );
not ( n10801 , n10800 );
not ( n10802 , n471 );
nor ( n10803 , n10802 , n472 );
not ( n10804 , n10803 );
or ( n10805 , n10801 , n10804 );
xor ( n10806 , n521 , n471 );
nand ( n10807 , n10806 , n472 );
nand ( n10808 , n10805 , n10807 );
and ( n10809 , n10795 , n10808 );
not ( n10810 , n10809 );
not ( n10811 , n10487 );
and ( n10812 , n523 , n469 );
not ( n10813 , n523 );
and ( n10814 , n10813 , n79958 );
nor ( n10815 , n10812 , n10814 );
nand ( n10816 , n10811 , n10815 );
and ( n10817 , n524 , n79958 );
not ( n10818 , n524 );
and ( n10819 , n10818 , n469 );
or ( n10820 , n10817 , n10819 );
nand ( n10821 , n10487 , n10489 , n10820 );
nor ( n10822 , n10292 , n10072 );
xor ( n10823 , n536 , n457 );
nand ( n10824 , n10822 , n10823 );
buf ( n10825 , n10066 );
not ( n10826 , n535 );
not ( n10827 , n10826 );
not ( n10828 , n457 );
or ( n10829 , n10827 , n10828 );
nand ( n10830 , n2714 , n535 );
nand ( n10831 , n10829 , n10830 );
nand ( n10832 , n10825 , n10831 );
nand ( n10833 , n10816 , n10821 , n10824 , n10832 );
xor ( n10834 , n528 , n465 );
and ( n10835 , n10141 , n10834 );
not ( n10836 , n10835 );
not ( n10837 , n10357 );
not ( n10838 , n10837 );
or ( n10839 , n10836 , n10838 );
xor ( n10840 , n527 , n465 );
nand ( n10841 , n10840 , n10357 );
nand ( n10842 , n10839 , n10841 );
nand ( n10843 , n10833 , n10842 );
nand ( n10844 , n10824 , n10832 );
nand ( n10845 , n10820 , n10489 );
not ( n10846 , n10845 );
not ( n10847 , n10563 );
and ( n10848 , n10846 , n10847 );
or ( n10849 , n10605 , n469 );
or ( n10850 , n79958 , n523 );
nand ( n10851 , n10849 , n10850 );
and ( n10852 , n10851 , n10486 );
nor ( n10853 , n10848 , n10852 );
not ( n10854 , n10853 );
nand ( n80649 , n10844 , n10854 );
nand ( n80650 , n10810 , n10843 , n80649 );
not ( n10857 , n80650 );
or ( n10858 , n10791 , n10857 );
nand ( n10859 , n10843 , n80649 );
nand ( n10860 , n10809 , n10859 );
nand ( n10861 , n10858 , n10860 );
xor ( n10862 , n10753 , n10861 );
xor ( n10863 , n534 , n459 );
not ( n10864 , n10863 );
not ( n10865 , n10087 );
or ( n10866 , n10864 , n10865 );
xor ( n10867 , n459 , n533 );
nand ( n10868 , n10094 , n10867 );
nand ( n10869 , n10866 , n10868 );
xor ( n10870 , n10795 , n10808 );
xor ( n10871 , n10869 , n10870 );
xor ( n10872 , n525 , n469 );
not ( n10873 , n10872 );
not ( n10874 , n10560 );
or ( n10875 , n10873 , n10874 );
nand ( n10876 , n10563 , n10820 );
nand ( n10877 , n10875 , n10876 );
not ( n10878 , n10877 );
and ( n10879 , n471 , n523 );
not ( n10880 , n471 );
and ( n10881 , n10880 , n10605 );
nor ( n10882 , n10879 , n10881 );
not ( n10883 , n10882 );
not ( n10884 , n471 );
nor ( n10885 , n10884 , n472 );
not ( n10886 , n10885 );
or ( n10887 , n10883 , n10886 );
nand ( n10888 , n10800 , n472 );
nand ( n10889 , n10887 , n10888 );
not ( n10890 , n10889 );
nand ( n10891 , n536 , n10066 );
nand ( n10892 , n10890 , n10891 );
not ( n10893 , n10892 );
or ( n10894 , n10878 , n10893 );
not ( n10895 , n10891 );
nand ( n10896 , n10895 , n10889 );
nand ( n10897 , n10894 , n10896 );
and ( n10898 , n10871 , n10897 );
and ( n10899 , n10869 , n10870 );
or ( n10900 , n10898 , n10899 );
xor ( n10901 , n10809 , n10859 );
xor ( n10902 , n10901 , n10790 );
xor ( n10903 , n10900 , n10902 );
not ( n10904 , n10785 );
xor ( n10905 , n10772 , n10904 );
xor ( n10906 , n10905 , n10764 );
not ( n10907 , n10906 );
not ( n10908 , n10907 );
not ( n10909 , n10842 );
not ( n10910 , n10844 );
and ( n10911 , n10910 , n10853 );
not ( n10912 , n10910 );
or ( n10913 , n10845 , n10811 );
nand ( n10914 , n10913 , n10816 );
and ( n10915 , n10912 , n10914 );
nor ( n10916 , n10911 , n10915 );
not ( n10917 , n10916 );
not ( n10918 , n10917 );
or ( n10919 , n10909 , n10918 );
not ( n10920 , n10842 );
nand ( n10921 , n10920 , n10916 );
nand ( n10922 , n10919 , n10921 );
not ( n10923 , n10922 );
or ( n10924 , n10908 , n10923 );
or ( n10925 , n10922 , n10907 );
xor ( n10926 , n531 , n463 );
not ( n10927 , n10926 );
not ( n10928 , n10480 );
or ( n80723 , n10927 , n10928 );
nand ( n10930 , n10112 , n10781 );
nand ( n10931 , n80723 , n10930 );
xor ( n10932 , n529 , n465 );
not ( n10933 , n10932 );
not ( n10934 , n10141 );
buf ( n10935 , n10356 );
nor ( n10936 , n10934 , n10935 );
not ( n10937 , n10936 );
or ( n10938 , n10933 , n10937 );
nand ( n80733 , n10935 , n10834 );
nand ( n10940 , n10938 , n80733 );
xor ( n10941 , n10931 , n10940 );
not ( n10942 , n10473 );
not ( n10943 , n10942 );
not ( n10944 , n10943 );
not ( n10945 , n10770 );
or ( n10946 , n10944 , n10945 );
xor ( n10947 , n467 , n527 );
nand ( n10948 , n10162 , n10947 );
nand ( n10949 , n10946 , n10948 );
and ( n10950 , n10941 , n10949 );
and ( n10951 , n10931 , n10940 );
or ( n10952 , n10950 , n10951 );
nand ( n10953 , n10925 , n10952 );
nand ( n10954 , n10924 , n10953 );
and ( n10955 , n10903 , n10954 );
and ( n10956 , n10900 , n10902 );
or ( n10957 , n10955 , n10956 );
not ( n10958 , n10957 );
xor ( n10959 , n10862 , n10958 );
xor ( n10960 , n461 , n530 );
not ( n10961 , n10960 );
not ( n10962 , n10253 );
or ( n10963 , n10961 , n10962 );
nand ( n10964 , n10244 , n10633 );
nand ( n10965 , n10963 , n10964 );
xor ( n10966 , n532 , n459 );
not ( n10967 , n10966 );
not ( n10968 , n10087 );
or ( n10969 , n10967 , n10968 );
nand ( n10970 , n10094 , n10640 );
nand ( n10971 , n10969 , n10970 );
xor ( n10972 , n10965 , n10971 );
and ( n10973 , n526 , n465 );
not ( n10974 , n526 );
and ( n10975 , n10974 , n10503 );
nor ( n10976 , n10973 , n10975 );
not ( n10977 , n10976 );
not ( n10978 , n10353 );
or ( n10979 , n10977 , n10978 );
nand ( n10980 , n10145 , n10629 );
nand ( n10981 , n10979 , n10980 );
not ( n10982 , n10981 );
xor ( n10983 , n10972 , n10982 );
not ( n10984 , n10815 );
not ( n10985 , n10714 );
or ( n10986 , n10984 , n10985 );
nand ( n10987 , n10563 , n10712 );
nand ( n10988 , n10986 , n10987 );
not ( n10989 , n10988 );
not ( n10990 , n10989 );
nand ( n10991 , n536 , n457 );
not ( n10992 , n10806 );
not ( n10993 , n10803 );
or ( n10994 , n10992 , n10993 );
nand ( n10995 , n471 , n472 );
nand ( n10996 , n10994 , n10995 );
and ( n10997 , n10991 , n10996 );
not ( n10998 , n10991 );
not ( n10999 , n10996 );
and ( n11000 , n10998 , n10999 );
nor ( n11001 , n10997 , n11000 );
not ( n11002 , n11001 );
and ( n11003 , n10990 , n11002 );
and ( n11004 , n10989 , n11001 );
nor ( n11005 , n11003 , n11004 );
not ( n11006 , n11005 );
not ( n11007 , n10067 );
not ( n11008 , n10724 );
and ( n11009 , n11007 , n11008 );
and ( n11010 , n10293 , n10831 );
nor ( n11011 , n11009 , n11010 );
not ( n11012 , n11011 );
not ( n11013 , n11012 );
nand ( n11014 , n10840 , n10141 );
not ( n11015 , n11014 );
not ( n11016 , n10139 );
and ( n11017 , n11015 , n11016 );
and ( n11018 , n10976 , n10356 );
nor ( n80813 , n11017 , n11018 );
not ( n11023 , n80813 );
not ( n80815 , n11023 );
or ( n11025 , n11013 , n80815 );
nand ( n11026 , n80813 , n11011 );
nand ( n11027 , n11025 , n11026 );
not ( n11028 , n10773 );
not ( n11029 , n10480 );
or ( n11030 , n11028 , n11029 );
nand ( n11031 , n10112 , n80499 );
nand ( n11032 , n11030 , n11031 );
buf ( n11033 , n11032 );
not ( n11034 , n11033 );
and ( n11035 , n11027 , n11034 );
not ( n11036 , n11027 );
and ( n11037 , n11036 , n11033 );
nor ( n11038 , n11035 , n11037 );
not ( n11039 , n11038 );
or ( n11040 , n11006 , n11039 );
not ( n11041 , n11038 );
not ( n11042 , n11041 );
not ( n11043 , n11005 );
not ( n11044 , n11043 );
or ( n11045 , n11042 , n11044 );
and ( n11046 , n460 , n461 );
not ( n11047 , n460 );
not ( n80839 , n461 );
and ( n11052 , n11047 , n80839 );
nor ( n11053 , n11046 , n11052 );
not ( n11054 , n11053 );
and ( n11055 , n459 , n460 );
not ( n11056 , n459 );
and ( n11057 , n11056 , n10082 );
nor ( n11058 , n11055 , n11057 );
nand ( n11059 , n11054 , n10867 , n11058 );
nand ( n11060 , n3088 , n460 );
not ( n11061 , n11060 );
nand ( n11062 , n10082 , n461 );
not ( n11063 , n11062 );
or ( n11064 , n11061 , n11063 );
nand ( n11065 , n11064 , n10966 );
nand ( n11066 , n11059 , n11065 );
not ( n11067 , n10700 );
not ( n11068 , n10767 );
or ( n11069 , n11067 , n11068 );
nand ( n11070 , n10473 , n10697 );
nand ( n11071 , n11069 , n11070 );
xor ( n11072 , n11066 , n11071 );
not ( n11073 , n10960 );
not ( n11074 , n80148 );
or ( n11075 , n11073 , n11074 );
nand ( n11076 , n10346 , n10340 , n10762 );
nand ( n11077 , n11075 , n11076 );
xor ( n11078 , n11072 , n11077 );
nand ( n11079 , n11045 , n11078 );
nand ( n11080 , n11040 , n11079 );
xor ( n11081 , n10983 , n11080 );
not ( n11082 , n11032 );
not ( n11083 , n11026 );
or ( n11084 , n11082 , n11083 );
nand ( n11085 , n11023 , n11012 );
nand ( n11086 , n11084 , n11085 );
not ( n11087 , n11086 );
not ( n11088 , n11087 );
xor ( n11089 , n11066 , n11071 );
and ( n11090 , n11089 , n11077 );
and ( n11091 , n11066 , n11071 );
or ( n11092 , n11090 , n11091 );
not ( n11093 , n11092 );
not ( n11094 , n11093 );
or ( n11095 , n11088 , n11094 );
nand ( n11096 , n11092 , n11086 );
nand ( n11097 , n11095 , n11096 );
not ( n11098 , n10991 );
not ( n11099 , n10999 );
or ( n11100 , n11098 , n11099 );
nand ( n11101 , n11100 , n10988 );
not ( n11102 , n10991 );
nand ( n11103 , n11102 , n10996 );
nand ( n11104 , n11101 , n11103 );
not ( n11105 , n11104 );
and ( n11106 , n11097 , n11105 );
not ( n11107 , n11097 );
and ( n11108 , n11107 , n11104 );
nor ( n11109 , n11106 , n11108 );
xnor ( n11110 , n11081 , n11109 );
xor ( n11111 , n10959 , n11110 );
xor ( n11112 , n11078 , n11043 );
xor ( n11113 , n11112 , n11041 );
xor ( n11114 , n461 , n533 );
not ( n11115 , n11114 );
nor ( n11116 , n10339 , n10345 );
not ( n11117 , n11116 );
or ( n11118 , n11115 , n11117 );
not ( n11119 , n10242 );
not ( n11120 , n10243 );
or ( n11121 , n11119 , n11120 );
nand ( n11122 , n11121 , n10754 );
nand ( n11123 , n11118 , n11122 );
not ( n11124 , n10863 );
not ( n11125 , n10093 );
or ( n11126 , n11124 , n11125 );
and ( n11127 , n459 , n535 );
not ( n11128 , n459 );
and ( n11129 , n11128 , n10826 );
nor ( n11130 , n11127 , n11129 );
nand ( n11131 , n10085 , n11130 );
nand ( n11132 , n11126 , n11131 );
or ( n11133 , n11123 , n11132 );
xor ( n11134 , n523 , n471 );
nand ( n11135 , n11134 , n472 );
not ( n11136 , n11135 );
nand ( n11137 , n10558 , n524 );
not ( n11138 , n11137 );
not ( n11139 , n524 );
nand ( n11140 , n11139 , n471 );
not ( n11141 , n11140 );
or ( n11142 , n11138 , n11141 );
nor ( n11143 , n10558 , n472 );
nand ( n11144 , n11142 , n11143 );
not ( n11145 , n11144 );
or ( n11146 , n11136 , n11145 );
and ( n11147 , n536 , n460 );
nor ( n11148 , n11147 , n2348 );
or ( n11149 , n536 , n460 );
nand ( n11150 , n11149 , n461 );
nand ( n11151 , n11148 , n11150 );
not ( n11152 , n11151 );
nand ( n11153 , n11146 , n11152 );
not ( n11154 , n11153 );
nand ( n11155 , n11133 , n11154 );
nand ( n11156 , n11123 , n11132 );
nand ( n11157 , n11155 , n11156 );
not ( n11158 , n11157 );
xor ( n11159 , n10869 , n10870 );
xor ( n11160 , n11159 , n10897 );
buf ( n80949 , n11160 );
not ( n80950 , n80949 );
or ( n11163 , n11158 , n80950 );
or ( n11164 , n11160 , n11157 );
nor ( n11165 , n10157 , n10947 );
not ( n11166 , n11165 );
xor ( n11167 , n467 , n528 );
not ( n11168 , n11167 );
not ( n11169 , n10160 );
or ( n11170 , n11168 , n11169 );
nand ( n11171 , n11170 , n10157 );
nand ( n11172 , n11166 , n11171 );
not ( n11173 , n80148 );
not ( n11174 , n11114 );
or ( n11175 , n11173 , n11174 );
not ( n11176 , n10250 );
xor ( n11177 , n461 , n534 );
nand ( n11178 , n11176 , n10183 , n11177 );
nand ( n11179 , n11175 , n11178 );
not ( n11180 , n11179 );
nand ( n11181 , n11172 , n11180 );
not ( n11182 , n11181 );
xor ( n11183 , n536 , n459 );
not ( n11184 , n11183 );
not ( n11185 , n10087 );
or ( n11186 , n11184 , n11185 );
nand ( n11187 , n10094 , n11130 );
nand ( n11188 , n11186 , n11187 );
not ( n11189 , n11188 );
or ( n11190 , n11182 , n11189 );
not ( n11191 , n11172 );
nand ( n11192 , n11191 , n11179 );
nand ( n11193 , n11190 , n11192 );
not ( n11194 , n11193 );
not ( n11195 , n11194 );
not ( n11196 , n10889 );
not ( n11197 , n10891 );
and ( n11198 , n11196 , n11197 );
and ( n11199 , n10889 , n10891 );
nor ( n11200 , n11198 , n11199 );
not ( n11201 , n11200 );
not ( n11202 , n11201 );
not ( n11203 , n10877 );
or ( n11204 , n11202 , n11203 );
not ( n11205 , n10877 );
nand ( n11206 , n11205 , n11200 );
nand ( n11207 , n11204 , n11206 );
not ( n11208 , n11207 );
or ( n11209 , n11195 , n11208 );
xor ( n11210 , n530 , n465 );
not ( n11211 , n11210 );
not ( n81000 , n10353 );
or ( n11213 , n11211 , n81000 );
nand ( n11214 , n10357 , n10932 );
nand ( n11215 , n11213 , n11214 );
and ( n11216 , n532 , n463 );
not ( n11217 , n532 );
and ( n11218 , n11217 , n2374 );
nor ( n11219 , n11216 , n11218 );
not ( n11220 , n11219 );
not ( n11221 , n10108 );
or ( n11222 , n11220 , n11221 );
nand ( n11223 , n10112 , n10926 );
nand ( n11224 , n11222 , n11223 );
xor ( n11225 , n11215 , n11224 );
xor ( n11226 , n526 , n469 );
not ( n11227 , n11226 );
not ( n11228 , n10714 );
or ( n11229 , n11227 , n11228 );
nand ( n11230 , n10811 , n10872 );
nand ( n11231 , n11229 , n11230 );
and ( n11232 , n11225 , n11231 );
and ( n11233 , n11215 , n11224 );
or ( n11234 , n11232 , n11233 );
nand ( n11235 , n11209 , n11234 );
not ( n11236 , n11207 );
nand ( n11237 , n11236 , n11193 );
nand ( n11238 , n11235 , n11237 );
nand ( n11239 , n11164 , n11238 );
nand ( n11240 , n11163 , n11239 );
xor ( n11241 , n11113 , n11240 );
xor ( n11242 , n10900 , n10902 );
xor ( n11243 , n11242 , n10954 );
and ( n11244 , n11241 , n11243 );
and ( n11245 , n11113 , n11240 );
or ( n11246 , n11244 , n11245 );
not ( n11247 , n11246 );
nand ( n11248 , n11111 , n11247 );
xor ( n11249 , n11193 , n11207 );
xor ( n11250 , n11249 , n11234 );
not ( n11251 , n11250 );
not ( n11252 , n11251 );
xor ( n11253 , n529 , n467 );
not ( n11254 , n11253 );
not ( n11255 , n10163 );
or ( n11256 , n11254 , n11255 );
nand ( n11257 , n10943 , n11167 );
nand ( n11258 , n11256 , n11257 );
not ( n11259 , n11258 );
nand ( n11260 , n536 , n462 );
or ( n11261 , n536 , n462 );
nand ( n11262 , n11261 , n463 );
nand ( n11263 , n11260 , n461 , n11262 );
not ( n11264 , n11263 );
xor ( n11265 , n528 , n469 );
not ( n11266 , n11265 );
not ( n11267 , n10714 );
or ( n11268 , n11266 , n11267 );
xor ( n11269 , n527 , n469 );
nand ( n11270 , n10563 , n11269 );
nand ( n11271 , n11268 , n11270 );
nand ( n11272 , n11264 , n11271 );
nand ( n11273 , n11259 , n11272 );
not ( n11274 , n11273 );
not ( n11275 , n10803 );
xor ( n11276 , n471 , n526 );
not ( n11277 , n11276 );
or ( n11278 , n11275 , n11277 );
and ( n11279 , n471 , n525 );
not ( n11280 , n471 );
not ( n11281 , n525 );
and ( n11282 , n11280 , n11281 );
nor ( n11283 , n11279 , n11282 );
nand ( n11284 , n11283 , n472 );
nand ( n11285 , n11278 , n11284 );
xor ( n11286 , n532 , n465 );
not ( n11287 , n11286 );
not ( n11288 , n10142 );
or ( n11289 , n11287 , n11288 );
and ( n11290 , n465 , n531 );
not ( n11291 , n465 );
and ( n11292 , n11291 , n10760 );
nor ( n81081 , n11290 , n11292 );
nand ( n81082 , n10145 , n81081 );
nand ( n11295 , n11289 , n81082 );
xor ( n11296 , n11285 , n11295 );
xor ( n11297 , n534 , n463 );
not ( n11298 , n11297 );
not ( n11299 , n10108 );
or ( n11300 , n11298 , n11299 );
xor ( n11301 , n533 , n463 );
nand ( n11302 , n10112 , n11301 );
nand ( n11303 , n11300 , n11302 );
and ( n11304 , n11296 , n11303 );
and ( n11305 , n11285 , n11295 );
or ( n11306 , n11304 , n11305 );
not ( n11307 , n11306 );
or ( n11308 , n11274 , n11307 );
not ( n11309 , n11272 );
nand ( n11310 , n11309 , n11258 );
nand ( n11311 , n11308 , n11310 );
not ( n11312 , n11311 );
xor ( n11313 , n11215 , n11224 );
xor ( n11314 , n11313 , n11231 );
not ( n11315 , n11314 );
xor ( n11316 , n11179 , n11172 );
xor ( n11317 , n11316 , n11188 );
nand ( n11318 , n11315 , n11317 );
not ( n11319 , n11318 );
or ( n11320 , n11312 , n11319 );
not ( n11321 , n11317 );
nand ( n11322 , n11321 , n11314 );
nand ( n11323 , n11320 , n11322 );
not ( n11324 , n11323 );
nand ( n11325 , n11252 , n11324 );
not ( n11326 , n11325 );
xor ( n11327 , n11153 , n11123 );
xnor ( n11328 , n11327 , n11132 );
xor ( n11329 , n10931 , n10940 );
xor ( n11330 , n11329 , n10949 );
xor ( n11331 , n11328 , n11330 );
buf ( n11332 , n11151 );
not ( n11333 , n11332 );
nand ( n11334 , n11144 , n11135 );
not ( n11335 , n11334 );
or ( n11336 , n11333 , n11335 );
or ( n11337 , n11334 , n11332 );
nand ( n11338 , n11336 , n11337 );
not ( n11339 , n11283 );
not ( n11340 , n10885 );
or ( n11341 , n11339 , n11340 );
not ( n11342 , n11137 );
not ( n11343 , n11140 );
or ( n11344 , n11342 , n11343 );
nand ( n11345 , n11344 , n472 );
nand ( n11346 , n11341 , n11345 );
not ( n11347 , n11346 );
nand ( n11348 , n11301 , n10783 , n10106 );
nand ( n11349 , n11219 , n10775 );
nand ( n11350 , n11348 , n11349 );
not ( n11351 , n11350 );
or ( n11352 , n11347 , n11351 );
not ( n11353 , n11346 );
nand ( n11354 , n11348 , n11349 , n11353 );
xor ( n11355 , n535 , n461 );
not ( n11356 , n11355 );
not ( n11357 , n10253 );
or ( n81146 , n11356 , n11357 );
nand ( n11359 , n80148 , n11177 );
nand ( n11360 , n81146 , n11359 );
nand ( n11361 , n11354 , n11360 );
nand ( n11362 , n11352 , n11361 );
xor ( n11363 , n11338 , n11362 );
not ( n11364 , n11210 );
not ( n11365 , n10935 );
or ( n11366 , n11364 , n11365 );
not ( n11367 , n10356 );
nand ( n11368 , n10141 , n11367 , n81081 );
nand ( n11369 , n11366 , n11368 );
not ( n11370 , n11369 );
nand ( n11371 , n11053 , n536 );
not ( n11372 , n11371 );
not ( n11373 , n11372 );
or ( n11374 , n11370 , n11373 );
or ( n11375 , n11369 , n11372 );
not ( n11376 , n11269 );
not ( n11377 , n10714 );
or ( n11378 , n11376 , n11377 );
nand ( n11379 , n10563 , n11226 );
nand ( n11380 , n11378 , n11379 );
nand ( n11381 , n11375 , n11380 );
nand ( n11382 , n11374 , n11381 );
and ( n11383 , n11363 , n11382 );
and ( n11384 , n11338 , n11362 );
or ( n11385 , n11383 , n11384 );
xor ( n11386 , n11331 , n11385 );
not ( n11387 , n11386 );
or ( n11388 , n11326 , n11387 );
nand ( n11389 , n11323 , n11251 );
nand ( n11390 , n11388 , n11389 );
xor ( n11391 , n11328 , n11330 );
and ( n11392 , n11391 , n11385 );
and ( n11393 , n11328 , n11330 );
or ( n11394 , n11392 , n11393 );
and ( n11395 , n10952 , n10906 );
not ( n11396 , n10952 );
and ( n81185 , n11396 , n10907 );
nor ( n11398 , n11395 , n81185 );
not ( n11399 , n10922 );
and ( n11400 , n11398 , n11399 );
not ( n11401 , n11398 );
and ( n11402 , n11401 , n10922 );
nor ( n11403 , n11400 , n11402 );
xor ( n11404 , n11394 , n11403 );
not ( n11405 , n11160 );
xor ( n11406 , n11157 , n11405 );
xnor ( n11407 , n11406 , n11238 );
xor ( n11408 , n11404 , n11407 );
nor ( n11409 , n11390 , n11408 );
not ( n11410 , n11409 );
xor ( n11411 , n11113 , n11240 );
xor ( n11412 , n11411 , n11243 );
not ( n11413 , n11412 );
xor ( n11414 , n11394 , n11403 );
and ( n11415 , n11414 , n11407 );
and ( n11416 , n11394 , n11403 );
or ( n11417 , n11415 , n11416 );
not ( n11418 , n11417 );
nand ( n11419 , n11413 , n11418 );
and ( n11420 , n11248 , n11410 , n11419 );
not ( n11421 , n11420 );
xor ( n11422 , n532 , n467 );
not ( n11423 , n11422 );
not ( n11424 , n10162 );
or ( n11425 , n11423 , n11424 );
xor ( n11426 , n531 , n467 );
nand ( n11427 , n10943 , n11426 );
nand ( n11428 , n11425 , n11427 );
not ( n11429 , n11428 );
not ( n11430 , n11429 );
xor ( n11431 , n530 , n469 );
not ( n11432 , n11431 );
not ( n11433 , n10492 );
or ( n11434 , n11432 , n11433 );
xor ( n11435 , n529 , n469 );
nand ( n11436 , n10563 , n11435 );
nand ( n11437 , n11434 , n11436 );
or ( n11438 , n536 , n464 );
nand ( n11439 , n11438 , n465 );
nand ( n11440 , n536 , n464 );
and ( n11441 , n11439 , n11440 , n463 );
nor ( n11442 , n11437 , n11441 );
not ( n11443 , n11442 );
nand ( n11444 , n11441 , n11437 );
nand ( n11445 , n11443 , n11444 );
not ( n81234 , n11445 );
or ( n11450 , n11430 , n81234 );
and ( n81236 , n10111 , n536 );
not ( n11452 , n472 );
xor ( n11453 , n471 , n528 );
not ( n11454 , n11453 );
or ( n11455 , n11452 , n11454 );
and ( n11456 , n471 , n529 );
not ( n11457 , n471 );
not ( n11458 , n529 );
and ( n11459 , n11457 , n11458 );
nor ( n11460 , n11456 , n11459 );
not ( n11461 , n471 );
nor ( n11462 , n11461 , n472 );
nand ( n11463 , n11460 , n11462 );
nand ( n11464 , n11455 , n11463 );
xor ( n11465 , n81236 , n11464 );
xor ( n11466 , n535 , n465 );
not ( n11467 , n11466 );
not ( n11468 , n10353 );
or ( n11469 , n11467 , n11468 );
xor ( n11470 , n534 , n465 );
nand ( n81256 , n11470 , n10145 );
nand ( n11475 , n11469 , n81256 );
and ( n11476 , n11465 , n11475 );
and ( n11477 , n81236 , n11464 );
or ( n11478 , n11476 , n11477 );
nand ( n11479 , n11450 , n11478 );
not ( n11480 , n11445 );
nand ( n11481 , n11480 , n11428 );
nand ( n11482 , n11479 , n11481 );
not ( n11483 , n11482 );
xor ( n11484 , n471 , n527 );
not ( n11485 , n11484 );
not ( n11486 , n10803 );
or ( n11487 , n11485 , n11486 );
nand ( n11488 , n11276 , n472 );
nand ( n11489 , n11487 , n11488 );
xor ( n11490 , n535 , n463 );
not ( n11491 , n11490 );
not ( n11492 , n10108 );
or ( n11493 , n11491 , n11492 );
nand ( n11494 , n10112 , n11297 );
nand ( n11495 , n11493 , n11494 );
xor ( n11496 , n11489 , n11495 );
not ( n11497 , n11426 );
not ( n11498 , n10162 );
or ( n11499 , n11497 , n11498 );
xor ( n11500 , n467 , n530 );
nand ( n11501 , n10473 , n11500 );
nand ( n11502 , n11499 , n11501 );
buf ( n11503 , n11502 );
xor ( n11504 , n11496 , n11503 );
not ( n11505 , n11504 );
or ( n11506 , n11483 , n11505 );
not ( n11507 , n11482 );
not ( n11508 , n11504 );
nand ( n11509 , n11507 , n11508 );
nand ( n11510 , n11506 , n11509 );
not ( n11511 , n11510 );
not ( n11512 , n11453 );
not ( n11513 , n11462 );
or ( n11514 , n11512 , n11513 );
nand ( n11515 , n11484 , n472 );
nand ( n11516 , n11514 , n11515 );
not ( n11517 , n11516 );
not ( n11518 , n11470 );
not ( n11519 , n10353 );
or ( n11520 , n11518 , n11519 );
xor ( n11521 , n533 , n465 );
nand ( n11522 , n10357 , n11521 );
nand ( n11523 , n11520 , n11522 );
not ( n11524 , n11523 );
or ( n11525 , n11517 , n11524 );
or ( n11526 , n11523 , n11516 );
xor ( n11527 , n536 , n463 );
not ( n11528 , n11527 );
not ( n11529 , n10108 );
or ( n11530 , n11528 , n11529 );
nand ( n11531 , n10112 , n11490 );
nand ( n11532 , n11530 , n11531 );
nand ( n11533 , n11526 , n11532 );
nand ( n11534 , n11525 , n11533 );
xor ( n11535 , n11444 , n11534 );
and ( n11536 , n80148 , n536 );
not ( n11537 , n11521 );
not ( n11538 , n10936 );
or ( n11539 , n11537 , n11538 );
nand ( n11540 , n10935 , n11286 );
nand ( n11541 , n11539 , n11540 );
not ( n11542 , n11541 );
xor ( n11543 , n11536 , n11542 );
not ( n11544 , n10714 );
not ( n11545 , n11435 );
or ( n11546 , n11544 , n11545 );
nand ( n11547 , n10563 , n11265 );
nand ( n11548 , n11546 , n11547 );
xnor ( n11549 , n11543 , n11548 );
xnor ( n11550 , n11535 , n11549 );
not ( n11551 , n11550 );
not ( n11552 , n11551 );
or ( n11553 , n11511 , n11552 );
or ( n11554 , n11510 , n11551 );
nand ( n11555 , n11553 , n11554 );
not ( n11556 , n11555 );
buf ( n11557 , n11445 );
xor ( n11558 , n11429 , n11557 );
xnor ( n11559 , n11558 , n11478 );
or ( n11560 , n536 , n466 );
nand ( n11561 , n11560 , n467 );
nand ( n11562 , n536 , n466 );
and ( n11563 , n11561 , n11562 , n465 );
nor ( n11564 , n530 , n472 );
nand ( n11565 , n11564 , n471 );
not ( n11566 , n471 );
nand ( n81349 , n11566 , n472 , n529 );
nand ( n81350 , n11458 , n471 , n472 );
nand ( n11569 , n11565 , n81349 , n81350 );
nand ( n11570 , n11563 , n11569 );
xor ( n11571 , n531 , n469 );
not ( n11572 , n11571 );
not ( n11573 , n10492 );
or ( n11574 , n11572 , n11573 );
nand ( n11575 , n11431 , n10563 );
nand ( n11576 , n11574 , n11575 );
not ( n11577 , n11576 );
xor ( n11578 , n11570 , n11577 );
xor ( n11579 , n533 , n467 );
not ( n11580 , n11579 );
not ( n11581 , n10162 );
or ( n11582 , n11580 , n11581 );
nand ( n11583 , n10329 , n11422 );
nand ( n11584 , n11582 , n11583 );
not ( n11585 , n11584 );
and ( n11586 , n11578 , n11585 );
and ( n11587 , n11570 , n11577 );
or ( n11588 , n11586 , n11587 );
xor ( n11589 , n11516 , n11532 );
xnor ( n11590 , n11589 , n11523 );
and ( n11591 , n11588 , n11590 );
or ( n11592 , n11559 , n11591 );
or ( n11593 , n11590 , n11588 );
nand ( n11594 , n11592 , n11593 );
nand ( n11595 , n11556 , n11594 );
not ( n11596 , n11595 );
xor ( n11597 , n81236 , n11464 );
xor ( n11598 , n11597 , n11475 );
not ( n11599 , n11598 );
xor ( n11600 , n11570 , n11577 );
xor ( n11601 , n11600 , n11585 );
or ( n11602 , n11599 , n11601 );
not ( n11603 , n11601 );
not ( n11604 , n11599 );
or ( n11605 , n11603 , n11604 );
xor ( n11606 , n536 , n465 );
not ( n11607 , n11606 );
not ( n11608 , n10142 );
or ( n11609 , n11607 , n11608 );
nand ( n11610 , n10145 , n11466 );
nand ( n11611 , n11609 , n11610 );
xor ( n11612 , n534 , n467 );
not ( n11613 , n11612 );
not ( n11614 , n10163 );
or ( n11615 , n11613 , n11614 );
nand ( n11616 , n10943 , n11579 );
nand ( n11617 , n11615 , n11616 );
xor ( n11618 , n11611 , n11617 );
xor ( n11619 , n532 , n469 );
not ( n11620 , n11619 );
not ( n11621 , n10714 );
or ( n11622 , n11620 , n11621 );
nand ( n11623 , n10563 , n11571 );
nand ( n11624 , n11622 , n11623 );
and ( n11625 , n11618 , n11624 );
and ( n11626 , n11611 , n11617 );
or ( n11627 , n11625 , n11626 );
nand ( n11628 , n11605 , n11627 );
nand ( n11629 , n11602 , n11628 );
not ( n11630 , n11629 );
xor ( n11631 , n11428 , n11478 );
xnor ( n81414 , n11631 , n11557 );
xor ( n11633 , n11588 , n11590 );
xnor ( n11634 , n81414 , n11633 );
nand ( n11635 , n11630 , n11634 );
not ( n11636 , n11599 );
not ( n11637 , n11601 );
not ( n11638 , n11637 );
or ( n11639 , n11636 , n11638 );
nand ( n11640 , n11601 , n11598 );
nand ( n11641 , n11639 , n11640 );
not ( n11642 , n11641 );
not ( n11643 , n11627 );
nand ( n11644 , n11642 , n11643 );
not ( n11645 , n11643 );
nand ( n11646 , n11645 , n11641 );
nand ( n11647 , n10357 , n536 );
not ( n11648 , n11647 );
not ( n11649 , n11648 );
xor ( n11650 , n531 , n471 );
not ( n11651 , n11650 );
not ( n11652 , n10803 );
or ( n11653 , n11651 , n11652 );
xor ( n11654 , n471 , n530 );
nand ( n11655 , n11654 , n472 );
nand ( n11656 , n11653 , n11655 );
not ( n11657 , n11656 );
or ( n11658 , n11649 , n11657 );
not ( n11659 , n11647 );
not ( n11660 , n11656 );
not ( n11661 , n11660 );
or ( n11662 , n11659 , n11661 );
xor ( n11663 , n533 , n469 );
not ( n11664 , n11663 );
not ( n11665 , n10714 );
or ( n11666 , n11664 , n11665 );
nand ( n11667 , n10563 , n11619 );
nand ( n11668 , n11666 , n11667 );
nand ( n11669 , n11662 , n11668 );
nand ( n11670 , n11658 , n11669 );
not ( n11671 , n11670 );
not ( n11672 , n11569 );
not ( n11673 , n11672 );
not ( n11674 , n11563 );
not ( n11675 , n11674 );
or ( n11676 , n11673 , n11675 );
nand ( n11677 , n11676 , n11570 );
nand ( n11678 , n11671 , n11677 );
not ( n11679 , n11678 );
xor ( n11680 , n11611 , n11617 );
xor ( n11681 , n11680 , n11624 );
not ( n11682 , n11681 );
or ( n11683 , n11679 , n11682 );
not ( n11684 , n11677 );
nand ( n11685 , n11684 , n11670 );
nand ( n11686 , n11683 , n11685 );
and ( n11687 , n11644 , n11646 , n11686 );
nand ( n11688 , n11635 , n11687 );
not ( n11689 , n11634 );
nand ( n11690 , n11689 , n11629 );
and ( n11691 , n11688 , n11690 );
xor ( n11692 , n536 , n467 );
nand ( n11693 , n10160 , n11692 );
not ( n11694 , n11693 );
not ( n11695 , n10329 );
and ( n11696 , n11694 , n11695 );
xor ( n11697 , n535 , n467 );
and ( n11698 , n10943 , n11697 );
nor ( n11699 , n11696 , n11698 );
not ( n81482 , n11699 );
xor ( n81483 , n534 , n469 );
not ( n11702 , n81483 );
not ( n11703 , n10714 );
or ( n11704 , n11702 , n11703 );
nand ( n11705 , n10563 , n11663 );
nand ( n11706 , n11704 , n11705 );
and ( n11707 , n81482 , n11706 );
not ( n11708 , n81482 );
not ( n11709 , n11706 );
and ( n11710 , n11708 , n11709 );
nor ( n11711 , n11707 , n11710 );
or ( n11712 , n536 , n468 );
nand ( n11713 , n11712 , n469 );
nand ( n11714 , n536 , n468 );
nand ( n11715 , n11713 , n11714 , n467 );
xor ( n11716 , n471 , n532 );
not ( n11717 , n11716 );
not ( n11718 , n11462 );
or ( n11719 , n11717 , n11718 );
nand ( n11720 , n11650 , n472 );
nand ( n11721 , n11719 , n11720 );
xor ( n11722 , n11715 , n11721 );
and ( n11723 , n11711 , n11722 );
not ( n11724 , n11711 );
not ( n11725 , n11722 );
and ( n11726 , n11724 , n11725 );
nor ( n11727 , n11723 , n11726 );
xor ( n11728 , n535 , n469 );
not ( n11729 , n11728 );
not ( n11730 , n10714 );
or ( n11731 , n11729 , n11730 );
nand ( n11732 , n10563 , n81483 );
nand ( n11733 , n11731 , n11732 );
not ( n11734 , n11733 );
xor ( n11735 , n471 , n533 );
not ( n11736 , n11735 );
not ( n11737 , n10803 );
or ( n11738 , n11736 , n11737 );
nand ( n11739 , n11716 , n472 );
nand ( n11740 , n11738 , n11739 );
not ( n11741 , n11740 );
not ( n11742 , n536 );
not ( n11743 , n11742 );
nand ( n11744 , n11743 , n10329 );
nand ( n11745 , n11741 , n11744 );
not ( n11746 , n11745 );
or ( n11747 , n11734 , n11746 );
not ( n11748 , n11744 );
nand ( n11749 , n11748 , n11740 );
nand ( n11750 , n11747 , n11749 );
not ( n11751 , n11750 );
nand ( n11752 , n11727 , n11751 );
not ( n11753 , n11752 );
not ( n11754 , n11462 );
xor ( n11755 , n534 , n471 );
not ( n11756 , n11755 );
or ( n11757 , n11754 , n11756 );
nand ( n11758 , n11735 , n472 );
nand ( n11759 , n11757 , n11758 );
not ( n11760 , n11759 );
or ( n11761 , n536 , n470 );
nand ( n11762 , n11761 , n471 );
nand ( n11763 , n536 , n470 );
nand ( n11764 , n11762 , n11763 , n469 );
not ( n11765 , n11764 );
and ( n11766 , n11760 , n11765 );
and ( n11767 , n11759 , n11764 );
nor ( n81550 , n11766 , n11767 );
xor ( n11769 , n536 , n469 );
not ( n11770 , n11769 );
not ( n11771 , n10714 );
or ( n11772 , n11770 , n11771 );
nand ( n11773 , n10563 , n11728 );
nand ( n11774 , n11772 , n11773 );
not ( n11775 , n11774 );
nand ( n11776 , n81550 , n11775 );
not ( n11777 , n11776 );
not ( n11778 , n11742 );
not ( n11779 , n11462 );
or ( n11780 , n11778 , n11779 );
xor ( n11781 , n471 , n535 );
nand ( n11782 , n11781 , n472 );
nand ( n81565 , n11780 , n11782 );
and ( n11784 , n536 , n472 );
nor ( n11785 , n11784 , n10558 );
nand ( n11786 , n81565 , n11785 );
nand ( n11787 , n10563 , n536 );
not ( n11788 , n11787 );
not ( n11789 , n11781 );
not ( n11790 , n10803 );
or ( n11791 , n11789 , n11790 );
nand ( n11792 , n11755 , n472 );
nand ( n11793 , n11791 , n11792 );
nor ( n11794 , n11788 , n11793 );
or ( n11795 , n11786 , n11794 );
not ( n11796 , n11787 );
nand ( n11797 , n11796 , n11793 );
nand ( n11798 , n11795 , n11797 );
not ( n11799 , n11798 );
or ( n11800 , n11777 , n11799 );
not ( n11801 , n81550 );
nand ( n11802 , n11801 , n11774 );
nand ( n11803 , n11800 , n11802 );
not ( n11804 , n11803 );
not ( n11805 , n11740 );
not ( n11806 , n11744 );
and ( n11807 , n11805 , n11806 );
and ( n11808 , n11740 , n11744 );
nor ( n11809 , n11807 , n11808 );
not ( n11810 , n11809 );
not ( n11811 , n11733 );
and ( n11812 , n11810 , n11811 );
and ( n11813 , n11733 , n11809 );
nor ( n11814 , n11812 , n11813 );
not ( n11815 , n11764 );
nand ( n11816 , n11815 , n11759 );
nand ( n11817 , n11814 , n11816 );
not ( n11818 , n11817 );
or ( n11819 , n11804 , n11818 );
not ( n11820 , n11814 );
not ( n11821 , n11816 );
nand ( n11822 , n11820 , n11821 );
nand ( n11823 , n11819 , n11822 );
not ( n11824 , n11823 );
or ( n11825 , n11753 , n11824 );
not ( n11826 , n11727 );
nand ( n11827 , n11826 , n11750 );
nand ( n11828 , n11825 , n11827 );
not ( n11829 , n11722 );
not ( n11830 , n11699 );
or ( n11831 , n11829 , n11830 );
nand ( n11832 , n11831 , n11706 );
nand ( n11833 , n11725 , n81482 );
nand ( n11834 , n11832 , n11833 );
not ( n11835 , n11834 );
not ( n11836 , n11656 );
not ( n11837 , n11647 );
or ( n11838 , n11836 , n11837 );
or ( n11839 , n11656 , n11647 );
nand ( n11840 , n11838 , n11839 );
xor ( n11841 , n11840 , n11668 );
not ( n11842 , n11841 );
not ( n11843 , n11721 );
nor ( n11844 , n11843 , n11715 );
not ( n11845 , n11844 );
not ( n11846 , n11697 );
not ( n11847 , n10162 );
or ( n11848 , n11846 , n11847 );
nand ( n11849 , n10943 , n11612 );
nand ( n11850 , n11848 , n11849 );
not ( n11851 , n11850 );
not ( n11852 , n11851 );
and ( n11853 , n11845 , n11852 );
and ( n11854 , n11844 , n11851 );
nor ( n11855 , n11853 , n11854 );
not ( n81638 , n11855 );
and ( n11860 , n11842 , n81638 );
and ( n81640 , n11841 , n11855 );
nor ( n11862 , n11860 , n81640 );
nand ( n11863 , n11835 , n11862 );
nand ( n11864 , n11828 , n11863 );
xor ( n11865 , n11677 , n11670 );
xnor ( n11866 , n11865 , n11681 );
or ( n11867 , n11844 , n11850 );
nand ( n11868 , n11867 , n11841 );
nand ( n11869 , n11844 , n11850 );
nand ( n11870 , n11868 , n11869 );
nand ( n11871 , n11866 , n11870 );
not ( n11872 , n11862 );
nand ( n11873 , n11872 , n11834 );
nand ( n11874 , n11864 , n11871 , n11873 );
nand ( n11875 , n11642 , n11643 );
and ( n11876 , n11875 , n11646 );
nor ( n11877 , n11876 , n11686 );
nor ( n11878 , n11866 , n11870 );
nor ( n11879 , n11877 , n11878 );
nand ( n11880 , n11635 , n11874 , n11879 );
nand ( n11881 , n11691 , n11880 );
not ( n11882 , n11594 );
nand ( n11883 , n11882 , n11555 );
nand ( n11884 , n11881 , n11883 );
not ( n81664 , n11884 );
or ( n11889 , n11596 , n81664 );
not ( n11890 , n11272 );
not ( n11891 , n11258 );
and ( n11892 , n11890 , n11891 );
and ( n11893 , n11272 , n11258 );
nor ( n11894 , n11892 , n11893 );
not ( n11895 , n11894 );
not ( n11896 , n11306 );
and ( n11897 , n11895 , n11896 );
and ( n11898 , n11306 , n11894 );
nor ( n11899 , n11897 , n11898 );
not ( n11900 , n11899 );
xor ( n11901 , n11346 , n11360 );
xor ( n11902 , n11901 , n11350 );
not ( n11903 , n11902 );
xor ( n11904 , n11372 , n11369 );
xnor ( n11905 , n11904 , n11380 );
nand ( n11906 , n11903 , n11905 );
not ( n11907 , n11906 );
not ( n11908 , n11253 );
not ( n11909 , n10943 );
or ( n11910 , n11908 , n11909 );
nand ( n11911 , n11500 , n10160 , n10602 );
nand ( n11912 , n11910 , n11911 );
buf ( n11913 , n11912 );
not ( n11914 , n11913 );
not ( n11915 , n10190 );
xnor ( n11916 , n536 , n461 );
not ( n11917 , n11916 );
and ( n11918 , n11915 , n11917 );
and ( n11919 , n10194 , n11355 );
nor ( n11920 , n11918 , n11919 );
nand ( n11921 , n11914 , n11920 );
not ( n11922 , n11263 );
not ( n11923 , n11922 );
not ( n11924 , n11271 );
not ( n11925 , n11924 );
or ( n11926 , n11923 , n11925 );
nand ( n11927 , n11271 , n11263 );
nand ( n11928 , n11926 , n11927 );
and ( n11929 , n11921 , n11928 );
not ( n11930 , n11920 );
and ( n11931 , n11930 , n11913 );
nor ( n11932 , n11929 , n11931 );
not ( n11933 , n11902 );
nor ( n11934 , n11933 , n11905 );
nor ( n11935 , n11932 , n11934 );
not ( n11936 , n11935 );
or ( n11937 , n11907 , n11936 );
not ( n11938 , n11905 );
nor ( n11939 , n11938 , n11902 );
or ( n11940 , n11939 , n11934 );
nand ( n11941 , n11940 , n11932 );
nand ( n11942 , n11937 , n11941 );
not ( n11943 , n11942 );
or ( n11944 , n11900 , n11943 );
not ( n11945 , n11489 );
not ( n11946 , n11495 );
or ( n11947 , n11945 , n11946 );
or ( n11948 , n11489 , n11495 );
nand ( n11949 , n11948 , n11502 );
nand ( n11950 , n11947 , n11949 );
not ( n11951 , n11950 );
xor ( n11952 , n11285 , n11295 );
xor ( n11953 , n11952 , n11303 );
not ( n11954 , n11953 );
or ( n11955 , n11951 , n11954 );
or ( n11956 , n11950 , n11953 );
not ( n11957 , n11536 );
not ( n11958 , n11541 );
or ( n11959 , n11957 , n11958 );
not ( n11960 , n11542 );
not ( n11961 , n11536 );
not ( n11962 , n11961 );
or ( n11963 , n11960 , n11962 );
nand ( n11964 , n11963 , n11548 );
nand ( n11965 , n11959 , n11964 );
nand ( n11966 , n11956 , n11965 );
nand ( n11967 , n11955 , n11966 );
nand ( n11968 , n11944 , n11967 );
not ( n11969 , n11899 );
not ( n11970 , n11942 );
nand ( n11971 , n11969 , n11970 );
nand ( n11972 , n11968 , n11971 );
not ( n11973 , n11972 );
xor ( n11974 , n11338 , n11362 );
xor ( n11975 , n11974 , n11382 );
not ( n11976 , n11975 );
not ( n11977 , n11902 );
not ( n11978 , n11938 );
or ( n11979 , n11977 , n11978 );
not ( n11980 , n11933 );
not ( n11981 , n11905 );
or ( n11982 , n11980 , n11981 );
not ( n11983 , n11932 );
nand ( n11984 , n11982 , n11983 );
nand ( n11985 , n11979 , n11984 );
xor ( n11986 , n11976 , n11985 );
and ( n81763 , n11314 , n11317 );
not ( n81764 , n11314 );
and ( n11989 , n81764 , n11321 );
nor ( n11990 , n81763 , n11989 );
and ( n11991 , n11990 , n11311 );
not ( n11992 , n11990 );
not ( n11993 , n11311 );
and ( n11994 , n11992 , n11993 );
nor ( n11995 , n11991 , n11994 );
xnor ( n11996 , n11986 , n11995 );
nand ( n11997 , n11973 , n11996 );
or ( n11998 , n11899 , n11967 );
nand ( n11999 , n11967 , n11899 );
nand ( n12000 , n11998 , n11999 );
xnor ( n12001 , n12000 , n11970 );
not ( n12002 , n11549 );
not ( n12003 , n11444 );
not ( n12004 , n12003 );
or ( n12005 , n12002 , n12004 );
or ( n12006 , n11549 , n12003 );
nand ( n12007 , n12006 , n11534 );
nand ( n12008 , n12005 , n12007 );
not ( n12009 , n12008 );
not ( n12010 , n12009 );
not ( n12011 , n11953 );
xor ( n12012 , n11950 , n11965 );
xor ( n12013 , n12011 , n12012 );
not ( n12014 , n12013 );
or ( n12015 , n12010 , n12014 );
xor ( n12016 , n11913 , n11930 );
xnor ( n12017 , n12016 , n11928 );
not ( n12018 , n12017 );
nand ( n12019 , n12015 , n12018 );
not ( n12020 , n12013 );
nand ( n12021 , n12020 , n12008 );
nand ( n12022 , n12019 , n12021 );
not ( n12023 , n12022 );
nand ( n12024 , n12001 , n12023 );
nor ( n12025 , n12008 , n12018 );
and ( n12026 , n12025 , n12013 );
nor ( n12027 , n12008 , n12017 );
not ( n12028 , n12013 );
and ( n12029 , n12027 , n12028 );
nor ( n12030 , n12026 , n12029 );
not ( n12031 , n12030 );
and ( n12032 , n12017 , n12013 );
not ( n12033 , n12017 );
and ( n12034 , n12033 , n12028 );
nor ( n12035 , n12032 , n12034 );
not ( n12036 , n12009 );
nand ( n12037 , n12035 , n12036 );
not ( n12038 , n12037 );
or ( n12039 , n12031 , n12038 );
not ( n12040 , n11550 );
nand ( n12041 , n11507 , n11508 );
not ( n81818 , n12041 );
or ( n12043 , n12040 , n81818 );
not ( n12044 , n11507 );
nand ( n12045 , n12044 , n11504 );
nand ( n12046 , n12043 , n12045 );
not ( n12047 , n12046 );
nand ( n12048 , n12039 , n12047 );
nand ( n12049 , n11997 , n12024 , n12048 );
not ( n12050 , n11995 );
not ( n12051 , n12050 );
not ( n12052 , n11976 );
not ( n12053 , n12052 );
or ( n12054 , n12051 , n12053 );
not ( n12055 , n11976 );
not ( n12056 , n11995 );
or ( n12057 , n12055 , n12056 );
buf ( n12058 , n11985 );
nand ( n12059 , n12057 , n12058 );
nand ( n12060 , n12054 , n12059 );
not ( n12061 , n12060 );
and ( n12062 , n11386 , n11251 );
not ( n12063 , n11386 );
and ( n12064 , n12063 , n11250 );
nor ( n12065 , n12062 , n12064 );
and ( n12066 , n12065 , n11324 );
not ( n12067 , n12065 );
and ( n12068 , n12067 , n11323 );
nor ( n12069 , n12066 , n12068 );
nand ( n12070 , n12061 , n12069 );
not ( n12071 , n12070 );
nor ( n12072 , n12049 , n12071 );
nand ( n12073 , n11889 , n12072 );
buf ( n12074 , n11997 );
nand ( n12075 , n12037 , n12030 );
nor ( n12076 , n12075 , n12047 );
not ( n12077 , n12076 );
not ( n12078 , n12024 );
or ( n12079 , n12077 , n12078 );
not ( n12080 , n12001 );
nand ( n12081 , n12080 , n12022 );
nand ( n12082 , n12079 , n12081 );
not ( n12083 , n12071 );
nand ( n12084 , n12074 , n12082 , n12083 );
not ( n12085 , n12070 );
nor ( n12086 , n11973 , n11996 );
not ( n12087 , n12086 );
or ( n12088 , n12085 , n12087 );
not ( n12089 , n12069 );
nand ( n12090 , n12089 , n12060 );
nand ( n12091 , n12088 , n12090 );
not ( n12092 , n12091 );
nand ( n12093 , n12073 , n12084 , n12092 );
not ( n12094 , n12093 );
or ( n12095 , n11421 , n12094 );
not ( n12096 , n11418 );
not ( n12097 , n11413 );
or ( n12098 , n12096 , n12097 );
nand ( n12099 , n11412 , n11417 );
nand ( n12100 , n11408 , n11390 );
nand ( n12101 , n12099 , n12100 );
nand ( n12102 , n12098 , n12101 );
not ( n12103 , n11248 );
or ( n12104 , n12102 , n12103 );
not ( n12105 , n11111 );
nand ( n12106 , n12105 , n11246 );
nand ( n12107 , n12104 , n12106 );
not ( n12108 , n12107 );
nand ( n12109 , n12095 , n12108 );
not ( n12110 , n12109 );
xor ( n12111 , n10625 , n10648 );
xor ( n12112 , n12111 , n10651 );
or ( n12113 , n10558 , n10733 );
nand ( n81890 , n12113 , n10731 );
nand ( n81891 , n10558 , n10733 );
nand ( n12116 , n81890 , n81891 );
xor ( n12117 , n10632 , n10638 );
xor ( n12118 , n12117 , n10645 );
xor ( n12119 , n12116 , n12118 );
xor ( n12120 , n80498 , n10710 );
and ( n12121 , n12120 , n10718 );
and ( n12122 , n80498 , n10710 );
or ( n12123 , n12121 , n12122 );
and ( n12124 , n12119 , n12123 );
and ( n12125 , n12116 , n12118 );
or ( n12126 , n12124 , n12125 );
xor ( n12127 , n12112 , n12126 );
or ( n12128 , n11092 , n11086 );
nand ( n12129 , n12128 , n11104 );
nand ( n12130 , n11092 , n11086 );
nand ( n12131 , n12129 , n12130 );
not ( n12132 , n12131 );
not ( n12133 , n10729 );
not ( n12134 , n10126 );
or ( n12135 , n12133 , n12134 );
nand ( n12136 , n10066 , n10538 );
nand ( n12137 , n12135 , n12136 );
not ( n12138 , n12137 );
not ( n12139 , n12138 );
not ( n12140 , n10565 );
not ( n12141 , n12140 );
or ( n12142 , n12139 , n12141 );
nand ( n12143 , n10565 , n12137 );
nand ( n12144 , n12142 , n12143 );
and ( n12145 , n12144 , n10982 );
not ( n12146 , n12144 );
and ( n12147 , n12146 , n10981 );
nor ( n12148 , n12145 , n12147 );
not ( n12149 , n10600 );
not ( n12150 , n10619 );
nand ( n12151 , n12150 , n10624 );
not ( n12152 , n12151 );
not ( n12153 , n12152 );
or ( n12154 , n12149 , n12153 );
not ( n12155 , n10600 );
nand ( n12156 , n12155 , n12151 );
nand ( n12157 , n12154 , n12156 );
nand ( n12158 , n12148 , n12157 );
not ( n12159 , n12158 );
or ( n12160 , n12132 , n12159 );
not ( n12161 , n12157 );
not ( n12162 , n12148 );
nand ( n12163 , n12161 , n12162 );
nand ( n12164 , n12160 , n12163 );
xor ( n12165 , n12127 , n12164 );
not ( n12166 , n12165 );
not ( n12167 , n10518 );
not ( n12168 , n10510 );
not ( n12169 , n10511 );
and ( n12170 , n12168 , n12169 );
and ( n12171 , n10510 , n10511 );
nor ( n12172 , n12170 , n12171 );
xor ( n12173 , n12167 , n12172 );
not ( n12174 , n12173 );
xor ( n12175 , n12140 , n10550 );
xnor ( n12176 , n12175 , n10543 );
not ( n12177 , n12176 );
xor ( n12178 , n12174 , n12177 );
not ( n12179 , n12138 );
not ( n12180 , n10982 );
or ( n81957 , n12179 , n12180 );
nand ( n12182 , n81957 , n12140 );
nand ( n12183 , n10981 , n12137 );
nand ( n12184 , n12182 , n12183 );
xor ( n12185 , n12178 , n12184 );
not ( n12186 , n12185 );
or ( n12187 , n12166 , n12186 );
not ( n12188 , n12165 );
not ( n12189 , n12176 );
not ( n12190 , n12184 );
not ( n12191 , n12173 );
or ( n12192 , n12190 , n12191 );
or ( n12193 , n12184 , n12173 );
nand ( n12194 , n12192 , n12193 );
not ( n12195 , n12194 );
not ( n12196 , n12195 );
or ( n12197 , n12189 , n12196 );
not ( n12198 , n12176 );
nand ( n12199 , n12198 , n12194 );
nand ( n12200 , n12197 , n12199 );
nand ( n12201 , n12188 , n12200 );
nand ( n12202 , n12187 , n12201 );
xor ( n12203 , n10965 , n10971 );
and ( n12204 , n12203 , n10982 );
and ( n12205 , n10965 , n10971 );
or ( n12206 , n12204 , n12205 );
not ( n12207 , n12206 );
xor ( n12208 , n12116 , n12118 );
xor ( n12209 , n12208 , n12123 );
not ( n12210 , n12209 );
or ( n12211 , n12207 , n12210 );
or ( n12212 , n12206 , n12209 );
not ( n12213 , n10751 );
not ( n12214 , n10861 );
or ( n12215 , n12213 , n12214 );
nand ( n81992 , n12215 , n10752 );
nand ( n12217 , n12212 , n81992 );
nand ( n12218 , n12211 , n12217 );
not ( n12219 , n12218 );
and ( n12220 , n12202 , n12219 );
not ( n12221 , n12202 );
and ( n12222 , n12221 , n12218 );
nor ( n12223 , n12220 , n12222 );
buf ( n12224 , n12131 );
and ( n12225 , n12162 , n12157 );
not ( n12226 , n12162 );
and ( n12227 , n12226 , n12161 );
nor ( n12228 , n12225 , n12227 );
xor ( n12229 , n12224 , n12228 );
not ( n12230 , n12229 );
xor ( n12231 , n12206 , n12209 );
xnor ( n12232 , n12231 , n81992 );
not ( n12233 , n12232 );
or ( n12234 , n12230 , n12233 );
not ( n12235 , n10983 );
not ( n12236 , n11109 );
or ( n12237 , n12235 , n12236 );
or ( n12238 , n11109 , n10983 );
nand ( n12239 , n12238 , n11080 );
nand ( n12240 , n12237 , n12239 );
nand ( n12241 , n12234 , n12240 );
not ( n12242 , n12232 );
not ( n12243 , n12229 );
nand ( n12244 , n12242 , n12243 );
nand ( n12245 , n12241 , n12244 );
not ( n12246 , n12245 );
nand ( n12247 , n12223 , n12246 );
and ( n12248 , n12240 , n12229 );
not ( n12249 , n12240 );
and ( n12250 , n12249 , n12243 );
nor ( n12251 , n12248 , n12250 );
and ( n12252 , n12251 , n12242 );
not ( n12253 , n12251 );
not ( n12254 , n12242 );
and ( n12255 , n12253 , n12254 );
nor ( n12256 , n12252 , n12255 );
xor ( n12257 , n10862 , n10958 );
and ( n12258 , n12257 , n11110 );
and ( n12259 , n10862 , n10958 );
or ( n12260 , n12258 , n12259 );
nand ( n12261 , n12256 , n12260 );
and ( n12262 , n12247 , n12261 );
not ( n12263 , n12262 );
not ( n12264 , n12173 );
not ( n12265 , n12177 );
or ( n12266 , n12264 , n12265 );
nand ( n12267 , n12266 , n12184 );
nand ( n12268 , n12176 , n12174 );
nand ( n82045 , n12267 , n12268 );
not ( n12273 , n82045 );
not ( n82047 , n12273 );
xor ( n12275 , n10654 , n10656 );
xor ( n12276 , n12275 , n10659 );
nand ( n12277 , n82047 , n12276 );
or ( n12278 , n12276 , n82045 );
xor ( n12279 , n12112 , n12126 );
and ( n12280 , n12279 , n12164 );
and ( n12281 , n12112 , n12126 );
or ( n12282 , n12280 , n12281 );
nand ( n12283 , n12278 , n12282 );
nand ( n12284 , n12277 , n12283 );
not ( n12285 , n12284 );
not ( n12286 , n12285 );
xor ( n12287 , n10585 , n10662 );
xor ( n12288 , n12287 , n10575 );
not ( n12289 , n12288 );
or ( n12290 , n12286 , n12289 );
not ( n12291 , n12282 );
not ( n12292 , n12273 );
not ( n12293 , n12276 );
or ( n82067 , n12292 , n12293 );
or ( n12298 , n12276 , n12273 );
nand ( n12299 , n82067 , n12298 );
xor ( n12300 , n12291 , n12299 );
not ( n12301 , n12200 );
not ( n12302 , n12188 );
not ( n12303 , n12302 );
or ( n12304 , n12301 , n12303 );
not ( n12305 , n12185 );
not ( n12306 , n12188 );
or ( n12307 , n12305 , n12306 );
nand ( n12308 , n12307 , n12218 );
nand ( n12309 , n12304 , n12308 );
not ( n12310 , n12309 );
nand ( n12311 , n12300 , n12310 );
nand ( n12312 , n12290 , n12311 );
nor ( n12313 , n12263 , n12312 );
not ( n12314 , n12313 );
or ( n12315 , n12110 , n12314 );
not ( n12316 , n12312 );
not ( n12317 , n12316 );
nor ( n12318 , n12256 , n12260 );
not ( n12319 , n12318 );
not ( n12320 , n12247 );
or ( n12321 , n12319 , n12320 );
not ( n12322 , n12223 );
nand ( n12323 , n12322 , n12245 );
nand ( n12324 , n12321 , n12323 );
not ( n12325 , n12324 );
not ( n12326 , n12325 );
not ( n12327 , n12326 );
or ( n12328 , n12317 , n12327 );
not ( n12329 , n12288 );
nand ( n12330 , n12329 , n12284 );
not ( n12331 , n12309 );
nor ( n12332 , n12331 , n12300 );
nand ( n12333 , n12285 , n12288 );
nand ( n12334 , n12332 , n12333 );
nand ( n12335 , n12330 , n12334 );
not ( n12336 , n12335 );
nand ( n12337 , n12328 , n12336 );
not ( n12338 , n12337 );
nand ( n12339 , n12315 , n12338 );
not ( n12340 , n12339 );
or ( n12341 , n10696 , n12340 );
not ( n12342 , n10467 );
nand ( n12343 , n10682 , n10664 );
or ( n12344 , n10691 , n12343 );
nand ( n12345 , n10688 , n10690 );
nand ( n12346 , n12344 , n12345 );
not ( n12347 , n12346 );
or ( n12348 , n12342 , n12347 );
not ( n12349 , n10387 );
nor ( n12350 , n12349 , n10466 );
not ( n12351 , n12350 );
nand ( n12352 , n12348 , n12351 );
not ( n12353 , n12352 );
nand ( n12354 , n12341 , n12353 );
not ( n12355 , n12354 );
not ( n12356 , n10428 );
nand ( n12357 , n12356 , n80235 );
not ( n12358 , n12357 );
not ( n12359 , n10451 );
or ( n12360 , n12358 , n12359 );
not ( n12361 , n80235 );
nand ( n12362 , n12361 , n10428 );
nand ( n12363 , n12360 , n12362 );
not ( n12364 , n12363 );
xor ( n12365 , n10408 , n10414 );
and ( n12366 , n12365 , n10420 );
and ( n12367 , n10408 , n10414 );
or ( n12368 , n12366 , n12367 );
and ( n12369 , n457 , n527 );
not ( n12370 , n80235 );
xor ( n12371 , n12369 , n12370 );
not ( n12372 , n10426 );
not ( n12373 , n10087 );
or ( n12374 , n12372 , n12373 );
xor ( n12375 , n523 , n459 );
nand ( n12376 , n10094 , n12375 );
nand ( n12377 , n12374 , n12376 );
xnor ( n12378 , n12371 , n12377 );
xor ( n12379 , n12368 , n12378 );
not ( n12380 , n10412 );
not ( n12381 , n10127 );
or ( n12382 , n12380 , n12381 );
xor ( n12383 , n457 , n525 );
nand ( n12384 , n10068 , n12383 );
nand ( n12385 , n12382 , n12384 );
not ( n12386 , n10433 );
not ( n12387 , n10191 );
or ( n12388 , n12386 , n12387 );
xor ( n12389 , n461 , n521 );
nand ( n82160 , n10194 , n12389 );
nand ( n82161 , n12388 , n82160 );
xor ( n12392 , n12385 , n82161 );
or ( n12393 , n10480 , n10112 );
nand ( n12394 , n12393 , n463 );
xor ( n12395 , n12392 , n12394 );
xor ( n12396 , n12379 , n12395 );
xor ( n12397 , n12364 , n12396 );
xor ( n12398 , n10407 , n10421 );
and ( n12399 , n12398 , n10455 );
and ( n12400 , n10407 , n10421 );
or ( n12401 , n12399 , n12400 );
xor ( n12402 , n12397 , n12401 );
not ( n12403 , n12402 );
nand ( n12404 , n10459 , n10402 );
not ( n12405 , n12404 );
not ( n12406 , n10395 );
or ( n12407 , n12405 , n12406 );
nand ( n12408 , n10456 , n10401 );
nand ( n12409 , n12407 , n12408 );
nand ( n12410 , n12403 , n12409 );
not ( n12411 , n12409 );
nand ( n12412 , n12411 , n12402 );
nand ( n12413 , n12410 , n12412 );
not ( n12414 , n12413 );
and ( n12415 , n12355 , n12414 );
and ( n12416 , n12354 , n12413 );
nor ( n12417 , n12415 , n12416 );
not ( n12418 , n12417 );
not ( n12419 , n12418 );
not ( n12420 , n12419 );
or ( n12421 , n10063 , n12420 );
not ( n12422 , n12419 );
not ( n12423 , n503 );
nand ( n12424 , n12422 , n12423 );
nand ( n12425 , n12421 , n12424 );
not ( n12426 , n12425 );
or ( n12427 , n10062 , n12426 );
not ( n12428 , n503 );
nor ( n12429 , n10694 , n12312 );
not ( n12430 , n12429 );
not ( n12431 , n12107 );
not ( n12432 , n12262 );
or ( n12433 , n12431 , n12432 );
nand ( n12434 , n12433 , n12325 );
not ( n12435 , n12434 );
not ( n12436 , n12103 );
and ( n12437 , n11410 , n11419 );
and ( n12438 , n12436 , n12437 , n12247 , n12261 );
nand ( n12439 , n12438 , n12093 );
nand ( n12440 , n12435 , n12439 );
not ( n12441 , n12440 );
or ( n12442 , n12430 , n12441 );
and ( n12443 , n10693 , n12335 );
nor ( n12444 , n12443 , n12346 );
nand ( n82215 , n12442 , n12444 );
not ( n12446 , n12350 );
nand ( n12447 , n12446 , n10467 );
not ( n12448 , n12447 );
and ( n12449 , n82215 , n12448 );
not ( n12450 , n82215 );
and ( n12451 , n12450 , n12447 );
nor ( n12452 , n12449 , n12451 );
not ( n12453 , n12452 );
not ( n12454 , n12453 );
or ( n12455 , n12428 , n12454 );
not ( n12456 , n12453 );
buf ( n12457 , n12423 );
nand ( n12458 , n12456 , n12457 );
nand ( n12459 , n12455 , n12458 );
not ( n12460 , n504 );
nand ( n12461 , n12460 , n503 );
not ( n12462 , n12461 );
nand ( n12463 , n12459 , n12462 );
nand ( n12464 , n12427 , n12463 );
and ( n12465 , n498 , n499 );
not ( n12466 , n498 );
not ( n12467 , n499 );
and ( n12468 , n12466 , n12467 );
or ( n12469 , n12465 , n12468 );
not ( n12470 , n12469 );
not ( n12471 , n12470 );
not ( n12472 , n497 );
or ( n12473 , n12260 , n12256 );
nand ( n12474 , n12261 , n12473 );
not ( n12475 , n12474 );
not ( n12476 , n12109 );
or ( n12477 , n12475 , n12476 );
not ( n12478 , n12109 );
not ( n12479 , n12474 );
nand ( n12480 , n12478 , n12479 );
nand ( n12481 , n12477 , n12480 );
not ( n12482 , n12481 );
buf ( n12483 , n12482 );
not ( n12484 , n12483 );
or ( n12485 , n12472 , n12484 );
not ( n12486 , n497 );
nand ( n12487 , n12481 , n12486 );
nand ( n12488 , n12485 , n12487 );
not ( n12489 , n12488 );
or ( n12490 , n12471 , n12489 );
not ( n12491 , n497 );
nand ( n12492 , n12436 , n12106 );
not ( n12493 , n12492 );
not ( n12494 , n12493 );
not ( n12495 , n12437 );
nand ( n12496 , n12092 , n12073 , n12084 );
not ( n12497 , n12496 );
or ( n12498 , n12495 , n12497 );
buf ( n12499 , n12102 );
nand ( n12500 , n12498 , n12499 );
not ( n12501 , n12500 );
not ( n12502 , n12501 );
or ( n12503 , n12494 , n12502 );
nand ( n12504 , n12500 , n12492 );
nand ( n12505 , n12503 , n12504 );
not ( n12506 , n12505 );
not ( n12507 , n12506 );
or ( n12508 , n12491 , n12507 );
buf ( n12509 , n12505 );
nand ( n12510 , n12509 , n12486 );
nand ( n12511 , n12508 , n12510 );
and ( n12512 , n498 , n497 );
not ( n12513 , n498 );
and ( n12514 , n12513 , n12486 );
nor ( n12515 , n12512 , n12514 );
and ( n12516 , n12469 , n12515 );
buf ( n12517 , n12516 );
nand ( n12518 , n12511 , n12517 );
nand ( n12519 , n12490 , n12518 );
not ( n12520 , n489 );
buf ( n12521 , n11877 );
not ( n12522 , n12521 );
buf ( n12523 , n11687 );
not ( n12524 , n12523 );
nand ( n82295 , n12522 , n12524 );
or ( n82296 , n11866 , n11870 );
not ( n12527 , n82296 );
not ( n12528 , n12527 );
buf ( n12529 , n11874 );
nand ( n12530 , n12528 , n12529 );
xor ( n12531 , n82295 , n12530 );
not ( n12532 , n12531 );
nor ( n12533 , n12520 , n12532 );
not ( n12534 , n12533 );
and ( n12535 , n490 , n491 );
not ( n12536 , n490 );
and ( n12537 , n12536 , n1693 );
nor ( n12538 , n12535 , n12537 );
not ( n12539 , n12538 );
xor ( n12540 , n489 , n490 );
nand ( n12541 , n12539 , n12540 );
not ( n12542 , n12541 );
not ( n12543 , n12542 );
not ( n12544 , n489 );
nand ( n12545 , n11690 , n11635 );
not ( n12546 , n12545 );
nor ( n12547 , n12521 , n12527 );
and ( n12548 , n12529 , n12547 );
nor ( n12549 , n12548 , n12523 );
not ( n12550 , n12549 );
not ( n12551 , n12550 );
or ( n12552 , n12546 , n12551 );
not ( n12553 , n12545 );
nand ( n12554 , n12553 , n12549 );
nand ( n12555 , n12552 , n12554 );
not ( n12556 , n12555 );
not ( n12557 , n12556 );
or ( n12558 , n12544 , n12557 );
buf ( n12559 , n12555 );
not ( n12560 , n489 );
nand ( n12561 , n12559 , n12560 );
nand ( n12562 , n12558 , n12561 );
not ( n12563 , n12562 );
or ( n12564 , n12543 , n12563 );
not ( n12565 , n11881 );
not ( n12566 , n12565 );
nand ( n12567 , n11595 , n11883 );
not ( n12568 , n12567 );
not ( n12569 , n12568 );
or ( n12570 , n12566 , n12569 );
nand ( n12571 , n12567 , n11881 );
nand ( n82342 , n12570 , n12571 );
buf ( n12573 , n82342 );
not ( n12574 , n12573 );
not ( n12575 , n12560 );
or ( n12576 , n12574 , n12575 );
not ( n12577 , n82342 );
nand ( n12578 , n12577 , n489 );
nand ( n12579 , n12576 , n12578 );
buf ( n12580 , n12538 );
nand ( n12581 , n12579 , n12580 );
nand ( n12582 , n12564 , n12581 );
not ( n12583 , n12582 );
or ( n12584 , n12534 , n12583 );
or ( n12585 , n12582 , n12533 );
nand ( n12586 , n12584 , n12585 );
and ( n12587 , n491 , n492 );
nor ( n12588 , n491 , n492 );
nor ( n12589 , n12587 , n12588 );
and ( n12590 , n492 , n493 );
not ( n12591 , n492 );
and ( n12592 , n12591 , n1976 );
or ( n12593 , n12590 , n12592 );
nand ( n12594 , n12589 , n12593 );
not ( n12595 , n12594 );
not ( n12596 , n12595 );
not ( n12597 , n491 );
not ( n12598 , n11883 );
not ( n12599 , n11881 );
or ( n12600 , n12598 , n12599 );
nand ( n12601 , n12600 , n11595 );
not ( n12602 , n12076 );
nand ( n12603 , n12047 , n12075 );
nand ( n12604 , n12602 , n12603 );
xnor ( n12605 , n12601 , n12604 );
buf ( n12606 , n12605 );
not ( n12607 , n12606 );
not ( n12608 , n12607 );
or ( n12609 , n12597 , n12608 );
not ( n12610 , n491 );
nand ( n82381 , n12606 , n12610 );
nand ( n12612 , n12609 , n82381 );
not ( n12613 , n12612 );
or ( n12614 , n12596 , n12613 );
not ( n12615 , n491 );
and ( n12616 , n12024 , n12081 );
not ( n12617 , n12616 );
not ( n12618 , n12603 );
nand ( n12619 , n11884 , n11595 );
not ( n12620 , n12619 );
or ( n12621 , n12618 , n12620 );
nand ( n12622 , n12621 , n12602 );
not ( n12623 , n12622 );
not ( n12624 , n12623 );
or ( n12625 , n12617 , n12624 );
not ( n12626 , n12616 );
nand ( n12627 , n12626 , n12622 );
nand ( n12628 , n12625 , n12627 );
not ( n12629 , n12628 );
not ( n12630 , n12629 );
or ( n12631 , n12615 , n12630 );
and ( n12632 , n12616 , n12623 );
not ( n12633 , n12616 );
and ( n12634 , n12633 , n12622 );
or ( n12635 , n12632 , n12634 );
nand ( n12636 , n12610 , n12635 );
nand ( n12637 , n12631 , n12636 );
not ( n12638 , n12593 );
nand ( n12639 , n12637 , n12638 );
nand ( n12640 , n12614 , n12639 );
and ( n12641 , n12586 , n12640 );
not ( n12642 , n12586 );
not ( n12643 , n12640 );
and ( n12644 , n12642 , n12643 );
or ( n12645 , n12641 , n12644 );
xor ( n12646 , n12519 , n12645 );
xor ( n12647 , n500 , n501 );
buf ( n12648 , n12647 );
not ( n12649 , n12648 );
not ( n12650 , n12649 );
not ( n12651 , n12650 );
not ( n12652 , n499 );
not ( n12653 , n12332 );
nand ( n12654 , n12300 , n12310 );
nand ( n12655 , n12653 , n12654 );
not ( n12656 , n12655 );
not ( n12657 , n12656 );
not ( n12658 , n12093 );
not ( n12659 , n12438 );
or ( n82430 , n12658 , n12659 );
not ( n12664 , n12434 );
nand ( n82432 , n82430 , n12664 );
not ( n12666 , n82432 );
not ( n12667 , n12666 );
or ( n12668 , n12657 , n12667 );
nand ( n12669 , n82432 , n12655 );
nand ( n12670 , n12668 , n12669 );
not ( n12671 , n12670 );
not ( n12672 , n12671 );
or ( n12673 , n12652 , n12672 );
not ( n12674 , n12671 );
nand ( n12675 , n12674 , n12467 );
nand ( n12676 , n12673 , n12675 );
not ( n12677 , n12676 );
or ( n12678 , n12651 , n12677 );
nand ( n12679 , n12323 , n12247 );
not ( n12680 , n12679 );
not ( n12681 , n12680 );
not ( n12682 , n12261 );
not ( n12683 , n12109 );
or ( n12684 , n12682 , n12683 );
nand ( n12685 , n12684 , n12473 );
not ( n12686 , n12685 );
not ( n12687 , n12686 );
or ( n12688 , n12681 , n12687 );
nand ( n82456 , n12685 , n12679 );
nand ( n12693 , n12688 , n82456 );
not ( n12694 , n12693 );
and ( n12695 , n12694 , n499 );
not ( n12696 , n12694 );
and ( n12697 , n12696 , n12467 );
or ( n12698 , n12695 , n12697 );
not ( n12699 , n12647 );
xor ( n12700 , n500 , n499 );
nand ( n12701 , n12699 , n12700 );
not ( n12702 , n12701 );
nand ( n12703 , n12698 , n12702 );
nand ( n12704 , n12678 , n12703 );
and ( n12705 , n12646 , n12704 );
and ( n12706 , n12519 , n12645 );
or ( n12707 , n12705 , n12706 );
xor ( n12708 , n12464 , n12707 );
not ( n12709 , n12580 );
and ( n12710 , n12532 , n489 );
not ( n12711 , n12532 );
and ( n12712 , n12711 , n12560 );
or ( n12713 , n12710 , n12712 );
not ( n12714 , n12713 );
or ( n12715 , n12709 , n12714 );
nand ( n12716 , n11864 , n11873 );
not ( n12717 , n12716 );
not ( n12718 , n12717 );
nand ( n12719 , n11871 , n82296 );
not ( n12720 , n12719 );
not ( n12721 , n12720 );
or ( n12722 , n12718 , n12721 );
nand ( n12723 , n12719 , n12716 );
nand ( n12724 , n12722 , n12723 );
buf ( n12725 , n12724 );
xor ( n12726 , n489 , n12725 );
nand ( n12727 , n12542 , n12726 );
nand ( n12728 , n12715 , n12727 );
not ( n12729 , n11834 );
not ( n12730 , n12729 );
not ( n12731 , n11862 );
or ( n12732 , n12730 , n12731 );
nand ( n12733 , n12732 , n11873 );
not ( n12734 , n11828 );
xor ( n12735 , n12733 , n12734 );
and ( n12736 , n489 , n12735 );
xor ( n12737 , n12728 , n12736 );
not ( n12738 , n12638 );
not ( n12739 , n491 );
not ( n12740 , n12577 );
or ( n12741 , n12739 , n12740 );
nand ( n12742 , n12573 , n12610 );
nand ( n12743 , n12741 , n12742 );
not ( n12744 , n12743 );
or ( n12745 , n12738 , n12744 );
not ( n12746 , n491 );
not ( n12747 , n12556 );
or ( n12748 , n12746 , n12747 );
nand ( n12749 , n12559 , n12610 );
nand ( n12750 , n12748 , n12749 );
nand ( n12751 , n12750 , n12595 );
nand ( n82516 , n12745 , n12751 );
and ( n82517 , n12737 , n82516 );
and ( n12754 , n12728 , n12736 );
or ( n12755 , n82517 , n12754 );
xor ( n12756 , n494 , n495 );
not ( n12757 , n12756 );
not ( n12758 , n12757 );
not ( n12759 , n12758 );
and ( n12760 , n12024 , n12048 );
not ( n12761 , n12760 );
not ( n12762 , n12619 );
or ( n12763 , n12761 , n12762 );
not ( n12764 , n12082 );
nand ( n12765 , n12763 , n12764 );
buf ( n12766 , n12765 );
not ( n12767 , n12086 );
nand ( n12768 , n12767 , n12074 );
not ( n12769 , n12768 );
and ( n12770 , n12766 , n12769 );
not ( n12771 , n12766 );
and ( n12772 , n12771 , n12768 );
nor ( n12773 , n12770 , n12772 );
buf ( n12774 , n12773 );
not ( n12775 , n493 );
and ( n12776 , n12774 , n12775 );
not ( n12777 , n12774 );
and ( n12778 , n12777 , n493 );
or ( n12779 , n12776 , n12778 );
not ( n12780 , n12779 );
or ( n12781 , n12759 , n12780 );
not ( n12782 , n493 );
buf ( n12783 , n12629 );
not ( n12784 , n12783 );
or ( n12785 , n12782 , n12784 );
nand ( n12786 , n12775 , n12635 );
nand ( n12787 , n12785 , n12786 );
and ( n12788 , n493 , n494 );
nor ( n12789 , n493 , n494 );
nor ( n12790 , n12788 , n12789 );
and ( n12791 , n12757 , n12790 );
nand ( n12792 , n12787 , n12791 );
nand ( n12793 , n12781 , n12792 );
xor ( n12794 , n12755 , n12793 );
buf ( n12795 , n12538 );
not ( n12796 , n12795 );
not ( n12797 , n12562 );
or ( n12798 , n12796 , n12797 );
nand ( n12799 , n12713 , n12542 );
nand ( n12800 , n12798 , n12799 );
and ( n12801 , n489 , n12725 );
xor ( n12802 , n12800 , n12801 );
not ( n12803 , n12638 );
not ( n12804 , n12612 );
or ( n12805 , n12803 , n12804 );
nand ( n12806 , n12743 , n12595 );
nand ( n12807 , n12805 , n12806 );
xor ( n12808 , n12802 , n12807 );
and ( n12809 , n12794 , n12808 );
and ( n12810 , n12755 , n12793 );
or ( n12811 , n12809 , n12810 );
not ( n12812 , n502 );
nand ( n12813 , n12812 , n501 );
not ( n12814 , n501 );
nand ( n12815 , n12814 , n502 );
and ( n12816 , n12813 , n12815 );
and ( n12817 , n502 , n3027 );
not ( n12818 , n502 );
and ( n12819 , n12818 , n503 );
or ( n12820 , n12817 , n12819 );
nor ( n12821 , n12816 , n12820 );
buf ( n12822 , n12821 );
not ( n12823 , n12822 );
nand ( n12824 , n12333 , n12330 );
not ( n12825 , n12824 );
not ( n12826 , n12654 );
not ( n12827 , n12440 );
or ( n12828 , n12826 , n12827 );
nand ( n12829 , n12828 , n12653 );
not ( n12830 , n12829 );
or ( n12831 , n12825 , n12830 );
not ( n12832 , n12824 );
nand ( n12833 , n12440 , n12654 );
nand ( n12834 , n12832 , n12833 , n12653 );
nand ( n12835 , n12831 , n12834 );
not ( n82600 , n12835 );
and ( n12837 , n70432 , n82600 );
not ( n12838 , n70432 );
and ( n12839 , n12838 , n12835 );
nor ( n12840 , n12837 , n12839 );
not ( n12841 , n12840 );
or ( n12842 , n12823 , n12841 );
buf ( n12843 , n12820 );
not ( n12844 , n501 );
or ( n12845 , n10682 , n10664 );
nand ( n12846 , n12343 , n12845 );
not ( n12847 , n12846 );
not ( n12848 , n12339 );
or ( n12849 , n12847 , n12848 );
or ( n12850 , n12846 , n12339 );
nand ( n12851 , n12849 , n12850 );
not ( n12852 , n12851 );
not ( n12853 , n12852 );
or ( n12854 , n12844 , n12853 );
not ( n12855 , n12852 );
not ( n12856 , n501 );
nand ( n12857 , n12855 , n12856 );
nand ( n12858 , n12854 , n12857 );
nand ( n12859 , n12843 , n12858 );
nand ( n12860 , n12842 , n12859 );
xor ( n12861 , n12811 , n12860 );
not ( n12862 , n12462 );
not ( n12863 , n10691 );
nand ( n12864 , n12863 , n12345 );
not ( n12865 , n12864 );
not ( n12866 , n12439 );
not ( n12867 , n12108 );
nand ( n12868 , n12867 , n12262 );
not ( n12869 , n12868 );
or ( n12870 , n12866 , n12869 );
and ( n12871 , n12316 , n12845 );
nand ( n12872 , n12870 , n12871 );
and ( n12873 , n12335 , n12845 );
not ( n12874 , n12343 );
nor ( n12875 , n12873 , n12874 );
nand ( n12876 , n12326 , n12845 );
not ( n12877 , n12876 );
nand ( n12878 , n12877 , n12316 );
nand ( n12879 , n12872 , n12875 , n12878 );
not ( n12880 , n12879 );
or ( n12881 , n12865 , n12880 );
not ( n12882 , n12873 );
nor ( n12883 , n12864 , n12874 );
nand ( n12884 , n12882 , n12872 , n12878 , n12883 );
nand ( n12885 , n12881 , n12884 );
not ( n12886 , n12885 );
not ( n12887 , n12886 );
or ( n12888 , n12862 , n12887 );
nand ( n12889 , n12459 , n504 );
nand ( n12890 , n12888 , n12889 );
and ( n12891 , n12861 , n12890 );
and ( n12892 , n12811 , n12860 );
or ( n82657 , n12891 , n12892 );
and ( n82658 , n12708 , n82657 );
and ( n12895 , n12464 , n12707 );
or ( n12896 , n82658 , n12895 );
and ( n12897 , n12582 , n12533 );
not ( n12898 , n12638 );
not ( n12899 , n491 );
not ( n12900 , n12774 );
not ( n12901 , n12900 );
or ( n12902 , n12899 , n12901 );
nand ( n12903 , n12774 , n12610 );
nand ( n12904 , n12902 , n12903 );
not ( n12905 , n12904 );
or ( n12906 , n12898 , n12905 );
nand ( n12907 , n12637 , n12595 );
nand ( n12908 , n12906 , n12907 );
xor ( n12909 , n12897 , n12908 );
and ( n12910 , n12559 , n489 );
not ( n12911 , n12795 );
not ( n12912 , n489 );
not ( n12913 , n12607 );
or ( n12914 , n12912 , n12913 );
nand ( n12915 , n12606 , n12560 );
nand ( n12916 , n12914 , n12915 );
not ( n12917 , n12916 );
or ( n12918 , n12911 , n12917 );
nand ( n12919 , n12579 , n12542 );
nand ( n12920 , n12918 , n12919 );
xor ( n12921 , n12910 , n12920 );
xor ( n12922 , n12909 , n12921 );
not ( n12923 , n12470 );
not ( n12924 , n497 );
not ( n12925 , n12694 );
or ( n12926 , n12924 , n12925 );
nand ( n12927 , n12693 , n12486 );
nand ( n12928 , n12926 , n12927 );
not ( n12929 , n12928 );
or ( n12930 , n12923 , n12929 );
nand ( n12931 , n12488 , n12517 );
nand ( n12932 , n12930 , n12931 );
xor ( n12933 , n12922 , n12932 );
not ( n12934 , n12791 );
not ( n12935 , n12779 );
or ( n12936 , n12934 , n12935 );
not ( n12937 , n493 );
not ( n12938 , n12074 );
not ( n12939 , n12765 );
or ( n12940 , n12938 , n12939 );
buf ( n12941 , n12767 );
nand ( n12942 , n12940 , n12941 );
nand ( n12943 , n12083 , n12090 );
not ( n12944 , n12943 );
and ( n12945 , n12942 , n12944 );
not ( n12946 , n12942 );
and ( n12947 , n12946 , n12943 );
nor ( n12948 , n12945 , n12947 );
buf ( n12949 , n12948 );
not ( n12950 , n12949 );
not ( n12951 , n12950 );
or ( n12952 , n12937 , n12951 );
nand ( n12953 , n12949 , n12775 );
nand ( n12954 , n12952 , n12953 );
nand ( n12955 , n12954 , n12758 );
nand ( n12956 , n12936 , n12955 );
xor ( n12957 , n12800 , n12801 );
and ( n12958 , n12957 , n12807 );
and ( n12959 , n12800 , n12801 );
or ( n12960 , n12958 , n12959 );
xor ( n12961 , n12956 , n12960 );
and ( n12962 , n496 , n497 );
not ( n12963 , n496 );
and ( n82728 , n12963 , n12486 );
or ( n12965 , n12962 , n82728 );
and ( n12966 , n496 , n495 );
nor ( n12967 , n495 , n496 );
nor ( n12968 , n12966 , n12967 );
and ( n12969 , n12965 , n12968 );
not ( n12970 , n12969 );
not ( n12971 , n495 );
nand ( n12972 , n12100 , n11410 );
not ( n12973 , n12972 );
buf ( n12974 , n12496 );
not ( n82739 , n12974 );
or ( n12976 , n12973 , n82739 );
not ( n12977 , n12974 );
not ( n12978 , n12972 );
nand ( n12979 , n12977 , n12978 );
nand ( n12980 , n12976 , n12979 );
not ( n12981 , n12980 );
not ( n12982 , n12981 );
or ( n12983 , n12971 , n12982 );
not ( n12984 , n495 );
buf ( n12985 , n12980 );
nand ( n12986 , n12984 , n12985 );
nand ( n12987 , n12983 , n12986 );
not ( n12988 , n12987 );
or ( n12989 , n12970 , n12988 );
not ( n12990 , n12765 );
not ( n12991 , n12071 );
nand ( n12992 , n12991 , n12074 );
nor ( n12993 , n12992 , n11409 );
not ( n12994 , n12993 );
or ( n12995 , n12990 , n12994 );
not ( n12996 , n12091 );
not ( n12997 , n11410 );
or ( n12998 , n12996 , n12997 );
nand ( n12999 , n12998 , n12100 );
not ( n13000 , n12999 );
nand ( n13001 , n12995 , n13000 );
nand ( n13002 , n11419 , n12099 );
not ( n13003 , n13002 );
and ( n13004 , n13001 , n13003 );
not ( n13005 , n13001 );
and ( n13006 , n13005 , n13002 );
nor ( n13007 , n13004 , n13006 );
buf ( n13008 , n13007 );
not ( n13009 , n13008 );
and ( n13010 , n495 , n13009 );
not ( n13011 , n495 );
and ( n13012 , n13011 , n13008 );
or ( n13013 , n13010 , n13012 );
not ( n13014 , n13013 );
or ( n13015 , n13014 , n12965 );
nand ( n13016 , n12989 , n13015 );
and ( n13017 , n12961 , n13016 );
and ( n13018 , n12956 , n12960 );
or ( n13019 , n13017 , n13018 );
xor ( n13020 , n12933 , n13019 );
nor ( n13021 , n12586 , n12643 );
not ( n13022 , n12758 );
and ( n13023 , n12985 , n493 );
not ( n13024 , n12985 );
and ( n13025 , n13024 , n1976 );
nor ( n13026 , n13023 , n13025 );
not ( n13027 , n13026 );
or ( n13028 , n13022 , n13027 );
nand ( n13029 , n12954 , n12791 );
nand ( n13030 , n13028 , n13029 );
xor ( n13031 , n13021 , n13030 );
not ( n13032 , n12965 );
not ( n13033 , n13032 );
and ( n13034 , n495 , n12506 );
not ( n13035 , n495 );
and ( n13036 , n13035 , n12505 );
or ( n13037 , n13034 , n13036 );
not ( n13038 , n13037 );
or ( n13039 , n13033 , n13038 );
nand ( n13040 , n13013 , n12969 );
nand ( n13041 , n13039 , n13040 );
xor ( n13042 , n13031 , n13041 );
not ( n13043 , n12843 );
and ( n13044 , n501 , n12886 );
not ( n13045 , n501 );
not ( n13046 , n12886 );
and ( n13047 , n13045 , n13046 );
or ( n13048 , n13044 , n13047 );
not ( n13049 , n13048 );
or ( n13050 , n13043 , n13049 );
nand ( n13051 , n12858 , n12821 );
nand ( n82816 , n13050 , n13051 );
xor ( n13056 , n13042 , n82816 );
not ( n82818 , n12650 );
and ( n13058 , n12835 , n12467 );
not ( n13059 , n12835 );
and ( n13060 , n13059 , n499 );
or ( n13061 , n13058 , n13060 );
not ( n13062 , n13061 );
or ( n13063 , n82818 , n13062 );
nand ( n13064 , n12676 , n12702 );
nand ( n13065 , n13063 , n13064 );
xor ( n13066 , n13056 , n13065 );
xor ( n13067 , n13020 , n13066 );
xor ( n13068 , n12956 , n12960 );
xor ( n13069 , n13068 , n13016 );
not ( n13070 , n13032 );
not ( n13071 , n12987 );
or ( n13072 , n13070 , n13071 );
not ( n13073 , n495 );
not ( n13074 , n12950 );
or ( n13075 , n13073 , n13074 );
not ( n82837 , n12949 );
not ( n13080 , n82837 );
nand ( n13081 , n13080 , n3325 );
nand ( n13082 , n13075 , n13081 );
nand ( n13083 , n13082 , n12969 );
nand ( n13084 , n13072 , n13083 );
not ( n13085 , n12470 );
not ( n13086 , n12511 );
or ( n13087 , n13085 , n13086 );
and ( n13088 , n12486 , n13009 );
not ( n13089 , n12486 );
and ( n13090 , n13089 , n13008 );
or ( n13091 , n13088 , n13090 );
not ( n13092 , n13091 );
nand ( n13093 , n13092 , n12517 );
nand ( n13094 , n13087 , n13093 );
xor ( n13095 , n13084 , n13094 );
not ( n13096 , n12758 );
not ( n13097 , n12787 );
or ( n13098 , n13096 , n13097 );
not ( n13099 , n493 );
not ( n13100 , n12605 );
not ( n13101 , n13100 );
or ( n13102 , n13099 , n13101 );
nand ( n13103 , n12775 , n12606 );
nand ( n13104 , n13102 , n13103 );
nand ( n13105 , n13104 , n12791 );
nand ( n13106 , n13098 , n13105 );
not ( n13107 , n12580 );
not ( n13108 , n12726 );
or ( n13109 , n13107 , n13108 );
xor ( n13110 , n489 , n12735 );
nand ( n13111 , n13110 , n12542 );
nand ( n13112 , n13109 , n13111 );
nand ( n13113 , n11827 , n11752 );
xnor ( n13114 , n11823 , n13113 );
and ( n13115 , n489 , n13114 );
xor ( n13116 , n13112 , n13115 );
not ( n13117 , n12638 );
not ( n13118 , n12750 );
or ( n13119 , n13117 , n13118 );
and ( n13120 , n12531 , n12610 );
not ( n13121 , n12531 );
and ( n13122 , n13121 , n491 );
or ( n13123 , n13120 , n13122 );
nand ( n13124 , n13123 , n12595 );
nand ( n13125 , n13119 , n13124 );
and ( n13126 , n13116 , n13125 );
and ( n13127 , n13112 , n13115 );
or ( n13128 , n13126 , n13127 );
xor ( n13129 , n13106 , n13128 );
not ( n13130 , n13032 );
not ( n13131 , n13082 );
or ( n13132 , n13130 , n13131 );
and ( n13133 , n495 , n12900 );
not ( n13134 , n495 );
and ( n13135 , n13134 , n12774 );
or ( n13136 , n13133 , n13135 );
nand ( n13137 , n13136 , n12969 );
nand ( n13138 , n13132 , n13137 );
and ( n13139 , n13129 , n13138 );
and ( n13140 , n13106 , n13128 );
or ( n13141 , n13139 , n13140 );
and ( n82900 , n13095 , n13141 );
and ( n82901 , n13084 , n13094 );
or ( n13144 , n82900 , n82901 );
xor ( n13145 , n13069 , n13144 );
xor ( n13146 , n12519 , n12645 );
xor ( n13147 , n13146 , n12704 );
and ( n13148 , n13145 , n13147 );
and ( n13149 , n13069 , n13144 );
or ( n13150 , n13148 , n13149 );
and ( n13151 , n13067 , n13150 );
and ( n13152 , n13020 , n13066 );
or ( n13153 , n13151 , n13152 );
xor ( n13154 , n12896 , n13153 );
xor ( n13155 , n13042 , n82816 );
and ( n13156 , n13155 , n13065 );
and ( n13157 , n13042 , n82816 );
or ( n13158 , n13156 , n13157 );
not ( n13159 , n12822 );
not ( n13160 , n13048 );
or ( n13161 , n13159 , n13160 );
not ( n13162 , n501 );
not ( n13163 , n12453 );
or ( n13164 , n13162 , n13163 );
nand ( n13165 , n12456 , n12856 );
nand ( n13166 , n13164 , n13165 );
nand ( n13167 , n13166 , n12843 );
nand ( n13168 , n13161 , n13167 );
not ( n13169 , n12702 );
not ( n13170 , n13061 );
or ( n13171 , n13169 , n13170 );
and ( n13172 , n499 , n12855 );
not ( n13173 , n499 );
and ( n13174 , n13173 , n12852 );
nor ( n13175 , n13172 , n13174 );
nand ( n13176 , n12650 , n13175 );
nand ( n13177 , n13171 , n13176 );
xor ( n13178 , n13168 , n13177 );
not ( n13179 , n12462 );
not ( n13180 , n12425 );
or ( n13181 , n13179 , n13180 );
not ( n13182 , n503 );
not ( n13183 , n10692 );
nand ( n13184 , n10467 , n12412 );
nor ( n13185 , n13183 , n13184 );
and ( n13186 , n13185 , n12316 );
not ( n13187 , n13186 );
not ( n13188 , n82432 );
or ( n13189 , n13187 , n13188 );
not ( n13190 , n12335 );
not ( n13191 , n13185 );
or ( n13192 , n13190 , n13191 );
nand ( n13193 , n13192 , n12410 );
nand ( n13194 , n12352 , n12412 );
not ( n13195 , n13194 );
nor ( n13196 , n13193 , n13195 );
nand ( n13197 , n13189 , n13196 );
not ( n13198 , n12369 );
not ( n13199 , n12377 );
or ( n13200 , n13198 , n13199 );
or ( n13201 , n12369 , n12377 );
nand ( n13202 , n13201 , n80235 );
nand ( n13203 , n13200 , n13202 );
xor ( n13204 , n12368 , n12378 );
and ( n13205 , n13204 , n12395 );
and ( n13206 , n12368 , n12378 );
or ( n13207 , n13205 , n13206 );
xor ( n13208 , n13203 , n13207 );
not ( n13209 , n12389 );
not ( n13210 , n10191 );
or ( n13211 , n13209 , n13210 );
nand ( n13212 , n10194 , n461 );
nand ( n13213 , n13211 , n13212 );
not ( n13214 , n13213 );
and ( n13215 , n457 , n526 );
not ( n13216 , n12383 );
not ( n82975 , n10127 );
or ( n13218 , n13216 , n82975 );
xor ( n13219 , n457 , n524 );
nand ( n13220 , n10068 , n13219 );
nand ( n13221 , n13218 , n13220 );
xor ( n13222 , n13215 , n13221 );
not ( n13223 , n12375 );
not ( n13224 , n10087 );
or ( n13225 , n13223 , n13224 );
xor ( n13226 , n459 , n522 );
nand ( n13227 , n10094 , n13226 );
nand ( n13228 , n13225 , n13227 );
xor ( n13229 , n13222 , n13228 );
xor ( n13230 , n13214 , n13229 );
xor ( n13231 , n12385 , n82161 );
and ( n13232 , n13231 , n12394 );
and ( n13233 , n12385 , n82161 );
or ( n13234 , n13232 , n13233 );
xor ( n13235 , n13230 , n13234 );
xor ( n13236 , n13208 , n13235 );
not ( n13237 , n12363 );
not ( n13238 , n12396 );
or ( n13239 , n13237 , n13238 );
not ( n13240 , n12364 );
not ( n13241 , n12396 );
not ( n13242 , n13241 );
or ( n13243 , n13240 , n13242 );
nand ( n13244 , n13243 , n12401 );
nand ( n13245 , n13239 , n13244 );
nor ( n13246 , n13236 , n13245 );
not ( n13247 , n13246 );
nand ( n13248 , n13245 , n13236 );
nand ( n13249 , n13247 , n13248 );
and ( n13250 , n13197 , n13249 );
not ( n13251 , n13197 );
not ( n13252 , n13249 );
and ( n13253 , n13251 , n13252 );
nor ( n13254 , n13250 , n13253 );
buf ( n13255 , n13254 );
not ( n13256 , n13255 );
or ( n13257 , n13182 , n13256 );
not ( n13258 , n13254 );
nand ( n13259 , n13258 , n12423 );
nand ( n13260 , n13257 , n13259 );
nand ( n13261 , n13260 , n504 );
nand ( n13262 , n13181 , n13261 );
xor ( n13263 , n13178 , n13262 );
xor ( n13264 , n13158 , n13263 );
not ( n13265 , n12791 );
not ( n13266 , n13026 );
or ( n13267 , n13265 , n13266 );
and ( n13268 , n493 , n13008 );
not ( n13269 , n493 );
and ( n13270 , n13269 , n13009 );
nor ( n13271 , n13268 , n13270 );
nand ( n13272 , n13271 , n12758 );
nand ( n13273 , n13267 , n13272 );
not ( n13274 , n12969 );
not ( n13275 , n13037 );
or ( n13276 , n13274 , n13275 );
and ( n13277 , n495 , n12481 );
not ( n13278 , n495 );
and ( n13279 , n13278 , n12482 );
nor ( n13280 , n13277 , n13279 );
nand ( n13281 , n13280 , n13032 );
nand ( n13282 , n13276 , n13281 );
xor ( n13283 , n13273 , n13282 );
xor ( n13284 , n12897 , n12908 );
and ( n13285 , n13284 , n12921 );
and ( n13286 , n12897 , n12908 );
or ( n13287 , n13285 , n13286 );
xor ( n13288 , n13283 , n13287 );
xor ( n13289 , n12922 , n12932 );
and ( n13290 , n13289 , n13019 );
and ( n13291 , n12922 , n12932 );
or ( n13292 , n13290 , n13291 );
xor ( n13293 , n13288 , n13292 );
not ( n13294 , n12517 );
not ( n13295 , n12928 );
or ( n13296 , n13294 , n13295 );
not ( n13297 , n497 );
not ( n13298 , n12671 );
or ( n13299 , n13297 , n13298 );
nand ( n13300 , n12674 , n12486 );
nand ( n13301 , n13299 , n13300 );
nand ( n13302 , n13301 , n12470 );
nand ( n13303 , n13296 , n13302 );
and ( n13304 , n12949 , n12610 );
not ( n13305 , n12949 );
and ( n13306 , n13305 , n491 );
or ( n13307 , n13304 , n13306 );
not ( n13308 , n13307 );
not ( n13309 , n12638 );
or ( n13310 , n13308 , n13309 );
nand ( n83069 , n12904 , n12595 );
nand ( n83070 , n13310 , n83069 );
and ( n13313 , n12910 , n12920 );
xor ( n13314 , n83070 , n13313 );
not ( n13315 , n12542 );
not ( n13316 , n12916 );
or ( n13317 , n13315 , n13316 );
not ( n13318 , n489 );
not ( n13319 , n12629 );
or ( n13320 , n13318 , n13319 );
nand ( n13321 , n12628 , n12560 );
nand ( n13322 , n13320 , n13321 );
nand ( n13323 , n13322 , n12795 );
nand ( n13324 , n13317 , n13323 );
and ( n13325 , n12573 , n489 );
xor ( n13326 , n13324 , n13325 );
xor ( n13327 , n13314 , n13326 );
xor ( n13328 , n13303 , n13327 );
xor ( n13329 , n13021 , n13030 );
and ( n13330 , n13329 , n13041 );
and ( n13331 , n13021 , n13030 );
or ( n13332 , n13330 , n13331 );
xor ( n13333 , n13328 , n13332 );
xor ( n83092 , n13293 , n13333 );
xor ( n13335 , n13264 , n83092 );
xor ( n13336 , n13154 , n13335 );
not ( n13337 , n13336 );
xor ( n13338 , n12464 , n12707 );
xor ( n13339 , n13338 , n82657 );
not ( n13340 , n12650 );
not ( n13341 , n12698 );
or ( n13342 , n13340 , n13341 );
and ( n13343 , n499 , n12482 );
not ( n13344 , n499 );
and ( n13345 , n13344 , n12481 );
nor ( n13346 , n13343 , n13345 );
not ( n13347 , n13346 );
nand ( n13348 , n13347 , n12702 );
nand ( n13349 , n13342 , n13348 );
xor ( n13350 , n12755 , n12793 );
xor ( n13351 , n13350 , n12808 );
xor ( n13352 , n13349 , n13351 );
not ( n13353 , n12843 );
not ( n13354 , n12840 );
or ( n13355 , n13353 , n13354 );
not ( n13356 , n501 );
not ( n13357 , n12670 );
not ( n13358 , n13357 );
or ( n13359 , n13356 , n13358 );
or ( n13360 , n13357 , n501 );
nand ( n13361 , n13359 , n13360 );
nand ( n13362 , n13361 , n12822 );
nand ( n13363 , n13355 , n13362 );
and ( n13364 , n13352 , n13363 );
and ( n13365 , n13349 , n13351 );
or ( n13366 , n13364 , n13365 );
not ( n13367 , n70376 );
nand ( n13368 , n13367 , n12886 );
buf ( n13369 , n12851 );
not ( n13370 , n13369 );
nand ( n13371 , n13370 , n12462 );
buf ( n13372 , n12885 );
nand ( n13373 , n13372 , n3971 );
nand ( n13374 , n13368 , n13371 , n13373 );
xor ( n13375 , n12728 , n12736 );
xor ( n13376 , n13375 , n82516 );
not ( n13377 , n497 );
not ( n13378 , n12985 );
not ( n13379 , n13378 );
or ( n13380 , n13377 , n13379 );
nand ( n13381 , n12985 , n12486 );
nand ( n13382 , n13380 , n13381 );
not ( n13383 , n13382 );
not ( n13384 , n12517 );
or ( n13385 , n13383 , n13384 );
or ( n13386 , n13091 , n12469 );
nand ( n13387 , n13385 , n13386 );
xor ( n13388 , n13376 , n13387 );
and ( n13389 , n12467 , n12509 );
not ( n13390 , n12467 );
and ( n13391 , n13390 , n12506 );
nor ( n13392 , n13389 , n13391 );
or ( n13393 , n13392 , n12701 );
or ( n13394 , n13346 , n12649 );
nand ( n13395 , n13393 , n13394 );
and ( n13396 , n13388 , n13395 );
and ( n13397 , n13376 , n13387 );
or ( n13398 , n13396 , n13397 );
xor ( n13399 , n13374 , n13398 );
xor ( n13400 , n13084 , n13094 );
xor ( n13401 , n13400 , n13141 );
and ( n13402 , n13399 , n13401 );
and ( n13403 , n13374 , n13398 );
or ( n13404 , n13402 , n13403 );
xor ( n13405 , n13366 , n13404 );
xor ( n13406 , n12811 , n12860 );
xor ( n13407 , n13406 , n12890 );
and ( n13408 , n13405 , n13407 );
and ( n13409 , n13366 , n13404 );
or ( n13410 , n13408 , n13409 );
xor ( n13411 , n13339 , n13410 );
xor ( n13412 , n13020 , n13066 );
xor ( n13413 , n13412 , n13150 );
and ( n13414 , n13411 , n13413 );
and ( n13415 , n13339 , n13410 );
or ( n13416 , n13414 , n13415 );
not ( n13417 , n13416 );
nand ( n83176 , n13337 , n13417 );
xor ( n13422 , n13339 , n13410 );
xor ( n83178 , n13422 , n13413 );
xor ( n13424 , n13069 , n13144 );
xor ( n13425 , n13424 , n13147 );
not ( n13426 , n12795 );
not ( n13427 , n13110 );
or ( n13428 , n13426 , n13427 );
xor ( n13429 , n489 , n13114 );
nand ( n13430 , n13429 , n12542 );
nand ( n13431 , n13428 , n13430 );
not ( n13432 , n11803 );
not ( n13433 , n11821 );
not ( n13434 , n11820 );
or ( n13435 , n13433 , n13434 );
nand ( n13436 , n13435 , n11817 );
not ( n13437 , n13436 );
or ( n13438 , n13432 , n13437 );
or ( n13439 , n13436 , n11803 );
nand ( n13440 , n13438 , n13439 );
buf ( n13441 , n13440 );
and ( n13442 , n489 , n13441 );
xor ( n13443 , n13431 , n13442 );
not ( n13444 , n12638 );
not ( n13445 , n13123 );
or ( n13446 , n13444 , n13445 );
not ( n83202 , n491 );
not ( n13451 , n12724 );
not ( n13452 , n13451 );
or ( n13453 , n83202 , n13452 );
nand ( n13454 , n12725 , n12610 );
nand ( n13455 , n13453 , n13454 );
nand ( n13456 , n13455 , n12595 );
nand ( n13457 , n13446 , n13456 );
and ( n13458 , n13443 , n13457 );
and ( n13459 , n13431 , n13442 );
or ( n13460 , n13458 , n13459 );
not ( n13461 , n12758 );
not ( n13462 , n13104 );
or ( n13463 , n13461 , n13462 );
not ( n13464 , n493 );
not ( n13465 , n82342 );
or ( n13466 , n13464 , n13465 );
or ( n13467 , n82342 , n493 );
nand ( n13468 , n13466 , n13467 );
not ( n13469 , n13468 );
nand ( n13470 , n13469 , n12791 );
nand ( n13471 , n13463 , n13470 );
xor ( n13472 , n13460 , n13471 );
xor ( n13473 , n13112 , n13115 );
xor ( n13474 , n13473 , n13125 );
and ( n13475 , n13472 , n13474 );
and ( n13476 , n13460 , n13471 );
or ( n13477 , n13475 , n13476 );
xor ( n13478 , n13106 , n13128 );
xor ( n13479 , n13478 , n13138 );
xor ( n13480 , n13477 , n13479 );
not ( n13481 , n12822 );
not ( n13482 , n501 );
buf ( n13483 , n12693 );
not ( n13484 , n13483 );
not ( n13485 , n13484 );
or ( n13486 , n13482 , n13485 );
nand ( n13487 , n13483 , n12856 );
nand ( n13488 , n13486 , n13487 );
not ( n13489 , n13488 );
or ( n13490 , n13481 , n13489 );
nand ( n13491 , n13361 , n12843 );
nand ( n13492 , n13490 , n13491 );
and ( n13493 , n13480 , n13492 );
and ( n13494 , n13477 , n13479 );
or ( n13495 , n13493 , n13494 );
not ( n13496 , n13032 );
not ( n13497 , n13136 );
or ( n13498 , n13496 , n13497 );
and ( n13499 , n495 , n12629 );
not ( n13500 , n495 );
and ( n13501 , n13500 , n12628 );
nor ( n13502 , n13499 , n13501 );
not ( n13503 , n13502 );
nand ( n83256 , n13503 , n12969 );
nand ( n83257 , n13498 , n83256 );
and ( n13506 , n11802 , n11776 );
buf ( n13507 , n11798 );
and ( n13508 , n13506 , n13507 );
not ( n13509 , n13506 );
not ( n13510 , n13507 );
and ( n13511 , n13509 , n13510 );
nor ( n13512 , n13508 , n13511 );
and ( n13513 , n489 , n13512 );
xor ( n13514 , n489 , n13441 );
not ( n13515 , n13514 );
not ( n13516 , n12542 );
or ( n13517 , n13515 , n13516 );
not ( n13518 , n13429 );
or ( n13519 , n13518 , n12539 );
nand ( n13520 , n13517 , n13519 );
xor ( n13521 , n13513 , n13520 );
not ( n13522 , n12595 );
not ( n13523 , n491 );
not ( n13524 , n12735 );
not ( n13525 , n13524 );
or ( n13526 , n13523 , n13525 );
nand ( n13527 , n12735 , n12610 );
nand ( n13528 , n13526 , n13527 );
not ( n13529 , n13528 );
or ( n13530 , n13522 , n13529 );
nand ( n13531 , n13455 , n12638 );
nand ( n13532 , n13530 , n13531 );
and ( n13533 , n13521 , n13532 );
and ( n13534 , n13513 , n13520 );
or ( n13535 , n13533 , n13534 );
and ( n13536 , n12775 , n12556 );
not ( n13537 , n12775 );
and ( n13538 , n13537 , n12559 );
or ( n13539 , n13536 , n13538 );
not ( n13540 , n12791 );
or ( n13541 , n13539 , n13540 );
or ( n13542 , n13468 , n12757 );
nand ( n13543 , n13541 , n13542 );
xor ( n13544 , n13535 , n13543 );
xor ( n13545 , n13431 , n13442 );
xor ( n13546 , n13545 , n13457 );
and ( n13547 , n13544 , n13546 );
and ( n13548 , n13535 , n13543 );
or ( n13549 , n13547 , n13548 );
xor ( n13550 , n83257 , n13549 );
not ( n13551 , n12470 );
not ( n13552 , n13382 );
or ( n13553 , n13551 , n13552 );
and ( n13554 , n12486 , n12949 );
not ( n13555 , n12486 );
and ( n13556 , n13555 , n82837 );
nor ( n13557 , n13554 , n13556 );
not ( n13558 , n13557 );
nand ( n13559 , n13558 , n12517 );
nand ( n13560 , n13553 , n13559 );
and ( n13561 , n13550 , n13560 );
and ( n13562 , n83257 , n13549 );
or ( n13563 , n13561 , n13562 );
not ( n13564 , n499 );
not ( n13565 , n13009 );
or ( n13566 , n13564 , n13565 );
nand ( n13567 , n13008 , n12467 );
nand ( n13568 , n13566 , n13567 );
nand ( n13569 , n13568 , n12702 );
nand ( n13570 , n12648 , n499 );
or ( n13571 , n12505 , n13570 );
nor ( n13572 , n12649 , n499 );
nand ( n13573 , n12505 , n13572 );
nand ( n13574 , n13569 , n13571 , n13573 );
xor ( n13575 , n13460 , n13471 );
xor ( n13576 , n13575 , n13474 );
xor ( n13577 , n13574 , n13576 );
and ( n13578 , n495 , n13100 );
not ( n13579 , n495 );
and ( n13580 , n13579 , n12606 );
nor ( n13581 , n13578 , n13580 );
not ( n13582 , n12969 );
or ( n83335 , n13581 , n13582 );
or ( n13584 , n13502 , n12965 );
nand ( n13585 , n83335 , n13584 );
xor ( n13586 , n12486 , n12774 );
or ( n13587 , n13586 , n13384 );
or ( n13588 , n13557 , n12469 );
nand ( n13589 , n13587 , n13588 );
xor ( n13590 , n13585 , n13589 );
not ( n13591 , n11786 );
not ( n13592 , n13591 );
not ( n13593 , n13592 );
not ( n13594 , n11794 );
nand ( n13595 , n13594 , n11797 );
not ( n13596 , n13595 );
not ( n13597 , n13596 );
or ( n13598 , n13593 , n13597 );
nand ( n13599 , n13595 , n13591 );
nand ( n13600 , n13598 , n13599 );
and ( n13601 , n13600 , n489 );
not ( n13602 , n12795 );
not ( n13603 , n13514 );
or ( n13604 , n13602 , n13603 );
xor ( n13605 , n489 , n13512 );
nand ( n13606 , n13605 , n12542 );
nand ( n13607 , n13604 , n13606 );
xor ( n13608 , n13601 , n13607 );
not ( n13609 , n12638 );
not ( n13610 , n13528 );
or ( n13611 , n13609 , n13610 );
not ( n13612 , n13114 );
not ( n13613 , n13612 );
and ( n13614 , n491 , n13613 );
not ( n13615 , n491 );
and ( n13616 , n13615 , n13612 );
nor ( n13617 , n13614 , n13616 );
nand ( n13618 , n13617 , n12595 );
nand ( n13619 , n13611 , n13618 );
and ( n13620 , n13608 , n13619 );
and ( n13621 , n13601 , n13607 );
or ( n13622 , n13620 , n13621 );
not ( n13623 , n493 );
not ( n13624 , n12532 );
or ( n13625 , n13623 , n13624 );
nand ( n13626 , n12531 , n12775 );
nand ( n13627 , n13625 , n13626 );
not ( n13628 , n13627 );
not ( n13629 , n12791 );
or ( n13630 , n13628 , n13629 );
or ( n13631 , n13539 , n12757 );
nand ( n13632 , n13630 , n13631 );
xor ( n13633 , n13622 , n13632 );
xor ( n13634 , n13513 , n13520 );
xor ( n13635 , n13634 , n13532 );
and ( n13636 , n13633 , n13635 );
and ( n13637 , n13622 , n13632 );
or ( n13638 , n13636 , n13637 );
and ( n13639 , n13590 , n13638 );
and ( n13640 , n13585 , n13589 );
or ( n13641 , n13639 , n13640 );
and ( n13642 , n13577 , n13641 );
and ( n13643 , n13574 , n13576 );
or ( n13644 , n13642 , n13643 );
xor ( n83397 , n13563 , n13644 );
not ( n83398 , n12462 );
not ( n13647 , n503 );
not ( n13648 , n82600 );
or ( n13649 , n13647 , n13648 );
not ( n13650 , n82600 );
nand ( n13651 , n13650 , n12457 );
nand ( n13652 , n13649 , n13651 );
not ( n13653 , n13652 );
or ( n13654 , n83398 , n13653 );
nand ( n13655 , n12855 , n12457 );
not ( n13656 , n13655 );
nand ( n13657 , n12852 , n503 );
not ( n13658 , n13657 );
or ( n13659 , n13656 , n13658 );
nand ( n13660 , n13659 , n504 );
nand ( n13661 , n13654 , n13660 );
and ( n13662 , n83397 , n13661 );
and ( n13663 , n13563 , n13644 );
or ( n13664 , n13662 , n13663 );
xor ( n13665 , n13495 , n13664 );
xor ( n13666 , n13349 , n13351 );
xor ( n13667 , n13666 , n13363 );
and ( n13668 , n13665 , n13667 );
and ( n13669 , n13495 , n13664 );
or ( n13670 , n13668 , n13669 );
xor ( n13671 , n13425 , n13670 );
xor ( n13672 , n13366 , n13404 );
xor ( n13673 , n13672 , n13407 );
and ( n13674 , n13671 , n13673 );
and ( n13675 , n13425 , n13670 );
or ( n13676 , n13674 , n13675 );
and ( n13677 , n83178 , n13676 );
and ( n13678 , n83176 , n13677 );
and ( n13679 , n13336 , n13416 );
nor ( n13680 , n13678 , n13679 );
not ( n13681 , n13680 );
xor ( n13682 , n13425 , n13670 );
xor ( n13683 , n13682 , n13673 );
xor ( n13684 , n13374 , n13398 );
xor ( n13685 , n13684 , n13401 );
xor ( n13686 , n13376 , n13387 );
xor ( n13687 , n13686 , n13395 );
xor ( n13688 , n13477 , n13479 );
xor ( n13689 , n13688 , n13492 );
xor ( n13690 , n13687 , n13689 );
xor ( n13691 , n83257 , n13549 );
xor ( n13692 , n13691 , n13560 );
not ( n13693 , n12843 );
not ( n13694 , n13488 );
or ( n13695 , n13693 , n13694 );
not ( n13696 , n501 );
not ( n13697 , n12483 );
or ( n13698 , n13696 , n13697 );
not ( n13699 , n12483 );
nand ( n13700 , n13699 , n12856 );
nand ( n83453 , n13698 , n13700 );
nand ( n13702 , n83453 , n12822 );
nand ( n13703 , n13695 , n13702 );
xor ( n13704 , n13692 , n13703 );
not ( n13705 , n13652 );
not ( n13706 , n504 );
or ( n13707 , n13705 , n13706 );
not ( n13708 , n503 );
not ( n13709 , n12671 );
or ( n13710 , n13708 , n13709 );
nand ( n13711 , n12674 , n12457 );
nand ( n13712 , n13710 , n13711 );
nand ( n13713 , n13712 , n12462 );
nand ( n13714 , n13707 , n13713 );
and ( n13715 , n13704 , n13714 );
and ( n13716 , n13692 , n13703 );
or ( n13717 , n13715 , n13716 );
and ( n13718 , n13690 , n13717 );
and ( n13719 , n13687 , n13689 );
or ( n13720 , n13718 , n13719 );
xor ( n13721 , n13685 , n13720 );
xor ( n13722 , n13495 , n13664 );
xor ( n13723 , n13722 , n13667 );
and ( n13724 , n13721 , n13723 );
and ( n13725 , n13685 , n13720 );
or ( n13726 , n13724 , n13725 );
nor ( n13727 , n13683 , n13726 );
not ( n13728 , n13727 );
not ( n13729 , n12758 );
not ( n13730 , n12735 );
not ( n13731 , n13730 );
and ( n13732 , n493 , n13731 );
not ( n13733 , n493 );
and ( n13734 , n13733 , n13524 );
nor ( n13735 , n13732 , n13734 );
not ( n13736 , n13735 );
or ( n13737 , n13729 , n13736 );
and ( n13738 , n493 , n13613 );
not ( n13739 , n493 );
and ( n13740 , n13739 , n13612 );
nor ( n13741 , n13738 , n13740 );
nand ( n13742 , n13741 , n12791 );
nand ( n13743 , n13737 , n13742 );
not ( n13744 , n13032 );
and ( n13745 , n495 , n12532 );
not ( n13746 , n495 );
and ( n13747 , n13746 , n12531 );
or ( n13748 , n13745 , n13747 );
not ( n13749 , n13748 );
or ( n13750 , n13744 , n13749 );
and ( n13751 , n495 , n12725 );
not ( n13752 , n495 );
and ( n13753 , n13752 , n13451 );
nor ( n13754 , n13751 , n13753 );
nand ( n13755 , n13754 , n12969 );
nand ( n13756 , n13750 , n13755 );
xor ( n13757 , n13743 , n13756 );
not ( n13758 , n12638 );
not ( n13759 , n491 );
not ( n13760 , n13441 );
not ( n13761 , n13760 );
or ( n13762 , n13759 , n13761 );
nand ( n13763 , n13441 , n12610 );
nand ( n13764 , n13762 , n13763 );
not ( n13765 , n13764 );
or ( n13766 , n13758 , n13765 );
buf ( n13767 , n13512 );
and ( n13768 , n491 , n13767 );
not ( n13769 , n491 );
not ( n13770 , n13512 );
and ( n13771 , n13769 , n13770 );
nor ( n13772 , n13768 , n13771 );
nand ( n13773 , n13772 , n12595 );
nand ( n13774 , n13766 , n13773 );
nand ( n13775 , n536 , n472 );
not ( n13776 , n13775 );
and ( n13777 , n489 , n13776 );
not ( n13778 , n12795 );
not ( n13779 , n489 );
not ( n13780 , n11786 );
not ( n13781 , n13595 );
or ( n13782 , n13780 , n13781 );
nand ( n83535 , n13596 , n13591 );
nand ( n13787 , n13782 , n83535 );
not ( n83537 , n13787 );
or ( n13789 , n13779 , n83537 );
or ( n13790 , n13787 , n489 );
nand ( n13791 , n13789 , n13790 );
not ( n13792 , n13791 );
or ( n13793 , n13778 , n13792 );
not ( n13794 , n11785 );
not ( n13795 , n81565 );
or ( n13796 , n13794 , n13795 );
or ( n13797 , n81565 , n11785 );
nand ( n13798 , n13796 , n13797 );
not ( n13799 , n13798 );
xor ( n13800 , n489 , n13799 );
nand ( n13801 , n13800 , n12542 );
nand ( n13802 , n13793 , n13801 );
xor ( n13803 , n13777 , n13802 );
or ( n13804 , n13776 , n490 );
nand ( n13805 , n13804 , n491 );
nand ( n13806 , n13776 , n490 );
and ( n83556 , n13805 , n13806 , n489 );
not ( n13811 , n12795 );
not ( n13812 , n13800 );
or ( n13813 , n13811 , n13812 );
xor ( n13814 , n489 , n13776 );
nand ( n13815 , n13814 , n12542 );
nand ( n13816 , n13813 , n13815 );
and ( n13817 , n83556 , n13816 );
xor ( n13818 , n13803 , n13817 );
xor ( n13819 , n13774 , n13818 );
xor ( n13820 , n83556 , n13816 );
not ( n13821 , n12638 );
not ( n13822 , n13772 );
or ( n13823 , n13821 , n13822 );
or ( n13824 , n13600 , n1693 );
nand ( n13825 , n13600 , n12610 );
nand ( n13826 , n13824 , n13825 );
nand ( n13827 , n12595 , n13826 );
nand ( n13828 , n13823 , n13827 );
xor ( n13829 , n13820 , n13828 );
nor ( n13830 , n13775 , n12539 );
not ( n13831 , n12638 );
not ( n13832 , n13826 );
or ( n13833 , n13831 , n13832 );
and ( n13834 , n491 , n13799 );
not ( n13835 , n491 );
and ( n13836 , n13835 , n13798 );
nor ( n13837 , n13834 , n13836 );
nand ( n13838 , n13837 , n12595 );
nand ( n13839 , n13833 , n13838 );
xor ( n13840 , n13830 , n13839 );
or ( n13841 , n13776 , n492 );
nand ( n13842 , n13841 , n493 );
and ( n13843 , n13776 , n492 );
nor ( n13844 , n13843 , n12610 );
and ( n13845 , n13842 , n13844 );
not ( n13846 , n12638 );
not ( n13847 , n13837 );
or ( n13848 , n13846 , n13847 );
or ( n13849 , n13775 , n491 );
or ( n13850 , n13776 , n12610 );
nand ( n13851 , n13849 , n13850 );
nand ( n13852 , n13851 , n12595 );
nand ( n13853 , n13848 , n13852 );
and ( n13854 , n13845 , n13853 );
and ( n13855 , n13840 , n13854 );
and ( n13856 , n13830 , n13839 );
or ( n13857 , n13855 , n13856 );
and ( n13858 , n13829 , n13857 );
and ( n13859 , n13820 , n13828 );
or ( n13860 , n13858 , n13859 );
xor ( n13861 , n13819 , n13860 );
and ( n13862 , n13757 , n13861 );
and ( n83609 , n13743 , n13756 );
or ( n83610 , n13862 , n83609 );
not ( n13865 , n12470 );
and ( n13866 , n497 , n12606 );
not ( n13867 , n497 );
and ( n13868 , n13867 , n12607 );
nor ( n13869 , n13866 , n13868 );
not ( n13870 , n13869 );
or ( n13871 , n13865 , n13870 );
not ( n13872 , n497 );
not ( n13873 , n12577 );
or ( n13874 , n13872 , n13873 );
nand ( n13875 , n12573 , n12486 );
nand ( n13876 , n13874 , n13875 );
nand ( n13877 , n12517 , n13876 );
nand ( n13878 , n13871 , n13877 );
xor ( n13879 , n83610 , n13878 );
not ( n13880 , n12650 );
not ( n13881 , n499 );
not ( n13882 , n12900 );
or ( n13883 , n13881 , n13882 );
nand ( n13884 , n12774 , n12467 );
nand ( n13885 , n13883 , n13884 );
not ( n13886 , n13885 );
or ( n13887 , n13880 , n13886 );
not ( n13888 , n499 );
not ( n13889 , n12629 );
or ( n13890 , n13888 , n13889 );
nand ( n13891 , n12467 , n12628 );
nand ( n13892 , n13890 , n13891 );
nand ( n13893 , n13892 , n12702 );
nand ( n13894 , n13887 , n13893 );
xor ( n13895 , n13879 , n13894 );
not ( n13896 , n12462 );
not ( n13897 , n503 );
not ( n13898 , n13009 );
or ( n13899 , n13897 , n13898 );
nand ( n13900 , n13008 , n12423 );
nand ( n13901 , n13899 , n13900 );
not ( n13902 , n13901 );
or ( n13903 , n13896 , n13902 );
and ( n13904 , n12506 , n503 );
not ( n13905 , n12506 );
and ( n13906 , n13905 , n12457 );
or ( n13907 , n13904 , n13906 );
nand ( n13908 , n13907 , n504 );
nand ( n13909 , n13903 , n13908 );
xor ( n13910 , n13895 , n13909 );
xor ( n13911 , n13743 , n13756 );
xor ( n13912 , n13911 , n13861 );
not ( n13913 , n12758 );
and ( n13914 , n12775 , n13760 );
not ( n13915 , n12775 );
and ( n13916 , n13915 , n13441 );
nor ( n13917 , n13914 , n13916 );
not ( n13918 , n13917 );
or ( n13919 , n13913 , n13918 );
and ( n13920 , n493 , n13512 );
not ( n13921 , n493 );
and ( n13922 , n13921 , n13770 );
nor ( n13923 , n13920 , n13922 );
nand ( n13924 , n13923 , n12791 );
nand ( n13925 , n13919 , n13924 );
xor ( n13926 , n13830 , n13839 );
xor ( n13927 , n13926 , n13854 );
xor ( n13928 , n13925 , n13927 );
xor ( n13929 , n13845 , n13853 );
not ( n13930 , n12758 );
not ( n13931 , n13923 );
or ( n13932 , n13930 , n13931 );
not ( n13933 , n493 );
not ( n13934 , n13787 );
or ( n13935 , n13933 , n13934 );
or ( n13936 , n13787 , n493 );
nand ( n13937 , n13935 , n13936 );
nand ( n13938 , n13937 , n12791 );
nand ( n13939 , n13932 , n13938 );
xor ( n83686 , n13929 , n13939 );
nor ( n13941 , n12593 , n13775 );
not ( n13942 , n12756 );
and ( n13943 , n493 , n13799 );
not ( n13944 , n493 );
and ( n13945 , n13944 , n13798 );
nor ( n13946 , n13943 , n13945 );
not ( n13947 , n13946 );
or ( n13948 , n13942 , n13947 );
or ( n13949 , n13775 , n493 );
or ( n13950 , n13776 , n12775 );
nand ( n13951 , n13949 , n13950 );
nand ( n13952 , n13951 , n12791 );
nand ( n13953 , n13948 , n13952 );
or ( n13954 , n13776 , n494 );
nand ( n13955 , n13954 , n495 );
and ( n13956 , n13776 , n494 );
nor ( n13957 , n13956 , n12775 );
nand ( n13958 , n13955 , n13957 );
not ( n13959 , n13958 );
and ( n13960 , n13953 , n13959 );
xor ( n13961 , n13941 , n13960 );
not ( n13962 , n12758 );
not ( n13963 , n13937 );
or ( n13964 , n13962 , n13963 );
nand ( n13965 , n13946 , n12791 );
nand ( n13966 , n13964 , n13965 );
and ( n13967 , n13961 , n13966 );
or ( n13969 , n13967 , C0 );
and ( n13970 , n83686 , n13969 );
and ( n13971 , n13929 , n13939 );
or ( n13972 , n13970 , n13971 );
and ( n13973 , n13928 , n13972 );
and ( n13974 , n13925 , n13927 );
or ( n13975 , n13973 , n13974 );
not ( n13976 , n12470 );
not ( n13977 , n497 );
not ( n13978 , n12556 );
or ( n13979 , n13977 , n13978 );
nand ( n13980 , n12559 , n12486 );
nand ( n13981 , n13979 , n13980 );
not ( n13982 , n13981 );
or ( n13983 , n13976 , n13982 );
and ( n13984 , n12531 , n12486 );
not ( n13985 , n12531 );
and ( n13986 , n13985 , n497 );
or ( n13987 , n13984 , n13986 );
nand ( n13988 , n13987 , n12517 );
nand ( n13989 , n13983 , n13988 );
xor ( n13990 , n13975 , n13989 );
not ( n13991 , n12758 );
not ( n13992 , n13741 );
or ( n13993 , n13991 , n13992 );
nand ( n13994 , n13917 , n12791 );
nand ( n13995 , n13993 , n13994 );
xor ( n13996 , n13820 , n13828 );
xor ( n13997 , n13996 , n13857 );
xor ( n13998 , n13995 , n13997 );
not ( n13999 , n13032 );
not ( n14000 , n13754 );
or ( n14001 , n13999 , n14000 );
and ( n14002 , n495 , n13730 );
not ( n14003 , n495 );
and ( n14004 , n14003 , n13731 );
or ( n14005 , n14002 , n14004 );
nand ( n14006 , n14005 , n12969 );
nand ( n14007 , n14001 , n14006 );
xor ( n14008 , n13998 , n14007 );
and ( n14009 , n13990 , n14008 );
and ( n14010 , n13975 , n13989 );
or ( n83756 , n14009 , n14010 );
xor ( n83757 , n13912 , n83756 );
not ( n14013 , n12843 );
not ( n14014 , n501 );
not ( n14015 , n12950 );
or ( n14016 , n14014 , n14015 );
nand ( n14017 , n13080 , n12856 );
nand ( n14018 , n14016 , n14017 );
not ( n14019 , n14018 );
or ( n14020 , n14013 , n14019 );
not ( n14021 , n501 );
not ( n14022 , n12900 );
or ( n14023 , n14021 , n14022 );
nand ( n14024 , n12774 , n12856 );
nand ( n14025 , n14023 , n14024 );
nand ( n14026 , n14025 , n12821 );
nand ( n14027 , n14020 , n14026 );
and ( n14028 , n83757 , n14027 );
and ( n14029 , n13912 , n83756 );
or ( n14030 , n14028 , n14029 );
and ( n14031 , n13910 , n14030 );
and ( n14032 , n13895 , n13909 );
or ( n14033 , n14031 , n14032 );
not ( n14034 , n12638 );
not ( n14035 , n13617 );
or ( n14036 , n14034 , n14035 );
nand ( n14037 , n13764 , n12595 );
nand ( n14038 , n14036 , n14037 );
and ( n14039 , n489 , n13799 );
not ( n14040 , n12542 );
not ( n14041 , n13791 );
or ( n14042 , n14040 , n14041 );
nand ( n14043 , n13605 , n12795 );
nand ( n14044 , n14042 , n14043 );
xor ( n14045 , n14039 , n14044 );
xor ( n14046 , n13777 , n13802 );
and ( n14047 , n14046 , n13817 );
and ( n14048 , n13777 , n13802 );
or ( n83794 , n14047 , n14048 );
xor ( n14050 , n14045 , n83794 );
xor ( n14051 , n14038 , n14050 );
not ( n14052 , n12791 );
not ( n14053 , n13735 );
or ( n14054 , n14052 , n14053 );
not ( n14055 , n493 );
not ( n14056 , n13451 );
or ( n14057 , n14055 , n14056 );
nand ( n14058 , n12725 , n12775 );
nand ( n14059 , n14057 , n14058 );
nand ( n14060 , n14059 , n12758 );
nand ( n14061 , n14054 , n14060 );
and ( n14062 , n14051 , n14061 );
and ( n14063 , n14038 , n14050 );
or ( n14064 , n14062 , n14063 );
not ( n14065 , n13032 );
and ( n14066 , n495 , n12577 );
not ( n14067 , n495 );
and ( n14068 , n14067 , n12573 );
or ( n14069 , n14066 , n14068 );
not ( n14070 , n14069 );
or ( n14071 , n14065 , n14070 );
not ( n14072 , n495 );
not ( n14073 , n12559 );
not ( n14074 , n14073 );
or ( n14075 , n14072 , n14074 );
not ( n14076 , n495 );
not ( n14077 , n12556 );
nand ( n14078 , n14076 , n14077 );
nand ( n14079 , n14075 , n14078 );
nand ( n14080 , n14079 , n12969 );
nand ( n14081 , n14071 , n14080 );
xor ( n14082 , n14064 , n14081 );
not ( n14083 , n12517 );
not ( n14084 , n13869 );
or ( n14085 , n14083 , n14084 );
not ( n14086 , n497 );
not ( n14087 , n12629 );
or ( n14088 , n14086 , n14087 );
not ( n14089 , n12783 );
nand ( n14090 , n14089 , n12486 );
nand ( n14091 , n14088 , n14090 );
nand ( n14092 , n14091 , n12470 );
nand ( n14093 , n14085 , n14092 );
xor ( n14094 , n14082 , n14093 );
not ( n14095 , n12821 );
not ( n14096 , n501 );
not ( n14097 , n12981 );
or ( n14098 , n14096 , n14097 );
not ( n14099 , n12981 );
nand ( n14100 , n14099 , n12856 );
nand ( n14101 , n14098 , n14100 );
not ( n14102 , n14101 );
or ( n14103 , n14095 , n14102 );
not ( n14104 , n501 );
not ( n14105 , n13009 );
or ( n14106 , n14104 , n14105 );
nand ( n14107 , n13008 , n12856 );
nand ( n14108 , n14106 , n14107 );
nand ( n14109 , n14108 , n12843 );
nand ( n14110 , n14103 , n14109 );
xor ( n14111 , n14094 , n14110 );
not ( n14112 , n504 );
not ( n14113 , n503 );
not ( n14114 , n12483 );
or ( n14115 , n14113 , n14114 );
nand ( n14116 , n13699 , n12457 );
nand ( n14117 , n14115 , n14116 );
not ( n14118 , n14117 );
or ( n14119 , n14112 , n14118 );
nand ( n14120 , n13907 , n12462 );
nand ( n14121 , n14119 , n14120 );
xor ( n14122 , n14111 , n14121 );
xor ( n14123 , n14033 , n14122 );
xor ( n14124 , n83610 , n13878 );
and ( n14125 , n14124 , n13894 );
and ( n14126 , n83610 , n13878 );
or ( n14127 , n14125 , n14126 );
xor ( n14128 , n14039 , n14044 );
and ( n83874 , n14128 , n83794 );
and ( n14133 , n14039 , n14044 );
or ( n83876 , n83874 , n14133 );
not ( n14135 , n12758 );
not ( n14136 , n13627 );
or ( n14137 , n14135 , n14136 );
nand ( n14138 , n14059 , n12791 );
nand ( n14139 , n14137 , n14138 );
xor ( n14140 , n83876 , n14139 );
xor ( n14141 , n13601 , n13607 );
xor ( n14142 , n14141 , n13619 );
xor ( n14143 , n14140 , n14142 );
not ( n14144 , n12702 );
not ( n14145 , n13885 );
or ( n14146 , n14144 , n14145 );
and ( n14147 , n12949 , n12467 );
not ( n14148 , n12949 );
and ( n14149 , n14148 , n499 );
or ( n14150 , n14147 , n14149 );
nand ( n14151 , n14150 , n12648 );
nand ( n14152 , n14146 , n14151 );
xor ( n14153 , n14143 , n14152 );
xor ( n14154 , n13774 , n13818 );
and ( n14155 , n14154 , n13860 );
and ( n14156 , n13774 , n13818 );
or ( n14157 , n14155 , n14156 );
not ( n83900 , n13032 );
not ( n14162 , n14079 );
or ( n14163 , n83900 , n14162 );
nand ( n14164 , n13748 , n12969 );
nand ( n14165 , n14163 , n14164 );
xor ( n14166 , n14157 , n14165 );
xor ( n14167 , n14038 , n14050 );
xor ( n14168 , n14167 , n14061 );
and ( n14169 , n14166 , n14168 );
and ( n14170 , n14157 , n14165 );
or ( n14171 , n14169 , n14170 );
xor ( n14172 , n14153 , n14171 );
xor ( n14173 , n14127 , n14172 );
xor ( n14174 , n14157 , n14165 );
xor ( n14175 , n14174 , n14168 );
not ( n14176 , n12517 );
not ( n14177 , n13981 );
or ( n14178 , n14176 , n14177 );
nand ( n14179 , n13876 , n12470 );
nand ( n14180 , n14178 , n14179 );
xor ( n14181 , n13995 , n13997 );
and ( n14182 , n14181 , n14007 );
and ( n14183 , n13995 , n13997 );
or ( n14184 , n14182 , n14183 );
xor ( n14185 , n14180 , n14184 );
not ( n14186 , n12702 );
not ( n14187 , n499 );
not ( n14188 , n13100 );
or ( n14189 , n14187 , n14188 );
nand ( n14190 , n12467 , n12606 );
nand ( n14191 , n14189 , n14190 );
not ( n14192 , n14191 );
or ( n14193 , n14186 , n14192 );
nand ( n14194 , n13892 , n12648 );
nand ( n14195 , n14193 , n14194 );
and ( n14196 , n14185 , n14195 );
and ( n14197 , n14180 , n14184 );
or ( n14198 , n14196 , n14197 );
xor ( n14199 , n14175 , n14198 );
not ( n14200 , n12843 );
not ( n14201 , n14101 );
or ( n14202 , n14200 , n14201 );
nand ( n14203 , n14018 , n12821 );
nand ( n14204 , n14202 , n14203 );
and ( n14205 , n14199 , n14204 );
and ( n14206 , n14175 , n14198 );
or ( n14207 , n14205 , n14206 );
xor ( n14208 , n14173 , n14207 );
xor ( n14209 , n14123 , n14208 );
xor ( n83949 , n14175 , n14198 );
xor ( n83950 , n83949 , n14204 );
xor ( n14212 , n14180 , n14184 );
xor ( n14213 , n14212 , n14195 );
not ( n14214 , n12462 );
not ( n14215 , n503 );
not ( n14216 , n13378 );
or ( n14217 , n14215 , n14216 );
not ( n14218 , n503 );
nand ( n14219 , n14218 , n14099 );
nand ( n14220 , n14217 , n14219 );
not ( n14221 , n14220 );
or ( n14222 , n14214 , n14221 );
nand ( n14223 , n13901 , n504 );
nand ( n14224 , n14222 , n14223 );
xor ( n14225 , n14213 , n14224 );
not ( n14226 , n13032 );
not ( n14227 , n14005 );
or ( n14228 , n14226 , n14227 );
and ( n14229 , n495 , n13114 );
not ( n14230 , n495 );
and ( n14231 , n14230 , n13612 );
nor ( n14232 , n14229 , n14231 );
nand ( n14233 , n14232 , n12969 );
nand ( n14234 , n14228 , n14233 );
not ( n14235 , n12470 );
not ( n14236 , n13987 );
or ( n14237 , n14235 , n14236 );
not ( n14238 , n497 );
not ( n14239 , n13451 );
or ( n14240 , n14238 , n14239 );
nand ( n14241 , n12725 , n12486 );
nand ( n14242 , n14240 , n14241 );
nand ( n14243 , n14242 , n12517 );
nand ( n14244 , n14237 , n14243 );
xor ( n14245 , n14234 , n14244 );
xor ( n14246 , n13925 , n13927 );
xor ( n14247 , n14246 , n13972 );
and ( n14248 , n14245 , n14247 );
and ( n14249 , n14234 , n14244 );
or ( n14250 , n14248 , n14249 );
not ( n14251 , n12650 );
not ( n14252 , n14191 );
or ( n14253 , n14251 , n14252 );
not ( n14254 , n499 );
not ( n14255 , n12577 );
or ( n14256 , n14254 , n14255 );
nand ( n14257 , n12573 , n12467 );
nand ( n14258 , n14256 , n14257 );
nand ( n14259 , n14258 , n12702 );
nand ( n14260 , n14253 , n14259 );
xor ( n14261 , n14250 , n14260 );
not ( n14262 , n12843 );
not ( n14263 , n14025 );
or ( n14264 , n14262 , n14263 );
and ( n14265 , n12629 , n501 );
not ( n14266 , n12629 );
and ( n14267 , n14266 , n12856 );
or ( n14268 , n14265 , n14267 );
nand ( n14269 , n14268 , n12821 );
nand ( n14270 , n14264 , n14269 );
and ( n14271 , n14261 , n14270 );
and ( n14272 , n14250 , n14260 );
or ( n14273 , n14271 , n14272 );
and ( n14274 , n14225 , n14273 );
and ( n14275 , n14213 , n14224 );
or ( n14276 , n14274 , n14275 );
xor ( n14277 , n83950 , n14276 );
xor ( n14278 , n13895 , n13909 );
xor ( n14279 , n14278 , n14030 );
and ( n14280 , n14277 , n14279 );
and ( n14281 , n83950 , n14276 );
or ( n14282 , n14280 , n14281 );
or ( n14283 , n14209 , n14282 );
not ( n14284 , n14283 );
xor ( n14285 , n83950 , n14276 );
xor ( n14286 , n14285 , n14279 );
xor ( n84026 , n13912 , n83756 );
xor ( n14288 , n84026 , n14027 );
xor ( n14289 , n13975 , n13989 );
xor ( n14290 , n14289 , n14008 );
not ( n14291 , n13032 );
not ( n14292 , n14232 );
or ( n14293 , n14291 , n14292 );
and ( n14294 , n495 , n13441 );
not ( n14295 , n495 );
and ( n14296 , n14295 , n13760 );
nor ( n14297 , n14294 , n14296 );
nand ( n14298 , n14297 , n12969 );
nand ( n14299 , n14293 , n14298 );
xor ( n14300 , n13929 , n13939 );
xor ( n14301 , n14300 , n13969 );
xor ( n14302 , n14299 , n14301 );
not ( n14303 , n12470 );
not ( n14304 , n14242 );
or ( n14305 , n14303 , n14304 );
buf ( n14306 , n12735 );
and ( n14307 , n497 , n14306 );
not ( n14308 , n497 );
and ( n14309 , n14308 , n13730 );
nor ( n14310 , n14307 , n14309 );
nand ( n14311 , n14310 , n12516 );
nand ( n14312 , n14305 , n14311 );
and ( n14313 , n14302 , n14312 );
and ( n14314 , n14299 , n14301 );
or ( n14315 , n14313 , n14314 );
not ( n14316 , n12702 );
and ( n14317 , n499 , n14077 );
not ( n14318 , n499 );
and ( n14319 , n14318 , n12556 );
nor ( n14320 , n14317 , n14319 );
not ( n14321 , n14320 );
or ( n14322 , n14316 , n14321 );
nand ( n14323 , n14258 , n12648 );
nand ( n14324 , n14322 , n14323 );
xor ( n14325 , n14315 , n14324 );
xor ( n14326 , n14234 , n14244 );
xor ( n14327 , n14326 , n14247 );
and ( n14328 , n14325 , n14327 );
and ( n14329 , n14315 , n14324 );
or ( n14330 , n14328 , n14329 );
xor ( n14331 , n14290 , n14330 );
not ( n14332 , n12462 );
not ( n14333 , n503 );
not ( n14334 , n82837 );
or ( n14335 , n14333 , n14334 );
nand ( n14336 , n13080 , n12423 );
nand ( n14337 , n14335 , n14336 );
not ( n14338 , n14337 );
or ( n14339 , n14332 , n14338 );
nand ( n14340 , n14220 , n504 );
nand ( n14341 , n14339 , n14340 );
and ( n14342 , n14331 , n14341 );
and ( n14343 , n14290 , n14330 );
or ( n14344 , n14342 , n14343 );
xor ( n14345 , n14288 , n14344 );
xor ( n14346 , n14213 , n14224 );
xor ( n14347 , n14346 , n14273 );
and ( n14348 , n14345 , n14347 );
and ( n14349 , n14288 , n14344 );
or ( n14350 , n14348 , n14349 );
or ( n14351 , n14286 , n14350 );
not ( n14352 , n14351 );
xor ( n14353 , n14288 , n14344 );
xor ( n14354 , n14353 , n14347 );
not ( n14355 , n14354 );
not ( n14356 , n12821 );
and ( n14357 , n501 , n12606 );
not ( n14358 , n501 );
and ( n14359 , n14358 , n12607 );
nor ( n14360 , n14357 , n14359 );
not ( n14361 , n14360 );
or ( n14362 , n14356 , n14361 );
nand ( n14363 , n14268 , n12843 );
nand ( n14364 , n14362 , n14363 );
not ( n14365 , n12969 );
and ( n14366 , n495 , n13767 );
not ( n14367 , n495 );
and ( n14368 , n14367 , n13770 );
nor ( n14369 , n14366 , n14368 );
not ( n14370 , n14369 );
or ( n14371 , n14365 , n14370 );
nand ( n14372 , n14297 , n13032 );
nand ( n14373 , n14371 , n14372 );
xor ( n14374 , n13941 , n13960 );
xor ( n84114 , n14374 , n13966 );
xor ( n14376 , n14373 , n84114 );
and ( n14377 , n13953 , n13959 );
not ( n14378 , n13953 );
and ( n14379 , n14378 , n13958 );
nor ( n14380 , n14377 , n14379 );
not ( n14381 , n13032 );
not ( n14382 , n14369 );
or ( n14383 , n14381 , n14382 );
not ( n14384 , n495 );
not ( n14385 , n13787 );
or ( n14386 , n14384 , n14385 );
or ( n14387 , n13787 , n495 );
nand ( n14388 , n14386 , n14387 );
nand ( n14389 , n14388 , n12969 );
nand ( n14390 , n14383 , n14389 );
xor ( n14391 , n14380 , n14390 );
nor ( n14392 , n13775 , n12757 );
not ( n14393 , n13032 );
not ( n14394 , n14388 );
or ( n14395 , n14393 , n14394 );
and ( n14396 , n495 , n13799 );
not ( n14397 , n495 );
and ( n14398 , n14397 , n13798 );
nor ( n14399 , n14396 , n14398 );
nand ( n14400 , n14399 , n12969 );
nand ( n14401 , n14395 , n14400 );
xor ( n14402 , n14392 , n14401 );
or ( n14403 , n13776 , n496 );
nand ( n14404 , n14403 , n497 );
and ( n14405 , n13776 , n496 );
nor ( n14406 , n14405 , n3325 );
and ( n14407 , n14404 , n14406 );
not ( n14408 , n12969 );
and ( n14409 , n495 , n13776 );
not ( n14410 , n495 );
and ( n14411 , n14410 , n13775 );
nor ( n14412 , n14409 , n14411 );
not ( n14413 , n14412 );
or ( n14414 , n14408 , n14413 );
nand ( n14415 , n14399 , n13032 );
nand ( n14416 , n14414 , n14415 );
and ( n14417 , n14407 , n14416 );
and ( n14418 , n14402 , n14417 );
and ( n14419 , n14392 , n14401 );
or ( n14420 , n14418 , n14419 );
and ( n14421 , n14391 , n14420 );
and ( n14422 , n14380 , n14390 );
or ( n14423 , n14421 , n14422 );
and ( n14424 , n14376 , n14423 );
and ( n14425 , n14373 , n84114 );
or ( n14426 , n14424 , n14425 );
xor ( n14427 , n14299 , n14301 );
xor ( n14428 , n14427 , n14312 );
xor ( n14429 , n14426 , n14428 );
not ( n14430 , n14320 );
or ( n14431 , n14430 , n12649 );
and ( n14432 , n12531 , n12467 );
not ( n14433 , n12531 );
and ( n14434 , n14433 , n499 );
or ( n14435 , n14432 , n14434 );
nand ( n14436 , n14435 , n12702 );
nand ( n14437 , n14431 , n14436 );
and ( n14438 , n14429 , n14437 );
and ( n14439 , n14426 , n14428 );
or ( n14440 , n14438 , n14439 );
xor ( n14441 , n14364 , n14440 );
not ( n14442 , n12462 );
not ( n14443 , n503 );
not ( n14444 , n12900 );
or ( n14445 , n14443 , n14444 );
nand ( n14446 , n12774 , n12423 );
nand ( n14447 , n14445 , n14446 );
not ( n14448 , n14447 );
or ( n14449 , n14442 , n14448 );
nand ( n14450 , n14337 , n504 );
nand ( n14451 , n14449 , n14450 );
and ( n14452 , n14441 , n14451 );
and ( n14453 , n14364 , n14440 );
or ( n14454 , n14452 , n14453 );
xor ( n84194 , n14250 , n14260 );
xor ( n14459 , n84194 , n14270 );
xor ( n84196 , n14454 , n14459 );
xor ( n14461 , n14290 , n14330 );
xor ( n14462 , n14461 , n14341 );
and ( n14463 , n84196 , n14462 );
and ( n14464 , n14454 , n14459 );
or ( n14465 , n14463 , n14464 );
not ( n14466 , n14465 );
and ( n14467 , n14355 , n14466 );
xor ( n14468 , n14454 , n14459 );
xor ( n14469 , n14468 , n14462 );
xor ( n14470 , n14315 , n14324 );
xor ( n14471 , n14470 , n14327 );
not ( n14472 , n12470 );
not ( n14473 , n14310 );
or ( n14474 , n14472 , n14473 );
and ( n14475 , n497 , n13613 );
not ( n14476 , n497 );
and ( n14477 , n14476 , n13612 );
nor ( n14478 , n14475 , n14477 );
nand ( n14479 , n14478 , n12516 );
nand ( n14480 , n14474 , n14479 );
not ( n14481 , n12648 );
not ( n14482 , n14435 );
or ( n14483 , n14481 , n14482 );
not ( n14484 , n499 );
not ( n14485 , n13451 );
or ( n84222 , n14484 , n14485 );
nand ( n14490 , n12725 , n12467 );
nand ( n14491 , n84222 , n14490 );
nand ( n14492 , n14491 , n12702 );
nand ( n14493 , n14483 , n14492 );
xor ( n14494 , n14480 , n14493 );
xor ( n14495 , n14373 , n84114 );
xor ( n14496 , n14495 , n14423 );
and ( n14497 , n14494 , n14496 );
and ( n14498 , n14480 , n14493 );
or ( n14499 , n14497 , n14498 );
not ( n14500 , n12843 );
not ( n14501 , n14360 );
or ( n14502 , n14500 , n14501 );
not ( n14503 , n501 );
not ( n14504 , n12577 );
or ( n14505 , n14503 , n14504 );
nand ( n14506 , n12573 , n12856 );
nand ( n14507 , n14505 , n14506 );
nand ( n14508 , n14507 , n12822 );
nand ( n14509 , n14502 , n14508 );
xor ( n14510 , n14499 , n14509 );
not ( n14511 , n504 );
not ( n14512 , n14447 );
or ( n14513 , n14511 , n14512 );
not ( n14514 , n503 );
not ( n14515 , n12783 );
or ( n14516 , n14514 , n14515 );
nand ( n14517 , n12457 , n12628 );
nand ( n14518 , n14516 , n14517 );
nand ( n14519 , n14518 , n12462 );
nand ( n14520 , n14513 , n14519 );
and ( n14521 , n14510 , n14520 );
and ( n14522 , n14499 , n14509 );
or ( n14523 , n14521 , n14522 );
xor ( n14524 , n14471 , n14523 );
xor ( n14525 , n14364 , n14440 );
xor ( n14526 , n14525 , n14451 );
and ( n14527 , n14524 , n14526 );
and ( n14528 , n14471 , n14523 );
or ( n14529 , n14527 , n14528 );
nor ( n14530 , n14469 , n14529 );
nor ( n14531 , n14467 , n14530 );
not ( n14532 , n14531 );
xor ( n14533 , n14471 , n14523 );
xor ( n14534 , n14533 , n14526 );
not ( n14535 , n14534 );
xor ( n14536 , n14426 , n14428 );
xor ( n14537 , n14536 , n14437 );
not ( n14538 , n12843 );
not ( n14539 , n14507 );
or ( n14540 , n14538 , n14539 );
and ( n14541 , n501 , n12559 );
not ( n14542 , n501 );
and ( n14543 , n14542 , n12556 );
nor ( n14544 , n14541 , n14543 );
nand ( n14545 , n14544 , n12821 );
nand ( n14546 , n14540 , n14545 );
not ( n14547 , n12516 );
and ( n14548 , n497 , n13441 );
not ( n14549 , n497 );
and ( n14550 , n14549 , n13760 );
nor ( n14551 , n14548 , n14550 );
not ( n14552 , n14551 );
or ( n14553 , n14547 , n14552 );
nand ( n14554 , n14478 , n12470 );
nand ( n14555 , n14553 , n14554 );
xor ( n84289 , n14380 , n14390 );
xor ( n84290 , n84289 , n14420 );
xor ( n14558 , n14555 , n84290 );
not ( n14559 , n12648 );
not ( n14560 , n14491 );
or ( n14561 , n14559 , n14560 );
and ( n14562 , n499 , n13731 );
not ( n14563 , n499 );
and ( n14564 , n14563 , n13524 );
nor ( n14565 , n14562 , n14564 );
nand ( n14566 , n14565 , n12702 );
nand ( n14567 , n14561 , n14566 );
and ( n14568 , n14558 , n14567 );
and ( n14569 , n14555 , n84290 );
or ( n14570 , n14568 , n14569 );
xor ( n14571 , n14546 , n14570 );
not ( n14572 , n504 );
not ( n14573 , n14518 );
or ( n14574 , n14572 , n14573 );
and ( n14575 , n503 , n12606 );
not ( n14576 , n503 );
and ( n14577 , n14576 , n12607 );
nor ( n14578 , n14575 , n14577 );
nand ( n14579 , n14578 , n12462 );
nand ( n14580 , n14574 , n14579 );
and ( n14581 , n14571 , n14580 );
and ( n14582 , n14546 , n14570 );
or ( n14583 , n14581 , n14582 );
xor ( n14584 , n14537 , n14583 );
xor ( n14585 , n14499 , n14509 );
xor ( n14586 , n14585 , n14520 );
and ( n14587 , n14584 , n14586 );
and ( n14588 , n14537 , n14583 );
or ( n14589 , n14587 , n14588 );
not ( n14590 , n14589 );
and ( n14591 , n14535 , n14590 );
xor ( n14592 , n14537 , n14583 );
xor ( n14593 , n14592 , n14586 );
xor ( n14594 , n14480 , n14493 );
xor ( n14595 , n14594 , n14496 );
not ( n14596 , n12470 );
not ( n14597 , n14551 );
or ( n14598 , n14596 , n14597 );
not ( n14599 , n497 );
not ( n14600 , n13770 );
or ( n14601 , n14599 , n14600 );
nand ( n14602 , n13767 , n12486 );
nand ( n14603 , n14601 , n14602 );
nand ( n14604 , n14603 , n12516 );
nand ( n14605 , n14598 , n14604 );
xor ( n14606 , n14392 , n14401 );
xor ( n14607 , n14606 , n14417 );
xor ( n14608 , n14605 , n14607 );
xor ( n84342 , n14407 , n14416 );
not ( n14610 , n12470 );
not ( n14611 , n14603 );
or ( n14612 , n14610 , n14611 );
not ( n14613 , n12486 );
not ( n14614 , n13600 );
or ( n14615 , n14613 , n14614 );
nand ( n14616 , n13787 , n497 );
nand ( n14617 , n14615 , n14616 );
nand ( n14618 , n14617 , n12516 );
nand ( n14619 , n14612 , n14618 );
xor ( n14620 , n84342 , n14619 );
nor ( n14621 , n13775 , n12965 );
not ( n14622 , n12470 );
not ( n14623 , n14617 );
or ( n14624 , n14622 , n14623 );
or ( n14625 , n13799 , n497 );
nand ( n14626 , n13799 , n497 );
nand ( n14627 , n14625 , n14626 );
not ( n14628 , n14627 );
nand ( n14629 , n14628 , n12516 );
nand ( n14630 , n14624 , n14629 );
xor ( n14631 , n14621 , n14630 );
or ( n14632 , n13776 , n498 );
nand ( n14633 , n14632 , n499 );
and ( n14634 , n13776 , n498 );
nor ( n14635 , n14634 , n12486 );
and ( n14636 , n14633 , n14635 );
not ( n14637 , n12516 );
or ( n14638 , n13775 , n497 );
or ( n14639 , n13776 , n12486 );
nand ( n14640 , n14638 , n14639 );
not ( n14641 , n14640 );
or ( n14642 , n14637 , n14641 );
or ( n14643 , n14627 , n12469 );
nand ( n14644 , n14642 , n14643 );
and ( n14645 , n14636 , n14644 );
and ( n14646 , n14631 , n14645 );
and ( n14647 , n14621 , n14630 );
or ( n14648 , n14646 , n14647 );
and ( n14649 , n14620 , n14648 );
and ( n14650 , n84342 , n14619 );
or ( n14651 , n14649 , n14650 );
and ( n14652 , n14608 , n14651 );
and ( n14653 , n14605 , n14607 );
or ( n14654 , n14652 , n14653 );
xor ( n14655 , n14555 , n84290 );
xor ( n14656 , n14655 , n14567 );
xor ( n14657 , n14654 , n14656 );
not ( n14658 , n12822 );
xor ( n14659 , n501 , n12531 );
not ( n14660 , n14659 );
or ( n14661 , n14658 , n14660 );
nand ( n14662 , n14544 , n12843 );
nand ( n14663 , n14661 , n14662 );
and ( n14664 , n14657 , n14663 );
and ( n14665 , n14654 , n14656 );
or ( n14666 , n14664 , n14665 );
xor ( n14667 , n14595 , n14666 );
xor ( n14668 , n14546 , n14570 );
xor ( n14669 , n14668 , n14580 );
and ( n14670 , n14667 , n14669 );
and ( n14671 , n14595 , n14666 );
or ( n14672 , n14670 , n14671 );
nor ( n14673 , n14593 , n14672 );
nor ( n14674 , n14591 , n14673 );
not ( n14675 , n14674 );
not ( n14676 , n12702 );
and ( n14677 , n499 , n13612 );
not ( n14678 , n499 );
and ( n14679 , n14678 , n13114 );
or ( n14680 , n14677 , n14679 );
not ( n14681 , n14680 );
or ( n14682 , n14676 , n14681 );
nand ( n14683 , n14565 , n12648 );
nand ( n14684 , n14682 , n14683 );
xor ( n14685 , n14605 , n14607 );
xor ( n14686 , n14685 , n14651 );
xor ( n14687 , n14684 , n14686 );
not ( n14688 , n12843 );
not ( n14689 , n14659 );
or ( n14690 , n14688 , n14689 );
and ( n14691 , n12821 , n12856 );
and ( n84425 , n12725 , n14691 );
not ( n14693 , n12725 );
not ( n14694 , n12423 );
nor ( n14695 , n14694 , n12813 );
and ( n14696 , n14693 , n14695 );
nor ( n14697 , n84425 , n14696 );
nand ( n14698 , n14690 , n14697 );
and ( n14699 , n14687 , n14698 );
and ( n14700 , n14684 , n14686 );
or ( n14701 , n14699 , n14700 );
not ( n14702 , n504 );
not ( n14703 , n14578 );
or ( n14704 , n14702 , n14703 );
and ( n14705 , n503 , n12573 );
not ( n14706 , n503 );
and ( n14707 , n14706 , n12577 );
nor ( n14708 , n14705 , n14707 );
nand ( n14709 , n14708 , n12462 );
nand ( n14710 , n14704 , n14709 );
xor ( n14711 , n14701 , n14710 );
xor ( n14712 , n14654 , n14656 );
xor ( n14713 , n14712 , n14663 );
and ( n14714 , n14711 , n14713 );
and ( n14715 , n14701 , n14710 );
or ( n14716 , n14714 , n14715 );
not ( n14717 , n14716 );
xor ( n14718 , n14595 , n14666 );
xor ( n14719 , n14718 , n14669 );
not ( n14720 , n14719 );
nand ( n14721 , n14717 , n14720 );
not ( n14722 , n14721 );
xor ( n14723 , n14701 , n14710 );
xor ( n14724 , n14723 , n14713 );
not ( n14725 , n12462 );
not ( n14726 , n503 );
not ( n14727 , n12556 );
or ( n14728 , n14726 , n14727 );
nand ( n14729 , n12559 , n12423 );
nand ( n14730 , n14728 , n14729 );
not ( n14731 , n14730 );
or ( n14732 , n14725 , n14731 );
nand ( n14733 , n14708 , n504 );
nand ( n14734 , n14732 , n14733 );
not ( n14735 , n12648 );
not ( n14736 , n14680 );
or ( n14737 , n14735 , n14736 );
and ( n14738 , n13760 , n1077 );
not ( n14739 , n13760 );
and ( n14740 , n14739 , n499 );
nor ( n14741 , n14738 , n14740 );
nand ( n14742 , n14741 , n12702 );
nand ( n14743 , n14737 , n14742 );
xor ( n14744 , n84342 , n14619 );
xor ( n14745 , n14744 , n14648 );
xor ( n14746 , n14743 , n14745 );
not ( n14747 , n501 );
not ( n14748 , n13451 );
or ( n14749 , n14747 , n14748 );
nand ( n14750 , n12725 , n12856 );
nand ( n14751 , n14749 , n14750 );
not ( n14752 , n14751 );
not ( n14753 , n12843 );
or ( n14754 , n14752 , n14753 );
not ( n14755 , n14306 );
not ( n14756 , n14695 );
not ( n14757 , n14756 );
and ( n14758 , n14755 , n14757 );
not ( n14759 , n13524 );
and ( n14760 , n14759 , n14691 );
nor ( n14761 , n14758 , n14760 );
nand ( n14762 , n14754 , n14761 );
and ( n14763 , n14746 , n14762 );
and ( n14764 , n14743 , n14745 );
or ( n14765 , n14763 , n14764 );
xor ( n14766 , n14734 , n14765 );
xor ( n14767 , n14684 , n14686 );
xor ( n84501 , n14767 , n14698 );
and ( n14772 , n14766 , n84501 );
and ( n84503 , n14734 , n14765 );
or ( n14774 , n14772 , n84503 );
or ( n14775 , n14724 , n14774 );
not ( n14776 , n14775 );
xor ( n14777 , n14636 , n14644 );
not ( n14778 , n12647 );
and ( n14779 , n499 , n13767 );
not ( n14780 , n499 );
and ( n14781 , n14780 , n13770 );
nor ( n14782 , n14779 , n14781 );
not ( n14783 , n14782 );
or ( n14784 , n14778 , n14783 );
not ( n14785 , n499 );
not ( n14786 , n13787 );
or ( n14787 , n14785 , n14786 );
nand ( n14788 , n13600 , n12467 );
nand ( n14789 , n14787 , n14788 );
nand ( n14790 , n14789 , n12702 );
nand ( n14791 , n14784 , n14790 );
xor ( n14792 , n14777 , n14791 );
nor ( n14793 , n13775 , n12469 );
not ( n14794 , n12647 );
not ( n14795 , n14789 );
or ( n14796 , n14794 , n14795 );
and ( n14797 , n499 , n13799 );
not ( n14798 , n499 );
and ( n14799 , n14798 , n13798 );
nor ( n14800 , n14797 , n14799 );
nand ( n84531 , n14800 , n12702 );
nand ( n14805 , n14796 , n84531 );
xor ( n14806 , n14793 , n14805 );
or ( n14807 , n13776 , n500 );
nand ( n14808 , n14807 , n501 );
and ( n14809 , n13776 , n500 );
nor ( n14810 , n14809 , n12467 );
and ( n14811 , n14808 , n14810 );
not ( n14812 , n12647 );
not ( n14813 , n14800 );
or ( n14814 , n14812 , n14813 );
or ( n14815 , n13775 , n499 );
or ( n14816 , n13776 , n12467 );
nand ( n14817 , n14815 , n14816 );
nand ( n14818 , n14817 , n12702 );
nand ( n14819 , n14814 , n14818 );
and ( n14820 , n14811 , n14819 );
and ( n14821 , n14806 , n14820 );
and ( n14822 , n14793 , n14805 );
or ( n14823 , n14821 , n14822 );
and ( n14824 , n14792 , n14823 );
and ( n14825 , n14777 , n14791 );
or ( n14826 , n14824 , n14825 );
not ( n14827 , n12648 );
not ( n14828 , n14741 );
or ( n14829 , n14827 , n14828 );
nand ( n14830 , n14782 , n12702 );
nand ( n14831 , n14829 , n14830 );
xor ( n14832 , n14621 , n14630 );
xor ( n14833 , n14832 , n14645 );
xor ( n14834 , n14831 , n14833 );
not ( n14835 , n12820 );
xor ( n14836 , n501 , n12735 );
not ( n14837 , n14836 );
or ( n14838 , n14835 , n14837 );
and ( n14839 , n501 , n13114 );
not ( n14840 , n501 );
and ( n14841 , n14840 , n13612 );
nor ( n14842 , n14839 , n14841 );
nand ( n14843 , n14842 , n12821 );
nand ( n14844 , n14838 , n14843 );
xor ( n14845 , n14834 , n14844 );
xor ( n14846 , n14826 , n14845 );
not ( n14847 , n70376 );
nand ( n14848 , n14847 , n12532 );
nand ( n14849 , n12531 , n3971 );
not ( n14850 , n503 );
not ( n14851 , n13451 );
or ( n14852 , n14850 , n14851 );
or ( n14853 , n13451 , n503 );
nand ( n14854 , n14852 , n14853 );
nand ( n14855 , n14854 , n12462 );
nand ( n14856 , n14848 , n14849 , n14855 );
xor ( n14857 , n14846 , n14856 );
not ( n14858 , n12821 );
or ( n14859 , n13441 , n12856 );
nand ( n14860 , n13441 , n3117 );
nand ( n14861 , n14859 , n14860 );
not ( n14862 , n14861 );
or ( n84590 , n14858 , n14862 );
nand ( n84591 , n14842 , n12820 );
nand ( n14865 , n84590 , n84591 );
xor ( n14866 , n14777 , n14791 );
xor ( n14867 , n14866 , n14823 );
xor ( n14868 , n14865 , n14867 );
not ( n14869 , n12462 );
xor ( n14870 , n503 , n12735 );
not ( n14871 , n14870 );
or ( n14872 , n14869 , n14871 );
nand ( n14873 , n14854 , n504 );
nand ( n14874 , n14872 , n14873 );
and ( n14875 , n14868 , n14874 );
and ( n14876 , n14865 , n14867 );
or ( n14877 , n14875 , n14876 );
or ( n14878 , n14857 , n14877 );
not ( n14879 , n14878 );
not ( n14880 , n12821 );
and ( n14881 , n13512 , n501 );
not ( n14882 , n13512 );
and ( n14883 , n14882 , n12856 );
nor ( n14884 , n14881 , n14883 );
not ( n14885 , n14884 );
or ( n14886 , n14880 , n14885 );
nand ( n14887 , n14861 , n12820 );
nand ( n14888 , n14886 , n14887 );
xor ( n14889 , n14793 , n14805 );
xor ( n14890 , n14889 , n14820 );
xor ( n14891 , n14888 , n14890 );
not ( n14892 , n12462 );
and ( n14893 , n13114 , n12423 );
not ( n14894 , n13114 );
and ( n14895 , n14894 , n503 );
or ( n14896 , n14893 , n14895 );
not ( n14897 , n14896 );
or ( n14898 , n14892 , n14897 );
nand ( n14899 , n14870 , n504 );
nand ( n14900 , n14898 , n14899 );
and ( n14901 , n14891 , n14900 );
and ( n14902 , n14888 , n14890 );
or ( n14903 , n14901 , n14902 );
xor ( n14904 , n14865 , n14867 );
xor ( n14905 , n14904 , n14874 );
xor ( n14906 , n14903 , n14905 );
xor ( n14907 , n14811 , n14819 );
not ( n14908 , n12820 );
not ( n14909 , n14884 );
or ( n14910 , n14908 , n14909 );
not ( n14911 , n501 );
not ( n14912 , n13787 );
or ( n14913 , n14911 , n14912 );
nand ( n14914 , n13600 , n12856 );
nand ( n14915 , n14913 , n14914 );
nand ( n14916 , n14915 , n12821 );
nand ( n14917 , n14910 , n14916 );
xor ( n14918 , n14907 , n14917 );
and ( n14919 , n13776 , n12647 );
and ( n84647 , n13798 , n3117 );
not ( n14921 , n13798 );
and ( n14922 , n14921 , n501 );
nor ( n14923 , n84647 , n14922 );
nand ( n14924 , n14923 , n12820 );
nand ( n14925 , n14691 , n13776 );
nand ( n14926 , n14695 , n13775 );
and ( n14927 , n14924 , n14925 , n14926 );
or ( n14928 , n13776 , n502 );
nand ( n14929 , n14928 , n503 );
and ( n14930 , n13776 , n502 );
nor ( n14931 , n14930 , n12856 );
nand ( n14932 , n14929 , n14931 );
nor ( n14933 , n14927 , n14932 );
xor ( n14934 , n14919 , n14933 );
not ( n14935 , n12820 );
not ( n14936 , n14915 );
or ( n14937 , n14935 , n14936 );
nand ( n14938 , n14923 , n12821 );
nand ( n14939 , n14937 , n14938 );
and ( n14940 , n14934 , n14939 );
or ( n14942 , n14940 , C0 );
and ( n14943 , n14918 , n14942 );
and ( n14944 , n14907 , n14917 );
or ( n14945 , n14943 , n14944 );
xor ( n14946 , n14907 , n14917 );
xor ( n14947 , n14946 , n14942 );
not ( n14948 , n14896 );
not ( n14949 , n504 );
or ( n14950 , n14948 , n14949 );
not ( n14951 , n13441 );
not ( n14952 , n503 );
and ( n14953 , n14951 , n14952 );
and ( n14954 , n13441 , n503 );
nor ( n14955 , n14953 , n14954 );
nand ( n14956 , n14955 , n12462 );
nand ( n14957 , n14950 , n14956 );
or ( n14958 , n14947 , n14957 );
xor ( n14959 , n14919 , n14933 );
xor ( n14960 , n14959 , n14939 );
not ( n14961 , n13512 );
not ( n14962 , n12423 );
or ( n14963 , n14961 , n14962 );
or ( n14964 , n13512 , n12423 );
nand ( n14965 , n14963 , n14964 );
not ( n14966 , n14965 );
not ( n14967 , n12462 );
or ( n14968 , n14966 , n14967 );
not ( n14969 , n14955 );
or ( n14970 , n14969 , n1636 );
nand ( n14971 , n14968 , n14970 );
nor ( n14972 , n14960 , n14971 );
not ( n14973 , n14932 );
nand ( n14974 , n14924 , n14925 , n14926 );
not ( n14975 , n14974 );
or ( n14976 , n14973 , n14975 );
or ( n14977 , n14974 , n14932 );
nand ( n14978 , n14976 , n14977 );
not ( n14979 , n504 );
not ( n14980 , n14965 );
or ( n14981 , n14979 , n14980 );
not ( n14982 , n13600 );
not ( n14983 , n503 );
and ( n14984 , n14982 , n14983 );
and ( n14985 , n13600 , n503 );
nor ( n14986 , n14984 , n14985 );
nand ( n14987 , n14986 , n12462 );
nand ( n14988 , n14981 , n14987 );
xor ( n14989 , n14978 , n14988 );
not ( n14990 , n504 );
or ( n14991 , n13799 , n12423 , n14990 );
nor ( n14992 , n503 , n14990 );
and ( n14993 , n13799 , n14992 );
and ( n14994 , n12462 , n13775 );
nor ( n14995 , n14993 , n14994 );
nand ( n14996 , n14991 , n14995 );
not ( n14997 , n504 );
nor ( n14998 , n14997 , n13775 );
nor ( n14999 , n14998 , n12423 );
nand ( n15000 , n14996 , n14999 );
not ( n15001 , n15000 );
not ( n15002 , n12820 );
nor ( n15003 , n15002 , n13775 );
nor ( n15004 , n15001 , n15003 );
not ( n15005 , n503 );
not ( n15006 , n13799 );
or ( n15007 , n15005 , n15006 );
or ( n84734 , n13799 , n503 );
nand ( n15009 , n15007 , n84734 );
not ( n15010 , n15009 );
not ( n15011 , n12461 );
and ( n15012 , n15010 , n15011 );
and ( n15013 , n14986 , n504 );
nor ( n15014 , n15012 , n15013 );
or ( n15015 , n15004 , n15014 );
nand ( n15017 , n15015 , C1 );
and ( n15018 , n14989 , n15017 );
and ( n15019 , n14978 , n14988 );
or ( n15020 , n15018 , n15019 );
not ( n15021 , n15020 );
or ( n15022 , n14972 , n15021 );
nand ( n15023 , n14971 , n14960 );
nand ( n15024 , n15022 , n15023 );
nand ( n15025 , n14958 , n15024 );
nand ( n15026 , n14947 , n14957 );
nand ( n15027 , n15025 , n15026 );
xor ( n15028 , n14945 , n15027 );
xor ( n15029 , n14888 , n14890 );
xor ( n15030 , n15029 , n14900 );
and ( n15031 , n15028 , n15030 );
and ( n15032 , n14945 , n15027 );
or ( n15033 , n15031 , n15032 );
and ( n15034 , n14906 , n15033 );
and ( n15035 , n14903 , n14905 );
or ( n15036 , n15034 , n15035 );
not ( n15037 , n15036 );
or ( n15038 , n14879 , n15037 );
nand ( n15039 , n14857 , n14877 );
nand ( n15040 , n15038 , n15039 );
not ( n15041 , n15040 );
xor ( n15042 , n14831 , n14833 );
and ( n15043 , n15042 , n14844 );
and ( n15044 , n14831 , n14833 );
or ( n15045 , n15043 , n15044 );
xor ( n15046 , n14743 , n14745 );
xor ( n15047 , n15046 , n14762 );
xor ( n15048 , n15045 , n15047 );
not ( n15049 , n504 );
not ( n15050 , n14730 );
or ( n15051 , n15049 , n15050 );
nand ( n15052 , n12532 , n12462 );
nand ( n15053 , n15051 , n15052 );
xor ( n15054 , n15048 , n15053 );
not ( n15055 , n15054 );
xor ( n15056 , n14826 , n14845 );
and ( n15057 , n15056 , n14856 );
and ( n15058 , n14826 , n14845 );
or ( n15059 , n15057 , n15058 );
not ( n15060 , n15059 );
nand ( n15061 , n15055 , n15060 );
not ( n15062 , n15061 );
or ( n15063 , n15041 , n15062 );
nand ( n15064 , n15054 , n15059 );
nand ( n15065 , n15063 , n15064 );
not ( n15066 , n15065 );
xor ( n15067 , n14734 , n14765 );
xor ( n15068 , n15067 , n84501 );
not ( n15069 , n15068 );
xor ( n15070 , n15045 , n15047 );
and ( n15071 , n15070 , n15053 );
and ( n15072 , n15045 , n15047 );
or ( n15073 , n15071 , n15072 );
not ( n15074 , n15073 );
nand ( n15075 , n15069 , n15074 );
not ( n84801 , n15075 );
or ( n15080 , n15066 , n84801 );
nand ( n84803 , n15068 , n15073 );
nand ( n15082 , n15080 , n84803 );
not ( n15083 , n15082 );
or ( n15084 , n14776 , n15083 );
nand ( n15085 , n14724 , n14774 );
nand ( n15086 , n15084 , n15085 );
not ( n15087 , n15086 );
or ( n15088 , n14722 , n15087 );
nand ( n15089 , n14719 , n14716 );
nand ( n15090 , n15088 , n15089 );
not ( n15091 , n15090 );
or ( n15092 , n14675 , n15091 );
or ( n15093 , n14589 , n14534 );
and ( n15094 , n14593 , n14672 );
and ( n15095 , n15093 , n15094 );
and ( n15096 , n14534 , n14589 );
nor ( n15097 , n15095 , n15096 );
nand ( n15098 , n15092 , n15097 );
not ( n15099 , n15098 );
or ( n15100 , n14532 , n15099 );
not ( n15101 , n14354 );
not ( n15102 , n14465 );
nand ( n84825 , n15101 , n15102 );
nand ( n15107 , n14469 , n14529 );
not ( n15108 , n15107 );
and ( n15109 , n84825 , n15108 );
nand ( n15110 , n14354 , n14465 );
not ( n15111 , n15110 );
nor ( n15112 , n15109 , n15111 );
nand ( n15113 , n15100 , n15112 );
not ( n15114 , n15113 );
or ( n15115 , n14352 , n15114 );
nand ( n15116 , n14286 , n14350 );
nand ( n15117 , n15115 , n15116 );
not ( n15118 , n15117 );
or ( n15119 , n14284 , n15118 );
nand ( n15120 , n14282 , n14209 );
nand ( n15121 , n15119 , n15120 );
not ( n15122 , n15121 );
xor ( n15123 , n83876 , n14139 );
and ( n15124 , n15123 , n14142 );
and ( n15125 , n83876 , n14139 );
or ( n15126 , n15124 , n15125 );
not ( n15127 , n13032 );
not ( n15128 , n13581 );
not ( n15129 , n15128 );
or ( n15130 , n15127 , n15129 );
nand ( n15131 , n14069 , n12969 );
nand ( n15132 , n15130 , n15131 );
xor ( n15133 , n15126 , n15132 );
not ( n15134 , n14091 );
not ( n15135 , n12517 );
or ( n15136 , n15134 , n15135 );
not ( n15137 , n13586 );
nand ( n15138 , n15137 , n12470 );
nand ( n15139 , n15136 , n15138 );
and ( n15140 , n15133 , n15139 );
and ( n15141 , n15126 , n15132 );
or ( n15142 , n15140 , n15141 );
xor ( n15143 , n13585 , n13589 );
xor ( n15144 , n15143 , n13638 );
xor ( n15145 , n15142 , n15144 );
xor ( n15146 , n13622 , n13632 );
xor ( n15147 , n15146 , n13635 );
not ( n15148 , n12650 );
not ( n15149 , n499 );
not ( n15150 , n13378 );
or ( n15151 , n15149 , n15150 );
not ( n15152 , n499 );
nand ( n15153 , n15152 , n14099 );
nand ( n15154 , n15151 , n15153 );
not ( n15155 , n15154 );
or ( n15156 , n15148 , n15155 );
nand ( n15157 , n12702 , n14150 );
nand ( n15158 , n15156 , n15157 );
xor ( n84878 , n15147 , n15158 );
xor ( n84879 , n14064 , n14081 );
and ( n15161 , n84879 , n14093 );
and ( n15162 , n14064 , n14081 );
or ( n15163 , n15161 , n15162 );
and ( n15164 , n84878 , n15163 );
and ( n15165 , n15147 , n15158 );
or ( n15166 , n15164 , n15165 );
xor ( n15167 , n15145 , n15166 );
not ( n15168 , n12462 );
not ( n15169 , n14117 );
or ( n15170 , n15168 , n15169 );
not ( n15171 , n503 );
not ( n15172 , n13484 );
or ( n15173 , n15171 , n15172 );
nand ( n15174 , n13483 , n12457 );
nand ( n15175 , n15173 , n15174 );
nand ( n15176 , n15175 , n504 );
nand ( n15177 , n15170 , n15176 );
xor ( n15178 , n15147 , n15158 );
xor ( n15179 , n15178 , n15163 );
xor ( n15180 , n15177 , n15179 );
xor ( n15181 , n14094 , n14110 );
and ( n15182 , n15181 , n14121 );
and ( n15183 , n14094 , n14110 );
or ( n15184 , n15182 , n15183 );
and ( n15185 , n15180 , n15184 );
and ( n15186 , n15177 , n15179 );
or ( n15187 , n15185 , n15186 );
xor ( n15188 , n15167 , n15187 );
not ( n15189 , n12462 );
not ( n15190 , n15175 );
or ( n15191 , n15189 , n15190 );
nand ( n15192 , n13712 , n504 );
nand ( n15193 , n15191 , n15192 );
xor ( n15194 , n14143 , n14152 );
and ( n15195 , n15194 , n14171 );
and ( n15196 , n14143 , n14152 );
or ( n15197 , n15195 , n15196 );
xor ( n15198 , n15126 , n15132 );
xor ( n15199 , n15198 , n15139 );
xor ( n15200 , n15197 , n15199 );
not ( n15201 , n14108 );
not ( n15202 , n12822 );
or ( n15203 , n15201 , n15202 );
not ( n15204 , n501 );
not ( n15205 , n12506 );
or ( n15206 , n15204 , n15205 );
nand ( n15207 , n12509 , n12856 );
nand ( n15208 , n15206 , n15207 );
not ( n15209 , n15208 );
not ( n15210 , n12843 );
or ( n15211 , n15209 , n15210 );
nand ( n15212 , n15203 , n15211 );
and ( n15213 , n15200 , n15212 );
and ( n15214 , n15197 , n15199 );
or ( n15215 , n15213 , n15214 );
xor ( n84935 , n15193 , n15215 );
xor ( n15217 , n13535 , n13543 );
xor ( n15218 , n15217 , n13546 );
not ( n15219 , n12702 );
not ( n15220 , n15154 );
or ( n15221 , n15219 , n15220 );
nand ( n15222 , n13568 , n12650 );
nand ( n15223 , n15221 , n15222 );
xor ( n15224 , n15218 , n15223 );
not ( n15225 , n12822 );
not ( n15226 , n15208 );
or ( n15227 , n15225 , n15226 );
nand ( n15228 , n83453 , n12843 );
nand ( n15229 , n15227 , n15228 );
xor ( n15230 , n15224 , n15229 );
xor ( n15231 , n84935 , n15230 );
xor ( n15232 , n15188 , n15231 );
xor ( n15233 , n15197 , n15199 );
xor ( n15234 , n15233 , n15212 );
xor ( n15235 , n14127 , n14172 );
and ( n15236 , n15235 , n14207 );
and ( n15237 , n14127 , n14172 );
or ( n15238 , n15236 , n15237 );
xor ( n15239 , n15234 , n15238 );
xor ( n15240 , n15177 , n15179 );
xor ( n15241 , n15240 , n15184 );
and ( n15242 , n15239 , n15241 );
and ( n15243 , n15234 , n15238 );
or ( n15244 , n15242 , n15243 );
nor ( n15245 , n15232 , n15244 );
xor ( n15246 , n15234 , n15238 );
xor ( n15247 , n15246 , n15241 );
xor ( n15248 , n14033 , n14122 );
and ( n15249 , n15248 , n14208 );
and ( n15250 , n14033 , n14122 );
or ( n15251 , n15249 , n15250 );
nor ( n15252 , n15247 , n15251 );
nor ( n15253 , n15245 , n15252 );
not ( n15254 , n15253 );
or ( n15255 , n15122 , n15254 );
not ( n15256 , n15245 );
nand ( n15257 , n15247 , n15251 );
not ( n15258 , n15257 );
and ( n15259 , n15256 , n15258 );
and ( n15260 , n15232 , n15244 );
nor ( n15261 , n15259 , n15260 );
nand ( n15262 , n15255 , n15261 );
xor ( n15263 , n15193 , n15215 );
and ( n15264 , n15263 , n15230 );
and ( n15265 , n15193 , n15215 );
or ( n15266 , n15264 , n15265 );
xor ( n15267 , n13692 , n13703 );
xor ( n15268 , n15267 , n13714 );
xor ( n15269 , n15266 , n15268 );
xor ( n15270 , n15218 , n15223 );
and ( n15271 , n15270 , n15229 );
and ( n15272 , n15218 , n15223 );
or ( n15273 , n15271 , n15272 );
xor ( n15274 , n13574 , n13576 );
xor ( n15275 , n15274 , n13641 );
xor ( n15276 , n15273 , n15275 );
xor ( n15277 , n15142 , n15144 );
and ( n15278 , n15277 , n15166 );
and ( n15279 , n15142 , n15144 );
or ( n15280 , n15278 , n15279 );
xor ( n15281 , n15276 , n15280 );
and ( n15282 , n15269 , n15281 );
and ( n15283 , n15266 , n15268 );
or ( n15284 , n15282 , n15283 );
xor ( n15285 , n13563 , n13644 );
xor ( n15286 , n15285 , n13661 );
xor ( n15287 , n15273 , n15275 );
and ( n15288 , n15287 , n15280 );
and ( n15289 , n15273 , n15275 );
or ( n15290 , n15288 , n15289 );
xor ( n15291 , n15286 , n15290 );
xor ( n15292 , n13687 , n13689 );
xor ( n15293 , n15292 , n13717 );
xor ( n15294 , n15291 , n15293 );
nor ( n15295 , n15284 , n15294 );
xor ( n15296 , n15266 , n15268 );
xor ( n15297 , n15296 , n15281 );
xor ( n15298 , n15167 , n15187 );
and ( n85018 , n15298 , n15231 );
and ( n15300 , n15167 , n15187 );
or ( n15301 , n85018 , n15300 );
nor ( n15302 , n15297 , n15301 );
nor ( n15303 , n15295 , n15302 );
xor ( n15304 , n13685 , n13720 );
xor ( n15305 , n15304 , n13723 );
xor ( n15306 , n15286 , n15290 );
and ( n15307 , n15306 , n15293 );
and ( n15308 , n15286 , n15290 );
or ( n15309 , n15307 , n15308 );
nor ( n15310 , n15305 , n15309 );
not ( n15311 , n15310 );
and ( n15312 , n13728 , n15262 , n15303 , n15311 );
nand ( n15313 , n15297 , n15301 );
or ( n15314 , n15295 , n15313 );
nand ( n15315 , n15284 , n15294 );
nand ( n15316 , n15314 , n15315 );
not ( n15317 , n15316 );
nor ( n15318 , n13727 , n15310 );
not ( n15319 , n15318 );
or ( n15320 , n15317 , n15319 );
not ( n15321 , n13727 );
nand ( n15322 , n15305 , n15309 );
not ( n15323 , n15322 );
and ( n15324 , n15321 , n15323 );
and ( n15325 , n13683 , n13726 );
nor ( n15326 , n15324 , n15325 );
nand ( n15327 , n15320 , n15326 );
or ( n15328 , n15312 , n15327 );
nand ( n15329 , n13337 , n13417 );
not ( n15330 , n83178 );
not ( n15331 , n13676 );
nand ( n15332 , n15330 , n15331 );
and ( n15333 , n15329 , n15332 );
nand ( n15334 , n15328 , n15333 );
not ( n15335 , n15334 );
or ( n15336 , n13681 , n15335 );
not ( n15337 , n12758 );
and ( n15338 , n493 , n12509 );
not ( n15339 , n493 );
and ( n15340 , n15339 , n12506 );
nor ( n15341 , n15338 , n15340 );
not ( n15342 , n15341 );
or ( n15343 , n15337 , n15342 );
buf ( n15344 , n12791 );
nand ( n15345 , n13271 , n15344 );
nand ( n15346 , n15343 , n15345 );
xor ( n15347 , n83070 , n13313 );
and ( n15348 , n15347 , n13326 );
and ( n15349 , n83070 , n13313 );
or ( n15350 , n15348 , n15349 );
xor ( n15351 , n15346 , n15350 );
and ( n15352 , n495 , n13484 );
not ( n15353 , n495 );
and ( n15354 , n15353 , n13483 );
or ( n15355 , n15352 , n15354 );
not ( n15356 , n15355 );
not ( n15357 , n13032 );
or ( n15358 , n15356 , n15357 );
nand ( n15359 , n13280 , n12969 );
nand ( n15360 , n15358 , n15359 );
xor ( n15361 , n15351 , n15360 );
xor ( n15362 , n13303 , n13327 );
and ( n85082 , n15362 , n13332 );
and ( n15367 , n13303 , n13327 );
or ( n85084 , n85082 , n15367 );
xor ( n15369 , n15361 , n85084 );
xor ( n15370 , n13168 , n13177 );
and ( n15371 , n15370 , n13262 );
and ( n15372 , n13168 , n13177 );
or ( n15373 , n15371 , n15372 );
and ( n15374 , n15369 , n15373 );
and ( n15375 , n15361 , n85084 );
or ( n15376 , n15374 , n15375 );
not ( n15377 , n12702 );
not ( n15378 , n13175 );
or ( n15379 , n15377 , n15378 );
not ( n15380 , n499 );
not ( n15381 , n12886 );
or ( n15382 , n15380 , n15381 );
nand ( n15383 , n13372 , n12467 );
nand ( n15384 , n15382 , n15383 );
nand ( n15385 , n15384 , n12650 );
nand ( n15386 , n15379 , n15385 );
not ( n15387 , n12470 );
not ( n15388 , n497 );
not ( n15389 , n82600 );
or ( n15390 , n15388 , n15389 );
nand ( n15391 , n13650 , n12486 );
nand ( n15392 , n15390 , n15391 );
not ( n85109 , n15392 );
or ( n15397 , n15387 , n85109 );
nand ( n15398 , n13301 , n12517 );
nand ( n15399 , n15397 , n15398 );
xor ( n15400 , n15386 , n15399 );
and ( n15401 , n13324 , n13325 );
not ( n15402 , n12638 );
not ( n15403 , n491 );
not ( n15404 , n12981 );
or ( n15405 , n15403 , n15404 );
not ( n15406 , n491 );
nand ( n15407 , n15406 , n12980 );
nand ( n15408 , n15405 , n15407 );
not ( n15409 , n15408 );
or ( n15410 , n15402 , n15409 );
nand ( n15411 , n13307 , n12595 );
nand ( n15412 , n15410 , n15411 );
xor ( n15413 , n15401 , n15412 );
nand ( n15414 , n12606 , n489 );
not ( n15415 , n15414 );
not ( n15416 , n15415 );
not ( n15417 , n12795 );
not ( n15418 , n489 );
not ( n15419 , n12900 );
or ( n15420 , n15418 , n15419 );
nand ( n15421 , n12774 , n12560 );
nand ( n15422 , n15420 , n15421 );
not ( n15423 , n15422 );
or ( n15424 , n15417 , n15423 );
nand ( n15425 , n13322 , n12542 );
nand ( n15426 , n15424 , n15425 );
not ( n15427 , n15426 );
not ( n15428 , n15427 );
or ( n15429 , n15416 , n15428 );
or ( n15430 , n15427 , n15415 );
nand ( n15431 , n15429 , n15430 );
xor ( n15432 , n15413 , n15431 );
xor ( n15433 , n15400 , n15432 );
not ( n15434 , n12820 );
not ( n15435 , n501 );
not ( n15436 , n12419 );
or ( n15437 , n15435 , n15436 );
not ( n15438 , n12418 );
not ( n15439 , n15438 );
nand ( n15440 , n15439 , n12856 );
nand ( n15441 , n15437 , n15440 );
not ( n15442 , n15441 );
or ( n15443 , n15434 , n15442 );
nand ( n15444 , n13166 , n12822 );
nand ( n15445 , n15443 , n15444 );
xor ( n15446 , n13273 , n13282 );
and ( n15447 , n15446 , n13287 );
and ( n15448 , n13273 , n13282 );
or ( n15449 , n15447 , n15448 );
xor ( n15450 , n15445 , n15449 );
not ( n15451 , n12462 );
not ( n15452 , n13260 );
or ( n15453 , n15451 , n15452 );
not ( n15454 , n503 );
not ( n15455 , n13248 );
xor ( n15456 , n13203 , n13207 );
and ( n15457 , n15456 , n13235 );
and ( n15458 , n13203 , n13207 );
or ( n15459 , n15457 , n15458 );
not ( n15460 , n15459 );
xor ( n15461 , n13214 , n13229 );
and ( n15462 , n15461 , n13234 );
and ( n15463 , n13214 , n13229 );
or ( n15464 , n15462 , n15463 );
not ( n15465 , n15464 );
nand ( n15466 , n525 , n457 );
not ( n15467 , n13226 );
not ( n15468 , n10087 );
or ( n15469 , n15467 , n15468 );
not ( n15470 , n459 );
nor ( n15471 , n15470 , n521 );
not ( n15472 , n521 );
nor ( n15473 , n15472 , n459 );
nor ( n15474 , n15471 , n15473 );
not ( n15475 , n15474 );
nand ( n15476 , n15475 , n10094 );
nand ( n15477 , n15469 , n15476 );
xor ( n15478 , n15466 , n15477 );
and ( n15479 , n462 , n463 );
not ( n15480 , n462 );
and ( n15481 , n15480 , n2374 );
nor ( n15482 , n15479 , n15481 );
or ( n15483 , n10184 , n15482 );
not ( n15484 , n10194 );
nand ( n85198 , n15483 , n15484 );
nand ( n15486 , n85198 , n461 );
xor ( n15487 , n15478 , n15486 );
not ( n15488 , n15487 );
not ( n15489 , n13219 );
not ( n15490 , n10127 );
or ( n15491 , n15489 , n15490 );
xor ( n15492 , n457 , n523 );
nand ( n15493 , n10068 , n15492 );
nand ( n15494 , n15491 , n15493 );
xor ( n15495 , n13213 , n15494 );
xor ( n15496 , n13215 , n13221 );
and ( n15497 , n15496 , n13228 );
and ( n15498 , n13215 , n13221 );
or ( n15499 , n15497 , n15498 );
xor ( n15500 , n15495 , n15499 );
not ( n15501 , n15500 );
or ( n15502 , n15488 , n15501 );
or ( n15503 , n15500 , n15487 );
nand ( n15504 , n15502 , n15503 );
not ( n15505 , n15504 );
or ( n15506 , n15465 , n15505 );
or ( n15507 , n15504 , n15464 );
nand ( n15508 , n15506 , n15507 );
nand ( n15509 , n15460 , n15508 );
not ( n15510 , n15509 );
not ( n15511 , n15510 );
not ( n15512 , n15508 );
nand ( n15513 , n15512 , n15459 );
nand ( n15514 , n15511 , n15513 );
nor ( n15515 , n15455 , n15514 );
not ( n15516 , n15515 );
nand ( n15517 , n12334 , n12330 , n12410 );
nor ( n15518 , n13195 , n15517 );
not ( n15519 , n15518 );
nand ( n15520 , n82432 , n12316 );
not ( n15521 , n15520 );
or ( n15522 , n15519 , n15521 );
not ( n15523 , n13184 );
not ( n15524 , n15523 );
not ( n15525 , n10692 );
or ( n15526 , n15524 , n15525 );
nand ( n15527 , n15526 , n12410 );
not ( n15528 , n15527 );
and ( n15529 , n15528 , n13194 );
nor ( n15530 , n15529 , n13246 );
nand ( n15531 , n15522 , n15530 );
not ( n15532 , n15531 );
or ( n15533 , n15516 , n15532 );
not ( n15534 , n13248 );
not ( n15535 , n15531 );
or ( n15536 , n15534 , n15535 );
nand ( n15537 , n15536 , n15514 );
nand ( n15538 , n15533 , n15537 );
buf ( n15539 , n15538 );
not ( n15540 , n15539 );
not ( n15541 , n15540 );
or ( n15542 , n15454 , n15541 );
not ( n15543 , n15538 );
not ( n15544 , n15543 );
nand ( n15545 , n15544 , n12423 );
nand ( n15546 , n15542 , n15545 );
nand ( n15547 , n15546 , n504 );
nand ( n15548 , n15453 , n15547 );
xor ( n15549 , n15450 , n15548 );
xor ( n15550 , n15433 , n15549 );
xor ( n15551 , n13288 , n13292 );
and ( n15552 , n15551 , n13333 );
and ( n15553 , n13288 , n13292 );
or ( n15554 , n15552 , n15553 );
and ( n15555 , n15550 , n15554 );
and ( n15556 , n15433 , n15549 );
or ( n15557 , n15555 , n15556 );
xor ( n15558 , n15376 , n15557 );
not ( n15559 , n12702 );
not ( n15560 , n15384 );
or ( n15561 , n15559 , n15560 );
not ( n15562 , n499 );
not ( n15563 , n12452 );
not ( n15564 , n15563 );
or ( n15565 , n15562 , n15564 );
buf ( n15566 , n12452 );
nand ( n15567 , n15566 , n12467 );
nand ( n85281 , n15565 , n15567 );
nand ( n15569 , n85281 , n12650 );
nand ( n15570 , n15561 , n15569 );
not ( n15571 , n12470 );
nand ( n15572 , n13369 , n12486 );
nand ( n15573 , n13370 , n497 );
nand ( n15574 , n15572 , n15573 );
not ( n15575 , n15574 );
or ( n15576 , n15571 , n15575 );
nand ( n15577 , n15392 , n12517 );
nand ( n15578 , n15576 , n15577 );
xor ( n15579 , n15570 , n15578 );
not ( n15580 , n15408 );
not ( n15581 , n12595 );
or ( n15582 , n15580 , n15581 );
not ( n15583 , n491 );
not ( n15584 , n13009 );
or ( n15585 , n15583 , n15584 );
or ( n15586 , n13009 , n491 );
nand ( n15587 , n15585 , n15586 );
nand ( n15588 , n15587 , n12638 );
nand ( n15589 , n15582 , n15588 );
not ( n15590 , n15426 );
nor ( n15591 , n15590 , n15414 );
xor ( n15592 , n15589 , n15591 );
not ( n15593 , n12629 );
and ( n15594 , n15593 , n489 );
not ( n15595 , n12542 );
not ( n15596 , n15422 );
or ( n15597 , n15595 , n15596 );
not ( n15598 , n489 );
not ( n15599 , n82837 );
or ( n15600 , n15598 , n15599 );
nand ( n15601 , n12949 , n12560 );
nand ( n15602 , n15600 , n15601 );
nand ( n15603 , n15602 , n12795 );
nand ( n15604 , n15597 , n15603 );
xor ( n15605 , n15594 , n15604 );
xor ( n15606 , n15592 , n15605 );
xor ( n15607 , n15579 , n15606 );
not ( n15608 , n12822 );
not ( n15609 , n15441 );
or ( n15610 , n15608 , n15609 );
not ( n15611 , n501 );
not ( n15612 , n13255 );
or ( n15613 , n15611 , n15612 );
nand ( n15614 , n13258 , n12856 );
nand ( n15615 , n15613 , n15614 );
nand ( n15616 , n15615 , n12843 );
nand ( n15617 , n15610 , n15616 );
not ( n15618 , n12462 );
not ( n15619 , n15546 );
or ( n15620 , n15618 , n15619 );
not ( n15621 , n15487 );
not ( n15622 , n15621 );
not ( n15623 , n15500 );
or ( n15624 , n15622 , n15623 );
not ( n15625 , n15500 );
nand ( n85339 , n15625 , n15487 );
nand ( n15630 , n15464 , n85339 );
nand ( n85341 , n15624 , n15630 );
not ( n15632 , n15466 );
or ( n15633 , n15477 , n15632 );
nand ( n15634 , n15633 , n15486 );
nand ( n15635 , n15477 , n15632 );
nand ( n15636 , n15634 , n15635 );
and ( n15637 , n457 , n524 );
not ( n15638 , n15492 );
not ( n15639 , n10127 );
or ( n15640 , n15638 , n15639 );
xnor ( n15641 , n457 , n522 );
not ( n15642 , n15641 );
nand ( n15643 , n15642 , n10068 );
nand ( n15644 , n15640 , n15643 );
xor ( n15645 , n15637 , n15644 );
not ( n15646 , n10086 );
not ( n15647 , n15474 );
and ( n15648 , n15646 , n15647 );
and ( n15649 , n10094 , n459 );
nor ( n85360 , n15648 , n15649 );
xor ( n15654 , n15645 , n85360 );
xor ( n15655 , n15636 , n15654 );
xor ( n15656 , n13213 , n15494 );
and ( n15657 , n15656 , n15499 );
and ( n15658 , n13213 , n15494 );
or ( n15659 , n15657 , n15658 );
xor ( n15660 , n15655 , n15659 );
or ( n15661 , n85341 , n15660 );
nand ( n15662 , n85341 , n15660 );
nand ( n15663 , n15661 , n15662 );
not ( n15664 , n15663 );
not ( n15665 , n15664 );
not ( n15666 , n12440 );
not ( n15667 , n13186 );
or ( n15668 , n15666 , n15667 );
buf ( n15669 , n13194 );
nand ( n15670 , n15668 , n15669 );
nor ( n15671 , n13245 , n13236 );
nor ( n15672 , n15510 , n15671 );
buf ( n15673 , n15672 );
nand ( n15674 , n15670 , n15673 );
and ( n15675 , n13193 , n15672 );
not ( n15676 , n15509 );
not ( n15677 , n13248 );
not ( n15678 , n15677 );
or ( n15679 , n15676 , n15678 );
nand ( n15680 , n15679 , n15513 );
nor ( n15681 , n15675 , n15680 );
nand ( n15682 , n15674 , n15681 );
not ( n15683 , n15682 );
not ( n15684 , n15683 );
or ( n15685 , n15665 , n15684 );
not ( n15686 , n15681 );
not ( n15687 , n15674 );
or ( n15688 , n15686 , n15687 );
nand ( n15689 , n15688 , n15663 );
nand ( n15690 , n15685 , n15689 );
and ( n15691 , n12457 , n15690 );
not ( n15692 , n12457 );
not ( n15693 , n15664 );
not ( n15694 , n15683 );
or ( n15695 , n15693 , n15694 );
nand ( n15696 , n15695 , n15689 );
not ( n15697 , n15696 );
and ( n15698 , n15692 , n15697 );
nor ( n15699 , n15691 , n15698 );
not ( n15700 , n15699 );
nand ( n15701 , n15700 , n504 );
nand ( n15702 , n15620 , n15701 );
xor ( n15703 , n15617 , n15702 );
xor ( n15704 , n15346 , n15350 );
and ( n15705 , n15704 , n15360 );
and ( n15706 , n15346 , n15350 );
or ( n15707 , n15705 , n15706 );
xor ( n15708 , n15703 , n15707 );
xor ( n15709 , n15607 , n15708 );
not ( n15710 , n15344 );
not ( n15711 , n15341 );
or ( n15712 , n15710 , n15711 );
and ( n15713 , n12482 , n493 );
not ( n15714 , n12482 );
and ( n15715 , n15714 , n12775 );
or ( n15716 , n15713 , n15715 );
nand ( n15717 , n15716 , n12758 );
nand ( n15718 , n15712 , n15717 );
xor ( n15719 , n15401 , n15412 );
and ( n15720 , n15719 , n15431 );
and ( n15721 , n15401 , n15412 );
or ( n15722 , n15720 , n15721 );
xor ( n15723 , n15718 , n15722 );
not ( n15724 , n12969 );
not ( n15725 , n15355 );
or ( n15726 , n15724 , n15725 );
not ( n15727 , n495 );
not ( n15728 , n12671 );
or ( n15729 , n15727 , n15728 );
not ( n15730 , n495 );
nand ( n15731 , n15730 , n12674 );
nand ( n15732 , n15729 , n15731 );
nand ( n15733 , n15732 , n13032 );
nand ( n15734 , n15726 , n15733 );
xor ( n15735 , n15723 , n15734 );
xor ( n15736 , n15386 , n15399 );
and ( n15737 , n15736 , n15432 );
and ( n15738 , n15386 , n15399 );
or ( n15739 , n15737 , n15738 );
xor ( n85447 , n15735 , n15739 );
xor ( n15741 , n15445 , n15449 );
and ( n15742 , n15741 , n15548 );
and ( n15743 , n15445 , n15449 );
or ( n15744 , n15742 , n15743 );
xor ( n15745 , n85447 , n15744 );
xor ( n15746 , n15709 , n15745 );
xor ( n15747 , n15558 , n15746 );
not ( n15748 , n15747 );
xor ( n15749 , n15361 , n85084 );
xor ( n15750 , n15749 , n15373 );
xor ( n15751 , n15433 , n15549 );
xor ( n15752 , n15751 , n15554 );
xor ( n15753 , n15750 , n15752 );
xor ( n15754 , n13158 , n13263 );
and ( n15755 , n15754 , n83092 );
and ( n15756 , n13158 , n13263 );
or ( n15757 , n15755 , n15756 );
and ( n15758 , n15753 , n15757 );
and ( n15759 , n15750 , n15752 );
or ( n15760 , n15758 , n15759 );
not ( n15761 , n15760 );
and ( n15762 , n15748 , n15761 );
xor ( n15763 , n15750 , n15752 );
xor ( n15764 , n15763 , n15757 );
xor ( n15765 , n12896 , n13153 );
and ( n15766 , n15765 , n13335 );
and ( n15767 , n12896 , n13153 );
or ( n15768 , n15766 , n15767 );
nor ( n15769 , n15764 , n15768 );
nor ( n15770 , n15762 , n15769 );
nand ( n15771 , n15336 , n15770 );
or ( n15772 , n15747 , n15760 );
nand ( n15773 , n15764 , n15768 );
not ( n15774 , n15773 );
and ( n15775 , n15772 , n15774 );
and ( n15776 , n15747 , n15760 );
nor ( n15777 , n15775 , n15776 );
nand ( n15778 , n15771 , n15777 );
xor ( n15779 , n15570 , n15578 );
and ( n15780 , n15779 , n15606 );
and ( n15781 , n15570 , n15578 );
or ( n15782 , n15780 , n15781 );
xor ( n15783 , n15589 , n15591 );
and ( n15784 , n15783 , n15605 );
and ( n15785 , n15589 , n15591 );
or ( n15786 , n15784 , n15785 );
not ( n15787 , n12758 );
and ( n15788 , n12694 , n493 );
not ( n15789 , n12694 );
and ( n15790 , n15789 , n12775 );
or ( n15791 , n15788 , n15790 );
not ( n15792 , n15791 );
or ( n15793 , n15787 , n15792 );
nand ( n15794 , n15716 , n15344 );
nand ( n15795 , n15793 , n15794 );
xor ( n15796 , n15786 , n15795 );
not ( n15797 , n13032 );
and ( n15798 , n495 , n12835 );
not ( n15799 , n495 );
and ( n15800 , n15799 , n82600 );
nor ( n15801 , n15798 , n15800 );
not ( n15802 , n15801 );
or ( n15803 , n15797 , n15802 );
nand ( n15804 , n15732 , n12969 );
nand ( n15805 , n15803 , n15804 );
xor ( n15806 , n15796 , n15805 );
xor ( n15807 , n15782 , n15806 );
not ( n15808 , n12650 );
not ( n15809 , n12467 );
not ( n15810 , n12422 );
or ( n15811 , n15809 , n15810 );
nand ( n85519 , n12419 , n499 );
nand ( n15813 , n15811 , n85519 );
not ( n15814 , n15813 );
or ( n15815 , n15808 , n15814 );
nand ( n15816 , n85281 , n12702 );
nand ( n15817 , n15815 , n15816 );
and ( n15818 , n15594 , n15604 );
not ( n15819 , n12638 );
xor ( n15820 , n491 , n12492 );
xnor ( n15821 , n15820 , n12500 );
not ( n15822 , n15821 );
or ( n15823 , n15819 , n15822 );
nand ( n15824 , n15587 , n12595 );
nand ( n15825 , n15823 , n15824 );
xor ( n15826 , n15818 , n15825 );
and ( n15827 , n12774 , n489 );
not ( n15828 , n12795 );
not ( n15829 , n489 );
not ( n15830 , n12981 );
or ( n15831 , n15829 , n15830 );
nand ( n15832 , n12980 , n12560 );
nand ( n15833 , n15831 , n15832 );
not ( n15834 , n15833 );
or ( n15835 , n15828 , n15834 );
nand ( n15836 , n15602 , n12542 );
nand ( n15837 , n15835 , n15836 );
xor ( n15838 , n15827 , n15837 );
xor ( n15839 , n15826 , n15838 );
xor ( n15840 , n15817 , n15839 );
xor ( n15841 , n15718 , n15722 );
and ( n15842 , n15841 , n15734 );
and ( n15843 , n15718 , n15722 );
or ( n15844 , n15842 , n15843 );
xor ( n15845 , n15840 , n15844 );
xor ( n15846 , n15807 , n15845 );
xor ( n15847 , n15617 , n15702 );
and ( n15848 , n15847 , n15707 );
and ( n15849 , n15617 , n15702 );
or ( n15850 , n15848 , n15849 );
not ( n15851 , n12470 );
not ( n15852 , n497 );
not ( n15853 , n13372 );
not ( n15854 , n15853 );
or ( n15855 , n15852 , n15854 );
nand ( n15856 , n13046 , n12486 );
nand ( n15857 , n15855 , n15856 );
not ( n15858 , n15857 );
or ( n15859 , n15851 , n15858 );
nand ( n15860 , n15574 , n12517 );
nand ( n15861 , n15859 , n15860 );
nand ( n15862 , n15539 , n12856 , n12843 );
nand ( n15863 , n15615 , n12822 );
nand ( n15864 , n15543 , n12843 , n501 );
nand ( n15865 , n15862 , n15863 , n15864 );
xor ( n85573 , n15861 , n15865 );
or ( n15870 , n15699 , n12461 );
xor ( n85575 , n15636 , n15654 );
and ( n15872 , n85575 , n15659 );
and ( n15873 , n15636 , n15654 );
or ( n15874 , n15872 , n15873 );
xor ( n15875 , n15637 , n15644 );
and ( n15876 , n15875 , n85360 );
and ( n15877 , n15637 , n15644 );
or ( n15878 , n15876 , n15877 );
not ( n15879 , n85360 );
xor ( n15880 , n15878 , n15879 );
not ( n15881 , n10127 );
or ( n15882 , n15881 , n15641 );
xnor ( n15883 , n457 , n521 );
or ( n15884 , n10067 , n15883 );
nand ( n15885 , n15882 , n15884 );
and ( n15886 , n457 , n523 );
xor ( n15887 , n15885 , n15886 );
not ( n15888 , n10094 );
not ( n15889 , n15888 );
not ( n15890 , n10086 );
or ( n15891 , n15889 , n15890 );
nand ( n15892 , n15891 , n459 );
xor ( n15893 , n15887 , n15892 );
xor ( n15894 , n15880 , n15893 );
nor ( n85599 , n15874 , n15894 );
not ( n15899 , n85599 );
nand ( n15900 , n15874 , n15894 );
nand ( n15901 , n15899 , n15900 );
nand ( n15902 , n15509 , n15661 );
nor ( n15903 , n15902 , n15671 );
nand ( n15904 , n12316 , n15903 );
not ( n15905 , n15904 );
buf ( n15906 , n12434 );
nand ( n15907 , n15905 , n15906 );
or ( n15908 , n15907 , n15528 );
not ( n15909 , n12412 );
not ( n15910 , n15903 );
nor ( n15911 , n15909 , n15910 );
and ( n15912 , n15911 , n12352 );
not ( n15913 , n15661 );
not ( n15914 , n15680 );
or ( n15915 , n15913 , n15914 );
nand ( n15916 , n15915 , n15662 );
nor ( n15917 , n15912 , n15916 );
nand ( n15918 , n15908 , n15917 );
not ( n15919 , n15527 );
nor ( n15920 , n12439 , n15904 );
not ( n15921 , n15920 );
or ( n15922 , n15919 , n15921 );
and ( n15923 , n12336 , n12410 );
nor ( n15924 , n15923 , n15910 );
nand ( n15925 , n15527 , n15924 );
nand ( n15926 , n15922 , n15925 );
nor ( n15927 , n15918 , n15926 );
xor ( n15928 , n15901 , n15927 );
and ( n15929 , n12457 , n15928 );
not ( n15930 , n12457 );
not ( n15931 , n15928 );
and ( n15932 , n15930 , n15931 );
nor ( n15933 , n15929 , n15932 );
or ( n15934 , n15933 , n14990 );
nand ( n15935 , n15870 , n15934 );
xor ( n15936 , n85573 , n15935 );
xor ( n15937 , n15850 , n15936 );
xor ( n15938 , n15735 , n15739 );
and ( n15939 , n15938 , n15744 );
and ( n15940 , n15735 , n15739 );
or ( n15941 , n15939 , n15940 );
xor ( n15942 , n15937 , n15941 );
xor ( n15943 , n15846 , n15942 );
xor ( n15944 , n15607 , n15708 );
and ( n15945 , n15944 , n15745 );
and ( n15946 , n15607 , n15708 );
or ( n15947 , n15945 , n15946 );
xor ( n15948 , n15943 , n15947 );
xor ( n15949 , n15376 , n15557 );
and ( n15950 , n15949 , n15746 );
and ( n15951 , n15376 , n15557 );
or ( n15952 , n15950 , n15951 );
or ( n15953 , n15948 , n15952 );
nand ( n15954 , n15948 , n15952 );
nand ( n15955 , n15953 , n15954 );
xnor ( n15956 , n15778 , n15955 );
nand ( n15957 , n10061 , n15956 );
nand ( n15958 , n10060 , n15957 );
and ( n15959 , n15958 , n471 );
not ( n15960 , n9263 );
not ( n15961 , n9911 );
buf ( n15962 , n9915 );
not ( n15963 , n15962 );
or ( n15964 , n15961 , n15963 );
nand ( n15965 , n15964 , n454 );
and ( n15966 , n15960 , n15965 );
not ( n15967 , n15960 );
nand ( n15968 , n454 , n9911 , n15962 );
and ( n15969 , n15967 , n15968 );
nor ( n15970 , n15966 , n15969 );
not ( n15971 , n15970 );
not ( n15972 , n15332 );
not ( n15973 , n15318 );
not ( n15974 , n15303 );
not ( n15975 , n15262 );
or ( n15976 , n15974 , n15975 );
not ( n15977 , n15316 );
nand ( n15978 , n15976 , n15977 );
not ( n15979 , n15978 );
or ( n85681 , n15973 , n15979 );
buf ( n15981 , n15326 );
nand ( n15982 , n85681 , n15981 );
not ( n15983 , n15982 );
or ( n15984 , n15972 , n15983 );
not ( n15985 , n13677 );
nand ( n15986 , n15984 , n15985 );
not ( n15987 , n13679 );
nand ( n15988 , n15987 , n83176 );
not ( n15989 , n15988 );
and ( n15990 , n15986 , n15989 );
not ( n15991 , n15986 );
and ( n15992 , n15991 , n15988 );
nor ( n15993 , n15990 , n15992 );
nand ( n15994 , n15993 , n10061 );
nand ( n15995 , n15971 , n15994 );
and ( n15996 , n15995 , n469 );
not ( n15997 , n10061 );
not ( n15998 , n15769 );
not ( n15999 , n15998 );
not ( n16000 , n15333 );
not ( n16001 , n15982 );
or ( n16002 , n16000 , n16001 );
nand ( n16003 , n16002 , n13680 );
not ( n16004 , n16003 );
or ( n16005 , n15999 , n16004 );
nand ( n16006 , n16005 , n15773 );
not ( n16007 , n15772 );
nor ( n16008 , n16007 , n15776 );
and ( n16009 , n16006 , n16008 );
not ( n16010 , n16006 );
not ( n16011 , n16008 );
and ( n16012 , n16010 , n16011 );
nor ( n16013 , n16009 , n16012 );
not ( n16014 , n16013 );
or ( n16015 , n15997 , n16014 );
buf ( n16016 , n9917 );
not ( n16017 , n16016 );
nor ( n16018 , n9667 , n9679 );
not ( n16019 , n16018 );
not ( n16020 , n16019 );
or ( n16021 , n16017 , n16020 );
not ( n16022 , n9911 );
nor ( n16023 , n16022 , n16018 );
nand ( n16024 , n15960 , n16023 );
nand ( n16025 , n16021 , n16024 );
nand ( n16026 , n9902 , n9919 );
not ( n16027 , n16026 );
and ( n16028 , n16025 , n16027 );
not ( n16029 , n16025 );
and ( n16030 , n16029 , n16026 );
nor ( n16031 , n16028 , n16030 );
nand ( n16032 , n16031 , n454 );
nand ( n16033 , n16015 , n16032 );
and ( n16034 , n16033 , n471 );
xor ( n16035 , n15996 , n16034 );
not ( n16036 , n454 );
not ( n16037 , n9911 );
not ( n16038 , n15960 );
or ( n16039 , n16037 , n16038 );
nand ( n16040 , n16039 , n15962 );
and ( n16041 , n16019 , n9916 );
xor ( n16042 , n16040 , n16041 );
not ( n16043 , n16042 );
or ( n16044 , n16036 , n16043 );
nand ( n16045 , n15998 , n15773 );
xnor ( n16046 , n16003 , n16045 );
nand ( n85748 , n16046 , n10061 );
nand ( n16048 , n16044 , n85748 );
and ( n16049 , n16048 , n470 );
and ( n16050 , n16035 , n16049 );
and ( n16051 , n15996 , n16034 );
or ( n16052 , n16050 , n16051 );
xor ( n16053 , n15959 , n16052 );
and ( n16054 , n16033 , n470 );
not ( n16055 , n16048 );
not ( n16056 , n469 );
nor ( n16057 , n16055 , n16056 );
xor ( n16058 , n16054 , n16057 );
buf ( n16059 , n10049 );
not ( n16060 , n16059 );
not ( n16061 , n16060 );
not ( n16062 , n9923 );
or ( n16063 , n16061 , n16062 );
nand ( n16064 , n16063 , n10052 );
xor ( n16065 , n79793 , n10038 );
and ( n16066 , n16065 , n10043 );
and ( n16067 , n79793 , n10038 );
or ( n16068 , n16066 , n16067 );
xor ( n16069 , n9940 , n9951 );
and ( n16070 , n16069 , n9958 );
and ( n16071 , n9940 , n9951 );
or ( n16072 , n16070 , n16071 );
not ( n16073 , n9595 );
and ( n16074 , n6440 , n4938 );
not ( n16075 , n6440 );
and ( n16076 , n16075 , n543 );
or ( n16077 , n16074 , n16076 );
not ( n16078 , n16077 );
or ( n16079 , n16073 , n16078 );
nand ( n16080 , n9965 , n4445 );
nand ( n16081 , n16079 , n16080 );
not ( n16082 , n541 );
not ( n16083 , n6847 );
or ( n16084 , n16082 , n16083 );
nand ( n16085 , n6843 , n5538 );
nand ( n16086 , n16084 , n16085 );
not ( n16087 , n16086 );
not ( n16088 , n5590 );
or ( n16089 , n16087 , n16088 );
nand ( n16090 , n9935 , n9938 );
nand ( n16091 , n16089 , n16090 );
xor ( n16092 , n16081 , n16091 );
xor ( n16093 , n10006 , n10008 );
and ( n16094 , n16093 , n10021 );
and ( n85796 , n10006 , n10008 );
or ( n16099 , n16094 , n85796 );
xor ( n85798 , n16092 , n16099 );
xor ( n16101 , n16072 , n85798 );
not ( n16102 , n4433 );
not ( n16103 , n539 );
not ( n16104 , n5265 );
or ( n16105 , n16103 , n16104 );
nand ( n16106 , n5264 , n4251 );
nand ( n16107 , n16105 , n16106 );
not ( n16108 , n16107 );
or ( n16109 , n16102 , n16108 );
nand ( n16110 , n9998 , n4224 );
nand ( n16111 , n16109 , n16110 );
not ( n16112 , n5399 );
not ( n16113 , n545 );
not ( n16114 , n9735 );
or ( n16115 , n16113 , n16114 );
nand ( n16116 , n9734 , n4440 );
nand ( n16117 , n16115 , n16116 );
not ( n16118 , n16117 );
or ( n16119 , n16112 , n16118 );
nand ( n16120 , n9949 , n5137 );
nand ( n16121 , n16119 , n16120 );
xor ( n16122 , n16111 , n16121 );
not ( n16123 , n6489 );
not ( n16124 , n9954 );
or ( n16125 , n16123 , n16124 );
not ( n85824 , n7018 );
not ( n16130 , n79653 );
or ( n16131 , n85824 , n16130 );
nand ( n16132 , n9848 , n549 );
nand ( n16133 , n16131 , n16132 );
nand ( n16134 , n16133 , n5905 );
nand ( n16135 , n16125 , n16134 );
xor ( n16136 , n16122 , n16135 );
xor ( n16137 , n16101 , n16136 );
not ( n16138 , n6811 );
and ( n16139 , n547 , n9557 );
not ( n16140 , n547 );
not ( n16141 , n9557 );
and ( n16142 , n16140 , n16141 );
or ( n16143 , n16139 , n16142 );
not ( n16144 , n16143 );
or ( n16145 , n16138 , n16144 );
nand ( n16146 , n9983 , n6854 );
nand ( n16147 , n16145 , n16146 );
not ( n16148 , n5501 );
and ( n16149 , n4937 , n5409 );
not ( n16150 , n4937 );
and ( n16151 , n16150 , n537 );
or ( n16152 , n16149 , n16151 );
not ( n16153 , n16152 );
or ( n16154 , n16148 , n16153 );
buf ( n16155 , n5413 );
nand ( n16156 , n10016 , n16155 );
nand ( n16157 , n16154 , n16156 );
and ( n16158 , n10010 , n10020 );
xor ( n16159 , n16157 , n16158 );
nand ( n16160 , n7786 , n537 );
nand ( n16161 , n8878 , n9991 );
or ( n16162 , n16160 , n16161 );
nand ( n16163 , n16160 , n16161 );
nand ( n16164 , n16162 , n16163 );
xor ( n16165 , n16159 , n16164 );
xor ( n16166 , n16147 , n16165 );
xor ( n16167 , n9970 , n9974 );
and ( n16168 , n16167 , n9985 );
and ( n16169 , n9970 , n9974 );
or ( n16170 , n16168 , n16169 );
xor ( n16171 , n16166 , n16170 );
xor ( n16172 , n9992 , n10022 );
and ( n16173 , n16172 , n10027 );
and ( n16174 , n9992 , n10022 );
or ( n16175 , n16173 , n16174 );
xor ( n16176 , n16171 , n16175 );
xor ( n16177 , n9928 , n9959 );
and ( n16178 , n16177 , n9986 );
and ( n16179 , n9928 , n9959 );
or ( n16180 , n16178 , n16179 );
xor ( n16181 , n16176 , n16180 );
xor ( n16182 , n16137 , n16181 );
xor ( n16183 , n10028 , n10032 );
and ( n16184 , n16183 , n10037 );
and ( n16185 , n10028 , n10032 );
or ( n16186 , n16184 , n16185 );
xor ( n16187 , n16182 , n16186 );
nand ( n16188 , n16068 , n16187 );
not ( n16189 , n16187 );
not ( n16190 , n16068 );
nand ( n16191 , n16189 , n16190 );
nand ( n16192 , n16188 , n16191 );
not ( n16193 , n16192 );
and ( n16194 , n16064 , n16193 );
not ( n16195 , n16064 );
and ( n16196 , n16195 , n16192 );
nor ( n16197 , n16194 , n16196 );
nand ( n16198 , n16197 , n454 );
not ( n16199 , n15953 );
not ( n16200 , n15778 );
or ( n16201 , n16199 , n16200 );
not ( n16202 , n15344 );
not ( n16203 , n15791 );
or ( n16204 , n16202 , n16203 );
not ( n16205 , n493 );
not ( n16206 , n13357 );
or ( n16207 , n16205 , n16206 );
nand ( n16208 , n12674 , n12775 );
nand ( n16209 , n16207 , n16208 );
nand ( n16210 , n16209 , n12758 );
nand ( n85906 , n16204 , n16210 );
not ( n16212 , n12969 );
not ( n16213 , n15801 );
or ( n16214 , n16212 , n16213 );
not ( n16215 , n495 );
nand ( n16216 , n16215 , n13369 );
not ( n16217 , n16216 );
nand ( n16218 , n13370 , n495 );
not ( n16219 , n16218 );
or ( n16220 , n16217 , n16219 );
nand ( n16221 , n16220 , n13032 );
nand ( n16222 , n16214 , n16221 );
xor ( n16223 , n85906 , n16222 );
not ( n16224 , n12517 );
not ( n16225 , n15857 );
or ( n16226 , n16224 , n16225 );
not ( n16227 , n12486 );
not ( n16228 , n15566 );
or ( n16229 , n16227 , n16228 );
nand ( n16230 , n15563 , n497 );
nand ( n16231 , n16229 , n16230 );
nand ( n16232 , n16231 , n12470 );
nand ( n16233 , n16226 , n16232 );
xor ( n16234 , n16223 , n16233 );
xor ( n16235 , n15861 , n15865 );
and ( n16236 , n16235 , n15935 );
and ( n16237 , n15861 , n15865 );
or ( n16238 , n16236 , n16237 );
xor ( n16239 , n16234 , n16238 );
xor ( n16240 , n15817 , n15839 );
and ( n16241 , n16240 , n15844 );
and ( n16242 , n15817 , n15839 );
or ( n16243 , n16241 , n16242 );
xor ( n16244 , n16239 , n16243 );
xor ( n16245 , n15850 , n15936 );
and ( n16246 , n16245 , n15941 );
and ( n16247 , n15850 , n15936 );
or ( n16248 , n16246 , n16247 );
xor ( n16249 , n16244 , n16248 );
not ( n16250 , n15664 );
not ( n16251 , n15683 );
or ( n16252 , n16250 , n16251 );
nand ( n16253 , n16252 , n15689 );
nand ( n16254 , n12843 , n501 );
or ( n16255 , n16253 , n16254 );
not ( n16256 , n15539 );
not ( n16257 , n12821 );
nor ( n16258 , n16257 , n12856 );
nand ( n16259 , n16256 , n16258 );
nor ( n16260 , n15210 , n501 );
nand ( n16261 , n15696 , n16260 );
nand ( n16262 , n15539 , n14691 );
nand ( n16263 , n16255 , n16259 , n16261 , n16262 );
xor ( n16264 , n15818 , n15825 );
and ( n16265 , n16264 , n15838 );
and ( n16266 , n15818 , n15825 );
or ( n16267 , n16265 , n16266 );
xor ( n16268 , n16263 , n16267 );
not ( n16269 , n12702 );
not ( n85965 , n15813 );
or ( n16271 , n16269 , n85965 );
and ( n16272 , n13258 , n12467 );
not ( n16273 , n13258 );
and ( n16274 , n16273 , n499 );
nor ( n16275 , n16272 , n16274 );
or ( n16276 , n16275 , n12649 );
nand ( n16277 , n16271 , n16276 );
xor ( n16278 , n16268 , n16277 );
not ( n16279 , n504 );
not ( n16280 , n503 );
or ( n16281 , n15918 , n15926 );
xor ( n16282 , n15878 , n15879 );
and ( n16283 , n16282 , n15893 );
and ( n16284 , n15878 , n15879 );
or ( n16285 , n16283 , n16284 );
or ( n16286 , n15881 , n15883 );
or ( n16287 , n10067 , n2714 );
nand ( n16288 , n16286 , n16287 );
nand ( n16289 , n522 , n457 );
xor ( n16290 , n16288 , n16289 );
xor ( n16291 , n15885 , n15886 );
and ( n16292 , n16291 , n15892 );
and ( n16293 , n15885 , n15886 );
or ( n16294 , n16292 , n16293 );
xor ( n16295 , n16290 , n16294 );
nor ( n16296 , n16285 , n16295 );
not ( n16297 , n16296 );
not ( n16298 , n16297 );
and ( n16299 , n16285 , n16295 );
nor ( n16300 , n16298 , n16299 );
not ( n16301 , n16300 );
not ( n16302 , n15900 );
and ( n16303 , n16301 , n16302 );
and ( n16304 , n16300 , n15900 , n85599 );
nor ( n16305 , n16303 , n16304 );
or ( n16306 , n16300 , n85599 );
nand ( n16307 , n16281 , n16305 , n16306 );
not ( n16308 , n15918 );
not ( n16309 , n15900 );
not ( n16310 , n16300 );
or ( n16311 , n16309 , n16310 );
nand ( n16312 , n16311 , n16305 );
nor ( n16313 , n15926 , n16312 );
nand ( n86009 , n16308 , n16313 );
nand ( n16318 , n16307 , n86009 );
not ( n86011 , n16318 );
or ( n16320 , n16280 , n86011 );
not ( n16321 , n16318 );
nand ( n16322 , n16321 , n12457 );
nand ( n16323 , n16320 , n16322 );
not ( n16324 , n16323 );
or ( n16325 , n16279 , n16324 );
not ( n16326 , n15933 );
nand ( n16327 , n16326 , n12462 );
nand ( n16328 , n16325 , n16327 );
not ( n16329 , n12595 );
not ( n16330 , n15821 );
or ( n16331 , n16329 , n16330 );
xor ( n16332 , n12481 , n12610 );
or ( n16333 , n16332 , n12593 );
nand ( n16334 , n16331 , n16333 );
and ( n16335 , n15837 , n15827 );
xor ( n16336 , n16334 , n16335 );
not ( n16337 , n489 );
nor ( n16338 , n16337 , n12950 );
not ( n16339 , n12795 );
xor ( n16340 , n13008 , n12560 );
not ( n16341 , n16340 );
not ( n16342 , n16341 );
or ( n16343 , n16339 , n16342 );
nand ( n16344 , n15833 , n12542 );
nand ( n16345 , n16343 , n16344 );
xor ( n16346 , n16338 , n16345 );
xor ( n86039 , n16336 , n16346 );
xor ( n16351 , n16328 , n86039 );
xor ( n16352 , n15786 , n15795 );
and ( n16353 , n16352 , n15805 );
and ( n16354 , n15786 , n15795 );
or ( n16355 , n16353 , n16354 );
xor ( n16356 , n16351 , n16355 );
xor ( n16357 , n16278 , n16356 );
xor ( n16358 , n15782 , n15806 );
and ( n16359 , n16358 , n15845 );
and ( n16360 , n15782 , n15806 );
or ( n16361 , n16359 , n16360 );
xor ( n16362 , n16357 , n16361 );
xor ( n16363 , n16249 , n16362 );
xor ( n16364 , n15846 , n15942 );
and ( n16365 , n16364 , n15947 );
and ( n16366 , n15846 , n15942 );
or ( n16367 , n16365 , n16366 );
nand ( n16368 , n16363 , n16367 );
buf ( n16369 , n16368 );
not ( n16370 , n16369 );
nor ( n16371 , n16363 , n16367 );
buf ( n16372 , n16371 );
nor ( n16373 , n16370 , n16372 );
not ( n16374 , n15954 );
nor ( n16375 , n16373 , n16374 );
nand ( n16376 , n16201 , n16375 );
and ( n16377 , n16373 , n16374 );
nor ( n16378 , n16377 , n454 );
nand ( n16379 , n15953 , n15778 , n16373 );
nand ( n16380 , n16376 , n16378 , n16379 );
nand ( n16381 , n16198 , n16380 );
not ( n16382 , n16381 );
not ( n16383 , n472 );
nor ( n16384 , n16382 , n16383 );
xor ( n16385 , n16058 , n16384 );
and ( n16386 , n16053 , n16385 );
and ( n16387 , n15959 , n16052 );
or ( n16388 , n16386 , n16387 );
not ( n16389 , n16388 );
nor ( n16390 , n16187 , n16068 );
nor ( n16391 , n16390 , n10049 );
not ( n16392 , n16391 );
not ( n16393 , n9923 );
or ( n16394 , n16392 , n16393 );
nand ( n16395 , n16188 , n10051 );
nand ( n16396 , n16395 , n16191 );
buf ( n16397 , n16396 );
nand ( n16398 , n16394 , n16397 );
xor ( n16399 , n16137 , n16181 );
and ( n16400 , n16399 , n16186 );
and ( n16401 , n16137 , n16181 );
or ( n16402 , n16400 , n16401 );
xor ( n16403 , n16111 , n16121 );
and ( n16404 , n16403 , n16135 );
and ( n16405 , n16111 , n16121 );
or ( n16406 , n16404 , n16405 );
not ( n16407 , n9938 );
not ( n16408 , n16086 );
or ( n16409 , n16407 , n16408 );
not ( n16410 , n541 );
not ( n16411 , n6479 );
or ( n16412 , n16410 , n16411 );
nand ( n16413 , n6478 , n5538 );
nand ( n16414 , n16412 , n16413 );
nand ( n16415 , n16414 , n5590 );
nand ( n16416 , n16409 , n16415 );
not ( n16417 , n5399 );
and ( n16418 , n9382 , n545 );
not ( n16419 , n9382 );
and ( n16420 , n16419 , n4440 );
or ( n16421 , n16418 , n16420 );
not ( n16422 , n16421 );
or ( n16423 , n16417 , n16422 );
nand ( n16424 , n16117 , n75018 );
nand ( n16425 , n16423 , n16424 );
xor ( n16426 , n16416 , n16425 );
not ( n16427 , n6489 );
not ( n86117 , n16133 );
or ( n16429 , n16427 , n86117 );
nand ( n16430 , n16429 , n7020 );
xor ( n16431 , n16426 , n16430 );
xor ( n16432 , n16406 , n16431 );
not ( n16433 , n4224 );
not ( n16434 , n16107 );
or ( n16435 , n16433 , n16434 );
nand ( n16436 , n539 , n9931 );
not ( n16437 , n16436 );
not ( n16438 , n9931 );
nand ( n16439 , n16438 , n4251 );
not ( n16440 , n16439 );
or ( n16441 , n16437 , n16440 );
nand ( n16442 , n16441 , n4221 );
nand ( n16443 , n16435 , n16442 );
not ( n16444 , n5128 );
not ( n16445 , n543 );
not ( n16446 , n6796 );
or ( n16447 , n16445 , n16446 );
nand ( n16448 , n76644 , n4938 );
nand ( n16449 , n16447 , n16448 );
not ( n16450 , n16449 );
or ( n16451 , n16444 , n16450 );
nand ( n16452 , n4445 , n16077 );
nand ( n16453 , n16451 , n16452 );
xor ( n16454 , n16443 , n16453 );
not ( n16455 , n6854 );
not ( n16456 , n16143 );
or ( n16457 , n16455 , n16456 );
xor ( n16458 , n547 , n9553 );
nand ( n16459 , n16458 , n6811 );
nand ( n16460 , n16457 , n16459 );
xor ( n16461 , n16454 , n16460 );
xor ( n16462 , n16432 , n16461 );
not ( n16463 , n16155 );
not ( n16464 , n16152 );
or ( n16465 , n16463 , n16464 );
not ( n16466 , n537 );
not ( n16467 , n7911 );
or ( n16468 , n16466 , n16467 );
nand ( n16469 , n6937 , n5409 );
nand ( n16470 , n16468 , n16469 );
nand ( n16471 , n16470 , n5501 );
nand ( n16472 , n16465 , n16471 );
nand ( n16473 , n77458 , n537 );
xor ( n16474 , n16472 , n16473 );
xor ( n16475 , n16474 , n16163 );
xor ( n16476 , n16157 , n16158 );
and ( n16477 , n16476 , n16164 );
and ( n16478 , n16157 , n16158 );
or ( n16479 , n16477 , n16478 );
xor ( n16480 , n16475 , n16479 );
xor ( n16481 , n16081 , n16091 );
and ( n16482 , n16481 , n16099 );
and ( n16483 , n16081 , n16091 );
or ( n16484 , n16482 , n16483 );
xor ( n86174 , n16480 , n16484 );
xor ( n16486 , n16147 , n16165 );
and ( n16487 , n16486 , n16170 );
and ( n16488 , n16147 , n16165 );
or ( n16489 , n16487 , n16488 );
xor ( n16490 , n86174 , n16489 );
xor ( n16491 , n16072 , n85798 );
and ( n16492 , n16491 , n16136 );
and ( n16493 , n16072 , n85798 );
or ( n16494 , n16492 , n16493 );
xor ( n16495 , n16490 , n16494 );
xor ( n16496 , n16462 , n16495 );
xor ( n16497 , n16171 , n16175 );
and ( n16498 , n16497 , n16180 );
and ( n16499 , n16171 , n16175 );
or ( n16500 , n16498 , n16499 );
xor ( n16501 , n16496 , n16500 );
nor ( n16502 , n16402 , n16501 );
buf ( n16503 , n16502 );
not ( n16504 , n16503 );
buf ( n16505 , n16501 );
nand ( n16506 , n16402 , n16505 );
nand ( n16507 , n16504 , n16506 );
not ( n16508 , n16507 );
and ( n16509 , n16398 , n16508 );
not ( n16510 , n16398 );
and ( n16511 , n16510 , n16507 );
nor ( n16512 , n16509 , n16511 );
not ( n16513 , n16512 );
not ( n16514 , n454 );
or ( n16515 , n16513 , n16514 );
not ( n16516 , n15953 );
nor ( n16517 , n16516 , n16372 );
not ( n16518 , n16517 );
not ( n16519 , n15778 );
or ( n16520 , n16518 , n16519 );
nor ( n16521 , n16371 , n15954 );
not ( n16522 , n16521 );
and ( n86212 , n16369 , n16522 );
nand ( n16527 , n16520 , n86212 );
not ( n86214 , n13032 );
and ( n16529 , n495 , n12886 );
not ( n16530 , n495 );
and ( n16531 , n16530 , n13372 );
or ( n16532 , n16529 , n16531 );
not ( n16533 , n16532 );
or ( n16534 , n86214 , n16533 );
not ( n16535 , n16218 );
not ( n16536 , n16216 );
or ( n16537 , n16535 , n16536 );
nand ( n16538 , n16537 , n12969 );
nand ( n16539 , n16534 , n16538 );
not ( n16540 , n12758 );
not ( n16541 , n493 );
not ( n16542 , n82600 );
or ( n16543 , n16541 , n16542 );
or ( n16544 , n82600 , n493 );
nand ( n16545 , n16543 , n16544 );
not ( n16546 , n16545 );
or ( n16547 , n16540 , n16546 );
nand ( n16548 , n16209 , n15344 );
nand ( n16549 , n16547 , n16548 );
xor ( n16550 , n16539 , n16549 );
not ( n16551 , n12822 );
and ( n16552 , n501 , n15690 );
not ( n16553 , n501 );
and ( n86240 , n16553 , n15697 );
nor ( n16558 , n16552 , n86240 );
not ( n16559 , n16558 );
or ( n16560 , n16551 , n16559 );
and ( n16561 , n15928 , n12856 );
not ( n16562 , n15928 );
and ( n16563 , n16562 , n501 );
or ( n16564 , n16561 , n16563 );
nand ( n16565 , n16564 , n12843 );
nand ( n16566 , n16560 , n16565 );
xor ( n16567 , n16550 , n16566 );
xor ( n16568 , n16263 , n16267 );
and ( n16569 , n16568 , n16277 );
and ( n16570 , n16263 , n16267 );
or ( n16571 , n16569 , n16570 );
xor ( n16572 , n16567 , n16571 );
not ( n16573 , n15438 );
nor ( n16574 , n12469 , n497 );
nand ( n16575 , n16573 , n16574 );
nand ( n16576 , n16231 , n12517 );
nand ( n16577 , n12470 , n497 );
or ( n16578 , n12418 , n16577 );
nand ( n16579 , n16575 , n16576 , n16578 );
xor ( n16580 , n16334 , n16335 );
and ( n16581 , n16580 , n16346 );
and ( n16582 , n16334 , n16335 );
or ( n16583 , n16581 , n16582 );
xor ( n16584 , n16579 , n16583 );
not ( n16585 , n12649 );
not ( n16586 , n499 );
not ( n16587 , n16256 );
or ( n16588 , n16586 , n16587 );
nand ( n16589 , n15539 , n1077 );
nand ( n16590 , n16588 , n16589 );
nand ( n16591 , n16585 , n16590 );
not ( n16592 , n16275 );
nand ( n16593 , n16592 , n12702 );
nand ( n16594 , n16591 , n16593 );
xor ( n16595 , n16584 , n16594 );
xor ( n16596 , n16572 , n16595 );
xor ( n16597 , n16328 , n86039 );
and ( n16598 , n16597 , n16355 );
and ( n16599 , n16328 , n86039 );
or ( n16600 , n16598 , n16599 );
not ( n16601 , n504 );
not ( n16602 , n503 );
or ( n16603 , n15662 , n85599 );
nand ( n16604 , n16603 , n15900 );
and ( n16605 , n16604 , n16297 );
nor ( n16606 , n16605 , n16299 );
not ( n16607 , n16606 );
xor ( n16608 , n16288 , n16289 );
and ( n16609 , n16608 , n16294 );
and ( n16610 , n16288 , n16289 );
or ( n16611 , n16609 , n16610 );
not ( n16612 , n16289 );
nand ( n16613 , n521 , n457 );
not ( n16614 , n16613 );
or ( n16615 , n10127 , n10068 );
nand ( n16616 , n16615 , n457 );
not ( n16617 , n16616 );
or ( n16618 , n16614 , n16617 );
or ( n16619 , n16616 , n16613 );
nand ( n16620 , n16618 , n16619 );
not ( n16621 , n16620 );
or ( n16622 , n16612 , n16621 );
or ( n16623 , n16620 , n16289 );
nand ( n16624 , n16622 , n16623 );
xnor ( n16625 , n16611 , n16624 );
nor ( n16626 , n16607 , n16625 );
not ( n16627 , n16626 );
not ( n16628 , n15681 );
not ( n16629 , n15674 );
or ( n86313 , n16628 , n16629 );
not ( n16631 , n15661 );
nor ( n16632 , n16631 , n16296 , n85599 );
nand ( n16633 , n86313 , n16632 );
not ( n16634 , n16633 );
or ( n16635 , n16627 , n16634 );
not ( n16636 , n16606 );
not ( n16637 , n16633 );
or ( n16638 , n16636 , n16637 );
xor ( n16639 , n16611 , n16289 );
xor ( n16640 , n16639 , n16620 );
nand ( n16641 , n16638 , n16640 );
nand ( n16642 , n16635 , n16641 );
not ( n16643 , n16642 );
not ( n16644 , n16643 );
or ( n16645 , n16602 , n16644 );
nand ( n16646 , n12423 , n16642 );
nand ( n16647 , n16645 , n16646 );
not ( n16648 , n16647 );
or ( n16649 , n16601 , n16648 );
nand ( n16650 , n16323 , n12462 );
nand ( n16651 , n16649 , n16650 );
xor ( n16652 , n85906 , n16222 );
and ( n16653 , n16652 , n16233 );
and ( n16654 , n85906 , n16222 );
or ( n16655 , n16653 , n16654 );
xor ( n16656 , n16651 , n16655 );
and ( n16657 , n16338 , n16345 );
xor ( n16658 , n491 , n12693 );
not ( n16659 , n16658 );
or ( n16660 , n16659 , n12593 );
not ( n16661 , n16332 );
nand ( n16662 , n16661 , n12595 );
nand ( n16663 , n16660 , n16662 );
xor ( n16664 , n16657 , n16663 );
and ( n16665 , n14099 , n489 );
not ( n16666 , n12580 );
and ( n16667 , n12505 , n12560 );
not ( n16668 , n12505 );
and ( n16669 , n16668 , n489 );
or ( n16670 , n16667 , n16669 );
not ( n16671 , n16670 );
or ( n16672 , n16666 , n16671 );
not ( n16673 , n16340 );
nand ( n16674 , n16673 , n12542 );
nand ( n16675 , n16672 , n16674 );
xor ( n16676 , n16665 , n16675 );
xor ( n16677 , n16664 , n16676 );
xor ( n16678 , n16656 , n16677 );
xor ( n16679 , n16600 , n16678 );
xor ( n16680 , n16234 , n16238 );
and ( n16681 , n16680 , n16243 );
and ( n16682 , n16234 , n16238 );
or ( n16683 , n16681 , n16682 );
xor ( n86367 , n16679 , n16683 );
xor ( n16685 , n16596 , n86367 );
xor ( n16686 , n16278 , n16356 );
and ( n16687 , n16686 , n16361 );
and ( n16688 , n16278 , n16356 );
or ( n16689 , n16687 , n16688 );
xor ( n16690 , n16685 , n16689 );
xor ( n16691 , n16244 , n16248 );
and ( n16692 , n16691 , n16362 );
and ( n16693 , n16244 , n16248 );
or ( n16694 , n16692 , n16693 );
or ( n16695 , n16690 , n16694 );
nand ( n16696 , n16690 , n16694 );
nand ( n16697 , n16695 , n16696 );
not ( n16698 , n16697 );
and ( n16699 , n16527 , n16698 );
not ( n16700 , n16527 );
and ( n16701 , n16700 , n16697 );
nor ( n16702 , n16699 , n16701 );
nand ( n16703 , n16702 , n10061 );
nand ( n16704 , n16515 , n16703 );
and ( n16705 , n16704 , n472 );
xor ( n16706 , n16054 , n16057 );
and ( n16707 , n16706 , n16384 );
and ( n16708 , n16054 , n16057 );
or ( n16709 , n16707 , n16708 );
xor ( n16710 , n16705 , n16709 );
and ( n16711 , n16033 , n469 );
nand ( n16712 , n16198 , n16380 );
and ( n16713 , n16712 , n471 );
xor ( n16714 , n16711 , n16713 );
and ( n16715 , n15958 , n470 );
xor ( n16716 , n16714 , n16715 );
xor ( n16717 , n16710 , n16716 );
not ( n86401 , n16717 );
and ( n16722 , n16389 , n86401 );
xor ( n86403 , n15959 , n16052 );
xor ( n16724 , n86403 , n16385 );
and ( n16725 , n15958 , n472 );
and ( n16726 , n15995 , n470 );
nor ( n16727 , n8169 , n8164 );
not ( n16728 , n454 );
nor ( n16729 , n16727 , n16728 );
or ( n16730 , n7374 , n7600 );
not ( n16731 , n16730 );
buf ( n16732 , n8150 );
not ( n16733 , n16732 );
not ( n16734 , n9261 );
not ( n16735 , n8185 );
not ( n16736 , n16735 );
or ( n16737 , n16734 , n16736 );
not ( n16738 , n8126 );
nand ( n16739 , n16737 , n16738 );
not ( n16740 , n16739 );
or ( n16741 , n16733 , n16740 );
buf ( n16742 , n8160 );
nand ( n16743 , n16741 , n16742 );
not ( n16744 , n16743 );
or ( n16745 , n16731 , n16744 );
nand ( n16746 , n16745 , n8166 );
and ( n86427 , n16729 , n16746 );
nand ( n16751 , n15985 , n15332 );
xnor ( n16752 , n15982 , n16751 );
and ( n16753 , n16752 , n10061 );
nor ( n16754 , n86427 , n16753 );
not ( n16755 , n16746 );
and ( n16756 , n16727 , n454 );
nand ( n16757 , n16755 , n16756 );
nand ( n16758 , n16754 , n16757 );
and ( n16759 , n16758 , n469 );
xor ( n16760 , n16726 , n16759 );
and ( n16761 , n16033 , n472 );
and ( n16762 , n16760 , n16761 );
and ( n16763 , n16726 , n16759 );
or ( n16764 , n16762 , n16763 );
xor ( n16765 , n16725 , n16764 );
xor ( n16766 , n15996 , n16034 );
xor ( n16767 , n16766 , n16049 );
and ( n16768 , n16765 , n16767 );
and ( n16769 , n16725 , n16764 );
or ( n16770 , n16768 , n16769 );
nor ( n16771 , n16724 , n16770 );
nor ( n16772 , n16722 , n16771 );
not ( n16773 , n15252 );
nand ( n16774 , n15257 , n16773 );
xnor ( n16775 , n15121 , n16774 );
nand ( n16776 , n16775 , n10061 );
buf ( n16777 , n9189 );
not ( n16778 , n9235 );
nand ( n16779 , n16777 , n16778 );
not ( n16780 , n9256 );
nand ( n16781 , n16779 , n16780 );
nand ( n16782 , n9258 , n9251 );
nand ( n16783 , n16781 , n16782 , n454 );
not ( n16784 , n16782 );
nand ( n16785 , n16784 , n16779 , n16780 , n454 );
nand ( n16786 , n16776 , n16783 , n16785 );
and ( n16787 , n16786 , n471 );
not ( n16788 , n8619 );
not ( n16789 , n16788 );
not ( n16790 , n8684 );
not ( n16791 , n9173 );
or ( n16792 , n16790 , n16791 );
nand ( n16793 , n16792 , n9177 );
buf ( n16794 , n16793 );
not ( n16795 , n16794 );
or ( n16796 , n16789 , n16795 );
buf ( n16797 , n9181 );
nand ( n16798 , n16796 , n16797 );
not ( n16799 , n16798 );
not ( n16800 , n454 );
not ( n16801 , n8526 );
nand ( n16802 , n16801 , n9186 );
nor ( n16803 , n16800 , n16802 );
nand ( n16804 , n16799 , n16803 );
and ( n16805 , n16802 , n454 );
and ( n16806 , n16798 , n16805 );
nand ( n16807 , n84825 , n15110 );
not ( n16808 , n14530 );
not ( n16809 , n16808 );
buf ( n16810 , n15098 );
not ( n16811 , n16810 );
or ( n16812 , n16809 , n16811 );
nand ( n16813 , n16812 , n15107 );
xnor ( n16814 , n16807 , n16813 );
and ( n16815 , n16814 , n10061 );
nor ( n16816 , n16806 , n16815 );
nand ( n16817 , n16804 , n16816 );
and ( n86495 , n16817 , n469 );
not ( n16819 , n9252 );
nand ( n16820 , n16819 , n9255 );
not ( n16821 , n16820 );
nor ( n16822 , n16821 , n16728 );
not ( n16823 , n16822 );
nand ( n16824 , n16777 , n9234 );
nand ( n16825 , n16824 , n9253 );
not ( n16826 , n16825 );
or ( n16827 , n16823 , n16826 );
nand ( n16828 , n9253 , n454 );
nor ( n16829 , n16820 , n16828 );
and ( n16830 , n16829 , n16824 );
nand ( n16831 , n14283 , n15120 );
xnor ( n16832 , n15117 , n16831 );
and ( n16833 , n16832 , n10061 );
nor ( n16834 , n16830 , n16833 );
nand ( n16835 , n16827 , n16834 );
and ( n16836 , n16835 , n471 );
xor ( n16837 , n86495 , n16836 );
not ( n16838 , n454 );
nand ( n16839 , n9234 , n9253 );
xnor ( n16840 , n16839 , n16777 );
not ( n16841 , n16840 );
or ( n16842 , n16838 , n16841 );
nand ( n16843 , n14351 , n15116 );
xnor ( n16844 , n15113 , n16843 );
nand ( n16845 , n16844 , n10061 );
nand ( n16846 , n16842 , n16845 );
and ( n16847 , n16846 , n470 );
and ( n16848 , n16837 , n16847 );
and ( n16849 , n86495 , n16836 );
or ( n16850 , n16848 , n16849 );
xor ( n16851 , n16787 , n16850 );
and ( n16852 , n16835 , n470 );
and ( n16853 , n16846 , n469 );
xor ( n16854 , n16852 , n16853 );
not ( n16855 , n15232 );
not ( n16856 , n15244 );
or ( n16857 , n16855 , n16856 );
or ( n16858 , n15244 , n15232 );
nand ( n16859 , n16857 , n16858 );
not ( n16860 , n16773 );
not ( n16861 , n15121 );
or ( n16862 , n16860 , n16861 );
nand ( n16863 , n16862 , n15257 );
xnor ( n16864 , n16859 , n16863 );
not ( n16865 , n16864 );
not ( n16866 , n10061 );
or ( n16867 , n16865 , n16866 );
buf ( n16868 , n8184 );
buf ( n16869 , n8123 );
nand ( n16870 , n16868 , n16869 );
not ( n16871 , n454 );
nor ( n86549 , n16870 , n16871 );
buf ( n16873 , n9261 );
or ( n16874 , n86549 , n16873 );
not ( n16875 , n454 );
not ( n16876 , n16870 );
or ( n16877 , n16875 , n16876 );
nand ( n16878 , n16877 , n16873 );
nand ( n16879 , n16874 , n16878 );
nand ( n16880 , n16867 , n16879 );
and ( n16881 , n16880 , n472 );
xor ( n16882 , n16854 , n16881 );
xor ( n16883 , n16851 , n16882 );
and ( n16884 , n16786 , n472 );
nand ( n16885 , n16788 , n16797 );
not ( n16886 , n16885 );
and ( n16887 , n16794 , n16886 );
not ( n16888 , n16794 );
and ( n16889 , n16888 , n16885 );
nor ( n16890 , n16887 , n16889 );
nand ( n16891 , n16890 , n454 );
nand ( n16892 , n16808 , n15107 );
xnor ( n16893 , n16810 , n16892 );
nand ( n16894 , n16893 , n10061 );
nand ( n16895 , n16891 , n16894 );
and ( n16896 , n16895 , n469 );
and ( n16897 , n16817 , n470 );
xor ( n16898 , n16896 , n16897 );
and ( n16899 , n16835 , n472 );
and ( n86577 , n16898 , n16899 );
and ( n16904 , n16896 , n16897 );
or ( n86579 , n86577 , n16904 );
xor ( n16906 , n16884 , n86579 );
xor ( n16907 , n86495 , n16836 );
xor ( n16908 , n16907 , n16847 );
and ( n16909 , n16906 , n16908 );
and ( n16910 , n16884 , n86579 );
or ( n16911 , n16909 , n16910 );
nor ( n16912 , n16883 , n16911 );
xor ( n16913 , n16884 , n86579 );
xor ( n16914 , n16913 , n16908 );
and ( n16915 , n16846 , n471 );
nand ( n16916 , n9177 , n8684 );
not ( n16917 , n16916 );
buf ( n16918 , n9173 );
not ( n16919 , n16918 );
or ( n16920 , n16917 , n16919 );
or ( n16921 , n16918 , n16916 );
nand ( n16922 , n16920 , n16921 );
nand ( n16923 , n16922 , n454 );
not ( n16924 , n15096 );
nand ( n86599 , n16924 , n15093 );
not ( n16929 , n86599 );
not ( n16930 , n14673 );
not ( n16931 , n16930 );
buf ( n16932 , n15090 );
not ( n16933 , n16932 );
or ( n16934 , n16931 , n16933 );
not ( n16935 , n15094 );
nand ( n16936 , n16934 , n16935 );
not ( n16937 , n16936 );
or ( n16938 , n16929 , n16937 );
or ( n16939 , n86599 , n16936 );
nand ( n16940 , n16938 , n16939 );
nand ( n16941 , n10061 , n16940 );
nand ( n16942 , n16923 , n16941 );
and ( n16943 , n16942 , n469 );
and ( n16944 , n16895 , n470 );
xor ( n16945 , n16943 , n16944 );
and ( n16946 , n16817 , n471 );
and ( n16947 , n16945 , n16946 );
and ( n16948 , n16943 , n16944 );
or ( n16949 , n16947 , n16948 );
xor ( n16950 , n16915 , n16949 );
xor ( n16951 , n16896 , n16897 );
xor ( n16952 , n16951 , n16899 );
and ( n16953 , n16950 , n16952 );
and ( n16954 , n16915 , n16949 );
or ( n16955 , n16953 , n16954 );
nor ( n16956 , n16914 , n16955 );
nor ( n16957 , n16912 , n16956 );
not ( n16958 , n16957 );
not ( n16959 , n16958 );
xor ( n16960 , n16915 , n16949 );
xor ( n16961 , n16960 , n16952 );
and ( n16962 , n16846 , n472 );
not ( n16963 , n8745 );
not ( n16964 , n8803 );
nand ( n16965 , n16963 , n16964 );
not ( n16966 , n16965 );
buf ( n16967 , n9162 );
not ( n16968 , n16967 );
or ( n16969 , n16966 , n16968 );
nand ( n16970 , n8745 , n8803 );
nand ( n16971 , n16969 , n16970 );
not ( n16972 , n16971 );
not ( n16973 , n9171 );
nand ( n16974 , n16973 , n9167 );
nor ( n16975 , n16974 , n16728 );
nand ( n16976 , n16972 , n16975 );
and ( n16977 , n16974 , n454 );
and ( n16978 , n16971 , n16977 );
nand ( n16979 , n16935 , n16930 );
xnor ( n16980 , n16932 , n16979 );
and ( n16981 , n16980 , n10061 );
nor ( n16982 , n16978 , n16981 );
nand ( n16983 , n16976 , n16982 );
and ( n16984 , n16983 , n469 );
and ( n16985 , n16942 , n470 );
xor ( n16986 , n16984 , n16985 );
and ( n16987 , n16895 , n471 );
and ( n16988 , n16986 , n16987 );
and ( n16989 , n16984 , n16985 );
or ( n86661 , n16988 , n16989 );
xor ( n16991 , n16962 , n86661 );
xor ( n16992 , n16943 , n16944 );
xor ( n16993 , n16992 , n16946 );
and ( n16994 , n16991 , n16993 );
and ( n16995 , n16962 , n86661 );
or ( n16996 , n16994 , n16995 );
or ( n16997 , n16961 , n16996 );
not ( n16998 , n16997 );
not ( n16999 , n10061 );
not ( n17000 , n14721 );
and ( n17001 , n15086 , n17000 );
not ( n17002 , n15089 );
and ( n17003 , n15086 , n17002 );
nor ( n17004 , n17001 , n17003 );
not ( n17005 , n14716 );
not ( n17006 , n15086 );
nand ( n17007 , n17005 , n17006 , n14719 );
not ( n17008 , n14719 );
nand ( n17009 , n17008 , n17006 , n14716 );
nand ( n17010 , n17004 , n17007 , n17009 );
not ( n17011 , n17010 );
or ( n17012 , n16999 , n17011 );
nand ( n17013 , n16965 , n16970 );
not ( n17014 , n9162 );
and ( n17015 , n17013 , n17014 );
not ( n17016 , n17013 );
and ( n17017 , n17016 , n16967 );
nor ( n17018 , n17015 , n17017 );
nand ( n17019 , n17018 , n454 );
nand ( n17020 , n17012 , n17019 );
and ( n17021 , n17020 , n469 );
and ( n17022 , n16983 , n470 );
xor ( n17023 , n17021 , n17022 );
and ( n17024 , n16942 , n471 );
and ( n17025 , n17023 , n17024 );
and ( n17026 , n17021 , n17022 );
or ( n17027 , n17025 , n17026 );
and ( n17028 , n16817 , n472 );
xor ( n17029 , n17027 , n17028 );
xor ( n17030 , n16984 , n16985 );
xor ( n17031 , n17030 , n16987 );
and ( n86703 , n17029 , n17031 );
and ( n17033 , n17027 , n17028 );
or ( n17034 , n86703 , n17033 );
not ( n17035 , n17034 );
xor ( n17036 , n16962 , n86661 );
xor ( n17037 , n17036 , n16993 );
not ( n17038 , n17037 );
nand ( n17039 , n17035 , n17038 );
not ( n17040 , n17039 );
xor ( n17041 , n17027 , n17028 );
xor ( n17042 , n17041 , n17031 );
and ( n17043 , n16895 , n472 );
nand ( n17044 , n9161 , n8871 );
buf ( n17045 , n9158 );
not ( n17046 , n17045 );
and ( n17047 , n17044 , n17046 );
not ( n17048 , n17044 );
and ( n17049 , n17048 , n17045 );
nor ( n17050 , n17047 , n17049 );
nand ( n17051 , n17050 , n454 );
nand ( n17052 , n14775 , n15085 );
xnor ( n17053 , n15082 , n17052 );
nand ( n17054 , n17053 , n10061 );
nand ( n17055 , n17051 , n17054 );
and ( n86727 , n17055 , n469 );
and ( n17060 , n17020 , n470 );
xor ( n86729 , n86727 , n17060 );
and ( n17062 , n16983 , n471 );
and ( n17063 , n86729 , n17062 );
and ( n17064 , n86727 , n17060 );
or ( n17065 , n17063 , n17064 );
xor ( n17066 , n17043 , n17065 );
xor ( n17067 , n17021 , n17022 );
xor ( n17068 , n17067 , n17024 );
and ( n17069 , n17066 , n17068 );
and ( n17070 , n17043 , n17065 );
or ( n17071 , n17069 , n17070 );
or ( n17072 , n17042 , n17071 );
not ( n17073 , n17072 );
and ( n17074 , n16942 , n472 );
not ( n17075 , n10061 );
nand ( n17076 , n15075 , n84803 );
xnor ( n17077 , n17076 , n15065 );
not ( n17078 , n17077 );
or ( n17079 , n17075 , n17078 );
not ( n17080 , n8874 );
not ( n17081 , n8910 );
nand ( n17082 , n17080 , n17081 );
nand ( n17083 , n17082 , n78975 );
not ( n17084 , n8974 );
not ( n86753 , n9151 );
or ( n17089 , n17084 , n86753 );
not ( n17090 , n9154 );
nand ( n17091 , n17089 , n17090 );
not ( n17092 , n17091 );
and ( n17093 , n17083 , n17092 );
not ( n17094 , n17083 );
and ( n17095 , n17094 , n17091 );
nor ( n17096 , n17093 , n17095 );
nand ( n17097 , n17096 , n454 );
nand ( n17098 , n17079 , n17097 );
and ( n17099 , n17098 , n469 );
and ( n17100 , n17055 , n470 );
xor ( n17101 , n17099 , n17100 );
and ( n17102 , n17020 , n471 );
and ( n17103 , n17101 , n17102 );
and ( n17104 , n17099 , n17100 );
or ( n17105 , n17103 , n17104 );
xor ( n17106 , n17074 , n17105 );
xor ( n17107 , n86727 , n17060 );
xor ( n17108 , n17107 , n17062 );
and ( n17109 , n17106 , n17108 );
and ( n17110 , n17074 , n17105 );
or ( n17111 , n17109 , n17110 );
not ( n17112 , n17111 );
xor ( n17113 , n17043 , n17065 );
xor ( n17114 , n17113 , n17068 );
not ( n17115 , n17114 );
nand ( n17116 , n17112 , n17115 );
not ( n17117 , n17116 );
xor ( n17118 , n17074 , n17105 );
xor ( n17119 , n17118 , n17108 );
not ( n17120 , n17119 );
and ( n17121 , n16983 , n472 );
nand ( n17122 , n8974 , n9153 );
not ( n17123 , n17122 );
xor ( n17124 , n9151 , n17123 );
not ( n17125 , n17124 );
not ( n17126 , n454 );
or ( n17127 , n17125 , n17126 );
not ( n17128 , n15040 );
nand ( n17129 , n15061 , n15064 );
not ( n17130 , n17129 );
or ( n17131 , n17128 , n17130 );
or ( n17132 , n17129 , n15040 );
nand ( n17133 , n17131 , n17132 );
nand ( n17134 , n17133 , n10061 );
nand ( n17135 , n17127 , n17134 );
and ( n17136 , n17135 , n469 );
and ( n17137 , n17098 , n470 );
xor ( n17138 , n17136 , n17137 );
and ( n17139 , n17055 , n471 );
and ( n17140 , n17138 , n17139 );
and ( n17141 , n17136 , n17137 );
or ( n17142 , n17140 , n17141 );
xor ( n17143 , n17121 , n17142 );
xor ( n86809 , n17099 , n17100 );
xor ( n17145 , n86809 , n17102 );
and ( n17146 , n17143 , n17145 );
and ( n17147 , n17121 , n17142 );
or ( n17148 , n17146 , n17147 );
not ( n17149 , n17148 );
nand ( n17150 , n17120 , n17149 );
not ( n17151 , n17150 );
xor ( n17152 , n17121 , n17142 );
xor ( n17153 , n17152 , n17145 );
not ( n17154 , n17153 );
and ( n17155 , n17020 , n472 );
not ( n17156 , n10061 );
not ( n17157 , n15036 );
nand ( n17158 , n14878 , n15039 );
not ( n17159 , n17158 );
or ( n17160 , n17157 , n17159 );
or ( n17161 , n17158 , n15036 );
nand ( n17162 , n17160 , n17161 );
not ( n17163 , n17162 );
or ( n17164 , n17156 , n17163 );
xnor ( n17165 , n8996 , n8976 );
buf ( n17166 , n9148 );
and ( n17167 , n17165 , n17166 );
not ( n17168 , n17165 );
not ( n17169 , n17166 );
and ( n17170 , n17168 , n17169 );
nor ( n17171 , n17167 , n17170 );
nand ( n17172 , n17171 , n454 );
nand ( n17173 , n17164 , n17172 );
and ( n17174 , n17173 , n469 );
and ( n17175 , n17135 , n470 );
xor ( n17176 , n17174 , n17175 );
and ( n17177 , n17098 , n471 );
and ( n17178 , n17176 , n17177 );
and ( n17179 , n17174 , n17175 );
or ( n17180 , n17178 , n17179 );
xor ( n17181 , n17155 , n17180 );
xor ( n17182 , n17136 , n17137 );
xor ( n17183 , n17182 , n17139 );
and ( n17184 , n17181 , n17183 );
and ( n17185 , n17155 , n17180 );
or ( n17186 , n17184 , n17185 );
not ( n86852 , n17186 );
nand ( n17188 , n17154 , n86852 );
not ( n17189 , n17188 );
xor ( n17190 , n17155 , n17180 );
xor ( n17191 , n17190 , n17183 );
not ( n17192 , n17191 );
and ( n17193 , n17055 , n472 );
not ( n17194 , n10061 );
xor ( n17195 , n14903 , n14905 );
xor ( n17196 , n17195 , n15033 );
not ( n17197 , n17196 );
or ( n17198 , n17194 , n17197 );
not ( n17199 , n9018 );
nand ( n17200 , n17199 , n9022 );
and ( n17201 , n17200 , n9146 );
and ( n17202 , n17201 , n9144 );
not ( n17203 , n17201 );
not ( n17204 , n9144 );
and ( n86870 , n17203 , n17204 );
nor ( n17209 , n17202 , n86870 );
nand ( n86872 , n454 , n17209 );
nand ( n17211 , n17198 , n86872 );
and ( n17212 , n17211 , n469 );
and ( n17213 , n17173 , n470 );
xor ( n17214 , n17212 , n17213 );
and ( n17215 , n17135 , n471 );
and ( n17216 , n17214 , n17215 );
and ( n17217 , n17212 , n17213 );
or ( n17218 , n17216 , n17217 );
xor ( n17219 , n17193 , n17218 );
xor ( n17220 , n17174 , n17175 );
xor ( n17221 , n17220 , n17177 );
and ( n17222 , n17219 , n17221 );
and ( n17223 , n17193 , n17218 );
or ( n17224 , n17222 , n17223 );
not ( n17225 , n17224 );
nand ( n17226 , n17192 , n17225 );
not ( n17227 , n17226 );
xor ( n17228 , n17193 , n17218 );
xor ( n86891 , n17228 , n17221 );
not ( n17233 , n86891 );
nand ( n17234 , n9140 , n9143 );
not ( n17235 , n9130 );
and ( n17236 , n17234 , n17235 );
not ( n17237 , n17234 );
and ( n17238 , n17237 , n9130 );
nor ( n17239 , n17236 , n17238 );
not ( n17240 , n17239 );
not ( n17241 , n454 );
or ( n17242 , n17240 , n17241 );
xor ( n17243 , n14945 , n15027 );
xor ( n17244 , n17243 , n15030 );
nand ( n17245 , n17244 , n10061 );
nand ( n17246 , n17242 , n17245 );
and ( n17247 , n17246 , n469 );
and ( n17248 , n17211 , n470 );
xor ( n17249 , n17247 , n17248 );
nand ( n17250 , n17246 , n470 );
not ( n17251 , n454 );
not ( n17252 , n9127 );
nand ( n17253 , n17252 , n9129 );
xor ( n17254 , n9110 , n17253 );
not ( n17255 , n17254 );
or ( n17256 , n17251 , n17255 );
not ( n17257 , n15024 );
or ( n17258 , n14947 , n14957 );
nand ( n17259 , n17258 , n15026 );
not ( n17260 , n17259 );
or ( n17261 , n17257 , n17260 );
or ( n17262 , n17259 , n15024 );
nand ( n17263 , n17261 , n17262 );
nand ( n17264 , n17263 , n10061 );
nand ( n17265 , n17256 , n17264 );
nand ( n17266 , n17265 , n469 );
nor ( n17267 , n17250 , n17266 );
and ( n17268 , n17249 , n17267 );
and ( n17269 , n17247 , n17248 );
or ( n17270 , n17268 , n17269 );
and ( n17271 , n17098 , n472 );
xor ( n17272 , n17270 , n17271 );
and ( n17273 , n17173 , n471 );
not ( n17274 , n17211 );
not ( n17275 , n471 );
nor ( n17276 , n17274 , n17275 );
not ( n17277 , n17266 );
not ( n17278 , n17277 );
not ( n17279 , n17250 );
or ( n17280 , n17278 , n17279 );
nand ( n17281 , n17266 , n470 , n17246 );
nand ( n17282 , n17280 , n17281 );
xor ( n17283 , n17276 , n17282 );
and ( n17284 , n17246 , n471 );
not ( n86944 , n17284 );
nand ( n17286 , n470 , n17265 );
nor ( n17287 , n86944 , n17286 );
and ( n17288 , n17283 , n17287 );
and ( n17289 , n17276 , n17282 );
or ( n17290 , n17288 , n17289 );
xor ( n17291 , n17273 , n17290 );
and ( n17292 , n17135 , n472 );
and ( n17293 , n17291 , n17292 );
and ( n17294 , n17273 , n17290 );
or ( n17295 , n17293 , n17294 );
and ( n17296 , n17272 , n17295 );
and ( n17297 , n17270 , n17271 );
or ( n17298 , n17296 , n17297 );
not ( n17299 , n17298 );
nand ( n17300 , n17233 , n17299 );
not ( n17301 , n17300 );
xor ( n17302 , n17270 , n17271 );
xor ( n17303 , n17302 , n17295 );
xor ( n17304 , n17212 , n17213 );
xor ( n17305 , n17304 , n17215 );
nor ( n17306 , n17303 , n17305 );
and ( n17307 , n17173 , n472 );
xor ( n17308 , n17276 , n17282 );
xor ( n17309 , n17308 , n17287 );
xor ( n17310 , n17307 , n17309 );
not ( n17311 , n17284 );
not ( n17312 , n17286 );
or ( n17313 , n17311 , n17312 );
or ( n17314 , n17286 , n17284 );
nand ( n17315 , n17313 , n17314 );
not ( n86975 , n17315 );
not ( n17320 , n472 );
nor ( n86977 , n17320 , n17274 );
not ( n17322 , n86977 );
nand ( n17323 , n17246 , n17265 , n471 , n472 );
nand ( n17324 , n17322 , n17323 );
not ( n17325 , n17324 );
or ( n17326 , n86975 , n17325 );
not ( n17327 , n17323 );
nand ( n17328 , n17327 , n86977 );
nand ( n17329 , n17326 , n17328 );
and ( n17330 , n17310 , n17329 );
and ( n17331 , n17307 , n17309 );
or ( n17332 , n17330 , n17331 );
xor ( n17333 , n17273 , n17290 );
xor ( n17334 , n17333 , n17292 );
not ( n17335 , n17334 );
xor ( n17336 , n17247 , n17248 );
xor ( n17337 , n17336 , n17267 );
not ( n17338 , n17337 );
nand ( n17339 , n17335 , n17338 );
and ( n17340 , n17332 , n17339 );
nor ( n17341 , n17335 , n17338 );
nor ( n17342 , n17340 , n17341 );
or ( n17343 , n17306 , n17342 );
nand ( n17344 , n17303 , n17305 );
nand ( n17345 , n17343 , n17344 );
not ( n17346 , n17345 );
or ( n87003 , n17301 , n17346 );
nand ( n17351 , n86891 , n17298 );
nand ( n17352 , n87003 , n17351 );
not ( n17353 , n17352 );
or ( n17354 , n17227 , n17353 );
nand ( n17355 , n17191 , n17224 );
nand ( n17356 , n17354 , n17355 );
not ( n17357 , n17356 );
or ( n17358 , n17189 , n17357 );
nand ( n17359 , n17153 , n17186 );
nand ( n17360 , n17358 , n17359 );
not ( n17361 , n17360 );
or ( n17362 , n17151 , n17361 );
nand ( n17363 , n17119 , n17148 );
nand ( n17364 , n17362 , n17363 );
not ( n17365 , n17364 );
or ( n17366 , n17117 , n17365 );
nand ( n17367 , n17114 , n17111 );
nand ( n17368 , n17366 , n17367 );
not ( n17369 , n17368 );
or ( n17370 , n17073 , n17369 );
nand ( n17371 , n17042 , n17071 );
nand ( n17372 , n17370 , n17371 );
not ( n17373 , n17372 );
or ( n17374 , n17040 , n17373 );
not ( n17375 , n17038 );
nand ( n17376 , n17375 , n17034 );
nand ( n17377 , n17374 , n17376 );
not ( n17378 , n17377 );
or ( n17379 , n16998 , n17378 );
nand ( n17380 , n16961 , n16996 );
nand ( n17381 , n17379 , n17380 );
and ( n17382 , n16758 , n472 );
buf ( n17383 , n8154 );
nand ( n17384 , n17383 , n8176 );
not ( n17385 , n17384 );
not ( n17386 , n9261 );
not ( n17387 , n16735 );
or ( n17388 , n17386 , n17387 );
nand ( n17389 , n17388 , n16738 );
not ( n17390 , n17389 );
or ( n17391 , n17385 , n17390 );
or ( n17392 , n17384 , n16739 );
nand ( n17393 , n17391 , n17392 );
nand ( n17394 , n17393 , n454 );
not ( n17395 , n15295 );
nand ( n17396 , n17395 , n15315 );
not ( n17397 , n17396 );
not ( n87051 , n17397 );
not ( n17399 , n15121 );
not ( n17400 , n15253 );
or ( n17401 , n17399 , n17400 );
not ( n17402 , n15245 );
not ( n17403 , n15257 );
and ( n17404 , n17402 , n17403 );
nor ( n17405 , n17404 , n15260 );
nand ( n17406 , n17401 , n17405 );
not ( n17407 , n17406 );
not ( n17408 , n15302 );
buf ( n17409 , n17408 );
not ( n17410 , n17409 );
or ( n17411 , n17407 , n17410 );
buf ( n17412 , n15313 );
nand ( n17413 , n17411 , n17412 );
not ( n17414 , n17413 );
or ( n17415 , n87051 , n17414 );
nand ( n17416 , n17406 , n17409 );
and ( n17417 , n17416 , n17396 , n17412 );
nor ( n17418 , n17417 , n454 );
nand ( n17419 , n17415 , n17418 );
and ( n17420 , n17394 , n17419 );
not ( n17421 , n470 );
nor ( n17422 , n17420 , n17421 );
nand ( n17423 , n17408 , n15313 );
not ( n17424 , n17423 );
not ( n17425 , n17406 );
or ( n17426 , n17424 , n17425 );
or ( n17427 , n17406 , n17423 );
nand ( n17428 , n17426 , n17427 );
nand ( n17429 , n17428 , n10061 );
not ( n17430 , n17429 );
nand ( n17431 , n8181 , n8125 );
not ( n17432 , n17431 );
not ( n87086 , n16868 );
not ( n17437 , n9261 );
or ( n87088 , n87086 , n17437 );
nand ( n17439 , n87088 , n16869 );
not ( n17440 , n17439 );
or ( n17441 , n17432 , n17440 );
or ( n17442 , n17431 , n17439 );
nand ( n17443 , n17441 , n17442 );
nand ( n17444 , n17443 , n454 );
not ( n17445 , n17444 );
or ( n17446 , n17430 , n17445 );
nand ( n17447 , n17446 , n469 );
not ( n17448 , n17447 );
xor ( n17449 , n17422 , n17448 );
buf ( n17450 , n8159 );
not ( n17451 , n8173 );
nor ( n17452 , n17450 , n17451 );
not ( n17453 , n17383 );
nor ( n17454 , n17452 , n17453 );
buf ( n17455 , n8176 );
nand ( n17456 , n17389 , n17455 );
and ( n87107 , n17454 , n17456 );
nor ( n17461 , n87107 , n16728 );
not ( n17462 , n17461 );
not ( n17463 , n17383 );
not ( n17464 , n17456 );
or ( n17465 , n17463 , n17464 );
buf ( n17466 , n17452 );
nand ( n17467 , n17465 , n17466 );
not ( n17468 , n17467 );
or ( n17469 , n17462 , n17468 );
nand ( n17470 , n15311 , n15322 );
not ( n17471 , n17470 );
not ( n17472 , n15978 );
or ( n17473 , n17471 , n17472 );
or ( n17474 , n15978 , n17470 );
nand ( n17475 , n17473 , n17474 );
nand ( n17476 , n17475 , n10061 );
nand ( n17477 , n17469 , n17476 );
and ( n17478 , n17477 , n471 );
and ( n17479 , n17449 , n17478 );
and ( n17480 , n17422 , n17448 );
or ( n17481 , n17479 , n17480 );
xor ( n17482 , n17382 , n17481 );
nand ( n17483 , n17394 , n17419 );
and ( n17484 , n17483 , n469 );
and ( n17485 , n17477 , n470 );
xor ( n17486 , n17484 , n17485 );
not ( n17487 , n454 );
nand ( n17488 , n16730 , n8166 );
not ( n17489 , n17488 );
and ( n17490 , n16743 , n17489 );
not ( n17491 , n16743 );
and ( n17492 , n17491 , n17488 );
nor ( n17493 , n17490 , n17492 );
not ( n17494 , n17493 );
or ( n17495 , n17487 , n17494 );
not ( n17496 , n15311 );
not ( n17497 , n15978 );
or ( n17498 , n17496 , n17497 );
nand ( n17499 , n17498 , n15322 );
not ( n17500 , n13728 );
nor ( n17501 , n17500 , n15325 );
xor ( n87149 , n17499 , n17501 );
nand ( n17503 , n87149 , n10061 );
nand ( n17504 , n17495 , n17503 );
and ( n17505 , n17504 , n471 );
xor ( n17506 , n17486 , n17505 );
xor ( n17507 , n17482 , n17506 );
not ( n17508 , n17507 );
and ( n17509 , n17504 , n472 );
and ( n17510 , n16880 , n469 );
not ( n17511 , n17483 );
nor ( n17512 , n17511 , n17275 );
xor ( n17513 , n17510 , n17512 );
nand ( n17514 , n17444 , n17429 );
and ( n17515 , n17514 , n470 );
and ( n17516 , n17513 , n17515 );
and ( n17517 , n17510 , n17512 );
or ( n17518 , n17516 , n17517 );
xor ( n17519 , n17509 , n17518 );
xor ( n17520 , n17422 , n17448 );
xor ( n17521 , n17520 , n17478 );
and ( n17522 , n17519 , n17521 );
and ( n17523 , n17509 , n17518 );
or ( n17524 , n17522 , n17523 );
not ( n17525 , n17524 );
nand ( n17526 , n17508 , n17525 );
and ( n17527 , n17514 , n471 );
and ( n17528 , n16835 , n469 );
and ( n17529 , n16880 , n471 );
xor ( n17530 , n17528 , n17529 );
not ( n17531 , n16786 );
nor ( n17532 , n17531 , n17421 );
and ( n17533 , n17530 , n17532 );
and ( n87181 , n17528 , n17529 );
or ( n17538 , n17533 , n87181 );
xor ( n87183 , n17527 , n17538 );
and ( n17540 , n16880 , n470 );
and ( n17541 , n16786 , n469 );
xor ( n17542 , n17540 , n17541 );
and ( n17543 , n17483 , n472 );
xor ( n17544 , n17542 , n17543 );
xor ( n17545 , n87183 , n17544 );
not ( n17546 , n17545 );
and ( n17547 , n17514 , n472 );
xor ( n17548 , n16852 , n16853 );
and ( n17549 , n17548 , n16881 );
and ( n17550 , n16852 , n16853 );
or ( n17551 , n17549 , n17550 );
xor ( n17552 , n17547 , n17551 );
xor ( n17553 , n17528 , n17529 );
xor ( n17554 , n17553 , n17532 );
and ( n17555 , n17552 , n17554 );
and ( n87200 , n17547 , n17551 );
or ( n17560 , n17555 , n87200 );
not ( n17561 , n17560 );
and ( n17562 , n17546 , n17561 );
xor ( n17563 , n17547 , n17551 );
xor ( n17564 , n17563 , n17554 );
xor ( n17565 , n16787 , n16850 );
and ( n17566 , n17565 , n16882 );
and ( n17567 , n16787 , n16850 );
or ( n17568 , n17566 , n17567 );
nor ( n17569 , n17564 , n17568 );
nor ( n17570 , n17562 , n17569 );
nand ( n17571 , n16959 , n17381 , n17526 , n17570 );
not ( n17572 , n17571 );
and ( n17573 , n16758 , n471 );
xor ( n17574 , n17484 , n17485 );
and ( n17575 , n17574 , n17505 );
and ( n17576 , n17484 , n17485 );
or ( n17577 , n17575 , n17576 );
xor ( n17578 , n17573 , n17577 );
not ( n17579 , n17461 );
not ( n17580 , n17467 );
or ( n17581 , n17579 , n17580 );
nand ( n17582 , n17581 , n17476 );
and ( n17583 , n17582 , n469 );
and ( n17584 , n17504 , n470 );
xor ( n17585 , n17583 , n17584 );
and ( n17586 , n15995 , n472 );
xor ( n17587 , n17585 , n17586 );
xor ( n17588 , n17578 , n17587 );
not ( n17589 , n17588 );
xor ( n17590 , n17382 , n17481 );
and ( n17591 , n17590 , n17506 );
and ( n17592 , n17382 , n17481 );
or ( n17593 , n17591 , n17592 );
not ( n17594 , n17593 );
and ( n17595 , n17589 , n17594 );
and ( n17596 , n17582 , n472 );
xor ( n87238 , n17540 , n17541 );
and ( n17598 , n87238 , n17543 );
and ( n17599 , n17540 , n17541 );
or ( n17600 , n17598 , n17599 );
xor ( n17601 , n17596 , n17600 );
xor ( n17602 , n17510 , n17512 );
xor ( n17603 , n17602 , n17515 );
and ( n17604 , n17601 , n17603 );
and ( n17605 , n17596 , n17600 );
or ( n17606 , n17604 , n17605 );
not ( n17607 , n17606 );
not ( n17608 , n17607 );
xor ( n17609 , n17509 , n17518 );
xor ( n17610 , n17609 , n17521 );
not ( n17611 , n17610 );
not ( n17612 , n17611 );
or ( n17613 , n17608 , n17612 );
xor ( n17614 , n17596 , n17600 );
xor ( n17615 , n17614 , n17603 );
not ( n17616 , n17615 );
xor ( n17617 , n17527 , n17538 );
and ( n17618 , n17617 , n17544 );
and ( n17619 , n17527 , n17538 );
or ( n17620 , n17618 , n17619 );
not ( n17621 , n17620 );
nand ( n17622 , n17616 , n17621 );
nand ( n87264 , n17613 , n17622 );
nor ( n17627 , n17595 , n87264 );
nand ( n17628 , n17572 , n17627 );
nand ( n17629 , n17589 , n17594 );
and ( n17630 , n17507 , n17524 );
nand ( n17631 , n17629 , n17630 );
buf ( n17632 , n17588 );
nand ( n17633 , n17632 , n17593 );
buf ( n17634 , n17526 );
not ( n17635 , n17607 );
not ( n17636 , n17611 );
or ( n17637 , n17635 , n17636 );
nand ( n17638 , n17637 , n17622 );
not ( n17639 , n17638 );
not ( n17640 , n17639 );
nand ( n17641 , n16914 , n16955 );
or ( n17642 , n16912 , n17641 );
nand ( n17643 , n16883 , n16911 );
nand ( n17644 , n17642 , n17643 );
not ( n17645 , n17644 );
not ( n17646 , n17570 );
or ( n17647 , n17645 , n17646 );
not ( n17648 , n17545 );
not ( n17649 , n17560 );
nand ( n17650 , n17648 , n17649 );
and ( n17651 , n17564 , n17568 );
and ( n17652 , n17650 , n17651 );
not ( n17653 , n17545 );
nor ( n17654 , n17653 , n17649 );
nor ( n17655 , n17652 , n17654 );
nand ( n17656 , n17647 , n17655 );
not ( n17657 , n17656 );
or ( n87296 , n17640 , n17657 );
nand ( n17659 , n17611 , n17607 );
and ( n17660 , n17615 , n17620 );
and ( n17661 , n17659 , n17660 );
and ( n17662 , n17610 , n17606 );
nor ( n17663 , n17661 , n17662 );
nand ( n17664 , n87296 , n17663 );
nand ( n17665 , n17634 , n17664 , n17629 );
nand ( n17666 , n17628 , n17631 , n17633 , n17665 );
xor ( n17667 , n16725 , n16764 );
xor ( n17668 , n17667 , n16767 );
not ( n17669 , n17668 );
and ( n17670 , n16048 , n471 );
and ( n17671 , n17504 , n469 );
not ( n17672 , n15995 );
nor ( n17673 , n17672 , n17275 );
xor ( n17674 , n17671 , n17673 );
and ( n17675 , n16758 , n470 );
and ( n17676 , n17674 , n17675 );
and ( n17677 , n17671 , n17673 );
or ( n87316 , n17676 , n17677 );
xor ( n17682 , n17670 , n87316 );
xor ( n17683 , n16726 , n16759 );
xor ( n17684 , n17683 , n16761 );
and ( n17685 , n17682 , n17684 );
and ( n17686 , n17670 , n87316 );
or ( n17687 , n17685 , n17686 );
not ( n17688 , n17687 );
nand ( n17689 , n17669 , n17688 );
not ( n17690 , n17689 );
xor ( n17691 , n17670 , n87316 );
xor ( n17692 , n17691 , n17684 );
and ( n17693 , n16048 , n472 );
xor ( n17694 , n17583 , n17584 );
and ( n17695 , n17694 , n17586 );
and ( n17696 , n17583 , n17584 );
or ( n17697 , n17695 , n17696 );
xor ( n17698 , n17693 , n17697 );
xor ( n17699 , n17671 , n17673 );
xor ( n17700 , n17699 , n17675 );
and ( n17701 , n17698 , n17700 );
and ( n17702 , n17693 , n17697 );
or ( n17703 , n17701 , n17702 );
nor ( n17704 , n17692 , n17703 );
xor ( n17705 , n17693 , n17697 );
xor ( n17706 , n17705 , n17700 );
xor ( n87342 , n17573 , n17577 );
and ( n17708 , n87342 , n17587 );
and ( n17709 , n17573 , n17577 );
or ( n17710 , n17708 , n17709 );
nor ( n17711 , n17706 , n17710 );
nor ( n17712 , n17704 , n17711 );
not ( n17713 , n17712 );
nor ( n17714 , n17690 , n17713 );
nand ( n17715 , n16772 , n17666 , n17714 );
nand ( n17716 , n17706 , n17710 );
or ( n17717 , n17704 , n17716 );
nand ( n17718 , n17692 , n17703 );
nand ( n17719 , n17717 , n17718 );
and ( n17720 , n17689 , n17719 );
not ( n17721 , n17668 );
nor ( n17722 , n17721 , n17688 );
nor ( n87358 , n17720 , n17722 );
not ( n17727 , n87358 );
nand ( n17728 , n17727 , n16772 );
nand ( n17729 , n16724 , n16770 );
not ( n17730 , n17729 );
not ( n17731 , n16717 );
not ( n17732 , n16388 );
nand ( n17733 , n17731 , n17732 );
and ( n17734 , n17730 , n17733 );
and ( n17735 , n16717 , n16388 );
nor ( n17736 , n17734 , n17735 );
nand ( n17737 , n17715 , n17728 , n17736 );
and ( n17738 , n16704 , n471 );
xor ( n17739 , n16711 , n16713 );
and ( n17740 , n17739 , n16715 );
and ( n17741 , n16711 , n16713 );
or ( n17742 , n17740 , n17741 );
xor ( n17743 , n17738 , n17742 );
not ( n17744 , n454 );
not ( n17745 , n15777 );
not ( n17746 , n15771 );
or ( n17747 , n17745 , n17746 );
or ( n17748 , n16363 , n16367 );
nand ( n87381 , n16695 , n15953 , n17748 );
not ( n17750 , n87381 );
nand ( n17751 , n17747 , n17750 );
nand ( n17752 , n16368 , n16696 );
or ( n17753 , n17752 , n16521 );
nand ( n17754 , n17753 , n16695 );
buf ( n17755 , n17754 );
nand ( n17756 , n17751 , n17755 );
not ( n17757 , n12969 );
not ( n87390 , n16532 );
or ( n17762 , n17757 , n87390 );
and ( n17763 , n495 , n15563 );
not ( n17764 , n495 );
and ( n17765 , n17764 , n15566 );
or ( n17766 , n17763 , n17765 );
nand ( n17767 , n17766 , n13032 );
nand ( n17768 , n17762 , n17767 );
not ( n17769 , n15344 );
not ( n17770 , n16545 );
or ( n17771 , n17769 , n17770 );
not ( n17772 , n493 );
not ( n17773 , n12852 );
or ( n17774 , n17772 , n17773 );
nand ( n17775 , n13369 , n12775 );
nand ( n17776 , n17774 , n17775 );
nand ( n87406 , n17776 , n12758 );
nand ( n17781 , n17771 , n87406 );
xor ( n87408 , n17768 , n17781 );
not ( n87409 , n12702 );
not ( n87410 , n16590 );
or ( n87411 , n87409 , n87410 );
not ( n87412 , n499 );
not ( n87413 , n15697 );
or ( n87414 , n87412 , n87413 );
nand ( n87415 , n15690 , n12467 );
nand ( n87416 , n87414 , n87415 );
nand ( n87417 , n87416 , n12650 );
nand ( n87418 , n87411 , n87417 );
xor ( n87419 , n87408 , n87418 );
xor ( n87420 , n16539 , n16549 );
and ( n87421 , n87420 , n16566 );
and ( n87422 , n16539 , n16549 );
or ( n87423 , n87421 , n87422 );
xor ( n87424 , n87419 , n87423 );
xor ( n87425 , n16651 , n16655 );
and ( n87426 , n87425 , n16677 );
and ( n87427 , n16651 , n16655 );
or ( n87428 , n87426 , n87427 );
xor ( n87429 , n87424 , n87428 );
not ( n87430 , n12517 );
not ( n87431 , n497 );
not ( n87432 , n15438 );
or ( n87433 , n87431 , n87432 );
nand ( n87434 , n12418 , n12486 );
nand ( n87435 , n87433 , n87434 );
not ( n87436 , n87435 );
or ( n87437 , n87430 , n87436 );
not ( n87438 , n13258 );
not ( n87439 , n16577 );
and ( n87440 , n87438 , n87439 );
not ( n87441 , n13255 );
and ( n87442 , n87441 , n16574 );
nor ( n87443 , n87440 , n87442 );
nand ( n87444 , n87437 , n87443 );
not ( n87445 , n12822 );
not ( n87446 , n16564 );
or ( n87447 , n87445 , n87446 );
and ( n87448 , n16321 , n16260 );
not ( n87449 , n16321 );
and ( n87450 , n12843 , n501 );
and ( n87451 , n87449 , n87450 );
nor ( n87452 , n87448 , n87451 );
nand ( n87453 , n87447 , n87452 );
xor ( n87454 , n87444 , n87453 );
xor ( n87455 , n16657 , n16663 );
and ( n87456 , n87455 , n16676 );
and ( n87457 , n16657 , n16663 );
or ( n87458 , n87456 , n87457 );
xor ( n87459 , n87454 , n87458 );
not ( n87460 , n12462 );
not ( n87461 , n16647 );
or ( n87462 , n87460 , n87461 );
nand ( n87463 , n87462 , n70376 );
not ( n87464 , n12595 );
not ( n87465 , n16658 );
or ( n87466 , n87464 , n87465 );
not ( n87467 , n491 );
not ( n87468 , n13357 );
or ( n87469 , n87467 , n87468 );
or ( n87470 , n491 , n13357 );
nand ( n87471 , n87469 , n87470 );
nand ( n87472 , n87471 , n12638 );
nand ( n87473 , n87466 , n87472 );
and ( n87474 , n16665 , n16675 );
xor ( n87475 , n87473 , n87474 );
nand ( n87476 , n489 , n13008 );
not ( n87477 , n87476 );
not ( n87478 , n12580 );
not ( n87479 , n489 );
not ( n87480 , n12482 );
or ( n87481 , n87479 , n87480 );
nand ( n87482 , n12481 , n12560 );
nand ( n87483 , n87481 , n87482 );
not ( n87484 , n87483 );
or ( n87485 , n87478 , n87484 );
nand ( n87486 , n16670 , n12542 );
nand ( n87487 , n87485 , n87486 );
not ( n87488 , n87487 );
or ( n87489 , n87477 , n87488 );
or ( n87490 , n87487 , n87476 );
nand ( n87491 , n87489 , n87490 );
xor ( n87492 , n87475 , n87491 );
xor ( n87493 , n87463 , n87492 );
xor ( n87494 , n16579 , n16583 );
and ( n87495 , n87494 , n16594 );
and ( n87496 , n16579 , n16583 );
or ( n87497 , n87495 , n87496 );
xor ( n87498 , n87493 , n87497 );
xor ( n87499 , n87459 , n87498 );
xor ( n87500 , n16567 , n16571 );
and ( n87501 , n87500 , n16595 );
and ( n87502 , n16567 , n16571 );
or ( n87503 , n87501 , n87502 );
xor ( n87504 , n87499 , n87503 );
xor ( n87505 , n87429 , n87504 );
xor ( n87506 , n16600 , n16678 );
and ( n87507 , n87506 , n16683 );
and ( n87508 , n16600 , n16678 );
or ( n87509 , n87507 , n87508 );
xor ( n87510 , n87505 , n87509 );
not ( n87511 , n87510 );
xor ( n87512 , n16596 , n86367 );
and ( n87513 , n87512 , n16689 );
and ( n87514 , n16596 , n86367 );
or ( n87515 , n87513 , n87514 );
not ( n87516 , n87515 );
nor ( n87517 , n87511 , n87516 );
not ( n87518 , n87517 );
not ( n87519 , n87510 );
nand ( n87520 , n87519 , n87516 );
buf ( n87521 , n87520 );
nand ( n87522 , n87518 , n87521 );
not ( n87523 , n87522 );
and ( n87524 , n17756 , n87523 );
not ( n87525 , n17756 );
and ( n87526 , n87525 , n87522 );
nor ( n87527 , n87524 , n87526 );
nand ( n87528 , n17744 , n87527 );
not ( n87529 , n16728 );
not ( n87530 , n16391 );
nor ( n87531 , n87530 , n16503 );
not ( n87532 , n87531 );
not ( n87533 , n9923 );
or ( n87534 , n87532 , n87533 );
buf ( n87535 , n16390 );
nor ( n87536 , n16503 , n87535 );
buf ( n87537 , n16395 );
and ( n87538 , n87536 , n87537 );
not ( n87539 , n16506 );
nor ( n87540 , n87538 , n87539 );
nand ( n87541 , n87534 , n87540 );
xor ( n87542 , n16416 , n16425 );
and ( n87543 , n87542 , n16430 );
and ( n87544 , n16416 , n16425 );
or ( n87545 , n87543 , n87544 );
not ( n87546 , n5590 );
not ( n87547 , n541 );
not ( n87548 , n7324 );
or ( n87549 , n87547 , n87548 );
nand ( n87550 , n6440 , n5538 );
nand ( n87551 , n87549 , n87550 );
not ( n87552 , n87551 );
or ( n87553 , n87546 , n87552 );
nand ( n87554 , n16414 , n9938 );
nand ( n87555 , n87553 , n87554 );
not ( n87556 , n4434 );
and ( n87557 , n6844 , n539 );
not ( n87558 , n6844 );
and ( n87559 , n87558 , n4251 );
or ( n87560 , n87557 , n87559 );
not ( n87561 , n87560 );
or ( n87562 , n87556 , n87561 );
and ( n87563 , n5392 , n4251 );
not ( n87564 , n5392 );
and ( n87565 , n87564 , n539 );
or ( n87566 , n87563 , n87565 );
nand ( n87567 , n87566 , n4224 );
nand ( n87568 , n87562 , n87567 );
xor ( n87569 , n87555 , n87568 );
not ( n87570 , n5399 );
not ( n87571 , n545 );
not ( n87572 , n9557 );
or ( n87573 , n87571 , n87572 );
nand ( n87574 , n16141 , n4440 );
nand ( n87575 , n87573 , n87574 );
not ( n87576 , n87575 );
or ( n87577 , n87570 , n87576 );
nand ( n87578 , n16421 , n75018 );
nand ( n87579 , n87577 , n87578 );
xor ( n87580 , n87569 , n87579 );
xor ( n87581 , n87545 , n87580 );
not ( n87582 , n5501 );
not ( n87583 , n537 );
not ( n87584 , n7378 );
or ( n87585 , n87583 , n87584 );
nand ( n87586 , n5264 , n5409 );
nand ( n87587 , n87585 , n87586 );
not ( n87588 , n87587 );
or ( n87589 , n87582 , n87588 );
nand ( n87590 , n16470 , n16155 );
nand ( n87591 , n87589 , n87590 );
not ( n87592 , n9595 );
not ( n87593 , n543 );
not ( n87594 , n9735 );
or ( n87595 , n87593 , n87594 );
nand ( n87596 , n9734 , n4938 );
nand ( n87597 , n87595 , n87596 );
not ( n87598 , n87597 );
or ( n87599 , n87592 , n87598 );
nand ( n87600 , n16449 , n4445 );
nand ( n87601 , n87599 , n87600 );
xor ( n87602 , n87591 , n87601 );
not ( n87603 , n6811 );
not ( n87604 , n547 );
not ( n87605 , n9848 );
or ( n87606 , n87604 , n87605 );
or ( n87607 , n9848 , n547 );
nand ( n87608 , n87606 , n87607 );
not ( n87609 , n87608 );
or ( n87610 , n87603 , n87609 );
nand ( n87611 , n16458 , n6854 );
nand ( n87612 , n87610 , n87611 );
xor ( n87613 , n87602 , n87612 );
xor ( n87614 , n87581 , n87613 );
or ( n87615 , n6489 , n5905 );
nand ( n87616 , n87615 , n549 );
and ( n87617 , n4937 , n537 );
xor ( n87618 , n87616 , n87617 );
not ( n87619 , n16473 );
xor ( n87620 , n87618 , n87619 );
xor ( n87621 , n16472 , n16473 );
and ( n87622 , n87621 , n16163 );
and ( n87623 , n16472 , n16473 );
or ( n87624 , n87622 , n87623 );
xor ( n87625 , n87620 , n87624 );
xor ( n87626 , n16443 , n16453 );
and ( n87627 , n87626 , n16460 );
and ( n87628 , n16443 , n16453 );
or ( n87629 , n87627 , n87628 );
xor ( n87630 , n87625 , n87629 );
xor ( n87631 , n16475 , n16479 );
and ( n87632 , n87631 , n16484 );
and ( n87633 , n16475 , n16479 );
or ( n87634 , n87632 , n87633 );
xor ( n87635 , n87630 , n87634 );
xor ( n87636 , n16406 , n16431 );
and ( n87637 , n87636 , n16461 );
and ( n87638 , n16406 , n16431 );
or ( n87639 , n87637 , n87638 );
xor ( n87640 , n87635 , n87639 );
xor ( n87641 , n87614 , n87640 );
xor ( n87642 , n86174 , n16489 );
and ( n87643 , n87642 , n16494 );
and ( n87644 , n86174 , n16489 );
or ( n87645 , n87643 , n87644 );
xor ( n87646 , n87641 , n87645 );
xor ( n87647 , n16462 , n16495 );
and ( n87648 , n87647 , n16500 );
and ( n87649 , n16462 , n16495 );
or ( n87650 , n87648 , n87649 );
nor ( n87651 , n87646 , n87650 );
not ( n87652 , n87651 );
buf ( n87653 , n87646 );
nand ( n87654 , n87653 , n87650 );
nand ( n87655 , n87652 , n87654 );
not ( n87656 , n87655 );
and ( n87657 , n87541 , n87656 );
not ( n87658 , n87541 );
and ( n87659 , n87658 , n87655 );
nor ( n87660 , n87657 , n87659 );
nand ( n87661 , n87529 , n87660 );
and ( n87662 , n87528 , n87661 );
nor ( n87663 , n87662 , n16383 );
and ( n87664 , n15958 , n469 );
xor ( n87665 , n87663 , n87664 );
nor ( n87666 , n16382 , n17421 );
xor ( n87667 , n87665 , n87666 );
xor ( n87668 , n17743 , n87667 );
xor ( n87669 , n16705 , n16709 );
and ( n87670 , n87669 , n16716 );
and ( n87671 , n16705 , n16709 );
or ( n87672 , n87670 , n87671 );
nor ( n87673 , n87668 , n87672 );
buf ( n87674 , n87673 );
not ( n87675 , n87674 );
nand ( n87676 , n87668 , n87672 );
nand ( n87677 , n87675 , n87676 );
not ( n87678 , n87677 );
and ( n87679 , n17737 , n87678 );
not ( n87680 , n17737 );
and ( n87681 , n87680 , n87677 );
or ( n87682 , n87679 , n87681 );
nor ( n87683 , n455 , n456 );
or ( n87684 , n87683 , n16871 );
or ( n87685 , n87682 , n87684 );
and ( n87686 , n536 , n6801 );
not ( n87687 , n536 );
and ( n87688 , n87687 , n552 );
or ( n87689 , n87686 , n87688 );
not ( n87690 , n87689 );
nand ( n87691 , n536 , n552 );
nand ( n87692 , n535 , n551 );
not ( n87693 , n87692 );
nor ( n87694 , n535 , n551 );
nor ( n87695 , n87693 , n87694 );
and ( n87696 , n87691 , n87695 );
not ( n87697 , n87691 );
not ( n87698 , n87695 );
and ( n87699 , n87697 , n87698 );
or ( n87700 , n87696 , n87699 );
nand ( n87701 , n87690 , n87700 );
not ( n87702 , n87701 );
not ( n87703 , n87702 );
not ( n87704 , n87700 );
buf ( n87705 , n87704 );
not ( n87706 , n87705 );
buf ( n87707 , n2088 );
xor ( n87708 , n1982 , n87707 );
not ( n87709 , n6022 );
not ( n87710 , n75980 );
or ( n87711 , n87709 , n87710 );
nand ( n87712 , n6120 , n1982 );
nand ( n87713 , n87711 , n87712 );
nor ( n87714 , n87708 , n87713 );
not ( n87715 , n87714 );
not ( n87716 , n87715 );
not ( n87717 , n87716 );
not ( n87718 , n75980 );
not ( n87719 , n87718 );
nor ( n87720 , n493 , n509 );
nor ( n87721 , n494 , n510 );
nor ( n87722 , n87720 , n87721 );
nor ( n87723 , n495 , n511 );
nor ( n87724 , n496 , n512 );
nor ( n87725 , n87723 , n87724 );
and ( n87726 , n87722 , n87725 );
not ( n87727 , n87726 );
nor ( n87728 , n498 , n514 );
not ( n87729 , n87728 );
not ( n87730 , n87729 );
or ( n87731 , n497 , n513 );
not ( n87732 , n87731 );
or ( n87733 , n87730 , n87732 );
nand ( n87734 , n497 , n513 );
nand ( n87735 , n87733 , n87734 );
not ( n87736 , n87735 );
nand ( n87737 , n500 , n516 );
nor ( n87738 , n499 , n515 );
or ( n87739 , n87737 , n87738 );
nand ( n87740 , n498 , n514 );
nand ( n87741 , n499 , n515 );
and ( n87742 , n87734 , n87740 , n87741 );
nand ( n87743 , n87739 , n87742 );
not ( n87744 , n87743 );
or ( n87745 , n87736 , n87744 );
nand ( n87746 , n501 , n517 );
nand ( n87747 , n502 , n518 );
and ( n87748 , n87746 , n87747 );
not ( n87749 , n87748 );
not ( n87750 , n504 );
not ( n87751 , n520 );
or ( n87752 , n87750 , n87751 );
nand ( n87753 , n503 , n519 );
nand ( n87754 , n87752 , n87753 );
nor ( n87755 , n503 , n519 );
not ( n87756 , n87755 );
not ( n87757 , n502 );
nand ( n87758 , n87757 , n70435 );
nand ( n87759 , n87754 , n87756 , n87758 );
not ( n87760 , n87759 );
or ( n87761 , n87749 , n87760 );
or ( n87762 , n501 , n517 );
nand ( n87763 , n87731 , n87762 , n87729 );
or ( n87764 , n500 , n516 );
or ( n87765 , n499 , n515 );
nand ( n87766 , n87764 , n87765 );
nor ( n87767 , n87763 , n87766 );
nand ( n87768 , n87761 , n87767 );
nand ( n87769 , n87745 , n87768 );
not ( n87770 , n87769 );
or ( n87771 , n87727 , n87770 );
nor ( n87772 , n495 , n511 );
nand ( n87773 , n496 , n512 );
or ( n87774 , n87772 , n87773 );
nand ( n87775 , n495 , n511 );
nand ( n87776 , n87774 , n87775 );
not ( n87777 , n87776 );
not ( n87778 , n87722 );
or ( n87779 , n87777 , n87778 );
not ( n87780 , n87720 );
nand ( n87781 , n494 , n510 );
not ( n87782 , n87781 );
and ( n87783 , n87780 , n87782 );
nand ( n87784 , n493 , n509 );
not ( n87785 , n87784 );
nor ( n87786 , n87783 , n87785 );
nand ( n87787 , n87779 , n87786 );
not ( n87788 , n87787 );
nand ( n87789 , n87771 , n87788 );
nor ( n87790 , n492 , n508 );
not ( n87791 , n87790 );
nand ( n87792 , n492 , n508 );
nand ( n87793 , n87791 , n87792 );
xnor ( n87794 , n87789 , n87793 );
buf ( n87795 , n87794 );
not ( n87796 , n87795 );
not ( n87797 , n87796 );
or ( n87798 , n87719 , n87797 );
not ( n87799 , n87718 );
nand ( n87800 , n87795 , n87799 );
nand ( n87801 , n87798 , n87800 );
not ( n87802 , n87801 );
or ( n87803 , n87717 , n87802 );
not ( n87804 , n87718 );
not ( n87805 , n87726 );
nor ( n87806 , n87805 , n87790 );
not ( n87807 , n87806 );
not ( n87808 , n87769 );
or ( n87809 , n87807 , n87808 );
and ( n87810 , n87787 , n87791 );
not ( n87811 , n87792 );
nor ( n87812 , n87810 , n87811 );
nand ( n87813 , n87809 , n87812 );
nor ( n87814 , n491 , n507 );
not ( n87815 , n87814 );
nand ( n87816 , n491 , n507 );
and ( n87817 , n87815 , n87816 );
xor ( n87818 , n87813 , n87817 );
not ( n87819 , n87818 );
not ( n87820 , n87819 );
or ( n87821 , n87804 , n87820 );
buf ( n87822 , n87818 );
nand ( n87823 , n87822 , n87799 );
nand ( n87824 , n87821 , n87823 );
not ( n87825 , n87824 );
buf ( n87826 , n87708 );
not ( n87827 , n87826 );
or ( n87828 , n87825 , n87827 );
nand ( n87829 , n87803 , n87828 );
buf ( n87830 , n1726 );
not ( n87831 , n87830 );
and ( n87832 , n87815 , n87791 );
nor ( n87833 , n490 , n506 );
nor ( n87834 , n489 , n505 );
nor ( n87835 , n87833 , n87834 );
nand ( n87836 , n87832 , n87835 );
nor ( n87837 , n87805 , n87836 );
not ( n87838 , n87837 );
not ( n87839 , n87769 );
or ( n87840 , n87838 , n87839 );
not ( n87841 , n87836 );
and ( n87842 , n87787 , n87841 );
not ( n87843 , n87835 );
or ( n87844 , n87814 , n87792 );
nand ( n87845 , n87844 , n87816 );
not ( n87846 , n87845 );
or ( n87847 , n87843 , n87846 );
nand ( n87848 , n490 , n506 );
not ( n87849 , n87848 );
not ( n87850 , n87834 );
and ( n87851 , n87849 , n87850 );
and ( n87852 , n489 , n505 );
nor ( n87853 , n87851 , n87852 );
nand ( n87854 , n87847 , n87853 );
nor ( n87855 , n87842 , n87854 );
nand ( n87856 , n87840 , n87855 );
not ( n87857 , n87856 );
xor ( n87858 , n87831 , n87857 );
not ( n87859 , n87858 );
buf ( n87860 , n1714 );
xnor ( n87861 , n87860 , n87830 );
not ( n87862 , n87860 );
buf ( n87863 , n2065 );
not ( n87864 , n87863 );
not ( n87865 , n87864 );
or ( n87866 , n87862 , n87865 );
not ( n87867 , n87860 );
nand ( n87868 , n87867 , n87863 );
nand ( n87869 , n87866 , n87868 );
nor ( n87870 , n87861 , n87869 );
buf ( n87871 , n87870 );
not ( n87872 , n87871 );
or ( n87873 , n87859 , n87872 );
not ( n87874 , n87869 );
not ( n87875 , n87830 );
or ( n87876 , n87874 , n87875 );
nand ( n87877 , n87873 , n87876 );
not ( n87878 , n87877 );
xor ( n87879 , n87829 , n87878 );
not ( n87880 , n87826 );
not ( n87881 , n87801 );
or ( n87882 , n87880 , n87881 );
not ( n87883 , n87718 );
not ( n87884 , n87721 );
and ( n87885 , n87725 , n87884 );
not ( n87886 , n87885 );
nand ( n87887 , n87743 , n87735 );
nand ( n87888 , n87768 , n87887 );
not ( n87889 , n87888 );
or ( n87890 , n87886 , n87889 );
and ( n87891 , n87776 , n87884 );
not ( n87892 , n87781 );
nor ( n87893 , n87891 , n87892 );
nand ( n87894 , n87890 , n87893 );
not ( n87895 , n87784 );
nor ( n87896 , n87895 , n87720 );
xor ( n87897 , n87894 , n87896 );
not ( n87898 , n87897 );
not ( n87899 , n87898 );
or ( n87900 , n87883 , n87899 );
not ( n87901 , n87898 );
nand ( n87902 , n87901 , n87799 );
nand ( n87903 , n87900 , n87902 );
nand ( n87904 , n87903 , n87716 );
nand ( n87905 , n87882 , n87904 );
not ( n87906 , n6039 );
not ( n87907 , n87906 );
not ( n87908 , n75980 );
or ( n87909 , n87907 , n87908 );
buf ( n87910 , n1881 );
not ( n87911 , n87910 );
and ( n87912 , n87911 , n6120 );
not ( n87913 , n2013 );
and ( n87914 , n87906 , n87913 );
and ( n87915 , n87911 , n2013 );
nor ( n87916 , n87914 , n87915 );
nor ( n87917 , n87912 , n87916 );
nand ( n87918 , n87909 , n87917 );
not ( n87919 , n87918 );
not ( n87920 , n87919 );
not ( n87921 , n2013 );
not ( n87922 , n87921 );
not ( n87923 , n87724 );
not ( n87924 , n87923 );
not ( n87925 , n87769 );
or ( n87926 , n87924 , n87925 );
nand ( n87927 , n87926 , n87773 );
not ( n87928 , n87723 );
nand ( n87929 , n87928 , n87775 );
not ( n87930 , n87929 );
and ( n87931 , n87927 , n87930 );
not ( n87932 , n87927 );
and ( n87933 , n87932 , n87929 );
nor ( n87934 , n87931 , n87933 );
not ( n87935 , n87934 );
not ( n87936 , n87935 );
xor ( n87937 , n87922 , n87936 );
not ( n87938 , n87937 );
or ( n87939 , n87920 , n87938 );
not ( n87940 , n87725 );
not ( n87941 , n87888 );
or ( n87942 , n87940 , n87941 );
not ( n87943 , n87776 );
nand ( n87944 , n87942 , n87943 );
not ( n87945 , n87781 );
nor ( n87946 , n87945 , n87721 );
buf ( n87947 , n87946 );
and ( n87948 , n87944 , n87947 );
not ( n87949 , n87944 );
not ( n87950 , n87946 );
and ( n87951 , n87949 , n87950 );
nor ( n87952 , n87948 , n87951 );
not ( n87953 , n87952 );
not ( n87954 , n87953 );
xor ( n87955 , n87922 , n87954 );
and ( n87956 , n456 , n1773 );
not ( n87957 , n456 );
and ( n87958 , n87957 , n1776 );
nor ( n87959 , n87956 , n87958 );
not ( n87960 , n87959 );
not ( n87961 , n6039 );
or ( n87962 , n87960 , n87961 );
not ( n87963 , n87959 );
nand ( n87964 , n87963 , n87906 );
nand ( n87965 , n87962 , n87964 );
not ( n87966 , n87965 );
not ( n87967 , n87966 );
nand ( n87968 , n87955 , n87967 );
nand ( n87969 , n87939 , n87968 );
xor ( n87970 , n87905 , n87969 );
not ( n87971 , n87830 );
not ( n87972 , n2910 );
or ( n87973 , n87971 , n87972 );
or ( n87974 , n2910 , n87830 );
nand ( n87975 , n87973 , n87974 );
not ( n87976 , n87975 );
buf ( n87977 , n87976 );
not ( n87978 , n87977 );
buf ( n87979 , n87707 );
not ( n87980 , n87832 );
nor ( n87981 , n87980 , n87805 );
not ( n87982 , n87981 );
not ( n87983 , n87769 );
or ( n87984 , n87982 , n87983 );
and ( n87985 , n87787 , n87832 );
nor ( n87986 , n87985 , n87845 );
nand ( n87987 , n87984 , n87986 );
not ( n87988 , n87833 );
nand ( n87989 , n87988 , n87848 );
not ( n87990 , n87989 );
and ( n87991 , n87987 , n87990 );
not ( n87992 , n87987 );
and ( n87993 , n87992 , n87989 );
nor ( n87994 , n87991 , n87993 );
buf ( n87995 , n87994 );
and ( n87996 , n87979 , n87995 );
not ( n87997 , n87979 );
not ( n87998 , n87994 );
and ( n87999 , n87997 , n87998 );
nor ( n88000 , n87996 , n87999 );
not ( n88001 , n88000 );
or ( n88002 , n87978 , n88001 );
not ( n88003 , n87979 );
and ( n88004 , n88003 , n87819 );
not ( n88005 , n88003 );
and ( n88006 , n88005 , n87822 );
nor ( n88007 , n88004 , n88006 );
not ( n88008 , n88007 );
not ( n88009 , n2176 );
not ( n88010 , n87707 );
or ( n88011 , n88009 , n88010 );
or ( n88012 , n87707 , n2176 );
nand ( n88013 , n88011 , n88012 );
nand ( n88014 , n88013 , n87975 );
not ( n88015 , n88014 );
not ( n88016 , n88015 );
or ( n88017 , n88008 , n88016 );
nand ( n88018 , n88002 , n88017 );
and ( n88019 , n87970 , n88018 );
and ( n88020 , n87905 , n87969 );
or ( n88021 , n88019 , n88020 );
xor ( n88022 , n87879 , n88021 );
not ( n88023 , n1971 );
buf ( n88024 , n2102 );
not ( n88025 , n88024 );
or ( n88026 , n88023 , n88025 );
nand ( n88027 , n88025 , n88023 );
nand ( n88028 , n88026 , n88027 );
not ( n88029 , n2065 );
and ( n88030 , n1971 , n88029 );
not ( n88031 , n1971 );
and ( n88032 , n88031 , n2065 );
or ( n88033 , n88030 , n88032 );
nand ( n88034 , n88028 , n88033 );
not ( n88035 , n88034 );
buf ( n88036 , n88035 );
not ( n88037 , n88025 );
not ( n88038 , n88023 );
and ( n88039 , n88037 , n88038 );
and ( n88040 , n88025 , n88023 );
nor ( n88041 , n88039 , n88040 );
buf ( n88042 , n88041 );
or ( n88043 , n88036 , n88042 );
not ( n88044 , n87863 );
buf ( n88045 , n88044 );
buf ( n88046 , n88045 );
not ( n88047 , n88046 );
buf ( n88048 , n88047 );
not ( n88049 , n88048 );
not ( n88050 , n88049 );
nand ( n88051 , n88043 , n88050 );
not ( n88052 , n87773 );
nor ( n88053 , n88052 , n87724 );
xor ( n88054 , n88053 , n87769 );
and ( n88055 , n87922 , n88054 );
xor ( n88056 , n88051 , n88055 );
not ( n88057 , n87871 );
not ( n88058 , n87875 );
not ( n88059 , n88058 );
nor ( n88060 , n87814 , n87790 );
nand ( n88061 , n88060 , n87988 );
nor ( n88062 , n87805 , n88061 );
not ( n88063 , n88062 );
not ( n88064 , n87769 );
or ( n88065 , n88063 , n88064 );
not ( n88066 , n88061 );
and ( n88067 , n87787 , n88066 );
not ( n88068 , n87988 );
not ( n88069 , n87845 );
or ( n88070 , n88068 , n88069 );
nand ( n88071 , n88070 , n87848 );
nor ( n88072 , n88067 , n88071 );
nand ( n88073 , n88065 , n88072 );
nor ( n88074 , n87834 , n87852 );
xor ( n88075 , n88073 , n88074 );
not ( n88076 , n88075 );
not ( n88077 , n88076 );
or ( n88078 , n88059 , n88077 );
not ( n88079 , n88076 );
nand ( n88080 , n87875 , n88079 );
nand ( n88081 , n88078 , n88080 );
not ( n88082 , n88081 );
or ( n88083 , n88057 , n88082 );
not ( n88084 , n87874 );
nand ( n88085 , n87858 , n88084 );
nand ( n88086 , n88083 , n88085 );
and ( n88087 , n88056 , n88086 );
and ( n88088 , n88051 , n88055 );
or ( n88089 , n88087 , n88088 );
not ( n88090 , n88015 );
not ( n88091 , n88000 );
or ( n88092 , n88090 , n88091 );
not ( n88093 , n87979 );
not ( n88094 , n88079 );
not ( n88095 , n88094 );
or ( n88096 , n88093 , n88095 );
nand ( n88097 , n88079 , n88003 );
nand ( n88098 , n88096 , n88097 );
nand ( n88099 , n88098 , n87977 );
nand ( n88100 , n88092 , n88099 );
xor ( n88101 , n87922 , n87901 );
not ( n88102 , n88101 );
not ( n88103 , n87967 );
or ( n88104 , n88102 , n88103 );
nand ( n88105 , n87955 , n87919 );
nand ( n88106 , n88104 , n88105 );
xor ( n88107 , n88100 , n88106 );
and ( n88108 , n87922 , n87936 );
xor ( n88109 , n88107 , n88108 );
xor ( n88110 , n88089 , n88109 );
not ( n88111 , n88046 );
not ( n88112 , n88111 );
and ( n88113 , n88112 , n87857 );
not ( n88114 , n88112 );
not ( n88115 , n87857 );
and ( n88116 , n88114 , n88115 );
nor ( n88117 , n88113 , n88116 );
not ( n88118 , n88117 );
not ( n88119 , n88036 );
or ( n88120 , n88118 , n88119 );
not ( n88121 , n88042 );
not ( n88122 , n88050 );
or ( n88123 , n88121 , n88122 );
nand ( n88124 , n88120 , n88123 );
buf ( n88125 , n2013 );
not ( n88126 , n87729 );
nor ( n88127 , n87766 , n88126 );
not ( n88128 , n88127 );
nor ( n88129 , n501 , n517 );
nor ( n88130 , n502 , n518 );
nor ( n88131 , n88129 , n88130 );
not ( n88132 , n88131 );
and ( n88133 , n504 , n520 );
not ( n88134 , n88133 );
not ( n88135 , n87756 );
or ( n88136 , n88134 , n88135 );
nand ( n88137 , n503 , n519 );
nand ( n88138 , n88136 , n88137 );
not ( n88139 , n88138 );
or ( n88140 , n88132 , n88139 );
or ( n88141 , n88129 , n87747 );
nand ( n88142 , n88141 , n87746 );
not ( n88143 , n88142 );
nand ( n88144 , n88140 , n88143 );
not ( n88145 , n88144 );
or ( n88146 , n88128 , n88145 );
not ( n88147 , n87740 );
not ( n88148 , n87729 );
not ( n88149 , n87738 );
not ( n88150 , n87737 );
and ( n88151 , n88149 , n88150 );
not ( n88152 , n87741 );
nor ( n88153 , n88151 , n88152 );
nor ( n88154 , n88148 , n88153 );
nor ( n88155 , n88147 , n88154 );
nand ( n88156 , n88146 , n88155 );
and ( n88157 , n87731 , n87734 );
xor ( n88158 , n88156 , n88157 );
buf ( n88159 , n88158 );
and ( n88160 , n88125 , n88159 );
not ( n88161 , n88084 );
not ( n88162 , n88081 );
or ( n88163 , n88161 , n88162 );
not ( n88164 , n88058 );
not ( n88165 , n87998 );
or ( n88166 , n88164 , n88165 );
nand ( n88167 , n87995 , n87875 );
nand ( n88168 , n88166 , n88167 );
nand ( n88169 , n88168 , n87871 );
nand ( n88170 , n88163 , n88169 );
xor ( n17782 , n88160 , n88170 );
not ( n88172 , n87716 );
not ( n17784 , n6120 );
not ( n88174 , n87953 );
or ( n17789 , n17784 , n88174 );
nand ( n17790 , n87954 , n87799 );
nand ( n88177 , n17789 , n17790 );
not ( n17792 , n88177 );
or ( n88179 , n88172 , n17792 );
nand ( n17797 , n87903 , n87826 );
nand ( n17798 , n88179 , n17797 );
and ( n88182 , n17782 , n17798 );
and ( n17800 , n88160 , n88170 );
or ( n88184 , n88182 , n17800 );
xor ( n17805 , n88124 , n88184 );
xor ( n17806 , n88051 , n88055 );
xor ( n88187 , n17806 , n88086 );
and ( n17808 , n17805 , n88187 );
and ( n88189 , n88124 , n88184 );
or ( n17813 , n17808 , n88189 );
xor ( n17814 , n88110 , n17813 );
xor ( n88192 , n88022 , n17814 );
not ( n17816 , n87967 );
not ( n88194 , n87937 );
or ( n17821 , n17816 , n88194 );
xor ( n88196 , n87922 , n88054 );
nand ( n88197 , n88196 , n87919 );
nand ( n88198 , n17821 , n88197 );
not ( n88199 , n88015 );
and ( n88200 , n87979 , n87795 );
not ( n88201 , n87979 );
and ( n88202 , n88201 , n87796 );
nor ( n88203 , n88200 , n88202 );
not ( n88204 , n88203 );
or ( n88205 , n88199 , n88204 );
nand ( n88206 , n88007 , n87977 );
nand ( n88207 , n88205 , n88206 );
xor ( n88208 , n88198 , n88207 );
not ( n88209 , n88124 );
and ( n88210 , n88208 , n88209 );
and ( n88211 , n88198 , n88207 );
or ( n88212 , n88210 , n88211 );
xor ( n88213 , n87905 , n87969 );
xor ( n88214 , n88213 , n88018 );
xor ( n88215 , n88212 , n88214 );
xor ( n88216 , n88124 , n88184 );
xor ( n88217 , n88216 , n88187 );
and ( n88218 , n88215 , n88217 );
and ( n88219 , n88212 , n88214 );
or ( n88220 , n88218 , n88219 );
and ( n88221 , n88192 , n88220 );
and ( n88222 , n88022 , n17814 );
or ( n88223 , n88221 , n88222 );
xor ( n88224 , n87829 , n87878 );
and ( n88225 , n88224 , n88021 );
and ( n88226 , n87829 , n87878 );
or ( n88227 , n88225 , n88226 );
xor ( n88228 , n88100 , n88106 );
and ( n88229 , n88228 , n88108 );
and ( n88230 , n88100 , n88106 );
or ( n88231 , n88229 , n88230 );
not ( n88232 , n87874 );
not ( n88233 , n87872 );
or ( n88234 , n88232 , n88233 );
nand ( n88235 , n88234 , n88058 );
not ( n88236 , n88098 );
or ( n88237 , n88236 , n88016 );
not ( n88238 , n87707 );
and ( n88239 , n88238 , n88115 );
not ( n88240 , n88238 );
and ( n88241 , n88240 , n87857 );
nor ( n88242 , n88239 , n88241 );
not ( n88243 , n87977 );
or ( n88244 , n88242 , n88243 );
nand ( n88245 , n88237 , n88244 );
xor ( n88246 , n88235 , n88245 );
not ( n88247 , n87967 );
xor ( n88248 , n87922 , n87795 );
not ( n88249 , n88248 );
or ( n88250 , n88247 , n88249 );
not ( n88251 , n88101 );
or ( n88252 , n88251 , n87918 );
nand ( n88253 , n88250 , n88252 );
xor ( n88254 , n88246 , n88253 );
xor ( n88255 , n88231 , n88254 );
and ( n88256 , n87922 , n87954 );
not ( n88257 , n87826 );
not ( n88258 , n87718 );
not ( n88259 , n87998 );
or ( n88260 , n88258 , n88259 );
nand ( n88261 , n87995 , n87799 );
nand ( n88262 , n88260 , n88261 );
not ( n88263 , n88262 );
or ( n88264 , n88257 , n88263 );
nand ( n88265 , n87824 , n87716 );
nand ( n88266 , n88264 , n88265 );
xor ( n88267 , n88256 , n88266 );
xor ( n88268 , n88267 , n87877 );
xor ( n88269 , n88255 , n88268 );
xor ( n88270 , n88227 , n88269 );
xor ( n88271 , n88089 , n88109 );
and ( n88272 , n88271 , n17813 );
and ( n88273 , n88089 , n88109 );
or ( n88274 , n88272 , n88273 );
xor ( n88275 , n88270 , n88274 );
or ( n88276 , n88223 , n88275 );
not ( n88277 , n88276 );
xor ( n88278 , n88227 , n88269 );
and ( n88279 , n88278 , n88274 );
and ( n88280 , n88227 , n88269 );
or ( n88281 , n88279 , n88280 );
and ( n88282 , n87922 , n87901 );
not ( n88283 , n87716 );
not ( n88284 , n88262 );
or ( n88285 , n88283 , n88284 );
not ( n88286 , n87718 );
not ( n88287 , n88094 );
or ( n88288 , n88286 , n88287 );
nand ( n88289 , n88079 , n87799 );
nand ( n88290 , n88288 , n88289 );
nand ( n88291 , n88290 , n87826 );
nand ( n88292 , n88285 , n88291 );
xor ( n88293 , n88282 , n88292 );
not ( n88294 , n87919 );
not ( n88295 , n88248 );
or ( n88296 , n88294 , n88295 );
xor ( n88297 , n87922 , n87822 );
nand ( n88298 , n88297 , n87967 );
nand ( n88299 , n88296 , n88298 );
xor ( n88300 , n88293 , n88299 );
or ( n88301 , n88242 , n88016 );
or ( n88302 , n88243 , n88003 );
nand ( n88303 , n88301 , n88302 );
not ( n88304 , n88303 );
xor ( n88305 , n88235 , n88245 );
and ( n88306 , n88305 , n88253 );
and ( n88307 , n88235 , n88245 );
or ( n88308 , n88306 , n88307 );
xor ( n88309 , n88304 , n88308 );
xor ( n88310 , n88256 , n88266 );
and ( n88311 , n88310 , n87877 );
and ( n88312 , n88256 , n88266 );
or ( n88313 , n88311 , n88312 );
xor ( n88314 , n88309 , n88313 );
xor ( n88315 , n88300 , n88314 );
xor ( n88316 , n88231 , n88254 );
and ( n88317 , n88316 , n88268 );
and ( n88318 , n88231 , n88254 );
or ( n88319 , n88317 , n88318 );
xor ( n88320 , n88315 , n88319 );
nor ( n88321 , n88281 , n88320 );
nor ( n88322 , n88277 , n88321 );
not ( n88323 , n88322 );
not ( n88324 , n87716 );
not ( n88325 , n87718 );
not ( n88326 , n88159 );
not ( n88327 , n88326 );
or ( n88328 , n88325 , n88327 );
nand ( n88329 , n88159 , n87799 );
nand ( n88330 , n88328 , n88329 );
not ( n88331 , n88330 );
or ( n88332 , n88324 , n88331 );
not ( n88333 , n88054 );
and ( n88334 , n88333 , n87718 );
not ( n88335 , n88333 );
and ( n88336 , n88335 , n87799 );
or ( n88337 , n88334 , n88336 );
nand ( n88338 , n88337 , n87826 );
nand ( n88339 , n88332 , n88338 );
not ( n88340 , n87919 );
not ( n88341 , n87738 );
nand ( n88342 , n88341 , n87741 );
not ( n88343 , n88342 );
not ( n88344 , n88343 );
not ( n88345 , n87748 );
not ( n88346 , n88138 );
not ( n88347 , n88346 );
or ( n88348 , n88345 , n88347 );
and ( n88349 , n87748 , n88130 );
not ( n88350 , n88129 );
or ( n88351 , n500 , n516 );
nand ( n88352 , n88350 , n88351 );
nor ( n88353 , n88349 , n88352 );
nand ( n88354 , n88348 , n88353 );
nand ( n88355 , n88354 , n87737 );
not ( n88356 , n88355 );
not ( n88357 , n88356 );
or ( n88358 , n88344 , n88357 );
nand ( n88359 , n88355 , n88342 );
nand ( n88360 , n88358 , n88359 );
not ( n88361 , n88360 );
not ( n88362 , n88361 );
xor ( n88363 , n87922 , n88362 );
not ( n88364 , n88363 );
or ( n88365 , n88340 , n88364 );
not ( n88366 , n87922 );
not ( n88367 , n87766 );
not ( n88368 , n88367 );
not ( n88369 , n88144 );
or ( n88370 , n88368 , n88369 );
nand ( n88371 , n88370 , n88153 );
not ( n88372 , n87740 );
nor ( n88373 , n88372 , n88126 );
xor ( n88374 , n88371 , n88373 );
not ( n88375 , n88374 );
not ( n88376 , n88375 );
or ( n88377 , n88366 , n88376 );
not ( n88378 , n88125 );
nand ( n88379 , n88378 , n88374 );
nand ( n88380 , n88377 , n88379 );
nand ( n88381 , n88380 , n87967 );
nand ( n88382 , n88365 , n88381 );
xor ( n88383 , n88339 , n88382 );
not ( n88384 , n87794 );
and ( n88385 , n87831 , n88384 );
not ( n88386 , n87831 );
and ( n88387 , n88386 , n87795 );
nor ( n88388 , n88385 , n88387 );
nand ( n88389 , n88388 , n88084 );
not ( n88390 , n87897 );
xor ( n88391 , n87875 , n88390 );
nand ( n88392 , n88391 , n87871 );
nand ( n88393 , n88389 , n88392 );
and ( n88394 , n88383 , n88393 );
and ( n88395 , n88339 , n88382 );
or ( n88396 , n88394 , n88395 );
not ( n88397 , n87967 );
xor ( n88398 , n88125 , n88159 );
not ( n88399 , n88398 );
or ( n88400 , n88397 , n88399 );
nand ( n88401 , n88380 , n87919 );
nand ( n88402 , n88400 , n88401 );
and ( n88403 , n87922 , n88362 );
xor ( n88404 , n88402 , n88403 );
not ( n88405 , n88042 );
and ( n88406 , n88048 , n88079 );
not ( n88407 , n88048 );
and ( n88408 , n88407 , n88076 );
nor ( n88409 , n88406 , n88408 );
not ( n88410 , n88409 );
or ( n88411 , n88405 , n88410 );
not ( n88412 , n88111 );
not ( n88413 , n87998 );
or ( n88414 , n88412 , n88413 );
not ( n88415 , n88111 );
nand ( n88416 , n87995 , n88415 );
nand ( n88417 , n88414 , n88416 );
nand ( n88418 , n88417 , n88036 );
nand ( n88419 , n88411 , n88418 );
xor ( n88420 , n88404 , n88419 );
xor ( n88421 , n88396 , n88420 );
not ( n88422 , n88015 );
and ( n88423 , n87953 , n87707 );
not ( n88424 , n87953 );
and ( n88425 , n88424 , n88238 );
or ( n88426 , n88423 , n88425 );
not ( n88427 , n88426 );
or ( n88428 , n88422 , n88427 );
not ( n88429 , n87707 );
not ( n88430 , n87898 );
or ( n88431 , n88429 , n88430 );
nand ( n88432 , n87901 , n88238 );
nand ( n88433 , n88431 , n88432 );
nand ( n88434 , n88433 , n87977 );
nand ( n88435 , n88428 , n88434 );
or ( n88436 , n2362 , n456 );
not ( n88437 , n17421 );
nand ( n88438 , n88437 , n456 );
and ( n88439 , n456 , n469 );
not ( n88440 , n456 );
and ( n88441 , n88440 , n485 );
nor ( n88442 , n88439 , n88441 );
not ( n88443 , n88442 );
nand ( n88444 , n88436 , n88438 , n88443 );
not ( n88445 , n88444 );
nand ( n88446 , n88436 , n88438 );
buf ( n88447 , n88446 );
or ( n88448 , n88445 , n88447 );
buf ( n88449 , n88442 );
not ( n88450 , n88449 );
buf ( n88451 , n88450 );
nand ( n88452 , n88448 , n88451 );
not ( n88453 , n88452 );
and ( n88454 , n88351 , n87737 );
xor ( n88455 , n88454 , n88144 );
buf ( n88456 , n88455 );
not ( n88457 , n88456 );
not ( n88458 , n88457 );
nand ( n88459 , n88458 , n87922 );
nand ( n88460 , n88453 , n88459 );
xor ( n88461 , n88435 , n88460 );
not ( n88462 , n87826 );
not ( n88463 , n87718 );
not ( n88464 , n87935 );
or ( n88465 , n88463 , n88464 );
nand ( n88466 , n87936 , n87799 );
nand ( n88467 , n88465 , n88466 );
not ( n88468 , n88467 );
or ( n88469 , n88462 , n88468 );
nand ( n88470 , n88337 , n87716 );
nand ( n88471 , n88469 , n88470 );
xor ( n88472 , n88461 , n88471 );
xor ( n88473 , n88421 , n88472 );
not ( n88474 , n88452 );
not ( n88475 , n88459 );
not ( n88476 , n88475 );
or ( n88477 , n88474 , n88476 );
nand ( n88478 , n88477 , n88460 );
nand ( n88479 , n87759 , n87747 );
not ( n88480 , n87746 );
nor ( n88481 , n88480 , n88129 );
and ( n88482 , n88479 , n88481 );
not ( n88483 , n88479 );
nand ( n88484 , n87762 , n87746 );
and ( n88485 , n88483 , n88484 );
nor ( n88486 , n88482 , n88485 );
buf ( n88487 , n88486 );
and ( n88488 , n88487 , n87922 );
not ( n88489 , n88445 );
not ( n88490 , n88451 );
not ( n88491 , n88490 );
not ( n88492 , n88115 );
or ( n88493 , n88491 , n88492 );
nand ( n88494 , n87857 , n88451 );
nand ( n88495 , n88493 , n88494 );
not ( n88496 , n88495 );
or ( n88497 , n88489 , n88496 );
nand ( n88498 , n88451 , n88447 );
nand ( n88499 , n88497 , n88498 );
and ( n88500 , n88488 , n88499 );
xor ( n88501 , n88478 , n88500 );
and ( n88502 , n88457 , n87922 );
not ( n88503 , n88457 );
and ( n88504 , n88503 , n87921 );
or ( n88505 , n88502 , n88504 );
and ( n88506 , n88505 , n87965 );
not ( n88507 , n88487 );
not ( n88508 , n87921 );
and ( n88509 , n88507 , n88508 );
and ( n88510 , n88487 , n87921 );
nor ( n88511 , n88509 , n88510 );
nor ( n88512 , n88511 , n87918 );
nor ( n88513 , n88506 , n88512 );
not ( n88514 , n88130 );
nand ( n88515 , n88514 , n87747 );
and ( n88516 , n88515 , n88346 );
not ( n88517 , n88515 );
not ( n88518 , n88346 );
and ( n88519 , n88517 , n88518 );
nor ( n88520 , n88516 , n88519 );
buf ( n88521 , n88520 );
not ( n88522 , n88521 );
or ( n88523 , n88522 , n87921 );
nor ( n88524 , n88513 , n88523 );
not ( n88525 , n87826 );
not ( n88526 , n88330 );
or ( n88527 , n88525 , n88526 );
not ( n88528 , n87718 );
not ( n88529 , n88375 );
or ( n88530 , n88528 , n88529 );
nand ( n88531 , n88374 , n87799 );
nand ( n88532 , n88530 , n88531 );
nand ( n88533 , n88532 , n87716 );
nand ( n88534 , n88527 , n88533 );
xor ( n88535 , n88524 , n88534 );
not ( n88536 , n87967 );
not ( n88537 , n88363 );
or ( n88538 , n88536 , n88537 );
nand ( n88539 , n88505 , n87919 );
nand ( n88540 , n88538 , n88539 );
and ( n88541 , n88535 , n88540 );
and ( n88542 , n88524 , n88534 );
or ( n88543 , n88541 , n88542 );
and ( n88544 , n88501 , n88543 );
and ( n88545 , n88478 , n88500 );
or ( n88546 , n88544 , n88545 );
not ( n88547 , n88084 );
not ( n88548 , n88058 );
not ( n88549 , n87819 );
or ( n88550 , n88548 , n88549 );
nand ( n88551 , n87822 , n87831 );
nand ( n88552 , n88550 , n88551 );
not ( n88553 , n88552 );
or ( n88554 , n88547 , n88553 );
nand ( n88555 , n88388 , n87871 );
nand ( n88556 , n88554 , n88555 );
not ( n88557 , n88024 );
not ( n88558 , n88557 );
and ( n88559 , n88558 , n87856 );
not ( n88560 , n88558 );
and ( n88561 , n88560 , n87857 );
nor ( n88562 , n88559 , n88561 );
not ( n88563 , n2578 );
and ( n88564 , n88024 , n88563 );
not ( n88565 , n88024 );
not ( n88566 , n88563 );
and ( n88567 , n88565 , n88566 );
nor ( n88568 , n88564 , n88567 );
not ( n88569 , n88563 );
not ( n88570 , n3052 );
or ( n88571 , n88569 , n88570 );
or ( n88572 , n3052 , n88563 );
nand ( n88573 , n88571 , n88572 );
nand ( n88574 , n88568 , n88573 );
not ( n88575 , n88574 );
and ( n88576 , n88562 , n88575 );
not ( n88577 , n88573 );
and ( n88578 , n88577 , n88558 );
nor ( n88579 , n88576 , n88578 );
xor ( n88580 , n88556 , n88579 );
not ( n88581 , n88575 );
not ( n88582 , n88025 );
xor ( n88583 , n88582 , n88075 );
not ( n88584 , n88583 );
or ( n88585 , n88581 , n88584 );
nand ( n88586 , n88562 , n88577 );
nand ( n88587 , n88585 , n88586 );
not ( n88588 , n87977 );
not ( n88589 , n88426 );
or ( n88590 , n88588 , n88589 );
not ( n88591 , n87707 );
not ( n88592 , n87935 );
or ( n88593 , n88591 , n88592 );
nand ( n88594 , n87934 , n88238 );
nand ( n88595 , n88593 , n88594 );
nand ( n88596 , n88595 , n88015 );
nand ( n88597 , n88590 , n88596 );
xor ( n88598 , n88587 , n88597 );
not ( n88599 , n88042 );
not ( n88600 , n88417 );
or ( n88601 , n88599 , n88600 );
not ( n88602 , n88045 );
buf ( n88603 , n88602 );
not ( n88604 , n88603 );
not ( n88605 , n88604 );
not ( n88606 , n88605 );
not ( n88607 , n87819 );
or ( n88608 , n88606 , n88607 );
nand ( n88609 , n87822 , n88049 );
nand ( n88610 , n88608 , n88609 );
nand ( n88611 , n88610 , n88036 );
nand ( n88612 , n88601 , n88611 );
and ( n88613 , n88598 , n88612 );
and ( n88614 , n88587 , n88597 );
or ( n88615 , n88613 , n88614 );
xor ( n88616 , n88580 , n88615 );
xor ( n88617 , n88546 , n88616 );
not ( n88618 , n87871 );
not ( n88619 , n88058 );
and ( n88620 , n87944 , n87947 );
not ( n88621 , n87944 );
and ( n88622 , n88621 , n87950 );
nor ( n88623 , n88620 , n88622 );
not ( n88624 , n88623 );
not ( n88625 , n88624 );
or ( n88626 , n88619 , n88625 );
not ( n88627 , n88623 );
or ( n88628 , n88627 , n87830 );
nand ( n88629 , n88626 , n88628 );
not ( n88630 , n88629 );
or ( n88631 , n88618 , n88630 );
nand ( n88632 , n88391 , n88084 );
nand ( n88633 , n88631 , n88632 );
not ( n88634 , n88577 );
not ( n88635 , n88583 );
or ( n88636 , n88634 , n88635 );
not ( n88637 , n88557 );
not ( n88638 , n87994 );
or ( n88639 , n88637 , n88638 );
not ( n88640 , n88558 );
or ( n88641 , n87994 , n88640 );
nand ( n88642 , n88639 , n88641 );
nand ( n88643 , n88642 , n88575 );
nand ( n88644 , n88636 , n88643 );
xor ( n88645 , n88633 , n88644 );
not ( n88646 , n88015 );
not ( n88647 , n87707 );
not ( n88648 , n88333 );
or ( n88649 , n88647 , n88648 );
nand ( n88650 , n88054 , n88238 );
nand ( n88651 , n88649 , n88650 );
not ( n88652 , n88651 );
or ( n88653 , n88646 , n88652 );
nand ( n88654 , n88595 , n87977 );
nand ( n88655 , n88653 , n88654 );
and ( n88656 , n88645 , n88655 );
and ( n88657 , n88633 , n88644 );
or ( n88658 , n88656 , n88657 );
xor ( n88659 , n88339 , n88382 );
xor ( n88660 , n88659 , n88393 );
xor ( n88661 , n88658 , n88660 );
xor ( n88662 , n88587 , n88597 );
xor ( n88663 , n88662 , n88612 );
and ( n88664 , n88661 , n88663 );
and ( n88665 , n88658 , n88660 );
or ( n88666 , n88664 , n88665 );
xor ( n88667 , n88617 , n88666 );
xor ( n88668 , n88473 , n88667 );
not ( n88669 , n88036 );
not ( n88670 , n88050 );
not ( n88671 , n87796 );
or ( n88672 , n88670 , n88671 );
nand ( n88673 , n87795 , n88049 );
nand ( n88674 , n88672 , n88673 );
not ( n88675 , n88674 );
or ( n88676 , n88669 , n88675 );
nand ( n88677 , n88610 , n88042 );
nand ( n88678 , n88676 , n88677 );
xor ( n88679 , n88488 , n88499 );
xor ( n88680 , n88678 , n88679 );
xor ( n88681 , n88513 , n88523 );
not ( n88682 , n88015 );
not ( n88683 , n87707 );
not ( n88684 , n88326 );
or ( n88685 , n88683 , n88684 );
nand ( n88686 , n88159 , n88238 );
nand ( n88687 , n88685 , n88686 );
not ( n88688 , n88687 );
or ( n88689 , n88682 , n88688 );
nand ( n88690 , n88651 , n87977 );
nand ( n88691 , n88689 , n88690 );
and ( n88692 , n88681 , n88691 );
and ( n88693 , n88680 , n88692 );
and ( n88694 , n88678 , n88679 );
or ( n88695 , n88693 , n88694 );
xor ( n88696 , n88478 , n88500 );
xor ( n88697 , n88696 , n88543 );
xor ( n88698 , n88695 , n88697 );
not ( n88699 , n87716 );
and ( n88700 , n88362 , n87799 );
not ( n88701 , n88362 );
and ( n88702 , n88701 , n87718 );
or ( n88703 , n88700 , n88702 );
not ( n88704 , n88703 );
or ( n88705 , n88699 , n88704 );
nand ( n88706 , n88532 , n87826 );
nand ( n88707 , n88705 , n88706 );
and ( n88708 , n87934 , n88058 );
not ( n88709 , n87934 );
and ( n88710 , n88709 , n87831 );
nor ( n88711 , n88708 , n88710 );
not ( n88712 , n88711 );
or ( n88713 , n88712 , n87872 );
not ( n88714 , n88629 );
or ( n88715 , n88714 , n87874 );
nand ( n88716 , n88713 , n88715 );
xor ( n88717 , n88707 , n88716 );
not ( n88718 , n88495 );
not ( n88719 , n88447 );
or ( n88720 , n88718 , n88719 );
and ( n88721 , n88075 , n88451 );
not ( n88722 , n88075 );
and ( n88723 , n88722 , n88490 );
or ( n88724 , n88721 , n88723 );
or ( n88725 , n88724 , n88444 );
nand ( n88726 , n88720 , n88725 );
and ( n88727 , n88717 , n88726 );
and ( n88728 , n88707 , n88716 );
or ( n88729 , n88727 , n88728 );
xor ( n88730 , n88524 , n88534 );
xor ( n88731 , n88730 , n88540 );
xor ( n88732 , n88729 , n88731 );
xor ( n88733 , n88633 , n88644 );
xor ( n88734 , n88733 , n88655 );
and ( n88735 , n88732 , n88734 );
and ( n88736 , n88729 , n88731 );
or ( n88737 , n88735 , n88736 );
and ( n88738 , n88698 , n88737 );
and ( n88739 , n88695 , n88697 );
or ( n88740 , n88738 , n88739 );
xor ( n88741 , n88668 , n88740 );
xor ( n88742 , n88658 , n88660 );
xor ( n88743 , n88742 , n88663 );
xor ( n88744 , n88678 , n88679 );
xor ( n88745 , n88744 , n88692 );
not ( n88746 , n88575 );
not ( n88747 , n88558 );
not ( n88748 , n87819 );
or ( n88749 , n88747 , n88748 );
not ( n88750 , n88582 );
nand ( n88751 , n87818 , n88750 );
nand ( n88752 , n88749 , n88751 );
not ( n88753 , n88752 );
or ( n88754 , n88746 , n88753 );
nand ( n88755 , n88642 , n88577 );
nand ( n88756 , n88754 , n88755 );
not ( n88757 , n88036 );
not ( n88758 , n88604 );
and ( n88759 , n88758 , n87901 );
not ( n88760 , n88758 );
and ( n88761 , n88760 , n87898 );
nor ( n88762 , n88759 , n88761 );
not ( n88763 , n88762 );
or ( n88764 , n88757 , n88763 );
nand ( n88765 , n88674 , n88042 );
nand ( n88766 , n88764 , n88765 );
xor ( n88767 , n88756 , n88766 );
not ( n88768 , n87965 );
not ( n88769 , n88511 );
not ( n88770 , n88769 );
or ( n88771 , n88768 , n88770 );
not ( n88772 , n88125 );
not ( n88773 , n88521 );
not ( n88774 , n88773 );
or ( n88775 , n88772 , n88774 );
nand ( n88776 , n88521 , n87921 );
nand ( n88777 , n88775 , n88776 );
nand ( n88778 , n88777 , n87919 );
nand ( n88779 , n88771 , n88778 );
nand ( n88780 , n504 , n520 );
not ( n88781 , n88780 );
nand ( n88782 , n87756 , n88137 );
not ( n88783 , n88782 );
not ( n88784 , n88783 );
or ( n88785 , n88781 , n88784 );
not ( n88786 , n88780 );
nand ( n88787 , n88786 , n88782 );
nand ( n88788 , n88785 , n88787 );
buf ( n88789 , n88788 );
and ( n88790 , n88125 , n88789 );
xor ( n88791 , n88779 , n88790 );
not ( n88792 , n87826 );
not ( n88793 , n88703 );
or ( n88794 , n88792 , n88793 );
not ( n88795 , n87718 );
not ( n88796 , n88457 );
or ( n88797 , n88795 , n88796 );
nand ( n88798 , n88456 , n87799 );
nand ( n88799 , n88797 , n88798 );
nand ( n88800 , n88799 , n87716 );
nand ( n88801 , n88794 , n88800 );
and ( n88802 , n88791 , n88801 );
and ( n88803 , n88779 , n88790 );
or ( n88804 , n88802 , n88803 );
and ( n88805 , n88767 , n88804 );
and ( n88806 , n88756 , n88766 );
or ( n88807 , n88805 , n88806 );
xor ( n88808 , n88745 , n88807 );
xor ( n88809 , n88681 , n88691 );
not ( n88810 , n87977 );
not ( n88811 , n88687 );
or ( n88812 , n88810 , n88811 );
not ( n88813 , n87707 );
not ( n88814 , n88375 );
or ( n88815 , n88813 , n88814 );
nand ( n88816 , n88374 , n88238 );
nand ( n88817 , n88815 , n88816 );
nand ( n88818 , n88817 , n88015 );
nand ( n88819 , n88812 , n88818 );
not ( n88820 , n88084 );
not ( n88821 , n88711 );
or ( n88822 , n88820 , n88821 );
and ( n88823 , n88333 , n88058 );
not ( n88824 , n88333 );
and ( n88825 , n88824 , n87875 );
or ( n88826 , n88823 , n88825 );
nand ( n88827 , n88826 , n87871 );
nand ( n88828 , n88822 , n88827 );
xor ( n88829 , n88819 , n88828 );
not ( n88830 , n87994 );
not ( n88831 , n88490 );
and ( n88832 , n88830 , n88831 );
and ( n88833 , n87995 , n88490 );
nor ( n88834 , n88832 , n88833 );
or ( n88835 , n88834 , n88444 );
not ( n88836 , n88447 );
or ( n88837 , n88724 , n88836 );
nand ( n88838 , n88835 , n88837 );
and ( n88839 , n88829 , n88838 );
and ( n88840 , n88819 , n88828 );
or ( n88841 , n88839 , n88840 );
xor ( n88842 , n88809 , n88841 );
not ( n88843 , n88577 );
not ( n88844 , n88752 );
or ( n88845 , n88843 , n88844 );
not ( n88846 , n88557 );
not ( n88847 , n87794 );
or ( n88848 , n88846 , n88847 );
or ( n88849 , n87794 , n88640 );
nand ( n88850 , n88848 , n88849 );
nand ( n88851 , n88850 , n88575 );
nand ( n88852 , n88845 , n88851 );
xor ( n88853 , n504 , n520 );
not ( n88854 , n88853 );
not ( n88855 , n88854 );
and ( n88856 , n88855 , n88125 );
not ( n88857 , n87919 );
xor ( n88858 , n88125 , n88789 );
not ( n88859 , n88858 );
or ( n88860 , n88857 , n88859 );
nand ( n88861 , n88777 , n87965 );
nand ( n88862 , n88860 , n88861 );
xor ( n88863 , n88856 , n88862 );
not ( n88864 , n87918 );
and ( n88865 , n88125 , n88854 );
not ( n88866 , n88125 );
buf ( n88867 , n88853 );
and ( n88868 , n88866 , n88867 );
nor ( n88869 , n88865 , n88868 );
not ( n88870 , n88869 );
and ( n88871 , n88864 , n88870 );
and ( n88872 , n87965 , n88858 );
nor ( n88873 , n88871 , n88872 );
and ( n88874 , n6120 , n87906 );
nor ( n88875 , n88874 , n87913 );
not ( n88876 , n87911 );
not ( n88877 , n75980 );
or ( n88878 , n88876 , n88877 );
nand ( n88879 , n88878 , n88855 );
nand ( n88880 , n88875 , n88879 );
nor ( n88881 , n88873 , n88880 );
and ( n88882 , n88863 , n88881 );
and ( n88883 , n88856 , n88862 );
or ( n88884 , n88882 , n88883 );
xor ( n88885 , n88852 , n88884 );
not ( n88886 , n88036 );
not ( n88887 , n88048 );
not ( n88888 , n87953 );
or ( n88889 , n88887 , n88888 );
nand ( n88890 , n87954 , n88604 );
nand ( n88891 , n88889 , n88890 );
not ( n88892 , n88891 );
or ( n88893 , n88886 , n88892 );
nand ( n88894 , n88762 , n88042 );
nand ( n88895 , n88893 , n88894 );
and ( n88896 , n88885 , n88895 );
and ( n88897 , n88852 , n88884 );
or ( n88898 , n88896 , n88897 );
and ( n88899 , n88842 , n88898 );
and ( n88900 , n88809 , n88841 );
or ( n88901 , n88899 , n88900 );
and ( n88902 , n88808 , n88901 );
and ( n88903 , n88745 , n88807 );
or ( n88904 , n88902 , n88903 );
xor ( n88905 , n88743 , n88904 );
xor ( n88906 , n88695 , n88697 );
xor ( n88907 , n88906 , n88737 );
and ( n88908 , n88905 , n88907 );
and ( n88909 , n88743 , n88904 );
or ( n88910 , n88908 , n88909 );
nor ( n88911 , n88741 , n88910 );
xor ( n88912 , n88729 , n88731 );
xor ( n88913 , n88912 , n88734 );
xor ( n88914 , n88745 , n88807 );
xor ( n88915 , n88914 , n88901 );
xor ( n88916 , n88913 , n88915 );
xor ( n88917 , n88707 , n88716 );
xor ( n88918 , n88917 , n88726 );
xor ( n88919 , n88756 , n88766 );
xor ( n88920 , n88919 , n88804 );
xor ( n88921 , n88918 , n88920 );
not ( n88922 , n87708 );
not ( n88923 , n88799 );
or ( n88924 , n88922 , n88923 );
and ( n88925 , n88487 , n87799 );
not ( n88926 , n88487 );
and ( n88927 , n88926 , n87718 );
or ( n88928 , n88925 , n88927 );
nand ( n88929 , n88928 , n87716 );
nand ( n88930 , n88924 , n88929 );
not ( n88931 , n88015 );
not ( n88932 , n88361 );
and ( n88933 , n87707 , n88932 );
not ( n88934 , n87707 );
and ( n88935 , n88934 , n88361 );
nor ( n88936 , n88933 , n88935 );
not ( n88937 , n88936 );
or ( n88938 , n88931 , n88937 );
nand ( n88939 , n88817 , n87977 );
nand ( n88940 , n88938 , n88939 );
xor ( n88941 , n88930 , n88940 );
not ( n88942 , n87871 );
not ( n88943 , n88058 );
not ( n88944 , n88326 );
or ( n88945 , n88943 , n88944 );
nand ( n88946 , n88159 , n87875 );
nand ( n88947 , n88945 , n88946 );
not ( n88948 , n88947 );
or ( n88949 , n88942 , n88948 );
nand ( n88950 , n88826 , n88084 );
nand ( n88951 , n88949 , n88950 );
and ( n88952 , n88941 , n88951 );
and ( n88953 , n88930 , n88940 );
or ( n88954 , n88952 , n88953 );
xor ( n88955 , n88779 , n88790 );
xor ( n88956 , n88955 , n88801 );
xor ( n88957 , n88954 , n88956 );
xor ( n88958 , n88856 , n88862 );
xor ( n88959 , n88958 , n88881 );
not ( n88960 , n88575 );
and ( n88961 , n88557 , n87898 );
not ( n88962 , n88557 );
and ( n88963 , n88962 , n87901 );
nor ( n88964 , n88961 , n88963 );
not ( n88965 , n88964 );
or ( n88966 , n88960 , n88965 );
nand ( n88967 , n88850 , n88577 );
nand ( n88968 , n88966 , n88967 );
xor ( n88969 , n88959 , n88968 );
not ( n88970 , n88490 );
not ( n88971 , n87818 );
or ( n88972 , n88970 , n88971 );
or ( n88973 , n87822 , n88490 );
nand ( n88974 , n88972 , n88973 );
not ( n88975 , n88974 );
not ( n88976 , n88445 );
or ( n88977 , n88975 , n88976 );
or ( n88978 , n88834 , n88836 );
nand ( n88979 , n88977 , n88978 );
and ( n88980 , n88969 , n88979 );
and ( n88981 , n88959 , n88968 );
or ( n88982 , n88980 , n88981 );
and ( n88983 , n88957 , n88982 );
and ( n88984 , n88954 , n88956 );
or ( n88985 , n88983 , n88984 );
and ( n88986 , n88921 , n88985 );
and ( n88987 , n88918 , n88920 );
or ( n88988 , n88986 , n88987 );
and ( n88989 , n88916 , n88988 );
and ( n88990 , n88913 , n88915 );
or ( n88991 , n88989 , n88990 );
xor ( n88992 , n88743 , n88904 );
xor ( n88993 , n88992 , n88907 );
nor ( n88994 , n88991 , n88993 );
nor ( n88995 , n88911 , n88994 );
xor ( n88996 , n88396 , n88420 );
and ( n88997 , n88996 , n88472 );
and ( n88998 , n88396 , n88420 );
or ( n88999 , n88997 , n88998 );
not ( n89000 , n88084 );
not ( n89001 , n88168 );
or ( n89002 , n89000 , n89001 );
nand ( n89003 , n88552 , n87871 );
nand ( n89004 , n89002 , n89003 );
not ( n89005 , n88579 );
xor ( n89006 , n89004 , n89005 );
xor ( n89007 , n88402 , n88403 );
and ( n89008 , n89007 , n88419 );
and ( n89009 , n88402 , n88403 );
or ( n89010 , n89008 , n89009 );
xor ( n89011 , n89006 , n89010 );
xor ( n89012 , n88556 , n88579 );
and ( n89013 , n89012 , n88615 );
and ( n89014 , n88556 , n88579 );
or ( n89015 , n89013 , n89014 );
xor ( n89016 , n89011 , n89015 );
xor ( n89017 , n88435 , n88460 );
and ( n89018 , n89017 , n88471 );
and ( n89019 , n88435 , n88460 );
or ( n89020 , n89018 , n89019 );
not ( n89021 , n88573 );
not ( n89022 , n88574 );
or ( n89023 , n89021 , n89022 );
nand ( n89024 , n89023 , n88558 );
not ( n89025 , n87919 );
not ( n89026 , n88398 );
or ( n89027 , n89025 , n89026 );
nand ( n89028 , n88196 , n87967 );
nand ( n89029 , n89027 , n89028 );
xor ( n89030 , n89024 , n89029 );
not ( n89031 , n87922 );
nor ( n89032 , n89031 , n88375 );
xor ( n89033 , n89030 , n89032 );
xor ( n89034 , n89020 , n89033 );
not ( n89035 , n88036 );
not ( n89036 , n88409 );
or ( n89037 , n89035 , n89036 );
nand ( n89038 , n88117 , n88042 );
nand ( n89039 , n89037 , n89038 );
not ( n89040 , n87977 );
not ( n89041 , n88203 );
or ( n89042 , n89040 , n89041 );
nand ( n89043 , n88433 , n88015 );
nand ( n89044 , n89042 , n89043 );
xor ( n89045 , n89039 , n89044 );
not ( n89046 , n87826 );
not ( n89047 , n88177 );
or ( n89048 , n89046 , n89047 );
nand ( n89049 , n88467 , n87716 );
nand ( n89050 , n89048 , n89049 );
xor ( n89051 , n89045 , n89050 );
xor ( n89052 , n89034 , n89051 );
xor ( n89053 , n89016 , n89052 );
xor ( n89054 , n88999 , n89053 );
xor ( n89055 , n88546 , n88616 );
and ( n89056 , n89055 , n88666 );
and ( n89057 , n88546 , n88616 );
or ( n89058 , n89056 , n89057 );
and ( n89059 , n89054 , n89058 );
and ( n89060 , n88999 , n89053 );
or ( n89061 , n89059 , n89060 );
not ( n89062 , n89061 );
xor ( n89063 , n89024 , n89029 );
and ( n89064 , n89063 , n89032 );
and ( n89065 , n89024 , n89029 );
or ( n89066 , n89064 , n89065 );
xor ( n89067 , n89039 , n89044 );
and ( n89068 , n89067 , n89050 );
and ( n89069 , n89039 , n89044 );
or ( n89070 , n89068 , n89069 );
xor ( n89071 , n89066 , n89070 );
xor ( n89072 , n88198 , n88207 );
xor ( n89073 , n89072 , n88209 );
xor ( n89074 , n89071 , n89073 );
xor ( n89075 , n88160 , n88170 );
xor ( n89076 , n89075 , n17798 );
xor ( n89077 , n89004 , n89005 );
and ( n89078 , n89077 , n89010 );
and ( n89079 , n89004 , n89005 );
or ( n89080 , n89078 , n89079 );
xor ( n89081 , n89076 , n89080 );
xor ( n89082 , n89020 , n89033 );
and ( n89083 , n89082 , n89051 );
and ( n89084 , n89020 , n89033 );
or ( n89085 , n89083 , n89084 );
xor ( n89086 , n89081 , n89085 );
xor ( n89087 , n89074 , n89086 );
xor ( n89088 , n89011 , n89015 );
and ( n89089 , n89088 , n89052 );
and ( n89090 , n89011 , n89015 );
or ( n89091 , n89089 , n89090 );
xor ( n89092 , n89087 , n89091 );
not ( n89093 , n89092 );
nand ( n89094 , n89062 , n89093 );
xor ( n89095 , n88999 , n89053 );
xor ( n89096 , n89095 , n89058 );
not ( n89097 , n89096 );
xor ( n89098 , n88473 , n88667 );
and ( n89099 , n89098 , n88740 );
and ( n89100 , n88473 , n88667 );
or ( n89101 , n89099 , n89100 );
not ( n89102 , n89101 );
nand ( n89103 , n89097 , n89102 );
and ( n89104 , n88995 , n89094 , n89103 );
not ( n89105 , n89104 );
xor ( n89106 , n88809 , n88841 );
xor ( n89107 , n89106 , n88898 );
xor ( n89108 , n88918 , n88920 );
xor ( n89109 , n89108 , n88985 );
xor ( n89110 , n89107 , n89109 );
xor ( n89111 , n88852 , n88884 );
xor ( n89112 , n89111 , n88895 );
xor ( n89113 , n88819 , n88828 );
xor ( n89114 , n89113 , n88838 );
xor ( n89115 , n89112 , n89114 );
xor ( n89116 , n88954 , n88956 );
xor ( n89117 , n89116 , n88982 );
and ( n89118 , n89115 , n89117 );
and ( n89119 , n89112 , n89114 );
or ( n89120 , n89118 , n89119 );
xor ( n89121 , n89110 , n89120 );
not ( n89122 , n89121 );
not ( n89123 , n88042 );
not ( n89124 , n88891 );
or ( n89125 , n89123 , n89124 );
not ( n89126 , n88605 );
not ( n89127 , n87935 );
or ( n89128 , n89126 , n89127 );
nand ( n89129 , n87936 , n88415 );
nand ( n89130 , n89128 , n89129 );
nand ( n89131 , n89130 , n88036 );
nand ( n89132 , n89125 , n89131 );
not ( n89133 , n87826 );
not ( n89134 , n88928 );
or ( n89135 , n89133 , n89134 );
not ( n89136 , n6120 );
not ( n89137 , n88522 );
or ( n89138 , n89136 , n89137 );
nand ( n89139 , n88521 , n87799 );
nand ( n89140 , n89138 , n89139 );
nand ( n89141 , n89140 , n87716 );
nand ( n89142 , n89135 , n89141 );
xor ( n89143 , n88873 , n88880 );
xor ( n89144 , n89142 , n89143 );
not ( n89145 , n87977 );
not ( n89146 , n88936 );
or ( n89147 , n89145 , n89146 );
not ( n89148 , n87707 );
not ( n89149 , n88457 );
or ( n89150 , n89148 , n89149 );
nand ( n89151 , n88456 , n88238 );
nand ( n89152 , n89150 , n89151 );
nand ( n89153 , n89152 , n88015 );
nand ( n89154 , n89147 , n89153 );
and ( n89155 , n89144 , n89154 );
and ( n89156 , n89142 , n89143 );
or ( n89157 , n89155 , n89156 );
xor ( n89158 , n89132 , n89157 );
xor ( n89159 , n88930 , n88940 );
xor ( n89160 , n89159 , n88951 );
and ( n89161 , n89158 , n89160 );
and ( n89162 , n89132 , n89157 );
or ( n89163 , n89161 , n89162 );
not ( n89164 , n88084 );
not ( n89165 , n88947 );
or ( n89166 , n89164 , n89165 );
not ( n89167 , n88058 );
not ( n89168 , n88375 );
or ( n89169 , n89167 , n89168 );
nand ( n89170 , n88374 , n87875 );
nand ( n89171 , n89169 , n89170 );
nand ( n89172 , n89171 , n87871 );
nand ( n89173 , n89166 , n89172 );
not ( n89174 , n88577 );
not ( n89175 , n88964 );
or ( n89176 , n89174 , n89175 );
not ( n89177 , n87953 );
not ( n89178 , n88558 );
or ( n89179 , n89177 , n89178 );
nand ( n89180 , n88623 , n88557 );
nand ( n89181 , n89179 , n89180 );
nand ( n89182 , n89181 , n88575 );
nand ( n89183 , n89176 , n89182 );
xor ( n89184 , n89173 , n89183 );
and ( n89185 , n87965 , n88855 );
not ( n89186 , n87708 );
not ( n89187 , n89140 );
or ( n89188 , n89186 , n89187 );
not ( n89189 , n6120 );
not ( n89190 , n88789 );
not ( n89191 , n89190 );
or ( n89192 , n89189 , n89191 );
nand ( n89193 , n88789 , n75980 );
nand ( n89194 , n89192 , n89193 );
nand ( n89195 , n89194 , n87714 );
nand ( n89196 , n89188 , n89195 );
xor ( n89197 , n89185 , n89196 );
nand ( n89198 , n88238 , n6022 );
and ( n89199 , n89198 , n88855 );
not ( n89200 , n1982 );
not ( n89201 , n87707 );
or ( n89202 , n89200 , n89201 );
nand ( n89203 , n89202 , n6120 );
nor ( n89204 , n89199 , n89203 );
not ( n89205 , n87708 );
not ( n89206 , n89194 );
or ( n89207 , n89205 , n89206 );
not ( n89208 , n6120 );
not ( n89209 , n88854 );
or ( n89210 , n89208 , n89209 );
nand ( n89211 , n75980 , n88855 );
nand ( n89212 , n89210 , n89211 );
nand ( n89213 , n87714 , n89212 );
nand ( n89214 , n89207 , n89213 );
and ( n89215 , n89204 , n89214 );
and ( n89216 , n89197 , n89215 );
and ( n89217 , n89185 , n89196 );
or ( n89218 , n89216 , n89217 );
and ( n89219 , n89184 , n89218 );
and ( n89220 , n89173 , n89183 );
or ( n89221 , n89219 , n89220 );
xor ( n89222 , n88959 , n88968 );
xor ( n89223 , n89222 , n88979 );
xor ( n89224 , n89221 , n89223 );
not ( n89225 , n88445 );
not ( n89226 , n88449 );
and ( n89227 , n89226 , n87795 );
not ( n89228 , n89226 );
and ( n89229 , n89228 , n88384 );
nor ( n89230 , n89227 , n89229 );
not ( n89231 , n89230 );
or ( n89232 , n89225 , n89231 );
nand ( n89233 , n88974 , n88447 );
nand ( n89234 , n89232 , n89233 );
not ( n89235 , n88042 );
not ( n89236 , n89130 );
or ( n89237 , n89235 , n89236 );
and ( n89238 , n88603 , n88054 );
not ( n89239 , n88603 );
and ( n89240 , n89239 , n88333 );
nor ( n89241 , n89238 , n89240 );
nand ( n89242 , n89241 , n88036 );
nand ( n89243 , n89237 , n89242 );
xor ( n89244 , n89234 , n89243 );
xor ( n89245 , n89142 , n89143 );
xor ( n89246 , n89245 , n89154 );
and ( n89247 , n89244 , n89246 );
and ( n89248 , n89234 , n89243 );
or ( n89249 , n89247 , n89248 );
and ( n89250 , n89224 , n89249 );
and ( n89251 , n89221 , n89223 );
or ( n89252 , n89250 , n89251 );
xor ( n89253 , n89163 , n89252 );
xor ( n89254 , n89112 , n89114 );
xor ( n89255 , n89254 , n89117 );
and ( n89256 , n89253 , n89255 );
and ( n89257 , n89163 , n89252 );
or ( n89258 , n89256 , n89257 );
not ( n89259 , n89258 );
and ( n89260 , n89122 , n89259 );
xor ( n89261 , n88913 , n88915 );
xor ( n89262 , n89261 , n88988 );
xor ( n89263 , n89107 , n89109 );
and ( n89264 , n89263 , n89120 );
and ( n89265 , n89107 , n89109 );
or ( n89266 , n89264 , n89265 );
nor ( n89267 , n89262 , n89266 );
nor ( n89268 , n89260 , n89267 );
not ( n89269 , n89268 );
xor ( n89270 , n89163 , n89252 );
xor ( n89271 , n89270 , n89255 );
not ( n89272 , n89271 );
xor ( n89273 , n89132 , n89157 );
xor ( n89274 , n89273 , n89160 );
not ( n89275 , n87977 );
not ( n89276 , n89152 );
or ( n89277 , n89275 , n89276 );
not ( n89278 , n87707 );
not ( n89279 , n88487 );
not ( n89280 , n89279 );
or ( n89281 , n89278 , n89280 );
nand ( n89282 , n88487 , n88238 );
nand ( n89283 , n89281 , n89282 );
nand ( n89284 , n89283 , n88015 );
nand ( n89285 , n89277 , n89284 );
not ( n89286 , n88036 );
and ( n89287 , n88159 , n88111 );
not ( n89288 , n88159 );
and ( n89289 , n89288 , n88604 );
nor ( n89290 , n89287 , n89289 );
not ( n89291 , n89290 );
or ( n89292 , n89286 , n89291 );
nand ( n89293 , n89241 , n88042 );
nand ( n89294 , n89292 , n89293 );
xor ( n89295 , n89285 , n89294 );
not ( n89296 , n88084 );
not ( n89297 , n89171 );
or ( n89298 , n89296 , n89297 );
not ( n89299 , n87830 );
not ( n89300 , n88361 );
or ( n89301 , n89299 , n89300 );
nand ( n89302 , n88360 , n87875 );
nand ( n89303 , n89301 , n89302 );
nand ( n89304 , n89303 , n87871 );
nand ( n89305 , n89298 , n89304 );
and ( n89306 , n89295 , n89305 );
and ( n89307 , n89285 , n89294 );
or ( n89308 , n89306 , n89307 );
not ( n89309 , n88575 );
and ( n89310 , n87934 , n88557 );
not ( n89311 , n87934 );
and ( n89312 , n89311 , n88558 );
or ( n89313 , n89310 , n89312 );
not ( n89314 , n89313 );
or ( n89315 , n89309 , n89314 );
nand ( n89316 , n89181 , n88577 );
nand ( n89317 , n89315 , n89316 );
xor ( n89318 , n89185 , n89196 );
xor ( n89319 , n89318 , n89215 );
xor ( n89320 , n89317 , n89319 );
not ( n89321 , n88445 );
not ( n89322 , n88451 );
not ( n89323 , n87898 );
or ( n89324 , n89322 , n89323 );
nand ( n89325 , n87901 , n88490 );
nand ( n89326 , n89324 , n89325 );
not ( n89327 , n89326 );
or ( n89328 , n89321 , n89327 );
nand ( n89329 , n89230 , n88447 );
nand ( n89330 , n89328 , n89329 );
and ( n89331 , n89320 , n89330 );
and ( n89332 , n89317 , n89319 );
or ( n89333 , n89331 , n89332 );
xor ( n89334 , n89308 , n89333 );
xor ( n89335 , n89173 , n89183 );
xor ( n89336 , n89335 , n89218 );
and ( n89337 , n89334 , n89336 );
and ( n89338 , n89308 , n89333 );
or ( n89339 , n89337 , n89338 );
xor ( n89340 , n89274 , n89339 );
xor ( n89341 , n89221 , n89223 );
xor ( n89342 , n89341 , n89249 );
and ( n89343 , n89340 , n89342 );
and ( n89344 , n89274 , n89339 );
or ( n89345 , n89343 , n89344 );
not ( n89346 , n89345 );
and ( n89347 , n89272 , n89346 );
xor ( n89348 , n89274 , n89339 );
xor ( n89349 , n89348 , n89342 );
xor ( n89350 , n89234 , n89243 );
xor ( n89351 , n89350 , n89246 );
not ( n89352 , n87976 );
not ( n89353 , n89283 );
or ( n89354 , n89352 , n89353 );
not ( n89355 , n87707 );
not ( n89356 , n88522 );
or ( n89357 , n89355 , n89356 );
nand ( n89358 , n88521 , n88238 );
nand ( n89359 , n89357 , n89358 );
nand ( n89360 , n89359 , n88015 );
nand ( n89361 , n89354 , n89360 );
xor ( n89362 , n89204 , n89214 );
xor ( n89363 , n89361 , n89362 );
not ( n89364 , n87869 );
not ( n89365 , n89303 );
or ( n89366 , n89364 , n89365 );
not ( n89367 , n87830 );
not ( n89368 , n88457 );
or ( n89369 , n89367 , n89368 );
nand ( n89370 , n88456 , n87875 );
nand ( n89371 , n89369 , n89370 );
nand ( n89372 , n89371 , n87871 );
nand ( n89373 , n89366 , n89372 );
and ( n89374 , n89363 , n89373 );
and ( n89375 , n89361 , n89362 );
or ( n89376 , n89374 , n89375 );
xor ( n89377 , n89285 , n89294 );
xor ( n89378 , n89377 , n89305 );
xor ( n89379 , n89376 , n89378 );
not ( n89380 , n88036 );
not ( n89381 , n88046 );
not ( n89382 , n89381 );
not ( n89383 , n88375 );
or ( n89384 , n89382 , n89383 );
not ( n89385 , n89381 );
nand ( n89386 , n88374 , n89385 );
nand ( n89387 , n89384 , n89386 );
not ( n89388 , n89387 );
or ( n89389 , n89380 , n89388 );
nand ( n89390 , n89290 , n88042 );
nand ( n89391 , n89389 , n89390 );
and ( n89392 , n87708 , n88855 );
not ( n89393 , n87976 );
not ( n89394 , n89359 );
or ( n89395 , n89393 , n89394 );
not ( n89396 , n87707 );
not ( n89397 , n89190 );
or ( n89398 , n89396 , n89397 );
nand ( n89399 , n88789 , n88238 );
nand ( n89400 , n89398 , n89399 );
nand ( n89401 , n89400 , n88015 );
nand ( n89402 , n89395 , n89401 );
xor ( n89403 , n89392 , n89402 );
not ( n89404 , n88084 );
not ( n89405 , n89371 );
or ( n89406 , n89404 , n89405 );
not ( n89407 , n87830 );
not ( n89408 , n89279 );
or ( n89409 , n89407 , n89408 );
nand ( n89410 , n88487 , n87831 );
nand ( n89411 , n89409 , n89410 );
nand ( n89412 , n89411 , n87870 );
nand ( n89413 , n89406 , n89412 );
and ( n89414 , n89403 , n89413 );
and ( n89415 , n89392 , n89402 );
or ( n89416 , n89414 , n89415 );
xor ( n89417 , n89391 , n89416 );
not ( n89418 , n88577 );
not ( n89419 , n89313 );
or ( n89420 , n89418 , n89419 );
and ( n89421 , n88054 , n88640 );
not ( n89422 , n88054 );
and ( n89423 , n89422 , n88558 );
or ( n89424 , n89421 , n89423 );
nand ( n89425 , n89424 , n88575 );
nand ( n89426 , n89420 , n89425 );
and ( n89427 , n89417 , n89426 );
and ( n89428 , n89391 , n89416 );
or ( n89429 , n89427 , n89428 );
and ( n89430 , n89379 , n89429 );
and ( n89431 , n89376 , n89378 );
or ( n89432 , n89430 , n89431 );
xor ( n89433 , n89351 , n89432 );
xor ( n89434 , n89308 , n89333 );
xor ( n89435 , n89434 , n89336 );
and ( n89436 , n89433 , n89435 );
and ( n89437 , n89351 , n89432 );
or ( n89438 , n89436 , n89437 );
nor ( n89439 , n89349 , n89438 );
nor ( n89440 , n89347 , n89439 );
not ( n89441 , n89440 );
xor ( n89442 , n89351 , n89432 );
xor ( n89443 , n89442 , n89435 );
xor ( n89444 , n89317 , n89319 );
xor ( n89445 , n89444 , n89330 );
not ( n89446 , n88447 );
not ( n89447 , n89326 );
or ( n89448 , n89446 , n89447 );
not ( n89449 , n89226 );
not ( n89450 , n87953 );
or ( n89451 , n89449 , n89450 );
not ( n89452 , n88451 );
nand ( n89453 , n89452 , n87952 );
nand ( n89454 , n89451 , n89453 );
nand ( n89455 , n89454 , n88445 );
nand ( n89456 , n89448 , n89455 );
xor ( n89457 , n89361 , n89362 );
xor ( n89458 , n89457 , n89373 );
xor ( n89459 , n89456 , n89458 );
nand ( n89460 , n87875 , n2176 );
and ( n89461 , n89460 , n88855 );
not ( n89462 , n2910 );
not ( n89463 , n87830 );
or ( n89464 , n89462 , n89463 );
nand ( n89465 , n89464 , n87707 );
nor ( n89466 , n89461 , n89465 );
not ( n89467 , n87976 );
not ( n89468 , n89400 );
or ( n89469 , n89467 , n89468 );
not ( n89470 , n88014 );
not ( n89471 , n87707 );
not ( n89472 , n88854 );
or ( n89473 , n89471 , n89472 );
nand ( n89474 , n88238 , n88855 );
nand ( n89475 , n89473 , n89474 );
nand ( n89476 , n89470 , n89475 );
nand ( n89477 , n89469 , n89476 );
and ( n89478 , n89466 , n89477 );
not ( n89479 , n89424 );
not ( n89480 , n88577 );
or ( n89481 , n89479 , n89480 );
not ( n89482 , n88582 );
not ( n89483 , n88326 );
or ( n89484 , n89482 , n89483 );
nand ( n89485 , n88159 , n88640 );
nand ( n89486 , n89484 , n89485 );
nand ( n89487 , n89486 , n88575 );
nand ( n89488 , n89481 , n89487 );
xor ( n89489 , n89478 , n89488 );
not ( n89490 , n88036 );
not ( n89491 , n88047 );
not ( n89492 , n88361 );
or ( n89493 , n89491 , n89492 );
nand ( n89494 , n88932 , n89385 );
nand ( n89495 , n89493 , n89494 );
not ( n89496 , n89495 );
or ( n89497 , n89490 , n89496 );
nand ( n89498 , n89387 , n88042 );
nand ( n89499 , n89497 , n89498 );
and ( n89500 , n89489 , n89499 );
and ( n89501 , n89478 , n89488 );
or ( n89502 , n89500 , n89501 );
and ( n89503 , n89459 , n89502 );
and ( n89504 , n89456 , n89458 );
or ( n89505 , n89503 , n89504 );
xor ( n89506 , n89445 , n89505 );
xor ( n89507 , n89376 , n89378 );
xor ( n89508 , n89507 , n89429 );
and ( n89509 , n89506 , n89508 );
and ( n89510 , n89445 , n89505 );
or ( n89511 , n89509 , n89510 );
nor ( n89512 , n89443 , n89511 );
xor ( n89513 , n89445 , n89505 );
xor ( n89514 , n89513 , n89508 );
xor ( n89515 , n89391 , n89416 );
xor ( n89516 , n89515 , n89426 );
xor ( n89517 , n89392 , n89402 );
xor ( n89518 , n89517 , n89413 );
not ( n89519 , n88445 );
not ( n89520 , n88451 );
not ( n89521 , n87935 );
or ( n89522 , n89520 , n89521 );
nand ( n89523 , n87934 , n88490 );
nand ( n89524 , n89522 , n89523 );
not ( n89525 , n89524 );
or ( n89526 , n89519 , n89525 );
nand ( n89527 , n89454 , n88447 );
nand ( n89528 , n89526 , n89527 );
xor ( n89529 , n89518 , n89528 );
not ( n89530 , n88084 );
not ( n89531 , n89411 );
or ( n89532 , n89530 , n89531 );
not ( n89533 , n87830 );
not ( n89534 , n88522 );
or ( n89535 , n89533 , n89534 );
nand ( n89536 , n88521 , n87831 );
nand ( n89537 , n89535 , n89536 );
nand ( n89538 , n89537 , n87870 );
nand ( n89539 , n89532 , n89538 );
xor ( n89540 , n89466 , n89477 );
xor ( n89541 , n89539 , n89540 );
not ( n89542 , n88577 );
not ( n89543 , n89486 );
or ( n89544 , n89542 , n89543 );
not ( n89545 , n88558 );
not ( n89546 , n88375 );
or ( n89547 , n89545 , n89546 );
not ( n89548 , n88582 );
nand ( n89549 , n89548 , n88374 );
nand ( n89550 , n89547 , n89549 );
nand ( n89551 , n89550 , n88575 );
nand ( n89552 , n89544 , n89551 );
and ( n89553 , n89541 , n89552 );
and ( n89554 , n89539 , n89540 );
or ( n89555 , n89553 , n89554 );
and ( n89556 , n89529 , n89555 );
and ( n89557 , n89518 , n89528 );
or ( n89558 , n89556 , n89557 );
xor ( n89559 , n89516 , n89558 );
xor ( n89560 , n89456 , n89458 );
xor ( n89561 , n89560 , n89502 );
and ( n89562 , n89559 , n89561 );
and ( n89563 , n89516 , n89558 );
or ( n89564 , n89562 , n89563 );
nor ( n89565 , n89514 , n89564 );
nor ( n89566 , n89512 , n89565 );
not ( n89567 , n89566 );
xor ( n89568 , n89516 , n89558 );
xor ( n89569 , n89568 , n89561 );
not ( n89570 , n89569 );
xor ( n89571 , n89478 , n89488 );
xor ( n89572 , n89571 , n89499 );
not ( n89573 , n88042 );
not ( n89574 , n89495 );
or ( n89575 , n89573 , n89574 );
not ( n89576 , n88602 );
not ( n89577 , n88457 );
or ( n89578 , n89576 , n89577 );
buf ( n89579 , n88044 );
nand ( n89580 , n88456 , n89579 );
nand ( n89581 , n89578 , n89580 );
nand ( n89582 , n89581 , n88036 );
nand ( n89583 , n89575 , n89582 );
and ( n89584 , n87976 , n88855 );
not ( n89585 , n88084 );
not ( n89586 , n89537 );
or ( n89587 , n89585 , n89586 );
not ( n89588 , n88788 );
and ( n89589 , n87830 , n89588 );
not ( n89590 , n87830 );
and ( n89591 , n89590 , n88789 );
or ( n89592 , n89589 , n89591 );
nand ( n89593 , n89592 , n87870 );
nand ( n89594 , n89587 , n89593 );
xor ( n89595 , n89584 , n89594 );
not ( n89596 , n88041 );
not ( n89597 , n89581 );
or ( n89598 , n89596 , n89597 );
and ( n89599 , n88487 , n88045 );
not ( n89600 , n88487 );
not ( n89601 , n89579 );
and ( n89602 , n89600 , n89601 );
or ( n89603 , n89599 , n89602 );
nand ( n89604 , n89603 , n88036 );
nand ( n89605 , n89598 , n89604 );
and ( n89606 , n89595 , n89605 );
and ( n89607 , n89584 , n89594 );
or ( n89608 , n89606 , n89607 );
xor ( n89609 , n89583 , n89608 );
not ( n89610 , n88447 );
not ( n89611 , n89524 );
or ( n89612 , n89610 , n89611 );
not ( n89613 , n88451 );
not ( n89614 , n88333 );
or ( n89615 , n89613 , n89614 );
not ( n89616 , n89226 );
nand ( n89617 , n89616 , n88054 );
nand ( n89618 , n89615 , n89617 );
nand ( n89619 , n89618 , n88445 );
nand ( n89620 , n89612 , n89619 );
and ( n89621 , n89609 , n89620 );
and ( n89622 , n89583 , n89608 );
or ( n89623 , n89621 , n89622 );
xor ( n89624 , n89572 , n89623 );
xor ( n89625 , n89518 , n89528 );
xor ( n89626 , n89625 , n89555 );
and ( n89627 , n89624 , n89626 );
and ( n89628 , n89572 , n89623 );
or ( n89629 , n89627 , n89628 );
not ( n89630 , n89629 );
and ( n89631 , n89570 , n89630 );
xor ( n89632 , n89572 , n89623 );
xor ( n89633 , n89632 , n89626 );
nand ( n89634 , n89579 , n87867 );
and ( n89635 , n89634 , n88855 );
not ( n89636 , n87860 );
not ( n89637 , n88044 );
not ( n89638 , n89637 );
or ( n89639 , n89636 , n89638 );
nand ( n89640 , n89639 , n87830 );
nor ( n89641 , n89635 , n89640 );
not ( n89642 , n87869 );
not ( n89643 , n89592 );
or ( n89644 , n89642 , n89643 );
nor ( n89645 , n87861 , n87869 );
not ( n89646 , n88855 );
not ( n89647 , n87875 );
or ( n89648 , n89646 , n89647 );
nand ( n89649 , n88854 , n87830 );
nand ( n89650 , n89648 , n89649 );
nand ( n89651 , n89645 , n89650 );
nand ( n89652 , n89644 , n89651 );
and ( n89653 , n89641 , n89652 );
not ( n89654 , n88575 );
and ( n89655 , n88582 , n88361 );
not ( n89656 , n88582 );
and ( n89657 , n89656 , n88360 );
or ( n89658 , n89655 , n89657 );
not ( n89659 , n89658 );
or ( n89660 , n89654 , n89659 );
nand ( n89661 , n89550 , n88577 );
nand ( n89662 , n89660 , n89661 );
xor ( n89663 , n89653 , n89662 );
not ( n89664 , n88447 );
not ( n89665 , n89618 );
or ( n89666 , n89664 , n89665 );
not ( n89667 , n88451 );
not ( n89668 , n88326 );
or ( n89669 , n89667 , n89668 );
not ( n89670 , n89226 );
nand ( n89671 , n89670 , n88159 );
nand ( n89672 , n89669 , n89671 );
nand ( n89673 , n89672 , n88445 );
nand ( n89674 , n89666 , n89673 );
and ( n89675 , n89663 , n89674 );
and ( n89676 , n89653 , n89662 );
or ( n89677 , n89675 , n89676 );
xor ( n89678 , n89539 , n89540 );
xor ( n89679 , n89678 , n89552 );
xor ( n89680 , n89677 , n89679 );
xor ( n89681 , n89583 , n89608 );
xor ( n89682 , n89681 , n89620 );
and ( n89683 , n89680 , n89682 );
and ( n89684 , n89677 , n89679 );
or ( n89685 , n89683 , n89684 );
nor ( n89686 , n89633 , n89685 );
nor ( n89687 , n89631 , n89686 );
not ( n89688 , n89687 );
xor ( n89689 , n89584 , n89594 );
xor ( n89690 , n89689 , n89605 );
not ( n89691 , n88041 );
not ( n89692 , n89603 );
or ( n89693 , n89691 , n89692 );
not ( n89694 , n88045 );
not ( n89695 , n89694 );
not ( n89696 , n88773 );
or ( n89697 , n89695 , n89696 );
nand ( n89698 , n88521 , n89579 );
nand ( n89699 , n89697 , n89698 );
nand ( n89700 , n89699 , n88035 );
nand ( n89701 , n89693 , n89700 );
xor ( n89702 , n89641 , n89652 );
xor ( n89703 , n89701 , n89702 );
not ( n89704 , n88577 );
not ( n89705 , n89658 );
or ( n89706 , n89704 , n89705 );
not ( n89707 , n88582 );
not ( n89708 , n88457 );
or ( n89709 , n89707 , n89708 );
nand ( n89710 , n88456 , n88750 );
nand ( n89711 , n89709 , n89710 );
nand ( n89712 , n89711 , n88575 );
nand ( n89713 , n89706 , n89712 );
and ( n89714 , n89703 , n89713 );
and ( n89715 , n89701 , n89702 );
or ( n89716 , n89714 , n89715 );
xor ( n89717 , n89690 , n89716 );
xor ( n89718 , n89653 , n89662 );
xor ( n89719 , n89718 , n89674 );
and ( n89720 , n89717 , n89719 );
and ( n89721 , n89690 , n89716 );
or ( n89722 , n89720 , n89721 );
not ( n89723 , n89722 );
xor ( n89724 , n89677 , n89679 );
xor ( n89725 , n89724 , n89682 );
not ( n89726 , n89725 );
nand ( n89727 , n89723 , n89726 );
not ( n89728 , n89727 );
xor ( n89729 , n89690 , n89716 );
xor ( n89730 , n89729 , n89719 );
not ( n89731 , n89730 );
not ( n89732 , n88447 );
not ( n89733 , n89672 );
or ( n89734 , n89732 , n89733 );
xor ( n89735 , n89226 , n88374 );
nand ( n89736 , n89735 , n88445 );
nand ( n89737 , n89734 , n89736 );
nor ( n89738 , n87874 , n88854 );
not ( n89739 , n88041 );
not ( n89740 , n89699 );
or ( n89741 , n89739 , n89740 );
not ( n89742 , n88044 );
not ( n89743 , n89742 );
not ( n89744 , n89588 );
or ( n89745 , n89743 , n89744 );
nand ( n89746 , n88788 , n88044 );
nand ( n89747 , n89745 , n89746 );
nand ( n89748 , n88035 , n89747 );
nand ( n89749 , n89741 , n89748 );
xor ( n89750 , n89738 , n89749 );
not ( n89751 , n1971 );
nand ( n89752 , n89751 , n88557 );
and ( n89753 , n89752 , n88867 );
not ( n89754 , n1971 );
not ( n89755 , n88582 );
or ( n89756 , n89754 , n89755 );
nand ( n89757 , n89756 , n89637 );
nor ( n89758 , n89753 , n89757 );
not ( n89759 , n88041 );
not ( n89760 , n89747 );
or ( n89761 , n89759 , n89760 );
not ( n89762 , n88034 );
not ( n89763 , n88855 );
not ( n89764 , n88044 );
or ( n89765 , n89763 , n89764 );
not ( n89766 , n88867 );
not ( n89767 , n88044 );
nand ( n89768 , n89766 , n89767 );
nand ( n89769 , n89765 , n89768 );
nand ( n89770 , n89762 , n89769 );
nand ( n89771 , n89761 , n89770 );
and ( n89772 , n89758 , n89771 );
and ( n89773 , n89750 , n89772 );
and ( n89774 , n89738 , n89749 );
or ( n89775 , n89773 , n89774 );
xor ( n89776 , n89737 , n89775 );
xor ( n89777 , n89701 , n89702 );
xor ( n89778 , n89777 , n89713 );
and ( n89779 , n89776 , n89778 );
and ( n89780 , n89737 , n89775 );
or ( n89781 , n89779 , n89780 );
not ( n89782 , n89781 );
nand ( n89783 , n89731 , n89782 );
not ( n89784 , n89783 );
nor ( n89785 , n88028 , n88854 );
not ( n89786 , n88577 );
and ( n89787 , n88521 , n88024 );
not ( n89788 , n88521 );
and ( n89789 , n89788 , n88025 );
nor ( n89790 , n89787 , n89789 );
not ( n89791 , n89790 );
or ( n89792 , n89786 , n89791 );
not ( n89793 , n88024 );
not ( n89794 , n89588 );
or ( n89795 , n89793 , n89794 );
nand ( n89796 , n88788 , n88025 );
nand ( n89797 , n89795 , n89796 );
nand ( n89798 , n89797 , n88575 );
nand ( n89799 , n89792 , n89798 );
xor ( n89800 , n89785 , n89799 );
not ( n89801 , n88574 );
and ( n89802 , n88853 , n88025 );
not ( n89803 , n88853 );
and ( n89804 , n89803 , n88582 );
nor ( n89805 , n89802 , n89804 );
not ( n89806 , n89805 );
and ( n89807 , n89801 , n89806 );
and ( n89808 , n88577 , n89797 );
nor ( n89809 , n89807 , n89808 );
not ( n89810 , n88566 );
and ( n89811 , n88450 , n89810 );
nor ( n89812 , n89811 , n88025 );
or ( n89813 , n89226 , n89810 );
nand ( n89814 , n89813 , n88867 );
nand ( n89815 , n89812 , n89814 );
nor ( n89816 , n89809 , n89815 );
xor ( n89817 , n89800 , n89816 );
not ( n89818 , n88447 );
not ( n89819 , n89226 );
not ( n89820 , n88457 );
or ( n89821 , n89819 , n89820 );
nand ( n89822 , n88456 , n88449 );
nand ( n89823 , n89821 , n89822 );
not ( n89824 , n89823 );
or ( n89825 , n89818 , n89824 );
not ( n89826 , n88449 );
not ( n89827 , n88487 );
not ( n89828 , n89827 );
or ( n89829 , n89826 , n89828 );
or ( n89830 , n89827 , n88449 );
nand ( n89831 , n89829 , n89830 );
not ( n89832 , n89831 );
nand ( n89833 , n89832 , n88445 );
nand ( n89834 , n89825 , n89833 );
or ( n89835 , n89817 , n89834 );
and ( n89836 , n88521 , n88450 );
not ( n89837 , n88521 );
and ( n89838 , n89837 , n88449 );
nor ( n89839 , n89836 , n89838 );
not ( n89840 , n89839 );
not ( n89841 , n88445 );
or ( n89842 , n89840 , n89841 );
or ( n89843 , n89831 , n88836 );
nand ( n89844 , n89842 , n89843 );
xor ( n89845 , n89815 , n89809 );
xor ( n89846 , n89844 , n89845 );
nor ( n89847 , n88573 , n88854 );
not ( n89848 , n88447 );
not ( n89849 , n89839 );
or ( n89850 , n89848 , n89849 );
not ( n89851 , n88450 );
not ( n89852 , n89588 );
or ( n89853 , n89851 , n89852 );
nand ( n89854 , n88788 , n88449 );
nand ( n89855 , n89853 , n89854 );
nand ( n89856 , n89855 , n88445 );
nand ( n89857 , n89850 , n89856 );
xor ( n89858 , n89847 , n89857 );
and ( n89859 , n89855 , n88447 );
nand ( n89860 , n89226 , n88854 );
nand ( n89861 , n88449 , n88867 );
and ( n89862 , n89860 , n89861 );
nor ( n89863 , n89862 , n88444 );
nor ( n89864 , n89859 , n89863 );
nand ( n89865 , n88855 , n88447 );
nand ( n89866 , n89865 , n88450 );
nor ( n89867 , n89864 , n89866 );
and ( n89868 , n89858 , n89867 );
and ( n89869 , n89847 , n89857 );
or ( n89870 , n89868 , n89869 );
and ( n89871 , n89846 , n89870 );
and ( n89872 , n89844 , n89845 );
or ( n89873 , n89871 , n89872 );
and ( n89874 , n89835 , n89873 );
nand ( n89875 , n89817 , n89834 );
not ( n89876 , n89875 );
nor ( n89877 , n89874 , n89876 );
not ( n89878 , n88577 );
not ( n89879 , n88582 );
not ( n89880 , n89279 );
or ( n89881 , n89879 , n89880 );
not ( n89882 , n88024 );
nand ( n89883 , n89882 , n88487 );
nand ( n89884 , n89881 , n89883 );
not ( n89885 , n89884 );
or ( n89886 , n89878 , n89885 );
nand ( n89887 , n89790 , n88575 );
nand ( n89888 , n89886 , n89887 );
xor ( n89889 , n89758 , n89771 );
xor ( n89890 , n89888 , n89889 );
not ( n89891 , n88447 );
not ( n89892 , n88361 );
xor ( n89893 , n88450 , n89892 );
not ( n89894 , n89893 );
or ( n89895 , n89891 , n89894 );
nand ( n89896 , n89823 , n88445 );
nand ( n89897 , n89895 , n89896 );
xor ( n89898 , n89890 , n89897 );
xor ( n89899 , n89785 , n89799 );
and ( n89900 , n89899 , n89816 );
and ( n89901 , n89785 , n89799 );
or ( n89902 , n89900 , n89901 );
nor ( n89903 , n89898 , n89902 );
or ( n89904 , n89877 , n89903 );
nand ( n89905 , n89898 , n89902 );
nand ( n89906 , n89904 , n89905 );
not ( n89907 , n88577 );
not ( n89908 , n89711 );
or ( n89909 , n89907 , n89908 );
nand ( n89910 , n89884 , n88575 );
nand ( n89911 , n89909 , n89910 );
not ( n89912 , n88445 );
not ( n89913 , n89893 );
or ( n89914 , n89912 , n89913 );
nand ( n89915 , n89735 , n88447 );
nand ( n89916 , n89914 , n89915 );
xor ( n89917 , n89911 , n89916 );
xor ( n89918 , n89738 , n89749 );
xor ( n89919 , n89918 , n89772 );
xor ( n89920 , n89917 , n89919 );
not ( n89921 , n89920 );
xor ( n89922 , n89888 , n89889 );
and ( n89923 , n89922 , n89897 );
and ( n89924 , n89888 , n89889 );
or ( n89925 , n89923 , n89924 );
not ( n89926 , n89925 );
nand ( n89927 , n89921 , n89926 );
and ( n89928 , n89906 , n89927 );
and ( n89929 , n89920 , n89925 );
nor ( n89930 , n89928 , n89929 );
xor ( n89931 , n89737 , n89775 );
xor ( n89932 , n89931 , n89778 );
xor ( n89933 , n89911 , n89916 );
and ( n89934 , n89933 , n89919 );
and ( n89935 , n89911 , n89916 );
or ( n89936 , n89934 , n89935 );
nor ( n89937 , n89932 , n89936 );
or ( n89938 , n89930 , n89937 );
nand ( n89939 , n89932 , n89936 );
nand ( n89940 , n89938 , n89939 );
not ( n89941 , n89940 );
or ( n89942 , n89784 , n89941 );
nand ( n89943 , n89730 , n89781 );
nand ( n89944 , n89942 , n89943 );
not ( n89945 , n89944 );
or ( n89946 , n89728 , n89945 );
not ( n89947 , n89726 );
nand ( n89948 , n89947 , n89722 );
nand ( n89949 , n89946 , n89948 );
not ( n89950 , n89949 );
or ( n89951 , n89688 , n89950 );
not ( n89952 , n89569 );
not ( n89953 , n89629 );
nand ( n89954 , n89952 , n89953 );
and ( n89955 , n89633 , n89685 );
and ( n89956 , n89954 , n89955 );
nor ( n89957 , n89952 , n89953 );
nor ( n89958 , n89956 , n89957 );
nand ( n89959 , n89951 , n89958 );
not ( n89960 , n89959 );
or ( n89961 , n89567 , n89960 );
nor ( n89962 , n89443 , n89511 );
not ( n89963 , n89962 );
nand ( n89964 , n89514 , n89564 );
not ( n89965 , n89964 );
and ( n89966 , n89963 , n89965 );
and ( n89967 , n89443 , n89511 );
nor ( n89968 , n89966 , n89967 );
nand ( n89969 , n89961 , n89968 );
not ( n89970 , n89969 );
or ( n89971 , n89441 , n89970 );
not ( n89972 , n89271 );
not ( n89973 , n89345 );
nand ( n89974 , n89972 , n89973 );
not ( n89975 , n89349 );
not ( n89976 , n89438 );
nor ( n89977 , n89975 , n89976 );
and ( n89978 , n89974 , n89977 );
and ( n89979 , n89271 , n89345 );
nor ( n89980 , n89978 , n89979 );
nand ( n89981 , n89971 , n89980 );
not ( n89982 , n89981 );
or ( n89983 , n89269 , n89982 );
not ( n89984 , n89267 );
nand ( n89985 , n89121 , n89258 );
not ( n89986 , n89985 );
and ( n89987 , n89984 , n89986 );
and ( n89988 , n89262 , n89266 );
nor ( n89989 , n89987 , n89988 );
nand ( n89990 , n89983 , n89989 );
not ( n89991 , n89990 );
or ( n89992 , n89105 , n89991 );
not ( n89993 , n89103 );
nand ( n89994 , n88991 , n88993 );
or ( n89995 , n88911 , n89994 );
nand ( n89996 , n88741 , n88910 );
nand ( n89997 , n89995 , n89996 );
not ( n89998 , n89997 );
or ( n89999 , n89993 , n89998 );
not ( n90000 , n89097 );
nand ( n90001 , n90000 , n89101 );
nand ( n90002 , n89999 , n90001 );
not ( n90003 , n89061 );
nand ( n90004 , n89093 , n90003 );
and ( n90005 , n90002 , n90004 );
nor ( n90006 , n89093 , n90003 );
nor ( n90007 , n90005 , n90006 );
nand ( n90008 , n89992 , n90007 );
not ( n90009 , n90008 );
xor ( n90010 , n89074 , n89086 );
and ( n90011 , n90010 , n89091 );
and ( n90012 , n89074 , n89086 );
or ( n90013 , n90011 , n90012 );
xor ( n90014 , n89066 , n89070 );
and ( n90015 , n90014 , n89073 );
and ( n90016 , n89066 , n89070 );
or ( n90017 , n90015 , n90016 );
xor ( n90018 , n88212 , n88214 );
xor ( n90019 , n90018 , n88217 );
xor ( n90020 , n90017 , n90019 );
xor ( n90021 , n89076 , n89080 );
and ( n90022 , n90021 , n89085 );
and ( n90023 , n89076 , n89080 );
or ( n90024 , n90022 , n90023 );
xor ( n90025 , n90020 , n90024 );
or ( n90026 , n90013 , n90025 );
xor ( n90027 , n88022 , n17814 );
xor ( n90028 , n90027 , n88220 );
xor ( n90029 , n90017 , n90019 );
and ( n90030 , n90029 , n90024 );
and ( n90031 , n90017 , n90019 );
or ( n90032 , n90030 , n90031 );
nor ( n90033 , n90028 , n90032 );
not ( n90034 , n90033 );
nand ( n90035 , n90026 , n90034 );
not ( n90036 , n90035 );
not ( n90037 , n90036 );
or ( n90038 , n90009 , n90037 );
nand ( n90039 , n90013 , n90025 );
not ( n90040 , n90039 );
not ( n90041 , n90033 );
and ( n90042 , n90040 , n90041 );
and ( n90043 , n90028 , n90032 );
nor ( n90044 , n90042 , n90043 );
nand ( n90045 , n90038 , n90044 );
not ( n90046 , n90045 );
or ( n90047 , n88323 , n90046 );
nand ( n90048 , n88223 , n88275 );
or ( n90049 , n88321 , n90048 );
nand ( n90050 , n88281 , n88320 );
nand ( n90051 , n90049 , n90050 );
not ( n90052 , n90051 );
nand ( n90053 , n90047 , n90052 );
or ( n90054 , n88015 , n87977 );
nand ( n90055 , n90054 , n87979 );
not ( n90056 , n87826 );
or ( n90057 , n88115 , n87799 );
or ( n90058 , n87857 , n87718 );
nand ( n90059 , n90057 , n90058 );
not ( n90060 , n90059 );
or ( n90061 , n90056 , n90060 );
nand ( n90062 , n88290 , n87716 );
nand ( n90063 , n90061 , n90062 );
xor ( n90064 , n90055 , n90063 );
and ( n90065 , n87922 , n87795 );
xor ( n90066 , n90064 , n90065 );
not ( n90067 , n87919 );
not ( n90068 , n88297 );
or ( n90069 , n90067 , n90068 );
and ( n90070 , n87921 , n87995 );
not ( n90071 , n87921 );
and ( n90072 , n90071 , n87998 );
nor ( n90073 , n90070 , n90072 );
or ( n90074 , n90073 , n87966 );
nand ( n90075 , n90069 , n90074 );
xor ( n90076 , n90075 , n88303 );
xor ( n90077 , n88282 , n88292 );
and ( n90078 , n90077 , n88299 );
and ( n90079 , n88282 , n88292 );
or ( n90080 , n90078 , n90079 );
xor ( n90081 , n90076 , n90080 );
xor ( n90082 , n90066 , n90081 );
xor ( n90083 , n88304 , n88308 );
and ( n90084 , n90083 , n88313 );
and ( n90085 , n88304 , n88308 );
or ( n90086 , n90084 , n90085 );
xor ( n90087 , n90082 , n90086 );
xor ( n90088 , n88300 , n88314 );
and ( n90089 , n90088 , n88319 );
and ( n90090 , n88300 , n88314 );
or ( n90091 , n90089 , n90090 );
or ( n90092 , n90087 , n90091 );
nand ( n90093 , n90091 , n90087 );
nand ( n90094 , n90092 , n90093 );
not ( n90095 , n90094 );
and ( n90096 , n90053 , n90095 );
not ( n90097 , n90053 );
and ( n90098 , n90097 , n90094 );
nor ( n90099 , n90096 , n90098 );
and ( n90100 , n87706 , n90099 );
not ( n90101 , n87706 );
not ( n90102 , n90099 );
and ( n90103 , n90101 , n90102 );
nor ( n90104 , n90100 , n90103 );
not ( n90105 , n90104 );
or ( n90106 , n87703 , n90105 );
and ( n90107 , n88322 , n90092 );
not ( n90108 , n90107 );
not ( n90109 , n90045 );
or ( n90110 , n90108 , n90109 );
and ( n90111 , n90051 , n90092 );
not ( n90112 , n90093 );
nor ( n90113 , n90111 , n90112 );
nand ( n90114 , n90110 , n90113 );
xor ( n90115 , n90066 , n90081 );
and ( n90116 , n90115 , n90086 );
and ( n90117 , n90066 , n90081 );
or ( n90118 , n90116 , n90117 );
xor ( n90119 , n90055 , n90063 );
and ( n90120 , n90119 , n90065 );
and ( n90121 , n90055 , n90063 );
or ( n90122 , n90120 , n90121 );
or ( n90123 , n90073 , n87918 );
not ( n90124 , n88079 );
not ( n90125 , n87921 );
and ( n90126 , n90124 , n90125 );
and ( n90127 , n88079 , n87921 );
nor ( n90128 , n90126 , n90127 );
or ( n90129 , n90128 , n87966 );
nand ( n90130 , n90123 , n90129 );
and ( n90131 , n87922 , n87822 );
xor ( n90132 , n90130 , n90131 );
and ( n90133 , n90059 , n87716 );
and ( n90134 , n87826 , n87718 );
nor ( n90135 , n90133 , n90134 );
xor ( n90136 , n90132 , n90135 );
xor ( n90137 , n90122 , n90136 );
xor ( n90138 , n90075 , n88303 );
and ( n90139 , n90138 , n90080 );
and ( n90140 , n90075 , n88303 );
or ( n90141 , n90139 , n90140 );
xor ( n90142 , n90137 , n90141 );
or ( n90143 , n90118 , n90142 );
nand ( n90144 , n90118 , n90142 );
nand ( n90145 , n90143 , n90144 );
and ( n90146 , n90114 , n90145 );
not ( n90147 , n90114 );
not ( n90148 , n90145 );
and ( n90149 , n90147 , n90148 );
nor ( n90150 , n90146 , n90149 );
not ( n90151 , n90150 );
and ( n90152 , n87706 , n90151 );
not ( n90153 , n87706 );
not ( n90154 , n90151 );
and ( n90155 , n90153 , n90154 );
nor ( n90156 , n90152 , n90155 );
nand ( n90157 , n90156 , n87689 );
nand ( n90158 , n90106 , n90157 );
nor ( n90159 , n524 , n540 );
not ( n90160 , n90159 );
nand ( n90161 , n524 , n540 );
and ( n90162 , n90160 , n90161 );
nand ( n90163 , n536 , n552 );
not ( n90164 , n90163 );
not ( n90165 , n87692 );
or ( n90166 , n90164 , n90165 );
nor ( n90167 , n534 , n550 );
nor ( n90168 , n87694 , n90167 );
nand ( n90169 , n90166 , n90168 );
nand ( n90170 , n533 , n549 );
nand ( n90171 , n534 , n550 );
nand ( n90172 , n90169 , n90170 , n90171 );
not ( n90173 , n90172 );
nor ( n90174 , n529 , n545 );
nor ( n90175 , n533 , n549 );
nor ( n90176 , n530 , n546 );
nor ( n90177 , n90174 , n90175 , n90176 );
nor ( n90178 , n531 , n547 );
nor ( n90179 , n532 , n548 );
nor ( n90180 , n90178 , n90179 );
and ( n90181 , n90177 , n90180 );
not ( n90182 , n90181 );
or ( n90183 , n90173 , n90182 );
nand ( n90184 , n530 , n546 );
nand ( n90185 , n529 , n545 );
nand ( n90186 , n531 , n547 );
and ( n90187 , n90184 , n90185 , n90186 );
not ( n90188 , n90187 );
not ( n90189 , n90178 );
nand ( n90190 , n532 , n548 );
not ( n90191 , n90190 );
nand ( n90192 , n90189 , n90191 );
not ( n90193 , n90192 );
or ( n90194 , n90188 , n90193 );
not ( n90195 , n90176 );
not ( n90196 , n90195 );
not ( n90197 , n90174 );
not ( n90198 , n90197 );
or ( n90199 , n90196 , n90198 );
nand ( n90200 , n90199 , n90185 );
nand ( n90201 , n90194 , n90200 );
nand ( n90202 , n90183 , n90201 );
not ( n90203 , n90202 );
nor ( n90204 , n525 , n541 );
nor ( n90205 , n526 , n542 );
nor ( n90206 , n90204 , n90205 );
nor ( n90207 , n527 , n543 );
nor ( n90208 , n528 , n544 );
nor ( n90209 , n90207 , n90208 );
nand ( n90210 , n90206 , n90209 );
not ( n90211 , n90210 );
not ( n90212 , n90211 );
or ( n90213 , n90203 , n90212 );
nand ( n90214 , n528 , n544 );
or ( n90215 , n90207 , n90214 );
nand ( n90216 , n527 , n543 );
nand ( n90217 , n90215 , n90216 );
not ( n90218 , n90217 );
not ( n90219 , n90206 );
or ( n90220 , n90218 , n90219 );
not ( n90221 , n90204 );
nand ( n90222 , n526 , n542 );
not ( n90223 , n90222 );
and ( n90224 , n90221 , n90223 );
and ( n90225 , n525 , n541 );
nor ( n90226 , n90224 , n90225 );
nand ( n90227 , n90220 , n90226 );
not ( n90228 , n90227 );
nand ( n90229 , n90213 , n90228 );
xor ( n90230 , n90162 , n90229 );
not ( n90231 , n90230 );
not ( n90232 , n90231 );
nor ( n90233 , n90204 , n90225 );
not ( n90234 , n90205 );
and ( n90235 , n90209 , n90234 );
not ( n90236 , n90235 );
not ( n90237 , n90202 );
or ( n90238 , n90236 , n90237 );
and ( n90239 , n90217 , n90234 );
not ( n90240 , n90222 );
nor ( n90241 , n90239 , n90240 );
nand ( n90242 , n90238 , n90241 );
xor ( n90243 , n90233 , n90242 );
not ( n90244 , n90243 );
or ( n90245 , n90232 , n90244 );
not ( n90246 , n90243 );
nand ( n90247 , n90246 , n90230 );
nand ( n90248 , n90245 , n90247 );
not ( n90249 , n90248 );
not ( n90250 , n90231 );
nor ( n90251 , n90210 , n90159 );
not ( n90252 , n90251 );
not ( n90253 , n90172 );
not ( n90254 , n90181 );
or ( n90255 , n90253 , n90254 );
nand ( n90256 , n90255 , n90201 );
not ( n90257 , n90256 );
or ( n90258 , n90252 , n90257 );
not ( n90259 , n90160 );
not ( n90260 , n90227 );
or ( n90261 , n90259 , n90260 );
nand ( n90262 , n90261 , n90161 );
not ( n90263 , n90262 );
nand ( n90264 , n90258 , n90263 );
nor ( n90265 , n523 , n539 );
not ( n90266 , n90265 );
nand ( n90267 , n523 , n539 );
nand ( n90268 , n90266 , n90267 );
not ( n90269 , n90268 );
and ( n90270 , n90264 , n90269 );
not ( n90271 , n90264 );
and ( n90272 , n90271 , n90268 );
nor ( n90273 , n90270 , n90272 );
not ( n90274 , n90273 );
or ( n90275 , n90250 , n90274 );
or ( n90276 , n90273 , n90231 );
nand ( n90277 , n90275 , n90276 );
nand ( n90278 , n90249 , n90277 );
not ( n90279 , n90278 );
not ( n90280 , n90279 );
not ( n90281 , n90269 );
not ( n90282 , n90264 );
not ( n90283 , n90282 );
or ( n90284 , n90281 , n90283 );
nand ( n90285 , n90264 , n90268 );
nand ( n90286 , n90284 , n90285 );
not ( n90287 , n89565 );
and ( n90288 , n89959 , n90287 );
not ( n90289 , n89964 );
nor ( n90290 , n90288 , n90289 );
xor ( n90291 , n89443 , n89511 );
and ( n90292 , n90290 , n90291 );
not ( n90293 , n90290 );
or ( n90294 , n89512 , n89967 );
and ( n90295 , n90293 , n90294 );
nor ( n90296 , n90292 , n90295 );
not ( n90297 , n90296 );
and ( n90298 , n90286 , n90297 );
not ( n90299 , n90286 );
not ( n90300 , n90297 );
and ( n90301 , n90299 , n90300 );
nor ( n90302 , n90298 , n90301 );
not ( n90303 , n90302 );
or ( n90304 , n90280 , n90303 );
buf ( n90305 , n90286 );
not ( n90306 , n90305 );
nand ( n90307 , n89349 , n89438 );
not ( n90308 , n89349 );
nand ( n90309 , n90308 , n89976 );
nand ( n90310 , n90307 , n90309 );
not ( n90311 , n90310 );
not ( n90312 , n90311 );
not ( n90313 , n89969 );
not ( n90314 , n90313 );
or ( n90315 , n90312 , n90314 );
nand ( n90316 , n89969 , n90310 );
nand ( n90317 , n90315 , n90316 );
not ( n90318 , n90317 );
not ( n90319 , n90318 );
or ( n90320 , n90306 , n90319 );
not ( n90321 , n90286 );
nand ( n90322 , n90317 , n90321 );
nand ( n90323 , n90320 , n90322 );
buf ( n90324 , n90248 );
nand ( n90325 , n90323 , n90324 );
nand ( n90326 , n90304 , n90325 );
nor ( n90327 , n90265 , n90159 );
nor ( n90328 , n522 , n538 );
nor ( n90329 , n521 , n537 );
nor ( n90330 , n90328 , n90329 );
and ( n90331 , n90327 , n90330 );
not ( n90332 , n90331 );
nor ( n90333 , n90332 , n90210 );
not ( n90334 , n90333 );
not ( n90335 , n90256 );
or ( n90336 , n90334 , n90335 );
and ( n90337 , n90331 , n90227 );
not ( n90338 , n90330 );
not ( n90339 , n90161 );
not ( n90340 , n90339 );
not ( n90341 , n90266 );
or ( n90342 , n90340 , n90341 );
nand ( n90343 , n90342 , n90267 );
not ( n90344 , n90343 );
or ( n90345 , n90338 , n90344 );
nand ( n90346 , n522 , n538 );
nor ( n90347 , n90346 , n90329 );
and ( n90348 , n521 , n537 );
nor ( n90349 , n90347 , n90348 );
nand ( n90350 , n90345 , n90349 );
nor ( n90351 , n90337 , n90350 );
nand ( n90352 , n90336 , n90351 );
nor ( n90353 , n90348 , n90329 );
not ( n90354 , n90328 );
and ( n90355 , n90327 , n90354 );
not ( n90356 , n90355 );
nor ( n90357 , n90356 , n90210 );
not ( n90358 , n90357 );
not ( n90359 , n90202 );
or ( n90360 , n90358 , n90359 );
and ( n90361 , n90355 , n90227 );
not ( n90362 , n90354 );
not ( n90363 , n90343 );
or ( n90364 , n90362 , n90363 );
nand ( n90365 , n90364 , n90346 );
nor ( n90366 , n90361 , n90365 );
nand ( n90367 , n90360 , n90366 );
xor ( n90368 , n90353 , n90367 );
xnor ( n90369 , n90352 , n90368 );
not ( n90370 , n90369 );
not ( n90371 , n90370 );
buf ( n90372 , n89944 );
xor ( n90373 , n89722 , n89725 );
not ( n90374 , n90373 );
and ( n90375 , n90372 , n90374 );
not ( n90376 , n90372 );
and ( n90377 , n90376 , n90373 );
nor ( n90378 , n90375 , n90377 );
buf ( n90379 , n90378 );
not ( n90380 , n90379 );
not ( n90381 , n90380 );
or ( n90382 , n90371 , n90381 );
and ( n90383 , n89943 , n89783 );
buf ( n90384 , n89940 );
xor ( n90385 , n90383 , n90384 );
not ( n90386 , n90385 );
nand ( n90387 , n90369 , n90352 );
or ( n90388 , n90386 , n90387 );
nand ( n90389 , n90382 , n90388 );
not ( n90390 , n90286 );
not ( n90391 , n90327 );
nor ( n90392 , n90391 , n90210 );
not ( n90393 , n90392 );
not ( n90394 , n90256 );
or ( n90395 , n90393 , n90394 );
and ( n90396 , n90327 , n90227 );
nor ( n90397 , n90396 , n90343 );
nand ( n90398 , n90395 , n90397 );
nand ( n90399 , n90354 , n90346 );
xnor ( n90400 , n90398 , n90399 );
not ( n90401 , n90400 );
or ( n90402 , n90390 , n90401 );
or ( n90403 , n90273 , n90400 );
nand ( n90404 , n90402 , n90403 );
not ( n90405 , n90404 );
not ( n90406 , n90405 );
buf ( n90407 , n90368 );
not ( n90408 , n90407 );
not ( n90409 , n89954 );
nor ( n90410 , n90409 , n89957 );
or ( n90411 , n89633 , n89685 );
not ( n90412 , n90411 );
not ( n90413 , n89949 );
or ( n90414 , n90412 , n90413 );
not ( n90415 , n89955 );
nand ( n90416 , n90414 , n90415 );
xor ( n90417 , n90410 , n90416 );
buf ( n90418 , n90417 );
not ( n90419 , n90418 );
not ( n90420 , n90419 );
or ( n90421 , n90408 , n90420 );
not ( n90422 , n90407 );
nand ( n90423 , n90418 , n90422 );
nand ( n90424 , n90421 , n90423 );
not ( n90425 , n90424 );
or ( n90426 , n90406 , n90425 );
nand ( n90427 , n90415 , n90411 );
xnor ( n90428 , n89949 , n90427 );
not ( n90429 , n90428 );
not ( n90430 , n90429 );
and ( n90431 , n90407 , n90430 );
not ( n90432 , n90407 );
and ( n90433 , n90432 , n90429 );
nor ( n90434 , n90431 , n90433 );
and ( n90435 , n90400 , n90368 );
not ( n90436 , n90400 );
not ( n90437 , n90368 );
and ( n90438 , n90436 , n90437 );
nor ( n90439 , n90435 , n90438 );
and ( n90440 , n90439 , n90404 );
not ( n90441 , n90440 );
not ( n90442 , n90441 );
nand ( n90443 , n90434 , n90442 );
nand ( n90444 , n90426 , n90443 );
and ( n90445 , n90389 , n90444 );
xor ( n90446 , n90326 , n90445 );
not ( n90447 , n90370 );
not ( n90448 , n90430 );
or ( n90449 , n90447 , n90448 );
or ( n90450 , n90379 , n90387 );
nand ( n90451 , n90449 , n90450 );
not ( n90452 , n90442 );
not ( n90453 , n90424 );
or ( n90454 , n90452 , n90453 );
not ( n90455 , n90407 );
nand ( n90456 , n90287 , n89964 );
not ( n90457 , n90456 );
buf ( n90458 , n89959 );
not ( n90459 , n90458 );
not ( n90460 , n90459 );
or ( n90461 , n90457 , n90460 );
not ( n90462 , n90456 );
nand ( n90463 , n90462 , n90458 );
nand ( n90464 , n90461 , n90463 );
not ( n90465 , n90464 );
or ( n90466 , n90455 , n90465 );
not ( n90467 , n90456 );
not ( n90468 , n90459 );
or ( n90469 , n90467 , n90468 );
nand ( n90470 , n90469 , n90463 );
not ( n90471 , n90470 );
nand ( n90472 , n90471 , n90422 );
nand ( n90473 , n90466 , n90472 );
nand ( n90474 , n90473 , n90405 );
nand ( n90475 , n90454 , n90474 );
xor ( n90476 , n90451 , n90475 );
xor ( n90477 , n90446 , n90476 );
not ( n90478 , n90180 );
nor ( n90479 , n90478 , n90176 );
not ( n90480 , n90479 );
nor ( n90481 , n90167 , n90175 );
not ( n90482 , n90481 );
or ( n90483 , n87694 , n90163 );
nand ( n90484 , n90483 , n87692 );
not ( n90485 , n90484 );
or ( n90486 , n90482 , n90485 );
nor ( n90487 , n533 , n549 );
or ( n90488 , n90487 , n90171 );
nand ( n90489 , n90488 , n90170 );
not ( n90490 , n90489 );
nand ( n90491 , n90486 , n90490 );
not ( n90492 , n90491 );
or ( n90493 , n90480 , n90492 );
nand ( n90494 , n90192 , n90186 );
and ( n90495 , n90494 , n90195 );
not ( n90496 , n90184 );
nor ( n90497 , n90495 , n90496 );
nand ( n90498 , n90493 , n90497 );
nand ( n90499 , n90197 , n90185 );
not ( n90500 , n90499 );
and ( n90501 , n90498 , n90500 );
not ( n90502 , n90498 );
and ( n90503 , n90502 , n90499 );
nor ( n90504 , n90501 , n90503 );
buf ( n90505 , n90504 );
nand ( n90506 , n90195 , n90184 );
not ( n90507 , n90180 );
not ( n90508 , n90491 );
or ( n90509 , n90507 , n90508 );
not ( n90510 , n90494 );
nand ( n90511 , n90509 , n90510 );
xnor ( n90512 , n90506 , n90511 );
and ( n90513 , n90505 , n90512 );
not ( n90514 , n90505 );
not ( n90515 , n90512 );
and ( n90516 , n90514 , n90515 );
nor ( n90517 , n90513 , n90516 );
not ( n90518 , n90517 );
not ( n90519 , n90515 );
not ( n90520 , n90179 );
not ( n90521 , n90520 );
not ( n90522 , n90491 );
or ( n90523 , n90521 , n90522 );
nand ( n90524 , n90523 , n90190 );
nand ( n90525 , n90189 , n90186 );
not ( n90526 , n90525 );
and ( n90527 , n90524 , n90526 );
not ( n90528 , n90524 );
and ( n90529 , n90528 , n90525 );
nor ( n90530 , n90527 , n90529 );
not ( n90531 , n90530 );
or ( n90532 , n90519 , n90531 );
not ( n90533 , n90530 );
nand ( n90534 , n90512 , n90533 );
nand ( n90535 , n90532 , n90534 );
nor ( n90536 , n90518 , n90535 );
buf ( n90537 , n90536 );
not ( n90538 , n90537 );
not ( n90539 , n90504 );
not ( n90540 , n90539 );
not ( n90541 , n90540 );
not ( n90542 , n88994 );
not ( n90543 , n90542 );
not ( n90544 , n89990 );
or ( n90545 , n90543 , n90544 );
nand ( n90546 , n90545 , n89994 );
not ( n90547 , n88911 );
nand ( n90548 , n90547 , n89996 );
nor ( n90549 , n90546 , n90548 );
and ( n90550 , n90546 , n90548 );
or ( n90551 , n90549 , n90550 );
not ( n90552 , n90551 );
not ( n90553 , n90552 );
or ( n90554 , n90541 , n90553 );
buf ( n90555 , n90551 );
nand ( n90556 , n90555 , n90539 );
nand ( n90557 , n90554 , n90556 );
not ( n90558 , n90557 );
or ( n90559 , n90538 , n90558 );
not ( n90560 , n90540 );
and ( n90561 , n89102 , n89096 );
not ( n90562 , n89102 );
and ( n90563 , n90562 , n89097 );
nor ( n90564 , n90561 , n90563 );
not ( n90565 , n90564 );
not ( n90566 , n90565 );
not ( n90567 , n89990 );
not ( n90568 , n88995 );
or ( n90569 , n90567 , n90568 );
not ( n90570 , n89997 );
nand ( n90571 , n90569 , n90570 );
not ( n90572 , n90571 );
not ( n90573 , n90572 );
or ( n90574 , n90566 , n90573 );
nand ( n90575 , n90571 , n90564 );
nand ( n90576 , n90574 , n90575 );
not ( n90577 , n90576 );
not ( n90578 , n90577 );
or ( n90579 , n90560 , n90578 );
nand ( n90580 , n90576 , n90539 );
nand ( n90581 , n90579 , n90580 );
buf ( n90582 , n90535 );
nand ( n90583 , n90581 , n90582 );
nand ( n90584 , n90559 , n90583 );
xor ( n90585 , n90477 , n90584 );
not ( n90586 , n90209 );
not ( n90587 , n90256 );
or ( n90588 , n90586 , n90587 );
not ( n90589 , n90217 );
nand ( n90590 , n90588 , n90589 );
nand ( n90591 , n90234 , n90222 );
xor ( n90592 , n90590 , n90591 );
not ( n90593 , n90208 );
not ( n90594 , n90593 );
not ( n90595 , n90202 );
or ( n90596 , n90594 , n90595 );
nand ( n90597 , n90596 , n90214 );
not ( n90598 , n90207 );
nand ( n90599 , n90598 , n90216 );
and ( n90600 , n90597 , n90599 );
not ( n90601 , n90597 );
not ( n90602 , n90599 );
and ( n90603 , n90601 , n90602 );
nor ( n90604 , n90600 , n90603 );
and ( n90605 , n90592 , n90604 );
not ( n90606 , n90592 );
not ( n90607 , n90604 );
and ( n90608 , n90606 , n90607 );
or ( n90609 , n90605 , n90608 );
not ( n90610 , n90609 );
not ( n90611 , n90610 );
buf ( n90612 , n90243 );
not ( n90613 , n90612 );
or ( n90614 , n89121 , n89258 );
nand ( n90615 , n90614 , n89985 );
not ( n90616 , n90615 );
not ( n90617 , n90616 );
not ( n90618 , n89981 );
not ( n90619 , n90618 );
or ( n90620 , n90617 , n90619 );
nand ( n90621 , n89981 , n90615 );
nand ( n90622 , n90620 , n90621 );
not ( n90623 , n90622 );
not ( n90624 , n90623 );
or ( n90625 , n90613 , n90624 );
not ( n90626 , n90616 );
not ( n90627 , n90618 );
or ( n90628 , n90626 , n90627 );
nand ( n90629 , n90628 , n90621 );
not ( n90630 , n90612 );
nand ( n90631 , n90629 , n90630 );
nand ( n90632 , n90625 , n90631 );
not ( n90633 , n90632 );
or ( n90634 , n90611 , n90633 );
not ( n90635 , n89979 );
nand ( n90636 , n90635 , n89974 );
not ( n90637 , n90309 );
not ( n90638 , n89969 );
or ( n90639 , n90637 , n90638 );
nand ( n90640 , n90639 , n90307 );
and ( n90641 , n90636 , n90640 );
not ( n90642 , n90636 );
not ( n90643 , n90640 );
and ( n90644 , n90642 , n90643 );
nor ( n90645 , n90641 , n90644 );
not ( n90646 , n90645 );
and ( n90647 , n90612 , n90646 );
not ( n90648 , n90612 );
buf ( n90649 , n90645 );
and ( n90650 , n90648 , n90649 );
nor ( n90651 , n90647 , n90650 );
and ( n90652 , n90592 , n90246 );
not ( n90653 , n90592 );
and ( n90654 , n90653 , n90243 );
nor ( n90655 , n90652 , n90654 );
and ( n90656 , n90655 , n90609 );
buf ( n90657 , n90656 );
nand ( n90658 , n90651 , n90657 );
nand ( n90659 , n90634 , n90658 );
buf ( n90660 , n90607 );
nor ( n90661 , n89267 , n89988 );
and ( n90662 , n89981 , n90614 );
not ( n90663 , n89985 );
nor ( n90664 , n90662 , n90663 );
and ( n90665 , n90661 , n90664 );
not ( n90666 , n90661 );
not ( n90667 , n90664 );
and ( n90668 , n90666 , n90667 );
or ( n90669 , n90665 , n90668 );
and ( n90670 , n90660 , n90669 );
not ( n90671 , n90660 );
not ( n90672 , n90669 );
and ( n90673 , n90671 , n90672 );
nor ( n90674 , n90670 , n90673 );
not ( n90675 , n90674 );
and ( n90676 , n90593 , n90214 );
xor ( n90677 , n90676 , n90256 );
xor ( n90678 , n90677 , n90607 );
xnor ( n90679 , n90677 , n90504 );
and ( n90680 , n90678 , n90679 );
not ( n90681 , n90680 );
or ( n90682 , n90675 , n90681 );
nand ( n90683 , n90542 , n89994 );
not ( n90684 , n89990 );
not ( n90685 , n90684 );
and ( n90686 , n90683 , n90685 );
not ( n90687 , n90683 );
and ( n90688 , n90687 , n90684 );
or ( n90689 , n90686 , n90688 );
buf ( n90690 , n90689 );
and ( n90691 , n90660 , n90690 );
not ( n90692 , n90660 );
not ( n90693 , n90689 );
and ( n90694 , n90692 , n90693 );
nor ( n90695 , n90691 , n90694 );
not ( n90696 , n90679 );
buf ( n90697 , n90696 );
nand ( n90698 , n90695 , n90697 );
nand ( n90699 , n90682 , n90698 );
xor ( n90700 , n90659 , n90699 );
not ( n90701 , n90405 );
not ( n90702 , n90434 );
or ( n90703 , n90701 , n90702 );
and ( n90704 , n90407 , n90379 );
not ( n90705 , n90407 );
and ( n90706 , n90705 , n90380 );
nor ( n90707 , n90704 , n90706 );
or ( n90708 , n90707 , n90441 );
nand ( n90709 , n90703 , n90708 );
not ( n90710 , n90709 );
not ( n90711 , n89930 );
not ( n90712 , n90711 );
or ( n90713 , n89932 , n89936 );
nand ( n90714 , n90713 , n89939 );
not ( n90715 , n90714 );
or ( n90716 , n90712 , n90715 );
not ( n90717 , n90714 );
not ( n90718 , n90711 );
nand ( n90719 , n90717 , n90718 );
nand ( n90720 , n90716 , n90719 );
buf ( n90721 , n90720 );
not ( n90722 , n90387 );
and ( n90723 , n90721 , n90722 );
not ( n90724 , n90386 );
and ( n90725 , n90724 , n90370 );
nor ( n90726 , n90723 , n90725 );
nor ( n90727 , n90710 , n90726 );
not ( n90728 , n90324 );
not ( n90729 , n90302 );
or ( n90730 , n90728 , n90729 );
and ( n90731 , n90305 , n90471 );
not ( n90732 , n90305 );
and ( n90733 , n90732 , n90464 );
nor ( n90734 , n90731 , n90733 );
nand ( n90735 , n90734 , n90279 );
nand ( n90736 , n90730 , n90735 );
xor ( n90737 , n90727 , n90736 );
xor ( n90738 , n90389 , n90444 );
and ( n90739 , n90737 , n90738 );
and ( n90740 , n90727 , n90736 );
or ( n90741 , n90739 , n90740 );
xor ( n90742 , n90700 , n90741 );
and ( n90743 , n90585 , n90742 );
and ( n90744 , n90477 , n90584 );
or ( n90745 , n90743 , n90744 );
xor ( n90746 , n90158 , n90745 );
not ( n90747 , n90726 );
not ( n90748 , n90709 );
or ( n90749 , n90747 , n90748 );
or ( n90750 , n90709 , n90726 );
nand ( n90751 , n90749 , n90750 );
not ( n90752 , n90324 );
not ( n90753 , n90734 );
or ( n90754 , n90752 , n90753 );
and ( n90755 , n90286 , n90418 );
not ( n90756 , n90286 );
and ( n90757 , n90756 , n90419 );
nor ( n90758 , n90755 , n90757 );
nand ( n90759 , n90758 , n90279 );
nand ( n90760 , n90754 , n90759 );
and ( n90761 , n90751 , n90760 );
not ( n90762 , n90610 );
not ( n90763 , n90651 );
or ( n90764 , n90762 , n90763 );
buf ( n90765 , n90317 );
and ( n90766 , n90612 , n90765 );
not ( n90767 , n90612 );
and ( n90768 , n90767 , n90318 );
nor ( n90769 , n90766 , n90768 );
nand ( n90770 , n90769 , n90657 );
nand ( n90771 , n90764 , n90770 );
xor ( n90772 , n90761 , n90771 );
xor ( n90773 , n90727 , n90736 );
xor ( n90774 , n90773 , n90738 );
and ( n90775 , n90772 , n90774 );
and ( n90776 , n90761 , n90771 );
or ( n90777 , n90775 , n90776 );
not ( n90778 , n90171 );
nor ( n90779 , n90778 , n90167 );
xor ( n90780 , n90779 , n90484 );
xor ( n90781 , n90780 , n87700 );
buf ( n90782 , n90781 );
not ( n90783 , n90782 );
and ( n90784 , n90169 , n90171 );
not ( n90785 , n90487 );
nand ( n90786 , n90785 , n90170 );
xor ( n90787 , n90784 , n90786 );
buf ( n90788 , n90787 );
not ( n90789 , n90788 );
nand ( n90790 , n88276 , n90048 );
not ( n90791 , n90790 );
and ( n90792 , n90045 , n90791 );
not ( n90793 , n90045 );
and ( n90794 , n90793 , n90790 );
nor ( n90795 , n90792 , n90794 );
not ( n90796 , n90795 );
not ( n90797 , n90796 );
or ( n90798 , n90789 , n90797 );
not ( n90799 , n90787 );
not ( n90800 , n90799 );
not ( n90801 , n90800 );
nand ( n90802 , n90795 , n90801 );
nand ( n90803 , n90798 , n90802 );
not ( n90804 , n90803 );
or ( n90805 , n90783 , n90804 );
not ( n90806 , n90788 );
not ( n90807 , n90026 );
not ( n90808 , n90008 );
or ( n90809 , n90807 , n90808 );
buf ( n90810 , n90039 );
nand ( n90811 , n90809 , n90810 );
not ( n90812 , n90034 );
nor ( n90813 , n90812 , n90043 );
xor ( n90814 , n90811 , n90813 );
not ( n90815 , n90814 );
not ( n90816 , n90815 );
or ( n90817 , n90806 , n90816 );
nand ( n90818 , n90814 , n90801 );
nand ( n90819 , n90817 , n90818 );
not ( n90820 , n90781 );
and ( n90821 , n90788 , n90780 );
nor ( n90822 , n90788 , n90780 );
nor ( n90823 , n90821 , n90822 );
and ( n90824 , n90820 , n90823 );
buf ( n90825 , n90824 );
nand ( n90826 , n90819 , n90825 );
nand ( n90827 , n90805 , n90826 );
xor ( n90828 , n90777 , n90827 );
nor ( n90829 , n90191 , n90179 );
xor ( n90830 , n90829 , n90491 );
xor ( n90831 , n90830 , n90530 );
not ( n90832 , n90787 );
not ( n90833 , n90832 );
not ( n90834 , n90830 );
not ( n90835 , n90834 );
or ( n90836 , n90833 , n90835 );
nand ( n90837 , n90830 , n90787 );
nand ( n90838 , n90836 , n90837 );
and ( n90839 , n90831 , n90838 );
buf ( n90840 , n90839 );
not ( n90841 , n90840 );
not ( n90842 , n90533 );
not ( n90843 , n90842 );
not ( n90844 , n90843 );
buf ( n90845 , n89103 );
nand ( n90846 , n90571 , n90845 );
and ( n90847 , n90846 , n90001 );
not ( n90848 , n90004 );
nor ( n90849 , n90848 , n90006 );
nor ( n90850 , n90847 , n90849 );
and ( n90851 , n90845 , n90571 );
nand ( n90852 , n90849 , n90001 );
nor ( n90853 , n90851 , n90852 );
nor ( n90854 , n90850 , n90853 );
not ( n90855 , n90854 );
and ( n90856 , n90844 , n90855 );
not ( n90857 , n90844 );
not ( n90858 , n90855 );
and ( n90859 , n90857 , n90858 );
nor ( n90860 , n90856 , n90859 );
not ( n90861 , n90860 );
or ( n90862 , n90841 , n90861 );
and ( n90863 , n90810 , n90026 );
buf ( n90864 , n90008 );
not ( n90865 , n90864 );
and ( n90866 , n90863 , n90865 );
not ( n90867 , n90863 );
and ( n90868 , n90867 , n90864 );
or ( n90869 , n90866 , n90868 );
buf ( n90870 , n90869 );
and ( n90871 , n90844 , n90870 );
not ( n90872 , n90844 );
not ( n90873 , n90869 );
and ( n90874 , n90872 , n90873 );
nor ( n90875 , n90871 , n90874 );
not ( n90876 , n90838 );
nand ( n90877 , n90875 , n90876 );
nand ( n90878 , n90862 , n90877 );
and ( n90879 , n90828 , n90878 );
and ( n90880 , n90777 , n90827 );
or ( n90881 , n90879 , n90880 );
xor ( n90882 , n90746 , n90881 );
xor ( n90883 , n90477 , n90584 );
xor ( n90884 , n90883 , n90742 );
xor ( n90885 , n90777 , n90827 );
xor ( n90886 , n90885 , n90878 );
xor ( n90887 , n90884 , n90886 );
xor ( n90888 , n90760 , n90751 );
not ( n90889 , n90582 );
not ( n90890 , n90539 );
and ( n90891 , n90890 , n90690 );
not ( n90892 , n90890 );
and ( n90893 , n90892 , n90693 );
nor ( n90894 , n90891 , n90893 );
not ( n90895 , n90894 );
or ( n90896 , n90889 , n90895 );
not ( n90897 , n90540 );
not ( n90898 , n90672 );
or ( n90899 , n90897 , n90898 );
nand ( n90900 , n90669 , n90539 );
nand ( n90901 , n90899 , n90900 );
nand ( n90902 , n90901 , n90537 );
nand ( n90903 , n90896 , n90902 );
xor ( n90904 , n90888 , n90903 );
not ( n90905 , n90442 );
not ( n90906 , n90407 );
not ( n90907 , n90721 );
or ( n90908 , n90906 , n90907 );
or ( n90909 , n90721 , n90407 );
nand ( n90910 , n90908 , n90909 );
not ( n90911 , n90910 );
not ( n90912 , n90911 );
or ( n90913 , n90905 , n90912 );
and ( n90914 , n90422 , n90724 );
not ( n90915 , n90422 );
and ( n90916 , n90915 , n90386 );
nor ( n90917 , n90914 , n90916 );
not ( n90918 , n90917 );
nand ( n90919 , n90918 , n90405 );
nand ( n90920 , n90913 , n90919 );
not ( n90921 , n90370 );
not ( n90922 , n89929 );
nand ( n90923 , n90922 , n89927 );
not ( n90924 , n89877 );
not ( n90925 , n89903 );
and ( n90926 , n90924 , n90925 );
not ( n90927 , n89905 );
nor ( n90928 , n90926 , n90927 );
and ( n90929 , n90923 , n90928 );
not ( n90930 , n90923 );
and ( n90931 , n90930 , n89906 );
nor ( n90932 , n90929 , n90931 );
not ( n90933 , n90932 );
not ( n90934 , n90933 );
not ( n90935 , n90934 );
or ( n90936 , n90921 , n90935 );
not ( n90937 , n89903 );
nand ( n90938 , n90937 , n89905 );
not ( n90939 , n90938 );
not ( n90940 , n90939 );
not ( n90941 , n89877 );
or ( n90942 , n90940 , n90941 );
not ( n90943 , n89877 );
nand ( n90944 , n90938 , n90943 );
nand ( n90945 , n90942 , n90944 );
not ( n90946 , n90945 );
or ( n90947 , n90946 , n90387 );
nand ( n90948 , n90936 , n90947 );
xor ( n90949 , n90920 , n90948 );
not ( n90950 , n90324 );
not ( n90951 , n90286 );
not ( n90952 , n90429 );
or ( n90953 , n90951 , n90952 );
nand ( n90954 , n90430 , n90321 );
nand ( n90955 , n90953 , n90954 );
not ( n90956 , n90955 );
or ( n90957 , n90950 , n90956 );
not ( n90958 , n90286 );
not ( n90959 , n90379 );
or ( n90960 , n90958 , n90959 );
nand ( n90961 , n90380 , n90321 );
nand ( n90962 , n90960 , n90961 );
nand ( n90963 , n90962 , n90279 );
nand ( n90964 , n90957 , n90963 );
and ( n90965 , n90949 , n90964 );
and ( n90966 , n90920 , n90948 );
or ( n90967 , n90965 , n90966 );
not ( n90968 , n90967 );
not ( n90969 , n90610 );
and ( n90970 , n90612 , n90297 );
not ( n90971 , n90612 );
and ( n90972 , n90971 , n90300 );
nor ( n90973 , n90970 , n90972 );
not ( n90974 , n90973 );
or ( n90975 , n90969 , n90974 );
and ( n90976 , n90612 , n90471 );
not ( n90977 , n90612 );
and ( n90978 , n90977 , n90464 );
nor ( n90979 , n90976 , n90978 );
nand ( n90980 , n90979 , n90656 );
nand ( n90981 , n90975 , n90980 );
not ( n90982 , n90981 );
or ( n90983 , n90968 , n90982 );
not ( n90984 , n90967 );
not ( n90985 , n90984 );
not ( n90986 , n90981 );
not ( n90987 , n90986 );
or ( n90988 , n90985 , n90987 );
buf ( n90989 , n90933 );
or ( n90990 , n90989 , n90387 );
not ( n90991 , n90720 );
or ( n90992 , n90991 , n90369 );
nand ( n90993 , n90990 , n90992 );
or ( n90994 , n90917 , n90441 );
not ( n90995 , n90405 );
or ( n90996 , n90707 , n90995 );
nand ( n90997 , n90994 , n90996 );
xor ( n90998 , n90993 , n90997 );
not ( n90999 , n90324 );
not ( n91000 , n90758 );
or ( n91001 , n90999 , n91000 );
nand ( n91002 , n90955 , n90279 );
nand ( n91003 , n91001 , n91002 );
xor ( n91004 , n90998 , n91003 );
nand ( n91005 , n90988 , n91004 );
nand ( n91006 , n90983 , n91005 );
and ( n91007 , n90904 , n91006 );
and ( n91008 , n90888 , n90903 );
or ( n91009 , n91007 , n91008 );
not ( n91010 , n90697 );
not ( n91011 , n91010 );
not ( n91012 , n91011 );
not ( n91013 , n90674 );
or ( n91014 , n91012 , n91013 );
and ( n91015 , n90660 , n90629 );
not ( n91016 , n90660 );
and ( n91017 , n91016 , n90623 );
nor ( n91018 , n91015 , n91017 );
nand ( n91019 , n91018 , n90680 );
nand ( n91020 , n91014 , n91019 );
not ( n91021 , n90656 );
not ( n91022 , n90973 );
or ( n91023 , n91021 , n91022 );
nand ( n91024 , n90769 , n90610 );
nand ( n91025 , n91023 , n91024 );
not ( n91026 , n91025 );
not ( n91027 , n91026 );
not ( n91028 , n90680 );
and ( n91029 , n90660 , n90646 );
not ( n91030 , n90660 );
and ( n91031 , n91030 , n90649 );
nor ( n91032 , n91029 , n91031 );
not ( n91033 , n91032 );
or ( n91034 , n91028 , n91033 );
nand ( n91035 , n91018 , n90697 );
nand ( n91036 , n91034 , n91035 );
not ( n91037 , n91036 );
not ( n91038 , n91037 );
or ( n91039 , n91027 , n91038 );
xor ( n91040 , n90993 , n90997 );
and ( n91041 , n91040 , n91003 );
and ( n91042 , n90993 , n90997 );
or ( n91043 , n91041 , n91042 );
nand ( n91044 , n91039 , n91043 );
not ( n91045 , n91026 );
nand ( n91046 , n91045 , n91036 );
nand ( n91047 , n91044 , n91046 );
xor ( n91048 , n91020 , n91047 );
not ( n91049 , n90582 );
not ( n91050 , n90557 );
or ( n91051 , n91049 , n91050 );
nand ( n91052 , n90894 , n90537 );
nand ( n91053 , n91051 , n91052 );
xor ( n91054 , n91048 , n91053 );
xor ( n91055 , n91009 , n91054 );
not ( n91056 , n87689 );
not ( n91057 , n87706 );
not ( n91058 , n88276 );
not ( n91059 , n90045 );
or ( n91060 , n91058 , n91059 );
nand ( n91061 , n91060 , n90048 );
not ( n91062 , n88321 );
nand ( n91063 , n91062 , n90050 );
and ( n91064 , n91061 , n91063 );
not ( n91065 , n91061 );
not ( n91066 , n91063 );
and ( n91067 , n91065 , n91066 );
nor ( n91068 , n91064 , n91067 );
not ( n91069 , n91068 );
or ( n91070 , n91057 , n91069 );
not ( n91071 , n91068 );
nand ( n91072 , n91071 , n87705 );
nand ( n91073 , n91070 , n91072 );
not ( n91074 , n91073 );
or ( n91075 , n91056 , n91074 );
and ( n91076 , n87705 , n90796 );
not ( n91077 , n87705 );
and ( n91078 , n91077 , n90795 );
nor ( n91079 , n91076 , n91078 );
nand ( n91080 , n91079 , n87702 );
nand ( n91081 , n91075 , n91080 );
and ( n91082 , n91055 , n91081 );
and ( n91083 , n91009 , n91054 );
or ( n91084 , n91082 , n91083 );
and ( n91085 , n90887 , n91084 );
and ( n91086 , n90884 , n90886 );
or ( n91087 , n91085 , n91086 );
xor ( n91088 , n90882 , n91087 );
and ( n91089 , n90451 , n90475 );
not ( n91090 , n90305 );
not ( n91091 , n90649 );
or ( n91092 , n91090 , n91091 );
nand ( n91093 , n90646 , n90321 );
nand ( n91094 , n91092 , n91093 );
not ( n91095 , n91094 );
or ( n91096 , n91095 , n90249 );
nand ( n91097 , n90323 , n90279 );
nand ( n91098 , n91096 , n91097 );
xor ( n91099 , n91089 , n91098 );
not ( n91100 , n90440 );
not ( n91101 , n90473 );
or ( n91102 , n91100 , n91101 );
not ( n91103 , n90995 );
not ( n91104 , n90407 );
not ( n91105 , n90300 );
or ( n91106 , n91104 , n91105 );
nand ( n91107 , n90297 , n90422 );
nand ( n91108 , n91106 , n91107 );
nand ( n91109 , n91103 , n91108 );
nand ( n91110 , n91102 , n91109 );
not ( n91111 , n90429 );
not ( n91112 , n90387 );
and ( n91113 , n91111 , n91112 );
and ( n91114 , n90418 , n90370 );
nor ( n91115 , n91113 , n91114 );
xnor ( n91116 , n91110 , n91115 );
xor ( n91117 , n91099 , n91116 );
not ( n91118 , n90840 );
not ( n91119 , n90875 );
or ( n91120 , n91118 , n91119 );
not ( n91121 , n90844 );
not ( n91122 , n90815 );
or ( n91123 , n91121 , n91122 );
nand ( n91124 , n90814 , n90843 );
nand ( n91125 , n91123 , n91124 );
nand ( n91126 , n91125 , n90876 );
nand ( n91127 , n91120 , n91126 );
xor ( n91128 , n91117 , n91127 );
not ( n91129 , n90582 );
and ( n91130 , n90890 , n90855 );
not ( n91131 , n90890 );
and ( n91132 , n91131 , n90858 );
nor ( n91133 , n91130 , n91132 );
not ( n91134 , n91133 );
or ( n91135 , n91129 , n91134 );
nand ( n91136 , n90581 , n90537 );
nand ( n91137 , n91135 , n91136 );
xor ( n91138 , n91128 , n91137 );
xor ( n91139 , n90659 , n90699 );
and ( n91140 , n91139 , n90741 );
and ( n91141 , n90659 , n90699 );
or ( n91142 , n91140 , n91141 );
xor ( n91143 , n90326 , n90445 );
and ( n91144 , n91143 , n90476 );
and ( n91145 , n90326 , n90445 );
or ( n91146 , n91144 , n91145 );
not ( n91147 , n90610 );
not ( n91148 , n90612 );
not ( n91149 , n90672 );
or ( n91150 , n91148 , n91149 );
nand ( n91151 , n90669 , n90630 );
nand ( n91152 , n91150 , n91151 );
not ( n91153 , n91152 );
or ( n91154 , n91147 , n91153 );
nand ( n91155 , n90632 , n90657 );
nand ( n91156 , n91154 , n91155 );
xor ( n91157 , n91146 , n91156 );
not ( n91158 , n90680 );
not ( n91159 , n90695 );
or ( n91160 , n91158 , n91159 );
not ( n91161 , n90660 );
not ( n91162 , n90552 );
or ( n91163 , n91161 , n91162 );
not ( n91164 , n90660 );
nand ( n91165 , n90555 , n91164 );
nand ( n91166 , n91163 , n91165 );
nand ( n91167 , n91166 , n91011 );
nand ( n91168 , n91160 , n91167 );
xor ( n91169 , n91157 , n91168 );
xor ( n91170 , n91142 , n91169 );
not ( n91171 , n90825 );
not ( n91172 , n90803 );
or ( n91173 , n91171 , n91172 );
not ( n91174 , n90788 );
not ( n91175 , n91068 );
or ( n91176 , n91174 , n91175 );
nand ( n91177 , n91071 , n90801 );
nand ( n91178 , n91176 , n91177 );
nand ( n91179 , n91178 , n90782 );
nand ( n91180 , n91173 , n91179 );
xor ( n91181 , n91170 , n91180 );
xor ( n91182 , n91138 , n91181 );
xor ( n91183 , n91020 , n91047 );
and ( n91184 , n91183 , n91053 );
and ( n91185 , n91020 , n91047 );
or ( n91186 , n91184 , n91185 );
not ( n91187 , n91186 );
not ( n91188 , n87702 );
not ( n91189 , n91073 );
or ( n91190 , n91188 , n91189 );
nand ( n91191 , n90104 , n87689 );
nand ( n91192 , n91190 , n91191 );
not ( n91193 , n91192 );
or ( n91194 , n91187 , n91193 );
not ( n91195 , n91186 );
not ( n91196 , n91195 );
not ( n91197 , n91192 );
not ( n91198 , n91197 );
or ( n91199 , n91196 , n91198 );
not ( n91200 , n90782 );
not ( n91201 , n90819 );
or ( n91202 , n91200 , n91201 );
not ( n91203 , n90788 );
not ( n91204 , n90873 );
or ( n91205 , n91203 , n91204 );
nand ( n91206 , n90870 , n90799 );
nand ( n91207 , n91205 , n91206 );
nand ( n91208 , n91207 , n90825 );
nand ( n91209 , n91202 , n91208 );
xor ( n91210 , n90761 , n90771 );
xor ( n91211 , n91210 , n90774 );
xor ( n91212 , n91209 , n91211 );
not ( n91213 , n90840 );
not ( n91214 , n90844 );
not ( n91215 , n90577 );
or ( n91216 , n91214 , n91215 );
nand ( n91217 , n90576 , n90843 );
nand ( n91218 , n91216 , n91217 );
not ( n91219 , n91218 );
or ( n91220 , n91213 , n91219 );
nand ( n91221 , n90860 , n90876 );
nand ( n91222 , n91220 , n91221 );
and ( n91223 , n91212 , n91222 );
and ( n91224 , n91209 , n91211 );
or ( n91225 , n91223 , n91224 );
nand ( n91226 , n91199 , n91225 );
nand ( n91227 , n91194 , n91226 );
xor ( n91228 , n91182 , n91227 );
xnor ( n91229 , n91088 , n91228 );
not ( n91230 , n91186 );
not ( n91231 , n91197 );
or ( n91232 , n91230 , n91231 );
nand ( n91233 , n91195 , n91192 );
nand ( n91234 , n91232 , n91233 );
xnor ( n91235 , n91234 , n91225 );
not ( n91236 , n91235 );
xor ( n91237 , n90884 , n90886 );
xor ( n91238 , n91237 , n91084 );
not ( n91239 , n91238 );
not ( n91240 , n91239 );
or ( n91241 , n91236 , n91240 );
not ( n91242 , n90840 );
not ( n91243 , n90844 );
not ( n91244 , n90552 );
or ( n91245 , n91243 , n91244 );
nand ( n91246 , n90555 , n90843 );
nand ( n91247 , n91245 , n91246 );
not ( n91248 , n91247 );
or ( n91249 , n91242 , n91248 );
nand ( n91250 , n91218 , n90876 );
nand ( n91251 , n91249 , n91250 );
nand ( n91252 , n91037 , n91043 , n91026 );
not ( n91253 , n91043 );
buf ( n91254 , n91025 );
nand ( n91255 , n91253 , n91037 , n91254 );
nand ( n91256 , n91036 , n91043 , n91254 );
nor ( n91257 , n91043 , n91254 );
nand ( n91258 , n91036 , n91257 );
nand ( n91259 , n91252 , n91255 , n91256 , n91258 );
xor ( n91260 , n91251 , n91259 );
not ( n91261 , n90825 );
not ( n91262 , n90788 );
not ( n91263 , n90858 );
or ( n91264 , n91262 , n91263 );
nand ( n91265 , n90855 , n90799 );
nand ( n91266 , n91264 , n91265 );
not ( n91267 , n91266 );
or ( n91268 , n91261 , n91267 );
nand ( n91269 , n91207 , n90782 );
nand ( n91270 , n91268 , n91269 );
and ( n91271 , n91260 , n91270 );
and ( n91272 , n91251 , n91259 );
or ( n91273 , n91271 , n91272 );
xor ( n91274 , n91209 , n91211 );
xor ( n91275 , n91274 , n91222 );
xor ( n91276 , n91273 , n91275 );
and ( n91277 , n90660 , n90765 );
not ( n91278 , n90660 );
and ( n91279 , n91278 , n90318 );
nor ( n91280 , n91277 , n91279 );
not ( n91281 , n91280 );
not ( n91282 , n90680 );
or ( n91283 , n91281 , n91282 );
not ( n91284 , n91032 );
or ( n91285 , n91284 , n91010 );
nand ( n91286 , n91283 , n91285 );
not ( n91287 , n90370 );
not ( n91288 , n90945 );
or ( n91289 , n91287 , n91288 );
and ( n91290 , n89835 , n89875 );
not ( n91291 , n91290 );
buf ( n91292 , n89873 );
nand ( n91293 , n91291 , n91292 );
not ( n91294 , n91292 );
nand ( n91295 , n91290 , n91294 );
nand ( n91296 , n91293 , n91295 );
not ( n91297 , n91296 );
not ( n91298 , n91297 );
not ( n91299 , n91298 );
or ( n91300 , n91299 , n90387 );
nand ( n91301 , n91289 , n91300 );
or ( n91302 , n90910 , n90404 );
and ( n91303 , n90407 , n90989 );
not ( n91304 , n90407 );
and ( n91305 , n91304 , n90934 );
nor ( n91306 , n91303 , n91305 );
or ( n91307 , n91306 , n90441 );
nand ( n91308 , n91302 , n91307 );
xor ( n91309 , n91301 , n91308 );
not ( n91310 , n90324 );
not ( n91311 , n90962 );
or ( n91312 , n91310 , n91311 );
not ( n91313 , n90305 );
not ( n91314 , n90386 );
or ( n91315 , n91313 , n91314 );
nand ( n91316 , n90724 , n90321 );
nand ( n91317 , n91315 , n91316 );
nand ( n91318 , n91317 , n90279 );
nand ( n91319 , n91312 , n91318 );
and ( n91320 , n91309 , n91319 );
and ( n91321 , n91301 , n91308 );
or ( n91322 , n91320 , n91321 );
not ( n91323 , n90610 );
not ( n91324 , n90979 );
or ( n91325 , n91323 , n91324 );
and ( n91326 , n90612 , n90418 );
not ( n91327 , n90612 );
and ( n91328 , n91327 , n90419 );
nor ( n91329 , n91326 , n91328 );
nand ( n91330 , n91329 , n90657 );
nand ( n91331 , n91325 , n91330 );
xor ( n91332 , n91322 , n91331 );
xor ( n91333 , n90920 , n90948 );
xor ( n91334 , n91333 , n90964 );
and ( n91335 , n91332 , n91334 );
and ( n91336 , n91322 , n91331 );
or ( n91337 , n91335 , n91336 );
xor ( n91338 , n91286 , n91337 );
not ( n91339 , n90582 );
not ( n91340 , n90901 );
or ( n91341 , n91339 , n91340 );
and ( n91342 , n90540 , n90622 );
not ( n91343 , n90540 );
and ( n91344 , n91343 , n90623 );
nor ( n91345 , n91342 , n91344 );
nand ( n91346 , n91345 , n90537 );
nand ( n91347 , n91341 , n91346 );
and ( n91348 , n91338 , n91347 );
and ( n91349 , n91286 , n91337 );
or ( n91350 , n91348 , n91349 );
not ( n91351 , n91350 );
not ( n91352 , n87689 );
not ( n91353 , n91079 );
or ( n91354 , n91352 , n91353 );
not ( n91355 , n87706 );
not ( n91356 , n90815 );
or ( n91357 , n91355 , n91356 );
nand ( n91358 , n90814 , n87705 );
nand ( n91359 , n91357 , n91358 );
nand ( n91360 , n91359 , n87702 );
nand ( n91361 , n91354 , n91360 );
not ( n91362 , n91361 );
or ( n91363 , n91351 , n91362 );
and ( n91364 , n90842 , n90690 );
not ( n91365 , n90842 );
and ( n91366 , n91365 , n90693 );
nor ( n91367 , n91364 , n91366 );
not ( n91368 , n91367 );
not ( n91369 , n90840 );
or ( n91370 , n91368 , n91369 );
not ( n91371 , n91247 );
or ( n91372 , n91371 , n90838 );
nand ( n91373 , n91370 , n91372 );
xor ( n91374 , n90967 , n90986 );
xnor ( n91375 , n91374 , n91004 );
or ( n91376 , n91373 , n91375 );
not ( n91377 , n90697 );
not ( n91378 , n91280 );
or ( n91379 , n91377 , n91378 );
and ( n91380 , n90660 , n90297 );
not ( n91381 , n90660 );
and ( n91382 , n91381 , n90300 );
nor ( n91383 , n91380 , n91382 );
nand ( n91384 , n91383 , n90680 );
nand ( n91385 , n91379 , n91384 );
xor ( n91386 , n91301 , n91308 );
xor ( n91387 , n91386 , n91319 );
not ( n91388 , n91387 );
not ( n91389 , n90370 );
not ( n91390 , n91297 );
not ( n91391 , n91390 );
or ( n91392 , n91389 , n91391 );
xor ( n91393 , n89844 , n89845 );
xor ( n91394 , n91393 , n89870 );
not ( n91395 , n91394 );
or ( n91396 , n91395 , n90387 );
nand ( n91397 , n91392 , n91396 );
nor ( n91398 , n91306 , n90995 );
nor ( n91399 , n90938 , n90943 );
not ( n91400 , n91399 );
nand ( n91401 , n91400 , n90944 );
and ( n91402 , n90407 , n91401 );
not ( n91403 , n90407 );
and ( n91404 , n91403 , n90946 );
nor ( n91405 , n91402 , n91404 );
not ( n91406 , n91405 );
nor ( n91407 , n91406 , n90441 );
or ( n91408 , n91398 , n91407 );
xor ( n91409 , n91397 , n91408 );
not ( n91410 , n90324 );
not ( n91411 , n91317 );
or ( n91412 , n91410 , n91411 );
not ( n91413 , n90286 );
not ( n91414 , n90991 );
or ( n91415 , n91413 , n91414 );
nand ( n91416 , n90721 , n90321 );
nand ( n91417 , n91415 , n91416 );
nand ( n91418 , n91417 , n90279 );
nand ( n91419 , n91412 , n91418 );
and ( n91420 , n91409 , n91419 );
and ( n91421 , n91397 , n91408 );
or ( n91422 , n91420 , n91421 );
not ( n91423 , n91422 );
nand ( n91424 , n91388 , n91423 );
not ( n91425 , n91424 );
not ( n91426 , n90656 );
and ( n91427 , n90612 , n90430 );
not ( n91428 , n90612 );
and ( n91429 , n91428 , n90429 );
nor ( n91430 , n91427 , n91429 );
not ( n91431 , n91430 );
or ( n91432 , n91426 , n91431 );
nand ( n91433 , n91329 , n90610 );
nand ( n91434 , n91432 , n91433 );
not ( n91435 , n91434 );
or ( n91436 , n91425 , n91435 );
not ( n91437 , n91423 );
nand ( n91438 , n91437 , n91387 );
nand ( n91439 , n91436 , n91438 );
xor ( n91440 , n91385 , n91439 );
nand ( n91441 , n91345 , n90582 );
and ( n91442 , n90540 , n90646 );
not ( n91443 , n90540 );
and ( n91444 , n91443 , n90649 );
nor ( n91445 , n91442 , n91444 );
nand ( n91446 , n90537 , n91445 );
nand ( n91447 , n91441 , n91446 );
and ( n91448 , n91440 , n91447 );
and ( n91449 , n91385 , n91439 );
or ( n91450 , n91448 , n91449 );
nand ( n91451 , n91376 , n91450 );
nand ( n91452 , n91375 , n91373 );
nand ( n91453 , n91451 , n91452 );
not ( n91454 , n91350 );
not ( n91455 , n91361 );
nand ( n91456 , n91454 , n91455 );
nand ( n91457 , n91453 , n91456 );
nand ( n91458 , n91363 , n91457 );
and ( n91459 , n91276 , n91458 );
and ( n91460 , n91273 , n91275 );
or ( n91461 , n91459 , n91460 );
nand ( n91462 , n91241 , n91461 );
not ( n91463 , n91235 );
nand ( n91464 , n91463 , n91238 );
and ( n91465 , n91462 , n91464 );
nor ( n91466 , n91229 , n91465 );
not ( n91467 , n91466 );
nand ( n91468 , n91229 , n91465 );
nand ( n91469 , n91467 , n91468 );
xor ( n91470 , n91461 , n91235 );
and ( n91471 , n91470 , n91238 );
not ( n91472 , n91470 );
and ( n91473 , n91472 , n91239 );
nor ( n91474 , n91471 , n91473 );
xor ( n91475 , n91273 , n91275 );
xor ( n91476 , n91475 , n91458 );
xor ( n91477 , n90888 , n90903 );
xor ( n91478 , n91477 , n91006 );
xor ( n91479 , n91251 , n91259 );
xor ( n91480 , n91479 , n91270 );
xor ( n91481 , n91478 , n91480 );
not ( n91482 , n87702 );
not ( n91483 , n87706 );
not ( n91484 , n90873 );
or ( n91485 , n91483 , n91484 );
nand ( n91486 , n90870 , n87705 );
nand ( n91487 , n91485 , n91486 );
not ( n91488 , n91487 );
or ( n91489 , n91482 , n91488 );
nand ( n91490 , n91359 , n87689 );
nand ( n91491 , n91489 , n91490 );
xor ( n91492 , n91286 , n91337 );
xor ( n91493 , n91492 , n91347 );
xor ( n91494 , n91491 , n91493 );
not ( n91495 , n90825 );
and ( n91496 , n90788 , n90576 );
not ( n91497 , n90788 );
and ( n91498 , n91497 , n90577 );
nor ( n91499 , n91496 , n91498 );
not ( n91500 , n91499 );
or ( n91501 , n91495 , n91500 );
nand ( n91502 , n91266 , n90782 );
nand ( n91503 , n91501 , n91502 );
and ( n91504 , n91494 , n91503 );
and ( n91505 , n91491 , n91493 );
or ( n91506 , n91504 , n91505 );
and ( n91507 , n91481 , n91506 );
and ( n91508 , n91478 , n91480 );
or ( n91509 , n91507 , n91508 );
not ( n91510 , n91509 );
xor ( n91511 , n91009 , n91054 );
xor ( n91512 , n91511 , n91081 );
not ( n91513 , n91512 );
nand ( n91514 , n91510 , n91513 );
and ( n91515 , n91476 , n91514 );
and ( n91516 , n91512 , n91509 );
nor ( n91517 , n91515 , n91516 );
nand ( n91518 , n91474 , n91517 );
not ( n91519 , n91509 );
not ( n91520 , n91513 );
or ( n91521 , n91519 , n91520 );
nand ( n91522 , n91510 , n91512 );
nand ( n91523 , n91521 , n91522 );
not ( n91524 , n91476 );
and ( n91525 , n91523 , n91524 );
not ( n91526 , n91523 );
and ( n91527 , n91526 , n91476 );
nor ( n91528 , n91525 , n91527 );
xor ( n91529 , n91478 , n91480 );
xor ( n91530 , n91529 , n91506 );
not ( n91531 , n91530 );
not ( n91532 , n91531 );
not ( n91533 , n91455 );
not ( n91534 , n91350 );
and ( n91535 , n91533 , n91534 );
and ( n91536 , n91350 , n91455 );
nor ( n91537 , n91535 , n91536 );
xor ( n91538 , n91537 , n91453 );
not ( n91539 , n91538 );
and ( n91540 , n91532 , n91539 );
nand ( n91541 , n91531 , n91538 );
xor ( n91542 , n91322 , n91331 );
xor ( n91543 , n91542 , n91334 );
not ( n91544 , n90876 );
not ( n91545 , n91367 );
or ( n91546 , n91544 , n91545 );
and ( n91547 , n90842 , n90669 );
not ( n91548 , n90842 );
and ( n91549 , n91548 , n90672 );
nor ( n91550 , n91547 , n91549 );
nand ( n91551 , n91550 , n90839 );
nand ( n91552 , n91546 , n91551 );
buf ( n91553 , n91552 );
xor ( n91554 , n91543 , n91553 );
not ( n91555 , n90782 );
not ( n91556 , n91499 );
or ( n91557 , n91555 , n91556 );
not ( n91558 , n90788 );
not ( n91559 , n90552 );
or ( n91560 , n91558 , n91559 );
nand ( n91561 , n90555 , n90799 );
nand ( n91562 , n91560 , n91561 );
nand ( n91563 , n91562 , n90825 );
nand ( n91564 , n91557 , n91563 );
and ( n91565 , n91554 , n91564 );
and ( n91566 , n91543 , n91553 );
or ( n91567 , n91565 , n91566 );
not ( n91568 , n91434 );
nand ( n91569 , n91568 , n91388 , n91422 );
nand ( n91570 , n91568 , n91387 , n91423 );
nand ( n91571 , n91434 , n91388 , n91423 );
nand ( n91572 , n91434 , n91387 , n91422 );
nand ( n91573 , n91569 , n91570 , n91571 , n91572 );
not ( n91574 , n91573 );
not ( n91575 , n90876 );
not ( n91576 , n91550 );
or ( n91577 , n91575 , n91576 );
and ( n91578 , n90842 , n90629 );
not ( n91579 , n90842 );
and ( n91580 , n91579 , n90623 );
nor ( n91581 , n91578 , n91580 );
nand ( n91582 , n91581 , n90839 );
nand ( n91583 , n91577 , n91582 );
not ( n91584 , n91583 );
not ( n91585 , n90370 );
xor ( n91586 , n89847 , n89857 );
xor ( n91587 , n91586 , n89867 );
not ( n91588 , n91587 );
not ( n91589 , n91588 );
not ( n91590 , n91589 );
or ( n91591 , n91585 , n91590 );
not ( n91592 , n89867 );
nand ( n91593 , n89864 , n89866 );
nand ( n91594 , n91592 , n91593 );
not ( n91595 , n91594 );
not ( n91596 , n91595 );
or ( n91597 , n90387 , n91596 );
nand ( n91598 , n91591 , n91597 );
not ( n91599 , n90440 );
and ( n91600 , n90407 , n91394 );
not ( n91601 , n90407 );
and ( n91602 , n91601 , n91395 );
nor ( n91603 , n91600 , n91602 );
not ( n91604 , n91603 );
or ( n91605 , n91599 , n91604 );
and ( n91606 , n90437 , n91299 );
not ( n91607 , n90437 );
and ( n91608 , n91607 , n91390 );
nor ( n91609 , n91606 , n91608 );
nand ( n91610 , n91609 , n90405 );
nand ( n91611 , n91605 , n91610 );
xor ( n91612 , n91598 , n91611 );
or ( n91613 , n90387 , n89865 );
or ( n91614 , n91596 , n90369 );
nand ( n91615 , n91613 , n91614 );
not ( n91616 , n90405 );
not ( n91617 , n91603 );
or ( n91618 , n91616 , n91617 );
not ( n91619 , n90407 );
not ( n91620 , n91588 );
or ( n91621 , n91619 , n91620 );
buf ( n91622 , n91587 );
nand ( n91623 , n91622 , n90437 );
nand ( n91624 , n91621 , n91623 );
not ( n91625 , n91624 );
or ( n91626 , n91625 , n90441 );
nand ( n91627 , n91618 , n91626 );
xor ( n91628 , n91615 , n91627 );
nor ( n91629 , n90369 , n89865 );
not ( n91630 , n90405 );
not ( n91631 , n91624 );
or ( n91632 , n91630 , n91631 );
not ( n91633 , n90368 );
not ( n91634 , n91596 );
or ( n91635 , n91633 , n91634 );
nand ( n91636 , n91595 , n90437 );
nand ( n91637 , n91635 , n91636 );
nand ( n91638 , n91637 , n90440 );
nand ( n91639 , n91632 , n91638 );
xor ( n91640 , n91629 , n91639 );
not ( n91641 , n89865 );
and ( n91642 , n90400 , n91641 );
nor ( n91643 , n91642 , n90437 );
or ( n91644 , n90400 , n91641 );
nand ( n91645 , n91644 , n90286 );
and ( n91646 , n91643 , n91645 );
not ( n91647 , n90405 );
not ( n91648 , n91637 );
or ( n91649 , n91647 , n91648 );
or ( n91650 , n90368 , n89865 );
or ( n91651 , n90437 , n91641 );
nand ( n91652 , n91650 , n91651 );
nand ( n91653 , n90440 , n91652 );
nand ( n91654 , n91649 , n91653 );
and ( n91655 , n91646 , n91654 );
and ( n91656 , n91640 , n91655 );
and ( n91657 , n91629 , n91639 );
or ( n91658 , n91656 , n91657 );
and ( n91659 , n91628 , n91658 );
and ( n91660 , n91615 , n91627 );
or ( n91661 , n91659 , n91660 );
and ( n91662 , n91612 , n91661 );
and ( n91663 , n91598 , n91611 );
or ( n91664 , n91662 , n91663 );
or ( n91665 , n91588 , n90387 );
or ( n91666 , n91395 , n90369 );
nand ( n91667 , n91665 , n91666 );
not ( n91668 , n90405 );
not ( n91669 , n91405 );
or ( n91670 , n91668 , n91669 );
not ( n91671 , n91609 );
or ( n91672 , n91671 , n90441 );
nand ( n91673 , n91670 , n91672 );
xor ( n91674 , n91667 , n91673 );
not ( n91675 , n90324 );
not ( n91676 , n91417 );
or ( n91677 , n91675 , n91676 );
and ( n91678 , n90932 , n90286 );
not ( n91679 , n90932 );
and ( n91680 , n91679 , n90321 );
nor ( n91681 , n91678 , n91680 );
nand ( n91682 , n91681 , n90279 );
nand ( n91683 , n91677 , n91682 );
xor ( n91684 , n91674 , n91683 );
xor ( n91685 , n91664 , n91684 );
not ( n91686 , n90610 );
not ( n91687 , n90612 );
not ( n91688 , n90379 );
or ( n91689 , n91687 , n91688 );
nand ( n91690 , n90380 , n90630 );
nand ( n91691 , n91689 , n91690 );
not ( n91692 , n91691 );
or ( n91693 , n91686 , n91692 );
not ( n91694 , n90612 );
not ( n91695 , n90386 );
or ( n91696 , n91694 , n91695 );
nand ( n91697 , n90724 , n90630 );
nand ( n91698 , n91696 , n91697 );
nand ( n91699 , n91698 , n90656 );
nand ( n91700 , n91693 , n91699 );
and ( n91701 , n91685 , n91700 );
and ( n91702 , n91664 , n91684 );
or ( n91703 , n91701 , n91702 );
not ( n91704 , n90697 );
not ( n91705 , n90660 );
not ( n91706 , n90470 );
or ( n91707 , n91705 , n91706 );
or ( n91708 , n90470 , n90660 );
nand ( n91709 , n91707 , n91708 );
not ( n91710 , n91709 );
or ( n91711 , n91704 , n91710 );
and ( n91712 , n90660 , n90418 );
not ( n91713 , n90660 );
and ( n91714 , n91713 , n90419 );
nor ( n91715 , n91712 , n91714 );
nand ( n91716 , n91715 , n90680 );
nand ( n91717 , n91711 , n91716 );
xor ( n91718 , n91703 , n91717 );
not ( n91719 , n90537 );
and ( n91720 , n90540 , n90297 );
not ( n91721 , n90540 );
and ( n91722 , n91721 , n90300 );
nor ( n91723 , n91720 , n91722 );
not ( n91724 , n91723 );
or ( n91725 , n91719 , n91724 );
not ( n91726 , n90540 );
not ( n91727 , n90318 );
or ( n91728 , n91726 , n91727 );
nand ( n91729 , n90317 , n90539 );
nand ( n91730 , n91728 , n91729 );
nand ( n91731 , n91730 , n90582 );
nand ( n91732 , n91725 , n91731 );
and ( n91733 , n91718 , n91732 );
and ( n91734 , n91703 , n91717 );
or ( n91735 , n91733 , n91734 );
not ( n91736 , n91735 );
nand ( n91737 , n91584 , n91736 );
not ( n91738 , n91737 );
or ( n91739 , n91574 , n91738 );
and ( n91740 , n91583 , n91735 );
not ( n91741 , n91740 );
nand ( n91742 , n91739 , n91741 );
not ( n91743 , n91742 );
xor ( n91744 , n91385 , n91439 );
xor ( n91745 , n91744 , n91447 );
not ( n91746 , n91745 );
not ( n91747 , n90697 );
not ( n91748 , n91383 );
or ( n91749 , n91747 , n91748 );
nand ( n91750 , n91709 , n90680 );
nand ( n91751 , n91749 , n91750 );
xor ( n91752 , n91667 , n91673 );
and ( n91753 , n91752 , n91683 );
and ( n91754 , n91667 , n91673 );
or ( n91755 , n91753 , n91754 );
xor ( n91756 , n91397 , n91408 );
xor ( n91757 , n91756 , n91419 );
xor ( n91758 , n91755 , n91757 );
not ( n91759 , n90656 );
not ( n91760 , n91691 );
or ( n91761 , n91759 , n91760 );
nand ( n91762 , n91430 , n90610 );
nand ( n91763 , n91761 , n91762 );
and ( n91764 , n91758 , n91763 );
and ( n91765 , n91755 , n91757 );
or ( n91766 , n91764 , n91765 );
xor ( n91767 , n91751 , n91766 );
not ( n91768 , n90582 );
not ( n91769 , n91445 );
or ( n91770 , n91768 , n91769 );
nand ( n91771 , n91730 , n90537 );
nand ( n91772 , n91770 , n91771 );
and ( n91773 , n91767 , n91772 );
and ( n91774 , n91751 , n91766 );
or ( n91775 , n91773 , n91774 );
not ( n91776 , n91775 );
nand ( n91777 , n91746 , n91776 );
not ( n91778 , n91777 );
or ( n91779 , n91743 , n91778 );
nand ( n91780 , n91745 , n91775 );
nand ( n91781 , n91779 , n91780 );
xor ( n91782 , n91567 , n91781 );
xor ( n91783 , n91450 , n91375 );
xor ( n91784 , n91783 , n91373 );
and ( n91785 , n91782 , n91784 );
and ( n91786 , n91567 , n91781 );
or ( n91787 , n91785 , n91786 );
and ( n91788 , n91541 , n91787 );
nor ( n91789 , n91540 , n91788 );
nand ( n91790 , n91528 , n91789 );
and ( n91791 , n91518 , n91790 );
not ( n91792 , n91791 );
not ( n91793 , n91538 );
not ( n91794 , n91787 );
or ( n91795 , n91793 , n91794 );
or ( n91796 , n91787 , n91538 );
nand ( n91797 , n91795 , n91796 );
and ( n91798 , n91797 , n91530 );
not ( n91799 , n91797 );
and ( n91800 , n91799 , n91531 );
nor ( n91801 , n91798 , n91800 );
xor ( n91802 , n91491 , n91493 );
xor ( n91803 , n91802 , n91503 );
nand ( n91804 , n91487 , n87689 );
not ( n91805 , n87706 );
not ( n91806 , n90858 );
or ( n91807 , n91805 , n91806 );
nand ( n91808 , n90855 , n87705 );
nand ( n91809 , n91807 , n91808 );
nand ( n91810 , n91809 , n87702 );
nand ( n91811 , n91804 , n91810 );
xor ( n91812 , n91543 , n91553 );
xor ( n91813 , n91812 , n91564 );
xor ( n91814 , n91811 , n91813 );
xor ( n91815 , n91751 , n91766 );
xor ( n91816 , n91815 , n91772 );
not ( n91817 , n91816 );
not ( n91818 , n90782 );
not ( n91819 , n91562 );
or ( n91820 , n91818 , n91819 );
not ( n91821 , n90788 );
not ( n91822 , n90693 );
or ( n91823 , n91821 , n91822 );
nand ( n91824 , n90690 , n90799 );
nand ( n91825 , n91823 , n91824 );
nand ( n91826 , n91825 , n90825 );
nand ( n91827 , n91820 , n91826 );
not ( n91828 , n91827 );
or ( n91829 , n91817 , n91828 );
or ( n91830 , n91827 , n91816 );
xor ( n91831 , n91755 , n91757 );
xor ( n91832 , n91831 , n91763 );
not ( n91833 , n90876 );
not ( n91834 , n91581 );
or ( n91835 , n91833 , n91834 );
and ( n91836 , n90842 , n90646 );
not ( n91837 , n90842 );
and ( n91838 , n91837 , n90649 );
nor ( n91839 , n91836 , n91838 );
nand ( n91840 , n91839 , n90839 );
nand ( n91841 , n91835 , n91840 );
xor ( n91842 , n91832 , n91841 );
xor ( n91843 , n91703 , n91717 );
xor ( n91844 , n91843 , n91732 );
and ( n91845 , n91842 , n91844 );
and ( n91846 , n91832 , n91841 );
or ( n91847 , n91845 , n91846 );
nand ( n91848 , n91830 , n91847 );
nand ( n91849 , n91829 , n91848 );
and ( n91850 , n91814 , n91849 );
and ( n91851 , n91811 , n91813 );
or ( n91852 , n91850 , n91851 );
xor ( n91853 , n91803 , n91852 );
xor ( n91854 , n91567 , n91781 );
xor ( n91855 , n91854 , n91784 );
and ( n91856 , n91853 , n91855 );
and ( n91857 , n91803 , n91852 );
or ( n91858 , n91856 , n91857 );
nor ( n91859 , n91801 , n91858 );
xor ( n91860 , n91803 , n91852 );
xor ( n91861 , n91860 , n91855 );
not ( n91862 , n87689 );
not ( n91863 , n91809 );
or ( n91864 , n91862 , n91863 );
and ( n91865 , n87706 , n90576 );
not ( n91866 , n87706 );
and ( n91867 , n91866 , n90577 );
nor ( n91868 , n91865 , n91867 );
nand ( n91869 , n91868 , n87702 );
nand ( n91870 , n91864 , n91869 );
not ( n91871 , n91573 );
and ( n91872 , n91871 , n91583 , n91736 );
not ( n91873 , n91872 );
not ( n91874 , n91871 );
nand ( n91875 , n91874 , n91740 );
nand ( n91876 , n91584 , n91573 , n91736 );
not ( n91877 , n91583 );
nand ( n91878 , n91877 , n91871 , n91735 );
nand ( n91879 , n91873 , n91875 , n91876 , n91878 );
xor ( n91880 , n91870 , n91879 );
not ( n91881 , n90324 );
not ( n91882 , n91681 );
or ( n91883 , n91881 , n91882 );
and ( n91884 , n90286 , n91401 );
not ( n91885 , n90286 );
and ( n91886 , n91885 , n90946 );
nor ( n91887 , n91884 , n91886 );
nand ( n91888 , n91887 , n90279 );
nand ( n91889 , n91883 , n91888 );
xor ( n91890 , n91598 , n91611 );
xor ( n91891 , n91890 , n91661 );
and ( n91892 , n91889 , n91891 );
not ( n91893 , n90610 );
not ( n91894 , n91698 );
or ( n91895 , n91893 , n91894 );
and ( n91896 , n90612 , n90721 );
not ( n91897 , n90612 );
and ( n91898 , n91897 , n90991 );
nor ( n91899 , n91896 , n91898 );
nand ( n91900 , n91899 , n90656 );
nand ( n91901 , n91895 , n91900 );
xor ( n91902 , n91598 , n91611 );
xor ( n91903 , n91902 , n91661 );
and ( n91904 , n91901 , n91903 );
and ( n91905 , n91889 , n91901 );
or ( n91906 , n91892 , n91904 , n91905 );
not ( n91907 , n90697 );
not ( n91908 , n91715 );
or ( n91909 , n91907 , n91908 );
and ( n91910 , n90660 , n90430 );
not ( n91911 , n90660 );
and ( n91912 , n91911 , n90429 );
nor ( n91913 , n91910 , n91912 );
nand ( n91914 , n91913 , n90680 );
nand ( n91915 , n91909 , n91914 );
xor ( n91916 , n91906 , n91915 );
not ( n91917 , n90582 );
not ( n91918 , n91723 );
or ( n91919 , n91917 , n91918 );
and ( n91920 , n90540 , n90471 );
not ( n91921 , n90540 );
not ( n91922 , n90456 );
not ( n91923 , n90459 );
or ( n91924 , n91922 , n91923 );
nand ( n91925 , n91924 , n90463 );
and ( n91926 , n91921 , n91925 );
nor ( n91927 , n91920 , n91926 );
nand ( n91928 , n91927 , n90537 );
nand ( n91929 , n91919 , n91928 );
and ( n91930 , n91916 , n91929 );
and ( n91931 , n91906 , n91915 );
or ( n91932 , n91930 , n91931 );
not ( n91933 , n91932 );
not ( n91934 , n90782 );
not ( n91935 , n91825 );
or ( n91936 , n91934 , n91935 );
not ( n91937 , n90788 );
not ( n91938 , n90672 );
or ( n91939 , n91937 , n91938 );
nand ( n91940 , n90801 , n90669 );
nand ( n91941 , n91939 , n91940 );
nand ( n91942 , n91941 , n90825 );
nand ( n91943 , n91936 , n91942 );
not ( n91944 , n91943 );
or ( n91945 , n91933 , n91944 );
or ( n91946 , n91943 , n91932 );
xor ( n91947 , n91664 , n91684 );
xor ( n91948 , n91947 , n91700 );
xor ( n91949 , n91615 , n91627 );
xor ( n91950 , n91949 , n91658 );
not ( n91951 , n90324 );
not ( n91952 , n91887 );
or ( n91953 , n91951 , n91952 );
nand ( n91954 , n91390 , n90321 );
not ( n91955 , n91298 );
nand ( n91956 , n91955 , n90286 );
nand ( n91957 , n91954 , n91956 );
nand ( n91958 , n91957 , n90279 );
nand ( n91959 , n91953 , n91958 );
xor ( n91960 , n91950 , n91959 );
xor ( n91961 , n91629 , n91639 );
xor ( n91962 , n91961 , n91655 );
not ( n91963 , n90248 );
not ( n91964 , n91957 );
or ( n91965 , n91963 , n91964 );
and ( n91966 , n90286 , n91394 );
not ( n91967 , n90286 );
and ( n91968 , n91967 , n91395 );
nor ( n91969 , n91966 , n91968 );
nand ( n91970 , n91969 , n90279 );
nand ( n91971 , n91965 , n91970 );
xor ( n91972 , n91962 , n91971 );
xor ( n91973 , n91646 , n91654 );
not ( n91974 , n90248 );
not ( n91975 , n91969 );
or ( n91976 , n91974 , n91975 );
not ( n91977 , n90286 );
not ( n91978 , n91622 );
not ( n91979 , n91978 );
or ( n91980 , n91977 , n91979 );
nand ( n91981 , n91589 , n90321 );
nand ( n91982 , n91980 , n91981 );
nand ( n91983 , n91982 , n90279 );
nand ( n91984 , n91976 , n91983 );
xor ( n91985 , n91973 , n91984 );
nor ( n91986 , n90404 , n89865 );
not ( n91987 , n90248 );
not ( n91988 , n91982 );
or ( n91989 , n91987 , n91988 );
not ( n91990 , n90286 );
not ( n91991 , n91595 );
not ( n91992 , n91991 );
or ( n91993 , n91990 , n91992 );
not ( n91994 , n91991 );
nand ( n91995 , n91994 , n90321 );
nand ( n91996 , n91993 , n91995 );
nand ( n91997 , n91996 , n90279 );
nand ( n91998 , n91989 , n91997 );
xor ( n91999 , n91986 , n91998 );
and ( n92000 , n90230 , n91641 );
and ( n92001 , n90231 , n89865 );
nor ( n92002 , n92001 , n90630 );
nor ( n92003 , n92000 , n92002 , n90321 );
not ( n92004 , n90248 );
not ( n92005 , n91996 );
or ( n92006 , n92004 , n92005 );
or ( n92007 , n90286 , n89865 );
or ( n92008 , n90321 , n91641 );
nand ( n92009 , n92007 , n92008 );
nand ( n92010 , n90279 , n92009 );
nand ( n92011 , n92006 , n92010 );
and ( n92012 , n92003 , n92011 );
and ( n92013 , n91999 , n92012 );
and ( n92014 , n91986 , n91998 );
or ( n92015 , n92013 , n92014 );
and ( n92016 , n91985 , n92015 );
and ( n92017 , n91973 , n91984 );
or ( n92018 , n92016 , n92017 );
and ( n92019 , n91972 , n92018 );
and ( n92020 , n91962 , n91971 );
or ( n92021 , n92019 , n92020 );
and ( n92022 , n91960 , n92021 );
and ( n92023 , n91950 , n91959 );
or ( n92024 , n92022 , n92023 );
not ( n92025 , n90697 );
not ( n92026 , n91913 );
or ( n92027 , n92025 , n92026 );
and ( n92028 , n90380 , n90660 );
not ( n92029 , n90380 );
and ( n92030 , n92029 , n91164 );
nor ( n92031 , n92028 , n92030 );
nand ( n92032 , n92031 , n90680 );
nand ( n92033 , n92027 , n92032 );
xor ( n92034 , n92024 , n92033 );
xor ( n92035 , n91598 , n91611 );
xor ( n92036 , n92035 , n91661 );
xor ( n92037 , n91889 , n91901 );
xor ( n92038 , n92036 , n92037 );
and ( n92039 , n92034 , n92038 );
and ( n92040 , n92024 , n92033 );
or ( n92041 , n92039 , n92040 );
xor ( n92042 , n91948 , n92041 );
not ( n92043 , n90876 );
not ( n92044 , n91839 );
or ( n92045 , n92043 , n92044 );
and ( n92046 , n90842 , n90765 );
not ( n92047 , n90842 );
and ( n92048 , n92047 , n90318 );
nor ( n92049 , n92046 , n92048 );
nand ( n92050 , n92049 , n90839 );
nand ( n92051 , n92045 , n92050 );
and ( n92052 , n92042 , n92051 );
and ( n92053 , n91948 , n92041 );
or ( n92054 , n92052 , n92053 );
nand ( n92055 , n91946 , n92054 );
nand ( n92056 , n91945 , n92055 );
and ( n92057 , n91880 , n92056 );
and ( n92058 , n91870 , n91879 );
or ( n92059 , n92057 , n92058 );
xor ( n92060 , n91776 , n91745 );
xnor ( n92061 , n92060 , n91742 );
xor ( n92062 , n92059 , n92061 );
xor ( n92063 , n91811 , n91813 );
xor ( n92064 , n92063 , n91849 );
and ( n92065 , n92062 , n92064 );
and ( n92066 , n92059 , n92061 );
or ( n92067 , n92065 , n92066 );
nor ( n92068 , n91861 , n92067 );
nor ( n92069 , n91859 , n92068 );
not ( n92070 , n92069 );
xor ( n92071 , n92059 , n92061 );
xor ( n92072 , n92071 , n92064 );
xor ( n92073 , n91870 , n91879 );
xor ( n92074 , n92073 , n92056 );
xor ( n92075 , n91816 , n91827 );
xnor ( n92076 , n92075 , n91847 );
not ( n92077 , n92076 );
or ( n92078 , n92074 , n92077 );
not ( n92079 , n87702 );
not ( n92080 , n87706 );
not ( n92081 , n90552 );
or ( n92082 , n92080 , n92081 );
nand ( n92083 , n90555 , n87705 );
nand ( n92084 , n92082 , n92083 );
not ( n92085 , n92084 );
or ( n92086 , n92079 , n92085 );
nand ( n92087 , n91868 , n87689 );
nand ( n92088 , n92086 , n92087 );
not ( n92089 , n92088 );
xor ( n92090 , n91832 , n91841 );
xor ( n92091 , n92090 , n91844 );
not ( n92092 , n92091 );
or ( n92093 , n92089 , n92092 );
or ( n92094 , n92088 , n92091 );
xor ( n92095 , n91906 , n91915 );
xor ( n92096 , n92095 , n91929 );
not ( n92097 , n90782 );
not ( n92098 , n91941 );
or ( n92099 , n92097 , n92098 );
and ( n92100 , n90788 , n90622 );
not ( n92101 , n90788 );
and ( n92102 , n92101 , n90623 );
nor ( n92103 , n92100 , n92102 );
nand ( n92104 , n92103 , n90825 );
nand ( n92105 , n92099 , n92104 );
xor ( n92106 , n92096 , n92105 );
not ( n92107 , n90582 );
not ( n92108 , n91927 );
or ( n92109 , n92107 , n92108 );
and ( n92110 , n90540 , n90418 );
not ( n92111 , n90540 );
and ( n92112 , n92111 , n90419 );
nor ( n92113 , n92110 , n92112 );
nand ( n92114 , n92113 , n90537 );
nand ( n92115 , n92109 , n92114 );
not ( n92116 , n90610 );
not ( n92117 , n91899 );
or ( n92118 , n92116 , n92117 );
and ( n92119 , n90612 , n90989 );
not ( n92120 , n90612 );
and ( n92121 , n92120 , n90934 );
nor ( n92122 , n92119 , n92121 );
not ( n92123 , n92122 );
nand ( n92124 , n92123 , n90656 );
nand ( n92125 , n92118 , n92124 );
xor ( n92126 , n91950 , n91959 );
xor ( n92127 , n92126 , n92021 );
xor ( n92128 , n92125 , n92127 );
not ( n92129 , n90680 );
and ( n92130 , n90660 , n90724 );
not ( n92131 , n90660 );
and ( n92132 , n92131 , n90386 );
nor ( n92133 , n92130 , n92132 );
not ( n92134 , n92133 );
or ( n92135 , n92129 , n92134 );
nand ( n92136 , n90697 , n92031 );
nand ( n92137 , n92135 , n92136 );
and ( n92138 , n92128 , n92137 );
and ( n92139 , n92125 , n92127 );
or ( n92140 , n92138 , n92139 );
xor ( n92141 , n92115 , n92140 );
not ( n92142 , n90876 );
not ( n92143 , n92049 );
or ( n92144 , n92142 , n92143 );
not ( n92145 , n90842 );
not ( n92146 , n90300 );
or ( n92147 , n92145 , n92146 );
nand ( n92148 , n90297 , n90843 );
nand ( n92149 , n92147 , n92148 );
nand ( n92150 , n92149 , n90839 );
nand ( n92151 , n92144 , n92150 );
and ( n92152 , n92141 , n92151 );
and ( n92153 , n92115 , n92140 );
or ( n92154 , n92152 , n92153 );
and ( n92155 , n92106 , n92154 );
and ( n92156 , n92096 , n92105 );
or ( n92157 , n92155 , n92156 );
nand ( n92158 , n92094 , n92157 );
nand ( n92159 , n92093 , n92158 );
nand ( n92160 , n92078 , n92159 );
nand ( n92161 , n92074 , n92077 );
nand ( n92162 , n92160 , n92161 );
xor ( n92163 , n92072 , n92162 );
xor ( n92164 , n91943 , n91932 );
xnor ( n92165 , n92164 , n92054 );
xor ( n92166 , n92024 , n92033 );
xor ( n92167 , n92166 , n92038 );
not ( n92168 , n92167 );
not ( n92169 , n90782 );
not ( n92170 , n92103 );
or ( n92171 , n92169 , n92170 );
and ( n92172 , n90646 , n90788 );
not ( n92173 , n90646 );
and ( n92174 , n92173 , n90799 );
nor ( n92175 , n92172 , n92174 );
nand ( n92176 , n92175 , n90825 );
nand ( n92177 , n92171 , n92176 );
not ( n92178 , n92177 );
or ( n92179 , n92168 , n92178 );
not ( n92180 , n92167 );
not ( n92181 , n92180 );
not ( n92182 , n92177 );
not ( n92183 , n92182 );
or ( n92184 , n92181 , n92183 );
not ( n92185 , n90657 );
not ( n92186 , n90612 );
not ( n92187 , n91401 );
not ( n92188 , n92187 );
or ( n92189 , n92186 , n92188 );
or ( n92190 , n92187 , n90612 );
nand ( n92191 , n92189 , n92190 );
not ( n92192 , n92191 );
or ( n92193 , n92185 , n92192 );
or ( n92194 , n92122 , n90609 );
nand ( n92195 , n92193 , n92194 );
xor ( n92196 , n91962 , n91971 );
xor ( n92197 , n92196 , n92018 );
xor ( n92198 , n92195 , n92197 );
not ( n92199 , n90697 );
not ( n92200 , n92133 );
or ( n92201 , n92199 , n92200 );
and ( n92202 , n90660 , n90991 );
not ( n92203 , n90660 );
and ( n92204 , n92203 , n90721 );
nor ( n92205 , n92202 , n92204 );
not ( n92206 , n92205 );
nand ( n92207 , n92206 , n90680 );
nand ( n92208 , n92201 , n92207 );
and ( n92209 , n92198 , n92208 );
and ( n92210 , n92195 , n92197 );
or ( n92211 , n92209 , n92210 );
not ( n92212 , n90582 );
not ( n92213 , n92113 );
or ( n92214 , n92212 , n92213 );
and ( n92215 , n90540 , n90430 );
not ( n92216 , n90540 );
and ( n92217 , n92216 , n90429 );
nor ( n92218 , n92215 , n92217 );
nand ( n92219 , n92218 , n90537 );
nand ( n92220 , n92214 , n92219 );
xor ( n92221 , n92211 , n92220 );
xor ( n92222 , n92125 , n92127 );
xor ( n92223 , n92222 , n92137 );
and ( n92224 , n92221 , n92223 );
and ( n92225 , n92211 , n92220 );
or ( n92226 , n92224 , n92225 );
nand ( n92227 , n92184 , n92226 );
nand ( n92228 , n92179 , n92227 );
xor ( n92229 , n91948 , n92041 );
xor ( n92230 , n92229 , n92051 );
xor ( n92231 , n92228 , n92230 );
not ( n92232 , n87702 );
not ( n92233 , n87706 );
not ( n92234 , n90693 );
or ( n92235 , n92233 , n92234 );
nand ( n92236 , n90690 , n87705 );
nand ( n92237 , n92235 , n92236 );
not ( n92238 , n92237 );
or ( n92239 , n92232 , n92238 );
nand ( n92240 , n92084 , n87689 );
nand ( n92241 , n92239 , n92240 );
and ( n92242 , n92231 , n92241 );
and ( n92243 , n92228 , n92230 );
or ( n92244 , n92242 , n92243 );
not ( n92245 , n92244 );
xor ( n92246 , n92165 , n92245 );
xor ( n92247 , n92088 , n92091 );
xnor ( n92248 , n92247 , n92157 );
xor ( n92249 , n92246 , n92248 );
xor ( n92250 , n92096 , n92105 );
xor ( n92251 , n92250 , n92154 );
not ( n92252 , n87689 );
not ( n92253 , n92237 );
or ( n92254 , n92252 , n92253 );
not ( n92255 , n87706 );
not ( n92256 , n90672 );
or ( n92257 , n92255 , n92256 );
nand ( n92258 , n90669 , n87705 );
nand ( n92259 , n92257 , n92258 );
nand ( n92260 , n92259 , n87702 );
nand ( n92261 , n92254 , n92260 );
xor ( n92262 , n92115 , n92140 );
xor ( n92263 , n92262 , n92151 );
xor ( n92264 , n92261 , n92263 );
not ( n92265 , n90876 );
not ( n92266 , n92149 );
or ( n92267 , n92265 , n92266 );
not ( n92268 , n90842 );
not ( n92269 , n90464 );
or ( n92270 , n92268 , n92269 );
nand ( n92271 , n90471 , n90843 );
nand ( n92272 , n92270 , n92271 );
nand ( n92273 , n92272 , n90839 );
nand ( n92274 , n92267 , n92273 );
not ( n92275 , n92274 );
not ( n92276 , n90782 );
not ( n92277 , n92175 );
or ( n92278 , n92276 , n92277 );
and ( n92279 , n90788 , n90765 );
not ( n92280 , n90788 );
and ( n92281 , n92280 , n90318 );
nor ( n92282 , n92279 , n92281 );
nand ( n92283 , n92282 , n90825 );
nand ( n92284 , n92278 , n92283 );
not ( n92285 , n92284 );
or ( n92286 , n92275 , n92285 );
or ( n92287 , n92284 , n92274 );
not ( n92288 , n90582 );
not ( n92289 , n92218 );
or ( n92290 , n92288 , n92289 );
not ( n92291 , n90540 );
not ( n92292 , n90379 );
or ( n92293 , n92291 , n92292 );
nand ( n92294 , n90380 , n90539 );
nand ( n92295 , n92293 , n92294 );
nand ( n92296 , n92295 , n90537 );
nand ( n92297 , n92290 , n92296 );
xor ( n92298 , n91973 , n91984 );
xor ( n92299 , n92298 , n92015 );
not ( n92300 , n92299 );
not ( n92301 , n90610 );
not ( n92302 , n92191 );
or ( n92303 , n92301 , n92302 );
and ( n92304 , n90612 , n91390 );
not ( n92305 , n90612 );
and ( n92306 , n92305 , n91955 );
nor ( n92307 , n92304 , n92306 );
nand ( n92308 , n92307 , n90656 );
nand ( n92309 , n92303 , n92308 );
not ( n92310 , n92309 );
or ( n92311 , n92300 , n92310 );
or ( n92312 , n92309 , n92299 );
xor ( n92313 , n91986 , n91998 );
xor ( n92314 , n92313 , n92012 );
not ( n92315 , n90610 );
not ( n92316 , n92307 );
or ( n92317 , n92315 , n92316 );
and ( n92318 , n90612 , n91394 );
not ( n92319 , n90612 );
and ( n92320 , n92319 , n91395 );
nor ( n92321 , n92318 , n92320 );
nand ( n92322 , n92321 , n90656 );
nand ( n92323 , n92317 , n92322 );
xor ( n92324 , n92314 , n92323 );
xor ( n92325 , n92003 , n92011 );
not ( n92326 , n90610 );
not ( n92327 , n92321 );
or ( n92328 , n92326 , n92327 );
and ( n92329 , n90612 , n91622 );
not ( n92330 , n90612 );
and ( n92331 , n92330 , n91978 );
nor ( n92332 , n92329 , n92331 );
nand ( n92333 , n92332 , n90656 );
nand ( n92334 , n92328 , n92333 );
xor ( n92335 , n92325 , n92334 );
and ( n92336 , n90248 , n91641 );
not ( n92337 , n90610 );
and ( n92338 , n90246 , n91596 );
not ( n92339 , n90246 );
and ( n92340 , n92339 , n91595 );
nor ( n92341 , n92338 , n92340 );
not ( n92342 , n92341 );
or ( n92343 , n92337 , n92342 );
and ( n92344 , n90246 , n91641 );
and ( n92345 , n90243 , n89865 );
nor ( n92346 , n92344 , n92345 );
not ( n92347 , n92346 );
nand ( n92348 , n92347 , n90656 );
nand ( n92349 , n92343 , n92348 );
not ( n92350 , n90592 );
and ( n92351 , n92350 , n91641 );
nor ( n92352 , n92351 , n90630 );
or ( n92353 , n91641 , n92350 );
nand ( n92354 , n92353 , n90660 );
and ( n92355 , n92352 , n92354 );
and ( n92356 , n92349 , n92355 );
xor ( n92357 , n92336 , n92356 );
not ( n92358 , n90610 );
not ( n92359 , n92332 );
or ( n92360 , n92358 , n92359 );
nand ( n92361 , n92341 , n90656 );
nand ( n92362 , n92360 , n92361 );
and ( n92363 , n92357 , n92362 );
or ( n92364 , n92363 , C0 );
and ( n92365 , n92335 , n92364 );
and ( n92366 , n92325 , n92334 );
or ( n92367 , n92365 , n92366 );
and ( n92368 , n92324 , n92367 );
and ( n92369 , n92314 , n92323 );
or ( n92370 , n92368 , n92369 );
nand ( n92371 , n92312 , n92370 );
nand ( n92372 , n92311 , n92371 );
or ( n92373 , n92297 , n92372 );
xor ( n92374 , n92195 , n92197 );
xor ( n92375 , n92374 , n92208 );
and ( n92376 , n92373 , n92375 );
and ( n92377 , n92372 , n92297 );
nor ( n92378 , n92376 , n92377 );
not ( n92379 , n92378 );
nand ( n92380 , n92287 , n92379 );
nand ( n92381 , n92286 , n92380 );
and ( n92382 , n92264 , n92381 );
and ( n92383 , n92261 , n92263 );
or ( n92384 , n92382 , n92383 );
xor ( n92385 , n92251 , n92384 );
xor ( n92386 , n92228 , n92230 );
xor ( n92387 , n92386 , n92241 );
and ( n92388 , n92385 , n92387 );
and ( n92389 , n92251 , n92384 );
nor ( n92390 , n92388 , n92389 );
and ( n92391 , n92249 , n92390 );
xnor ( n92392 , n92159 , n92076 );
not ( n92393 , n92074 );
and ( n92394 , n92392 , n92393 );
not ( n92395 , n92392 );
and ( n92396 , n92395 , n92074 );
nor ( n92397 , n92394 , n92396 );
xor ( n92398 , n92165 , n92245 );
and ( n92399 , n92398 , n92248 );
and ( n92400 , n92165 , n92245 );
or ( n92401 , n92399 , n92400 );
and ( n92402 , n92397 , n92401 );
nor ( n92403 , n92391 , n92402 );
not ( n92404 , n92403 );
xor ( n92405 , n92261 , n92263 );
xor ( n92406 , n92405 , n92381 );
not ( n92407 , n92406 );
xor ( n92408 , n92211 , n92220 );
xor ( n92409 , n92408 , n92223 );
not ( n92410 , n92409 );
not ( n92411 , n92205 );
not ( n92412 , n91010 );
and ( n92413 , n92411 , n92412 );
not ( n92414 , n90660 );
not ( n92415 , n90989 );
or ( n92416 , n92414 , n92415 );
nand ( n92417 , n90934 , n91164 );
nand ( n92418 , n92416 , n92417 );
and ( n92419 , n92418 , n90680 );
nor ( n92420 , n92413 , n92419 );
not ( n92421 , n92420 );
not ( n92422 , n92421 );
xor ( n92423 , n92309 , n92299 );
xnor ( n92424 , n92423 , n92370 );
not ( n92425 , n92424 );
not ( n92426 , n92425 );
or ( n92427 , n92422 , n92426 );
and ( n92428 , n92295 , n90582 );
and ( n92429 , n90540 , n90386 );
not ( n92430 , n90540 );
and ( n92431 , n92430 , n90724 );
or ( n92432 , n92429 , n92431 );
and ( n92433 , n92432 , n90537 );
nor ( n92434 , n92428 , n92433 );
nand ( n92435 , n92427 , n92434 );
nand ( n92436 , n92424 , n92420 );
nand ( n92437 , n92435 , n92436 );
not ( n92438 , n92437 );
and ( n92439 , n90843 , n90418 );
not ( n92440 , n90843 );
and ( n92441 , n92440 , n90419 );
nor ( n92442 , n92439 , n92441 );
not ( n92443 , n92442 );
not ( n92444 , n90839 );
not ( n92445 , n92444 );
and ( n92446 , n92443 , n92445 );
and ( n92447 , n92272 , n90876 );
nor ( n92448 , n92446 , n92447 );
not ( n92449 , n92448 );
or ( n92450 , n92438 , n92449 );
xor ( n92451 , n92372 , n92297 );
xor ( n92452 , n92451 , n92375 );
nand ( n92453 , n92450 , n92452 );
not ( n92454 , n92448 );
not ( n92455 , n92437 );
nand ( n92456 , n92454 , n92455 );
and ( n92457 , n92453 , n92456 );
not ( n92458 , n92457 );
not ( n92459 , n92458 );
or ( n92460 , n92410 , n92459 );
not ( n92461 , n92409 );
not ( n92462 , n92461 );
not ( n92463 , n92457 );
or ( n92464 , n92462 , n92463 );
and ( n92465 , n87706 , n90629 );
not ( n92466 , n87706 );
and ( n92467 , n92466 , n90623 );
nor ( n92468 , n92465 , n92467 );
not ( n92469 , n92468 );
not ( n92470 , n87702 );
or ( n92471 , n92469 , n92470 );
not ( n92472 , n87689 );
not ( n92473 , n92472 );
nand ( n92474 , n92473 , n92259 );
nand ( n92475 , n92471 , n92474 );
nand ( n92476 , n92464 , n92475 );
nand ( n92477 , n92460 , n92476 );
not ( n92478 , n92477 );
and ( n92479 , n92177 , n92180 );
not ( n92480 , n92177 );
and ( n92481 , n92480 , n92167 );
or ( n92482 , n92479 , n92481 );
not ( n92483 , n92226 );
and ( n92484 , n92482 , n92483 );
not ( n92485 , n92482 );
and ( n92486 , n92485 , n92226 );
nor ( n92487 , n92484 , n92486 );
nand ( n92488 , n92478 , n92487 );
not ( n92489 , n92488 );
or ( n92490 , n92407 , n92489 );
not ( n92491 , n92487 );
nand ( n92492 , n92477 , n92491 );
nand ( n92493 , n92490 , n92492 );
xor ( n92494 , n92251 , n92384 );
xor ( n92495 , n92494 , n92387 );
xor ( n92496 , n92493 , n92495 );
not ( n92497 , n90537 );
not ( n92498 , n90539 );
and ( n92499 , n92498 , n90934 );
not ( n92500 , n92498 );
and ( n92501 , n92500 , n90989 );
nor ( n92502 , n92499 , n92501 );
not ( n92503 , n92502 );
or ( n92504 , n92497 , n92503 );
and ( n92505 , n90539 , n90721 );
not ( n92506 , n90539 );
and ( n92507 , n92506 , n90991 );
nor ( n92508 , n92505 , n92507 );
not ( n92509 , n90582 );
or ( n92510 , n92508 , n92509 );
nand ( n92511 , n92504 , n92510 );
xor ( n92512 , n92325 , n92334 );
xor ( n92513 , n92512 , n92364 );
not ( n92514 , n90697 );
and ( n92515 , n90660 , n90945 );
not ( n92516 , n90660 );
and ( n92517 , n92516 , n92187 );
nor ( n92518 , n92515 , n92517 );
not ( n92519 , n92518 );
or ( n92520 , n92514 , n92519 );
and ( n92521 , n90660 , n91390 );
not ( n92522 , n90660 );
and ( n92523 , n92522 , n91299 );
nor ( n92524 , n92521 , n92523 );
nand ( n92525 , n92524 , n90680 );
nand ( n92526 , n92520 , n92525 );
xor ( n92527 , n92513 , n92526 );
xor ( n92528 , n92336 , n92356 );
xor ( n92529 , n92528 , n92362 );
not ( n92530 , n90697 );
not ( n92531 , n92524 );
or ( n92532 , n92530 , n92531 );
and ( n92533 , n90660 , n91394 );
not ( n92534 , n90660 );
and ( n92535 , n92534 , n91395 );
nor ( n92536 , n92533 , n92535 );
nand ( n92537 , n92536 , n90680 );
nand ( n92538 , n92532 , n92537 );
xor ( n92539 , n92529 , n92538 );
xor ( n92540 , n92349 , n92355 );
not ( n92541 , n90697 );
not ( n92542 , n92536 );
or ( n92543 , n92541 , n92542 );
and ( n92544 , n90660 , n91622 );
not ( n92545 , n90660 );
and ( n92546 , n92545 , n91588 );
nor ( n92547 , n92544 , n92546 );
nand ( n92548 , n92547 , n90680 );
nand ( n92549 , n92543 , n92548 );
xor ( n92550 , n92540 , n92549 );
and ( n92551 , n90610 , n91641 );
not ( n92552 , n90697 );
not ( n92553 , n92547 );
or ( n92554 , n92552 , n92553 );
and ( n92555 , n90660 , n91994 );
not ( n92556 , n90660 );
and ( n92557 , n92556 , n91991 );
nor ( n92558 , n92555 , n92557 );
nand ( n92559 , n92558 , n90680 );
nand ( n92560 , n92554 , n92559 );
xor ( n92561 , n92551 , n92560 );
or ( n92562 , n90677 , n91641 );
nand ( n92563 , n92562 , n92498 );
nand ( n92564 , n90677 , n91641 );
and ( n92565 , n92563 , n90660 , n92564 );
not ( n92566 , n90697 );
not ( n92567 , n92558 );
or ( n92568 , n92566 , n92567 );
or ( n92569 , n90660 , n89865 );
or ( n92570 , n91164 , n91641 );
nand ( n92571 , n92569 , n92570 );
nand ( n92572 , n90680 , n92571 );
nand ( n92573 , n92568 , n92572 );
and ( n92574 , n92565 , n92573 );
and ( n92575 , n92561 , n92574 );
and ( n92576 , n92551 , n92560 );
or ( n92577 , n92575 , n92576 );
and ( n92578 , n92550 , n92577 );
and ( n92579 , n92540 , n92549 );
or ( n92580 , n92578 , n92579 );
and ( n92581 , n92539 , n92580 );
and ( n92582 , n92529 , n92538 );
or ( n92583 , n92581 , n92582 );
xor ( n92584 , n92527 , n92583 );
xor ( n92585 , n92511 , n92584 );
not ( n92586 , n90839 );
and ( n92587 , n90842 , n90724 );
not ( n92588 , n90842 );
and ( n92589 , n92588 , n90386 );
nor ( n92590 , n92587 , n92589 );
not ( n92591 , n92590 );
or ( n92592 , n92586 , n92591 );
not ( n92593 , n90842 );
not ( n92594 , n90379 );
or ( n92595 , n92593 , n92594 );
nand ( n92596 , n90380 , n90843 );
nand ( n92597 , n92595 , n92596 );
nand ( n92598 , n92597 , n90876 );
nand ( n92599 , n92592 , n92598 );
and ( n92600 , n92585 , n92599 );
and ( n92601 , n92511 , n92584 );
or ( n92602 , n92600 , n92601 );
not ( n92603 , n90782 );
not ( n92604 , n91925 );
and ( n92605 , n92604 , n90788 );
not ( n92606 , n92604 );
and ( n92607 , n92606 , n90801 );
nor ( n92608 , n92605 , n92607 );
not ( n92609 , n92608 );
or ( n92610 , n92603 , n92609 );
and ( n92611 , n90417 , n90799 );
not ( n92612 , n90417 );
and ( n92613 , n92612 , n90788 );
or ( n92614 , n92611 , n92613 );
nand ( n92615 , n92614 , n90825 );
nand ( n92616 , n92610 , n92615 );
xor ( n92617 , n92602 , n92616 );
and ( n92618 , n87705 , n90318 );
not ( n92619 , n87705 );
and ( n92620 , n92619 , n90317 );
nor ( n92621 , n92618 , n92620 );
not ( n92622 , n92621 );
not ( n92623 , n87689 );
or ( n92624 , n92622 , n92623 );
and ( n92625 , n87706 , n90297 );
not ( n92626 , n87706 );
and ( n92627 , n92626 , n90300 );
nor ( n92628 , n92625 , n92627 );
nand ( n92629 , n92628 , n87702 );
nand ( n92630 , n92624 , n92629 );
and ( n92631 , n92617 , n92630 );
and ( n92632 , n92602 , n92616 );
or ( n92633 , n92631 , n92632 );
xor ( n92634 , n92314 , n92323 );
xor ( n92635 , n92634 , n92367 );
not ( n92636 , n90697 );
not ( n92637 , n92418 );
or ( n92638 , n92636 , n92637 );
nand ( n92639 , n92518 , n90680 );
nand ( n92640 , n92638 , n92639 );
xor ( n92641 , n92635 , n92640 );
not ( n92642 , n90582 );
not ( n92643 , n92432 );
or ( n92644 , n92642 , n92643 );
not ( n92645 , n92508 );
nand ( n92646 , n92645 , n90537 );
nand ( n92647 , n92644 , n92646 );
and ( n92648 , n92641 , n92647 );
and ( n92649 , n92635 , n92640 );
or ( n92650 , n92648 , n92649 );
not ( n92651 , n90876 );
not ( n92652 , n92442 );
not ( n92653 , n92652 );
or ( n92654 , n92651 , n92653 );
and ( n92655 , n90842 , n90430 );
not ( n92656 , n90842 );
and ( n92657 , n92656 , n90429 );
or ( n92658 , n92655 , n92657 );
not ( n92659 , n92658 );
nand ( n92660 , n92659 , n90839 );
nand ( n92661 , n92654 , n92660 );
xor ( n92662 , n92650 , n92661 );
not ( n92663 , n90782 );
not ( n92664 , n90788 );
not ( n92665 , n90300 );
or ( n92666 , n92664 , n92665 );
nand ( n92667 , n90297 , n90801 );
nand ( n92668 , n92666 , n92667 );
not ( n92669 , n92668 );
or ( n92670 , n92663 , n92669 );
nand ( n92671 , n92608 , n90825 );
nand ( n92672 , n92670 , n92671 );
xor ( n92673 , n92662 , n92672 );
xor ( n92674 , n92633 , n92673 );
xor ( n92675 , n92420 , n92425 );
xnor ( n92676 , n92675 , n92434 );
xor ( n92677 , n92513 , n92526 );
and ( n92678 , n92677 , n92583 );
and ( n92679 , n92513 , n92526 );
or ( n92680 , n92678 , n92679 );
not ( n92681 , n92597 );
not ( n92682 , n90839 );
or ( n92683 , n92681 , n92682 );
or ( n92684 , n92658 , n90838 );
nand ( n92685 , n92683 , n92684 );
xor ( n92686 , n92680 , n92685 );
xor ( n92687 , n92635 , n92640 );
xor ( n92688 , n92687 , n92647 );
and ( n92689 , n92686 , n92688 );
and ( n92690 , n92680 , n92685 );
or ( n92691 , n92689 , n92690 );
xor ( n92692 , n92676 , n92691 );
xor ( n92693 , n87706 , n90636 );
xor ( n92694 , n92693 , n90643 );
not ( n92695 , n92694 );
not ( n92696 , n87689 );
or ( n92697 , n92695 , n92696 );
nand ( n92698 , n92621 , n87702 );
nand ( n92699 , n92697 , n92698 );
not ( n92700 , n92699 );
and ( n92701 , n92692 , n92700 );
not ( n92702 , n92692 );
and ( n92703 , n92702 , n92699 );
nor ( n92704 , n92701 , n92703 );
and ( n92705 , n92674 , n92704 );
and ( n92706 , n92633 , n92673 );
or ( n92707 , n92705 , n92706 );
not ( n92708 , n92707 );
xor ( n92709 , n92454 , n92455 );
xnor ( n92710 , n92709 , n92452 );
not ( n92711 , n92676 );
not ( n92712 , n92700 );
or ( n92713 , n92711 , n92712 );
nand ( n92714 , n92713 , n92691 );
not ( n92715 , n92676 );
nand ( n92716 , n92715 , n92699 );
and ( n92717 , n92714 , n92716 );
xor ( n92718 , n92710 , n92717 );
not ( n92719 , n90782 );
not ( n92720 , n92282 );
or ( n92721 , n92719 , n92720 );
nand ( n92722 , n92668 , n90825 );
nand ( n92723 , n92721 , n92722 );
not ( n92724 , n87689 );
not ( n92725 , n92468 );
or ( n92726 , n92724 , n92725 );
nand ( n92727 , n92694 , n87702 );
nand ( n92728 , n92726 , n92727 );
xor ( n92729 , n92723 , n92728 );
xor ( n92730 , n92650 , n92661 );
and ( n92731 , n92730 , n92672 );
and ( n92732 , n92650 , n92661 );
or ( n92733 , n92731 , n92732 );
xnor ( n92734 , n92729 , n92733 );
xor ( n92735 , n92718 , n92734 );
nand ( n92736 , n92708 , n92735 );
not ( n92737 , n92736 );
xor ( n92738 , n92680 , n92685 );
xor ( n92739 , n92738 , n92688 );
not ( n92740 , n92739 );
xor ( n92741 , n92602 , n92616 );
xor ( n92742 , n92741 , n92630 );
not ( n92743 , n92742 );
or ( n92744 , n92740 , n92743 );
not ( n92745 , n92739 );
not ( n92746 , n92745 );
not ( n92747 , n92742 );
not ( n92748 , n92747 );
or ( n92749 , n92746 , n92748 );
not ( n92750 , n90782 );
not ( n92751 , n92614 );
or ( n92752 , n92750 , n92751 );
not ( n92753 , n90788 );
not ( n92754 , n90429 );
or ( n92755 , n92753 , n92754 );
nand ( n92756 , n90428 , n90799 );
nand ( n92757 , n92755 , n92756 );
nand ( n92758 , n92757 , n90825 );
nand ( n92759 , n92752 , n92758 );
not ( n92760 , n90582 );
not ( n92761 , n92502 );
or ( n92762 , n92760 , n92761 );
and ( n92763 , n92498 , n90945 );
not ( n92764 , n92498 );
and ( n92765 , n92764 , n90946 );
nor ( n92766 , n92763 , n92765 );
nand ( n92767 , n92766 , n90537 );
nand ( n92768 , n92762 , n92767 );
xor ( n92769 , n92529 , n92538 );
xor ( n92770 , n92769 , n92580 );
xor ( n92771 , n92768 , n92770 );
not ( n92772 , n90876 );
not ( n92773 , n92590 );
or ( n92774 , n92772 , n92773 );
and ( n92775 , n90842 , n90721 );
not ( n92776 , n90842 );
and ( n92777 , n92776 , n90991 );
nor ( n92778 , n92775 , n92777 );
nand ( n92779 , n92778 , n90839 );
nand ( n92780 , n92774 , n92779 );
and ( n92781 , n92771 , n92780 );
and ( n92782 , n92768 , n92770 );
or ( n92783 , n92781 , n92782 );
or ( n92784 , n92759 , n92783 );
not ( n92785 , n92784 );
xor ( n92786 , n92540 , n92549 );
xor ( n92787 , n92786 , n92577 );
not ( n92788 , n90582 );
not ( n92789 , n92766 );
or ( n92790 , n92788 , n92789 );
xor ( n92791 , n92498 , n91390 );
nand ( n92792 , n92791 , n90537 );
nand ( n92793 , n92790 , n92792 );
xor ( n92794 , n92787 , n92793 );
xor ( n92795 , n92551 , n92560 );
xor ( n92796 , n92795 , n92574 );
not ( n92797 , n90582 );
not ( n92798 , n92791 );
or ( n92799 , n92797 , n92798 );
not ( n92800 , n92498 );
not ( n92801 , n91395 );
or ( n92802 , n92800 , n92801 );
nand ( n92803 , n91394 , n90539 );
nand ( n92804 , n92802 , n92803 );
nand ( n92805 , n92804 , n90537 );
nand ( n92806 , n92799 , n92805 );
xor ( n92807 , n92796 , n92806 );
xor ( n92808 , n92565 , n92573 );
not ( n92809 , n90582 );
not ( n92810 , n92804 );
or ( n92811 , n92809 , n92810 );
and ( n92812 , n91587 , n90539 );
not ( n92813 , n91587 );
and ( n92814 , n92813 , n92498 );
or ( n92815 , n92812 , n92814 );
nand ( n92816 , n92815 , n90536 );
nand ( n92817 , n92811 , n92816 );
xor ( n92818 , n92808 , n92817 );
not ( n92819 , n90582 );
not ( n92820 , n92815 );
or ( n92821 , n92819 , n92820 );
not ( n92822 , n90539 );
not ( n92823 , n92822 );
not ( n92824 , n91596 );
or ( n92825 , n92823 , n92824 );
nand ( n92826 , n91595 , n90539 );
nand ( n92827 , n92825 , n92826 );
nand ( n92828 , n92827 , n90536 );
nand ( n92829 , n92821 , n92828 );
nand ( n92830 , n90696 , n91641 );
not ( n92831 , n92830 );
or ( n92832 , n92829 , n92831 );
not ( n92833 , n90535 );
not ( n92834 , n92827 );
or ( n92835 , n92833 , n92834 );
or ( n92836 , n92822 , n89865 );
or ( n92837 , n90539 , n91641 );
nand ( n92838 , n92836 , n92837 );
nand ( n92839 , n90536 , n92838 );
nand ( n92840 , n92835 , n92839 );
or ( n92841 , n90512 , n91641 );
nand ( n92842 , n92841 , n90842 );
nand ( n92843 , n90512 , n91641 );
and ( n92844 , n92842 , n92498 , n92843 );
nand ( n92845 , n92832 , n92840 , n92844 );
nand ( n92846 , n92829 , n92831 );
nand ( n92847 , n92845 , n92846 );
and ( n92848 , n92818 , n92847 );
and ( n92849 , n92808 , n92817 );
or ( n92850 , n92848 , n92849 );
and ( n92851 , n92807 , n92850 );
and ( n92852 , n92796 , n92806 );
or ( n92853 , n92851 , n92852 );
and ( n92854 , n92794 , n92853 );
and ( n92855 , n92787 , n92793 );
or ( n92856 , n92854 , n92855 );
not ( n92857 , n92856 );
not ( n92858 , n90782 );
not ( n92859 , n92757 );
or ( n92860 , n92858 , n92859 );
and ( n92861 , n90378 , n90788 );
not ( n92862 , n90378 );
and ( n92863 , n92862 , n90799 );
or ( n92864 , n92861 , n92863 );
nand ( n92865 , n92864 , n90825 );
nand ( n92866 , n92860 , n92865 );
not ( n92867 , n92866 );
nand ( n92868 , n92857 , n92867 );
not ( n92869 , n92868 );
xor ( n92870 , n92768 , n92770 );
xor ( n92871 , n92870 , n92780 );
not ( n92872 , n92871 );
or ( n92873 , n92869 , n92872 );
nand ( n92874 , n92866 , n92856 );
nand ( n92875 , n92873 , n92874 );
not ( n92876 , n92875 );
or ( n92877 , n92785 , n92876 );
nand ( n92878 , n92759 , n92783 );
nand ( n92879 , n92877 , n92878 );
nand ( n92880 , n92749 , n92879 );
nand ( n92881 , n92744 , n92880 );
xor ( n92882 , n92633 , n92673 );
xor ( n92883 , n92882 , n92704 );
xor ( n92884 , n92881 , n92883 );
xor ( n92885 , n92511 , n92584 );
xor ( n92886 , n92885 , n92599 );
not ( n92887 , n87689 );
not ( n92888 , n92628 );
or ( n92889 , n92887 , n92888 );
not ( n92890 , n91925 );
not ( n92891 , n87706 );
or ( n92892 , n92890 , n92891 );
nand ( n92893 , n92604 , n87705 );
nand ( n92894 , n92892 , n92893 );
nand ( n92895 , n92894 , n87702 );
nand ( n92896 , n92889 , n92895 );
xor ( n92897 , n92886 , n92896 );
not ( n92898 , n92875 );
not ( n92899 , n92783 );
not ( n92900 , n92759 );
or ( n92901 , n92899 , n92900 );
or ( n92902 , n92759 , n92783 );
nand ( n92903 , n92901 , n92902 );
not ( n92904 , n92903 );
or ( n92905 , n92898 , n92904 );
or ( n92906 , n92903 , n92875 );
nand ( n92907 , n92905 , n92906 );
and ( n92908 , n92897 , n92907 );
and ( n92909 , n92886 , n92896 );
or ( n92910 , n92908 , n92909 );
xor ( n92911 , n92879 , n92745 );
xnor ( n92912 , n92911 , n92742 );
xor ( n92913 , n92910 , n92912 );
not ( n92914 , n90876 );
nand ( n92915 , n92187 , n90842 );
nand ( n92916 , n91401 , n90843 );
nand ( n92917 , n92915 , n92916 );
not ( n92918 , n92917 );
or ( n92919 , n92914 , n92918 );
or ( n92920 , n90842 , n91299 );
nand ( n92921 , n91297 , n90842 );
nand ( n92922 , n92920 , n92921 );
nand ( n92923 , n92922 , n90839 );
nand ( n92924 , n92919 , n92923 );
xor ( n92925 , n92808 , n92817 );
xor ( n92926 , n92925 , n92847 );
xor ( n92927 , n92924 , n92926 );
and ( n92928 , n92829 , n92830 );
not ( n92929 , n92829 );
and ( n92930 , n92929 , n92831 );
or ( n92931 , n92928 , n92930 );
and ( n92932 , n92844 , n92840 );
xnor ( n92933 , n92931 , n92932 );
not ( n92934 , n92933 );
not ( n92935 , n90842 );
nand ( n92936 , n92935 , n90876 );
or ( n92937 , n91299 , n92936 );
not ( n92938 , n92921 );
nand ( n92939 , n92938 , n90876 );
not ( n92940 , n90842 );
not ( n92941 , n91395 );
or ( n92942 , n92940 , n92941 );
nand ( n92943 , n91394 , n90533 );
nand ( n92944 , n92942 , n92943 );
nand ( n92945 , n92944 , n90839 );
nand ( n92946 , n92937 , n92939 , n92945 );
not ( n92947 , n92946 );
not ( n92948 , n92947 );
or ( n92949 , n92934 , n92948 );
xor ( n92950 , n92844 , n92840 );
not ( n92951 , n90876 );
not ( n92952 , n92944 );
or ( n92953 , n92951 , n92952 );
and ( n92954 , n91587 , n90533 );
not ( n92955 , n91587 );
and ( n92956 , n92955 , n90842 );
or ( n92957 , n92954 , n92956 );
nand ( n92958 , n92957 , n90839 );
nand ( n92959 , n92953 , n92958 );
xor ( n92960 , n92950 , n92959 );
nand ( n92961 , n90535 , n91641 );
not ( n92962 , n92961 );
not ( n92963 , n90876 );
not ( n92964 , n92957 );
or ( n92965 , n92963 , n92964 );
not ( n92966 , n90842 );
not ( n92967 , n91991 );
or ( n92968 , n92966 , n92967 );
nand ( n92969 , n91595 , n90533 );
nand ( n92970 , n92968 , n92969 );
nand ( n92971 , n92970 , n90839 );
nand ( n92972 , n92965 , n92971 );
not ( n92973 , n92972 );
not ( n92974 , n92973 );
or ( n92975 , n92962 , n92974 );
not ( n92976 , n90876 );
not ( n92977 , n92970 );
or ( n92978 , n92976 , n92977 );
or ( n92979 , n90842 , n89865 );
or ( n92980 , n90533 , n91641 );
nand ( n92981 , n92979 , n92980 );
nand ( n92982 , n90839 , n92981 );
nand ( n92983 , n92978 , n92982 );
or ( n92984 , n90830 , n91641 );
nand ( n92985 , n92984 , n90788 );
nand ( n92986 , n90830 , n91641 );
and ( n92987 , n90842 , n92985 , n92986 );
and ( n92988 , n92983 , n92987 );
nand ( n92989 , n92975 , n92988 );
not ( n92990 , n92961 );
nand ( n92991 , n92972 , n92990 );
nand ( n92992 , n92989 , n92991 );
and ( n92993 , n92960 , n92992 );
and ( n92994 , n92950 , n92959 );
or ( n92995 , n92993 , n92994 );
nand ( n92996 , n92949 , n92995 );
not ( n92997 , n92933 );
nand ( n92998 , n92997 , n92946 );
nand ( n92999 , n92996 , n92998 );
and ( n93000 , n92927 , n92999 );
and ( n93001 , n92924 , n92926 );
or ( n93002 , n93000 , n93001 );
not ( n93003 , n87689 );
not ( n93004 , n87706 );
not ( n93005 , n90429 );
or ( n93006 , n93004 , n93005 );
nand ( n93007 , n90428 , n87705 );
nand ( n93008 , n93006 , n93007 );
not ( n93009 , n93008 );
or ( n93010 , n93003 , n93009 );
not ( n93011 , n87706 );
not ( n93012 , n90378 );
or ( n93013 , n93011 , n93012 );
or ( n93014 , n90378 , n87706 );
nand ( n93015 , n93013 , n93014 );
nand ( n93016 , n93015 , n87702 );
nand ( n93017 , n93010 , n93016 );
xor ( n93018 , n93002 , n93017 );
not ( n93019 , n90782 );
not ( n93020 , n90788 );
not ( n93021 , n90386 );
or ( n93022 , n93020 , n93021 );
nand ( n93023 , n90385 , n90799 );
nand ( n93024 , n93022 , n93023 );
not ( n93025 , n93024 );
or ( n93026 , n93019 , n93025 );
not ( n93027 , n90788 );
not ( n93028 , n90991 );
or ( n93029 , n93027 , n93028 );
nand ( n93030 , n90721 , n90799 );
nand ( n93031 , n93029 , n93030 );
nand ( n93032 , n93031 , n90825 );
nand ( n93033 , n93026 , n93032 );
not ( n93034 , n90842 );
not ( n93035 , n90989 );
or ( n93036 , n93034 , n93035 );
nand ( n93037 , n90934 , n90843 );
nand ( n93038 , n93036 , n93037 );
and ( n93039 , n93038 , n90876 );
and ( n93040 , n92917 , n90839 );
nor ( n93041 , n93039 , n93040 );
not ( n93042 , n93041 );
xor ( n93043 , n92796 , n92806 );
xor ( n93044 , n93043 , n92850 );
not ( n93045 , n93044 );
or ( n93046 , n93042 , n93045 );
or ( n93047 , n93044 , n93041 );
nand ( n93048 , n93046 , n93047 );
xor ( n93049 , n93033 , n93048 );
and ( n93050 , n93018 , n93049 );
and ( n93051 , n93002 , n93017 );
or ( n93052 , n93050 , n93051 );
not ( n93053 , n93052 );
not ( n93054 , n87689 );
xor ( n93055 , n87706 , n90417 );
not ( n93056 , n93055 );
or ( n93057 , n93054 , n93056 );
nand ( n93058 , n93008 , n87702 );
nand ( n93059 , n93057 , n93058 );
not ( n93060 , n93033 );
not ( n93061 , n93060 );
not ( n93062 , n93041 );
and ( n93063 , n93061 , n93062 );
nand ( n93064 , n93060 , n93041 );
and ( n93065 , n93064 , n93044 );
nor ( n93066 , n93063 , n93065 );
xor ( n93067 , n93059 , n93066 );
not ( n93068 , n93067 );
and ( n93069 , n93053 , n93068 );
and ( n93070 , n93052 , n93067 );
nor ( n93071 , n93069 , n93070 );
not ( n93072 , n93071 );
not ( n93073 , n90782 );
not ( n93074 , n92864 );
or ( n93075 , n93073 , n93074 );
nand ( n93076 , n93024 , n90825 );
nand ( n93077 , n93075 , n93076 );
not ( n93078 , n93077 );
xor ( n93079 , n92787 , n92793 );
xor ( n93080 , n93079 , n92853 );
not ( n93081 , n90876 );
not ( n93082 , n92778 );
or ( n93083 , n93081 , n93082 );
nand ( n93084 , n93038 , n90839 );
nand ( n93085 , n93083 , n93084 );
xnor ( n93086 , n93080 , n93085 );
not ( n93087 , n93086 );
or ( n93088 , n93078 , n93087 );
or ( n93089 , n93086 , n93077 );
nand ( n93090 , n93088 , n93089 );
nand ( n93091 , n93072 , n93090 );
not ( n93092 , n90782 );
not ( n93093 , n93031 );
or ( n93094 , n93092 , n93093 );
xor ( n93095 , n90788 , n90932 );
nand ( n93096 , n93095 , n90825 );
nand ( n93097 , n93094 , n93096 );
xor ( n93098 , n92924 , n92926 );
xor ( n93099 , n93098 , n92999 );
xor ( n93100 , n93097 , n93099 );
not ( n93101 , n87702 );
xor ( n93102 , n87700 , n90385 );
not ( n93103 , n93102 );
or ( n93104 , n93101 , n93103 );
nand ( n93105 , n93015 , n87689 );
nand ( n93106 , n93104 , n93105 );
and ( n93107 , n93100 , n93106 );
and ( n93108 , n93097 , n93099 );
or ( n93109 , n93107 , n93108 );
xor ( n93110 , n93002 , n93017 );
xor ( n93111 , n93110 , n93049 );
xor ( n93112 , n93109 , n93111 );
not ( n93113 , n87689 );
not ( n93114 , n93102 );
or ( n93115 , n93113 , n93114 );
not ( n93116 , n87706 );
not ( n93117 , n90991 );
or ( n93118 , n93116 , n93117 );
nand ( n93119 , n90721 , n87705 );
nand ( n93120 , n93118 , n93119 );
nand ( n93121 , n93120 , n87702 );
nand ( n93122 , n93115 , n93121 );
not ( n93123 , n93122 );
not ( n93124 , n93123 );
not ( n93125 , n90782 );
not ( n93126 , n93095 );
or ( n93127 , n93125 , n93126 );
not ( n93128 , n90799 );
not ( n93129 , n91401 );
or ( n93130 , n93128 , n93129 );
or ( n93131 , n90799 , n91401 );
nand ( n93132 , n93130 , n93131 );
nand ( n93133 , n93132 , n90824 );
nand ( n93134 , n93127 , n93133 );
not ( n93135 , n93134 );
not ( n93136 , n93135 );
or ( n93137 , n93124 , n93136 );
buf ( n93138 , n92933 );
and ( n93139 , n92947 , n93138 );
not ( n93140 , n92947 );
not ( n93141 , n92933 );
and ( n93142 , n93140 , n93141 );
nor ( n93143 , n93139 , n93142 );
not ( n93144 , n92995 );
and ( n93145 , n93143 , n93144 );
not ( n93146 , n93143 );
and ( n93147 , n93146 , n92995 );
nor ( n93148 , n93145 , n93147 );
not ( n93149 , n93148 );
nand ( n93150 , n93137 , n93149 );
nand ( n93151 , n93122 , n93134 );
nand ( n93152 , n93150 , n93151 );
xor ( n93153 , n93097 , n93099 );
xor ( n93154 , n93153 , n93106 );
xor ( n93155 , n93152 , n93154 );
xor ( n93156 , n92950 , n92959 );
xor ( n93157 , n93156 , n92992 );
not ( n93158 , n90782 );
not ( n93159 , n93132 );
or ( n93160 , n93158 , n93159 );
not ( n93161 , n90788 );
not ( n93162 , n91955 );
or ( n93163 , n93161 , n93162 );
not ( n93164 , n90787 );
nand ( n93165 , n93164 , n91296 );
nand ( n93166 , n93163 , n93165 );
nand ( n93167 , n93166 , n90824 );
nand ( n93168 , n93160 , n93167 );
or ( n93169 , n93157 , n93168 );
not ( n93170 , n93169 );
not ( n93171 , n92990 );
not ( n93172 , n92973 );
or ( n93173 , n93171 , n93172 );
nand ( n93174 , n92972 , n92961 );
nand ( n93175 , n93173 , n93174 );
xnor ( n93176 , n93175 , n92988 );
not ( n93177 , n93176 );
not ( n93178 , n93177 );
not ( n93179 , n90782 );
not ( n93180 , n93166 );
or ( n93181 , n93179 , n93180 );
and ( n93182 , n90788 , n91394 );
not ( n93183 , n90788 );
and ( n93184 , n93183 , n91395 );
nor ( n93185 , n93182 , n93184 );
nand ( n93186 , n93185 , n90824 );
nand ( n93187 , n93181 , n93186 );
not ( n93188 , n93187 );
or ( n93189 , n93178 , n93188 );
or ( n93190 , n93187 , n93177 );
xor ( n93191 , n92987 , n92983 );
not ( n93192 , n90782 );
not ( n93193 , n93185 );
or ( n93194 , n93192 , n93193 );
and ( n93195 , n90788 , n91622 );
not ( n93196 , n90788 );
and ( n93197 , n93196 , n91588 );
nor ( n93198 , n93195 , n93197 );
nand ( n93199 , n93198 , n90824 );
nand ( n93200 , n93194 , n93199 );
xor ( n93201 , n93191 , n93200 );
and ( n93202 , n90876 , n91641 );
not ( n93203 , n90781 );
not ( n93204 , n93198 );
or ( n93205 , n93203 , n93204 );
not ( n93206 , n90788 );
not ( n93207 , n91991 );
or ( n93208 , n93206 , n93207 );
nand ( n93209 , n91595 , n90799 );
nand ( n93210 , n93208 , n93209 );
nand ( n93211 , n93210 , n90824 );
nand ( n93212 , n93205 , n93211 );
xor ( n93213 , n93202 , n93212 );
not ( n93214 , n90781 );
not ( n93215 , n93210 );
or ( n93216 , n93214 , n93215 );
or ( n93217 , n90788 , n89865 );
or ( n93218 , n90799 , n91641 );
nand ( n93219 , n93217 , n93218 );
nand ( n93220 , n90824 , n93219 );
nand ( n93221 , n93216 , n93220 );
not ( n93222 , n93221 );
or ( n93223 , n91641 , n90780 );
nand ( n93224 , n93223 , n87700 );
nand ( n93225 , n91641 , n90780 );
nand ( n93226 , n93224 , n90788 , n93225 );
nor ( n93227 , n93222 , n93226 );
and ( n93228 , n93213 , n93227 );
and ( n93229 , n93202 , n93212 );
or ( n93230 , n93228 , n93229 );
and ( n93231 , n93201 , n93230 );
and ( n93232 , n93191 , n93200 );
or ( n93233 , n93231 , n93232 );
nand ( n93234 , n93190 , n93233 );
nand ( n93235 , n93189 , n93234 );
not ( n93236 , n93235 );
or ( n93237 , n93170 , n93236 );
nand ( n93238 , n93168 , n93157 );
nand ( n93239 , n93237 , n93238 );
not ( n93240 , n93239 );
not ( n93241 , n93149 );
not ( n93242 , n93135 );
or ( n93243 , n93241 , n93242 );
nand ( n93244 , n93148 , n93134 );
nand ( n93245 , n93243 , n93244 );
and ( n93246 , n93245 , n93123 );
not ( n93247 , n93245 );
and ( n93248 , n93247 , n93122 );
nor ( n93249 , n93246 , n93248 );
nand ( n93250 , n93240 , n93249 );
not ( n93251 , n93250 );
not ( n93252 , n93120 );
or ( n93253 , n93252 , n92472 );
and ( n93254 , n90989 , n87706 );
not ( n93255 , n90989 );
and ( n93256 , n93255 , n87705 );
nor ( n93257 , n93254 , n93256 );
or ( n93258 , n93257 , n87701 );
nand ( n93259 , n93253 , n93258 );
not ( n93260 , n93259 );
or ( n93261 , n93157 , n93168 );
nand ( n93262 , n93157 , n93168 );
nand ( n93263 , n93261 , n93262 );
xor ( n93264 , n93263 , n93235 );
nand ( n93265 , n93260 , n93264 );
not ( n93266 , n93265 );
not ( n93267 , n87704 );
not ( n93268 , n91390 );
or ( n93269 , n93267 , n93268 );
nand ( n93270 , n91293 , n91295 , n87700 );
nand ( n93271 , n93269 , n93270 );
not ( n93272 , n93271 );
not ( n93273 , n87702 );
or ( n93274 , n93272 , n93273 );
not ( n93275 , n91401 );
not ( n93276 , n87704 );
and ( n93277 , n93275 , n93276 );
and ( n93278 , n90945 , n87704 );
nor ( n93279 , n93277 , n93278 );
or ( n93280 , n93279 , n92472 );
nand ( n93281 , n93274 , n93280 );
xor ( n93282 , n93191 , n93200 );
xor ( n93283 , n93282 , n93230 );
nor ( n93284 , n93281 , n93283 );
xor ( n93285 , n93202 , n93212 );
xor ( n93286 , n93285 , n93227 );
not ( n93287 , n87689 );
not ( n93288 , n93271 );
or ( n93289 , n93287 , n93288 );
and ( n93290 , n87704 , n91394 );
not ( n93291 , n87704 );
and ( n93292 , n93291 , n91395 );
nor ( n93293 , n93290 , n93292 );
or ( n93294 , n93293 , n87701 );
nand ( n93295 , n93289 , n93294 );
xor ( n93296 , n93286 , n93295 );
not ( n93297 , n93226 );
not ( n93298 , n93221 );
or ( n93299 , n93297 , n93298 );
or ( n93300 , n93221 , n93226 );
nand ( n93301 , n93299 , n93300 );
or ( n93302 , n93293 , n92472 );
and ( n93303 , n87700 , n91588 );
not ( n93304 , n87700 );
and ( n93305 , n93304 , n91622 );
nor ( n93306 , n93303 , n93305 );
or ( n93307 , n93306 , n87701 );
nand ( n93308 , n93302 , n93307 );
xor ( n93309 , n93301 , n93308 );
nor ( n93310 , n90820 , n89865 );
not ( n93311 , n91641 );
not ( n93312 , n87701 );
and ( n93313 , n93311 , n93312 );
not ( n93314 , n87700 );
not ( n93315 , n91991 );
or ( n93316 , n93314 , n93315 );
nand ( n93317 , n91595 , n87704 );
nand ( n93318 , n93316 , n93317 );
and ( n93319 , n93318 , n87689 );
nor ( n93320 , n93313 , n93319 );
nand ( n93321 , n91641 , n87689 );
nand ( n93322 , n93321 , n87700 );
nor ( n93323 , n93320 , n93322 );
xor ( n93324 , n93310 , n93323 );
not ( n93325 , n87702 );
not ( n93326 , n93318 );
or ( n93327 , n93325 , n93326 );
or ( n93328 , n93306 , n92472 );
nand ( n93329 , n93327 , n93328 );
and ( n93330 , n93324 , n93329 );
or ( n93331 , n93330 , C0 );
and ( n93332 , n93309 , n93331 );
and ( n93333 , n93301 , n93308 );
or ( n93334 , n93332 , n93333 );
and ( n93335 , n93296 , n93334 );
and ( n93336 , n93286 , n93295 );
or ( n93337 , n93335 , n93336 );
not ( n93338 , n93337 );
or ( n93339 , n93284 , n93338 );
nand ( n93340 , n93281 , n93283 );
nand ( n93341 , n93339 , n93340 );
not ( n93342 , n93341 );
xor ( n93343 , n93176 , n93187 );
xor ( n93344 , n93343 , n93233 );
not ( n93345 , n93257 );
not ( n93346 , n92472 );
and ( n93347 , n93345 , n93346 );
not ( n93348 , n93279 );
and ( n93349 , n93348 , n87702 );
nor ( n93350 , n93347 , n93349 );
nand ( n93351 , n93344 , n93350 );
not ( n93352 , n93351 );
or ( n93353 , n93342 , n93352 );
or ( n93354 , n93344 , n93350 );
nand ( n93355 , n93353 , n93354 );
not ( n93356 , n93355 );
or ( n93357 , n93266 , n93356 );
not ( n93358 , n93264 );
nand ( n93359 , n93358 , n93259 );
nand ( n93360 , n93357 , n93359 );
not ( n93361 , n93360 );
or ( n93362 , n93251 , n93361 );
not ( n93363 , n93249 );
nand ( n93364 , n93363 , n93239 );
nand ( n93365 , n93362 , n93364 );
and ( n93366 , n93155 , n93365 );
and ( n93367 , n93152 , n93154 );
or ( n93368 , n93366 , n93367 );
and ( n93369 , n93112 , n93368 );
and ( n93370 , n93109 , n93111 );
or ( n93371 , n93369 , n93370 );
not ( n93372 , n93090 );
nand ( n93373 , n93372 , n93071 );
nand ( n93374 , n93371 , n93373 );
nand ( n93375 , n93091 , n93374 );
and ( n93376 , n92856 , n92867 );
not ( n93377 , n92856 );
and ( n93378 , n93377 , n92866 );
or ( n93379 , n93376 , n93378 );
xnor ( n93380 , n92871 , n93379 );
not ( n93381 , n93380 );
or ( n93382 , n93077 , n93085 );
nand ( n93383 , n93382 , n93080 );
nand ( n93384 , n93077 , n93085 );
and ( n93385 , n93383 , n93384 );
and ( n93386 , n92894 , n87689 );
not ( n93387 , n93055 );
nor ( n93388 , n93387 , n87701 );
nor ( n93389 , n93386 , n93388 );
xor ( n93390 , n93385 , n93389 );
not ( n93391 , n93390 );
and ( n93392 , n93381 , n93391 );
and ( n93393 , n93380 , n93390 );
nor ( n93394 , n93392 , n93393 );
not ( n93395 , n93059 );
not ( n93396 , n93395 );
not ( n93397 , n93066 );
and ( n93398 , n93396 , n93397 );
nand ( n93399 , n93395 , n93066 );
and ( n93400 , n93052 , n93399 );
nor ( n93401 , n93398 , n93400 );
and ( n93402 , n93394 , n93401 );
not ( n93403 , n93402 );
and ( n93404 , n93375 , n93403 );
or ( n93405 , n93394 , n93401 );
not ( n93406 , n93405 );
nor ( n93407 , n93404 , n93406 );
xor ( n93408 , n92886 , n92896 );
xor ( n93409 , n93408 , n92907 );
and ( n93410 , n93385 , n93389 );
or ( n93411 , n93380 , n93410 );
or ( n93412 , n93389 , n93385 );
nand ( n93413 , n93411 , n93412 );
buf ( n93414 , n93413 );
nor ( n93415 , n93409 , n93414 );
or ( n93416 , n93407 , n93415 );
nand ( n93417 , n93409 , n93414 );
nand ( n93418 , n93416 , n93417 );
and ( n93419 , n92913 , n93418 );
and ( n93420 , n92910 , n92912 );
or ( n93421 , n93419 , n93420 );
and ( n93422 , n92884 , n93421 );
and ( n93423 , n92881 , n92883 );
or ( n93424 , n93422 , n93423 );
not ( n93425 , n93424 );
or ( n93426 , n92737 , n93425 );
not ( n93427 , n92735 );
nand ( n93428 , n93427 , n92707 );
nand ( n93429 , n93426 , n93428 );
not ( n93430 , n93429 );
not ( n93431 , n92491 );
not ( n93432 , n92478 );
or ( n93433 , n93431 , n93432 );
nand ( n93434 , n92477 , n92487 );
nand ( n93435 , n93433 , n93434 );
not ( n93436 , n92406 );
and ( n93437 , n93435 , n93436 );
not ( n93438 , n93435 );
and ( n93439 , n93438 , n92406 );
nor ( n93440 , n93437 , n93439 );
xor ( n93441 , n92274 , n92378 );
xor ( n93442 , n93441 , n92284 );
not ( n93443 , n93442 );
not ( n93444 , n92723 );
not ( n93445 , n92728 );
or ( n93446 , n93444 , n93445 );
or ( n93447 , n92728 , n92723 );
nand ( n93448 , n93447 , n92733 );
nand ( n93449 , n93446 , n93448 );
not ( n93450 , n93449 );
not ( n93451 , n93450 );
or ( n93452 , n93443 , n93451 );
xor ( n93453 , n92409 , n92457 );
xnor ( n93454 , n93453 , n92475 );
nand ( n93455 , n93452 , n93454 );
not ( n93456 , n93442 );
nand ( n93457 , n93449 , n93456 );
and ( n93458 , n93455 , n93457 );
nand ( n93459 , n93440 , n93458 );
not ( n93460 , n93456 );
not ( n93461 , n93450 );
or ( n93462 , n93460 , n93461 );
nand ( n93463 , n93449 , n93442 );
nand ( n93464 , n93462 , n93463 );
not ( n93465 , n93454 );
and ( n93466 , n93464 , n93465 );
not ( n93467 , n93464 );
buf ( n93468 , n93454 );
and ( n93469 , n93467 , n93468 );
nor ( n93470 , n93466 , n93469 );
xor ( n93471 , n92710 , n92717 );
and ( n93472 , n93471 , n92734 );
and ( n93473 , n92710 , n92717 );
or ( n93474 , n93472 , n93473 );
nand ( n93475 , n93470 , n93474 );
and ( n93476 , n93459 , n93475 );
not ( n93477 , n93476 );
or ( n93478 , n93430 , n93477 );
nor ( n93479 , n93470 , n93474 );
and ( n93480 , n93479 , n93459 );
nor ( n93481 , n93440 , n93458 );
nor ( n93482 , n93480 , n93481 );
nand ( n93483 , n93478 , n93482 );
and ( n93484 , n92496 , n93483 );
and ( n93485 , n92493 , n92495 );
or ( n93486 , n93484 , n93485 );
not ( n93487 , n93486 );
or ( n93488 , n92404 , n93487 );
nand ( n93489 , n92397 , n92401 );
nor ( n93490 , n92249 , n92390 );
and ( n93491 , n93489 , n93490 );
nor ( n93492 , n92397 , n92401 );
nor ( n93493 , n93491 , n93492 );
nand ( n93494 , n93488 , n93493 );
and ( n93495 , n92163 , n93494 );
and ( n93496 , n92072 , n92162 );
or ( n93497 , n93495 , n93496 );
not ( n93498 , n93497 );
or ( n93499 , n92070 , n93498 );
not ( n93500 , n91859 );
and ( n93501 , n91861 , n92067 );
and ( n93502 , n93500 , n93501 );
and ( n93503 , n91858 , n91801 );
nor ( n93504 , n93502 , n93503 );
nand ( n93505 , n93499 , n93504 );
not ( n93506 , n93505 );
or ( n93507 , n91792 , n93506 );
nor ( n93508 , n91528 , n91789 );
and ( n93509 , n91518 , n93508 );
nor ( n93510 , n91474 , n91517 );
nor ( n93511 , n93509 , n93510 );
nand ( n93512 , n93507 , n93511 );
xor ( n93513 , n91469 , n93512 );
not ( n93514 , n87684 );
or ( n93515 , n93513 , n93514 );
nand ( n93516 , n87685 , n93515 );
and ( n93517 , n17246 , n472 );
and ( n93518 , n17265 , n471 );
nor ( n93519 , n93517 , n93518 );
nor ( n93520 , n17327 , n93519 );
buf ( n93521 , n87684 );
not ( n93522 , n93521 );
and ( n93523 , n93520 , n93522 );
and ( n93524 , n93320 , n93322 );
nor ( n93525 , n93524 , n93323 );
and ( n93526 , n93525 , n93521 );
nor ( n93527 , n93523 , n93526 );
or ( n93528 , n17690 , n17722 );
not ( n93529 , n93528 );
not ( n93530 , n93529 );
buf ( n93531 , n17704 );
not ( n93532 , n93531 );
not ( n93533 , n93532 );
not ( n93534 , n17711 );
not ( n93535 , n93534 );
not ( n93536 , n17666 );
or ( n93537 , n93535 , n93536 );
buf ( n93538 , n17716 );
nand ( n93539 , n93537 , n93538 );
not ( n93540 , n93539 );
or ( n93541 , n93533 , n93540 );
buf ( n93542 , n17718 );
nand ( n93543 , n93541 , n93542 );
not ( n93544 , n93543 );
or ( n93545 , n93530 , n93544 );
not ( n93546 , n93528 );
or ( n93547 , n93543 , n93546 );
nand ( n93548 , n93545 , n93547 );
or ( n93549 , n93548 , n87684 );
not ( n93550 , n93503 );
nand ( n93551 , n93550 , n93500 );
not ( n93552 , n92068 );
not ( n93553 , n93552 );
not ( n93554 , n93497 );
or ( n93555 , n93553 , n93554 );
not ( n93556 , n93501 );
nand ( n93557 , n93555 , n93556 );
xor ( n93558 , n93551 , n93557 );
or ( n93559 , n93558 , n93514 );
nand ( n93560 , n93549 , n93559 );
nand ( n93561 , n93532 , n93542 );
and ( n93562 , n93539 , n93561 );
not ( n93563 , n93539 );
not ( n93564 , n93561 );
and ( n93565 , n93563 , n93564 );
nor ( n93566 , n93562 , n93565 );
or ( n93567 , n93566 , n87684 );
nand ( n93568 , n93556 , n93552 );
xor ( n93569 , n93568 , n93497 );
or ( n93570 , n93569 , n93514 );
nand ( n93571 , n93567 , n93570 );
nand ( n93572 , n93534 , n93538 );
not ( n93573 , n93572 );
and ( n93574 , n17666 , n93573 );
not ( n93575 , n17666 );
and ( n93576 , n93575 , n93572 );
or ( n93577 , n93574 , n93576 );
or ( n93578 , n93577 , n87684 );
xor ( n93579 , n92072 , n92162 );
xor ( n93580 , n93579 , n93494 );
not ( n93581 , n93580 );
or ( n93582 , n93581 , n93514 );
nand ( n93583 , n93578 , n93582 );
not ( n93584 , n17639 );
not ( n93585 , n17570 );
not ( n93586 , n16957 );
not ( n93587 , n17381 );
or ( n93588 , n93586 , n93587 );
not ( n93589 , n17644 );
nand ( n93590 , n93588 , n93589 );
not ( n93591 , n93590 );
or ( n93592 , n93585 , n93591 );
nand ( n93593 , n93592 , n17655 );
not ( n93594 , n93593 );
or ( n93595 , n93584 , n93594 );
nand ( n93596 , n93595 , n17663 );
not ( n93597 , n93596 );
not ( n93598 , n17630 );
and ( n93599 , n93598 , n17634 );
not ( n93600 , n93599 );
or ( n93601 , n93597 , n93600 );
or ( n93602 , n93599 , n93596 );
nand ( n93603 , n93601 , n93602 );
or ( n93604 , n93603 , n87684 );
not ( n93605 , n93490 );
nand ( n93606 , n92249 , n92390 );
nand ( n93607 , n93605 , n93606 );
xor ( n93608 , n93607 , n93486 );
or ( n93609 , n93608 , n93514 );
nand ( n93610 , n93604 , n93609 );
not ( n93611 , n17660 );
nand ( n93612 , n93611 , n17622 );
xor ( n93613 , n93593 , n93612 );
or ( n93614 , n93613 , n93521 );
not ( n93615 , n93481 );
nand ( n93616 , n93615 , n93459 );
and ( n93617 , n93424 , n92736 );
not ( n93618 , n93428 );
nor ( n93619 , n93617 , n93618 );
not ( n93620 , n93475 );
or ( n93621 , n93619 , n93620 );
not ( n93622 , n93479 );
nand ( n93623 , n93621 , n93622 );
xor ( n93624 , n93616 , n93623 );
not ( n93625 , n93521 );
or ( n93626 , n93624 , n93625 );
nand ( n93627 , n93614 , n93626 );
not ( n93628 , n10061 );
or ( n93629 , n12702 , n12650 );
nand ( n93630 , n93629 , n499 );
not ( n93631 , n12795 );
xor ( n93632 , n489 , n13046 );
not ( n93633 , n93632 );
or ( n93634 , n93631 , n93633 );
xor ( n93635 , n489 , n13369 );
nand ( n93636 , n93635 , n12542 );
nand ( n93637 , n93634 , n93636 );
xor ( n93638 , n93630 , n93637 );
and ( n93639 , n12835 , n489 );
and ( n93640 , n93638 , n93639 );
and ( n93641 , n93630 , n93637 );
or ( n93642 , n93640 , n93641 );
not ( n93643 , n12758 );
not ( n93644 , n493 );
not ( n93645 , n15540 );
or ( n93646 , n93644 , n93645 );
nand ( n93647 , n15539 , n12775 );
nand ( n93648 , n93646 , n93647 );
not ( n93649 , n93648 );
or ( n93650 , n93643 , n93649 );
not ( n93651 , n493 );
not ( n93652 , n13255 );
or ( n93653 , n93651 , n93652 );
nand ( n93654 , n13258 , n12775 );
nand ( n93655 , n93653 , n93654 );
nand ( n93656 , n93655 , n15344 );
nand ( n93657 , n93650 , n93656 );
and ( n93658 , n12674 , n489 );
xor ( n93659 , n93657 , n93658 );
not ( n93660 , n12638 );
not ( n93661 , n491 );
not ( n93662 , n12419 );
or ( n93663 , n93661 , n93662 );
nand ( n93664 , n12422 , n12610 );
nand ( n93665 , n93663 , n93664 );
not ( n93666 , n93665 );
or ( n93667 , n93660 , n93666 );
not ( n93668 , n491 );
not ( n93669 , n12453 );
or ( n93670 , n93668 , n93669 );
nand ( n93671 , n12456 , n12610 );
nand ( n93672 , n93670 , n93671 );
nand ( n93673 , n93672 , n12595 );
nand ( n93674 , n93667 , n93673 );
and ( n93675 , n93659 , n93674 );
and ( n93676 , n93657 , n93658 );
or ( n93677 , n93675 , n93676 );
xor ( n93678 , n93642 , n93677 );
and ( n93679 , n489 , n13369 );
not ( n93680 , n12758 );
not ( n93681 , n15697 );
and ( n93682 , n93681 , n12775 );
not ( n93683 , n93681 );
and ( n93684 , n93683 , n493 );
or ( n93685 , n93682 , n93684 );
not ( n93686 , n93685 );
or ( n93687 , n93680 , n93686 );
nand ( n93688 , n93648 , n15344 );
nand ( n93689 , n93687 , n93688 );
xor ( n93690 , n93679 , n93689 );
not ( n93691 , n12595 );
not ( n93692 , n93665 );
or ( n93693 , n93691 , n93692 );
not ( n93694 , n491 );
not ( n93695 , n13255 );
or ( n93696 , n93694 , n93695 );
nand ( n93697 , n87441 , n12610 );
nand ( n93698 , n93696 , n93697 );
nand ( n93699 , n93698 , n12638 );
nand ( n93700 , n93693 , n93699 );
xor ( n93701 , n93690 , n93700 );
xor ( n93702 , n93678 , n93701 );
not ( n93703 , n13032 );
not ( n93704 , n16321 );
and ( n93705 , n495 , n93704 );
not ( n93706 , n495 );
and ( n93707 , n93706 , n16321 );
or ( n93708 , n93705 , n93707 );
not ( n93709 , n93708 );
or ( n93710 , n93703 , n93709 );
not ( n93711 , n15928 );
and ( n93712 , n495 , n93711 );
not ( n93713 , n495 );
not ( n93714 , n93711 );
and ( n93715 , n93713 , n93714 );
or ( n93716 , n93712 , n93715 );
nand ( n93717 , n93716 , n12969 );
nand ( n93718 , n93710 , n93717 );
not ( n93719 , n12517 );
buf ( n93720 , n16642 );
and ( n93721 , n497 , n93720 );
not ( n93722 , n497 );
not ( n93723 , n93720 );
and ( n93724 , n93722 , n93723 );
nor ( n93725 , n93721 , n93724 );
not ( n93726 , n93725 );
or ( n93727 , n93719 , n93726 );
nand ( n93728 , n93727 , n16577 );
xor ( n93729 , n93718 , n93728 );
not ( n93730 , n12542 );
not ( n93731 , n93632 );
or ( n93732 , n93730 , n93731 );
xor ( n93733 , n489 , n15566 );
nand ( n93734 , n93733 , n12580 );
nand ( n93735 , n93732 , n93734 );
not ( n93736 , n93735 );
xor ( n93737 , n93729 , n93736 );
not ( n93738 , n12969 );
not ( n93739 , n15697 );
xor ( n93740 , n495 , n93739 );
not ( n93741 , n93740 );
or ( n93742 , n93738 , n93741 );
nand ( n93743 , n93716 , n13032 );
nand ( n93744 , n93742 , n93743 );
not ( n93745 , n12470 );
not ( n93746 , n93725 );
or ( n93747 , n93745 , n93746 );
and ( n93748 , n497 , n16321 );
not ( n93749 , n497 );
and ( n93750 , n93749 , n93704 );
nor ( n93751 , n93748 , n93750 );
nand ( n93752 , n93751 , n12517 );
nand ( n93753 , n93747 , n93752 );
xor ( n93754 , n93744 , n93753 );
not ( n93755 , n12595 );
not ( n93756 , n491 );
not ( n93757 , n15853 );
or ( n93758 , n93756 , n93757 );
nand ( n93759 , n13046 , n12610 );
nand ( n93760 , n93758 , n93759 );
not ( n93761 , n93760 );
or ( n93762 , n93755 , n93761 );
nand ( n93763 , n93672 , n12638 );
nand ( n93764 , n93762 , n93763 );
not ( n93765 , n12580 );
not ( n93766 , n93635 );
or ( n93767 , n93765 , n93766 );
not ( n93768 , n489 );
not ( n93769 , n82600 );
or ( n93770 , n93768 , n93769 );
nand ( n93771 , n12835 , n12560 );
nand ( n93772 , n93770 , n93771 );
nand ( n93773 , n93772 , n12542 );
nand ( n93774 , n93767 , n93773 );
xor ( n93775 , n93764 , n93774 );
not ( n93776 , n12969 );
and ( n93777 , n495 , n15539 );
not ( n93778 , n495 );
and ( n93779 , n93778 , n15543 );
nor ( n93780 , n93777 , n93779 );
not ( n93781 , n93780 );
or ( n93782 , n93776 , n93781 );
nand ( n93783 , n93740 , n13032 );
nand ( n93784 , n93782 , n93783 );
and ( n93785 , n93775 , n93784 );
and ( n93786 , n93764 , n93774 );
or ( n93787 , n93785 , n93786 );
and ( n93788 , n93754 , n93787 );
and ( n93789 , n93744 , n93753 );
or ( n93790 , n93788 , n93789 );
xor ( n93791 , n93737 , n93790 );
xor ( n93792 , n93630 , n93637 );
xor ( n93793 , n93792 , n93639 );
xor ( n93794 , n93657 , n93658 );
xor ( n93795 , n93794 , n93674 );
xor ( n93796 , n93793 , n93795 );
not ( n93797 , n12758 );
not ( n93798 , n93655 );
or ( n93799 , n93797 , n93798 );
not ( n93800 , n493 );
not ( n93801 , n12419 );
or ( n93802 , n93800 , n93801 );
nand ( n93803 , n12775 , n12418 );
nand ( n93804 , n93802 , n93803 );
nand ( n93805 , n93804 , n15344 );
nand ( n93806 , n93799 , n93805 );
not ( n93807 , n93658 );
xor ( n93808 , n93806 , n93807 );
not ( n93809 , n12517 );
xnor ( n93810 , n497 , n15931 );
not ( n93811 , n93810 );
or ( n93812 , n93809 , n93811 );
nand ( n93813 , n93751 , n12470 );
nand ( n93814 , n93812 , n93813 );
and ( n93815 , n93808 , n93814 );
and ( n93816 , n93806 , n93807 );
or ( n93817 , n93815 , n93816 );
and ( n93818 , n93796 , n93817 );
and ( n93819 , n93793 , n93795 );
or ( n93820 , n93818 , n93819 );
xor ( n93821 , n93791 , n93820 );
xor ( n93822 , n93702 , n93821 );
or ( n93823 , n12822 , n12843 );
nand ( n93824 , n93823 , n501 );
and ( n93825 , n13483 , n489 );
xor ( n93826 , n93824 , n93825 );
nand ( n93827 , n13699 , n489 );
not ( n93828 , n93827 );
and ( n93829 , n93826 , n93828 );
and ( n93830 , n93824 , n93825 );
or ( n93831 , n93829 , n93830 );
not ( n93832 , n12702 );
and ( n93833 , n499 , n16643 );
not ( n93834 , n499 );
and ( n93835 , n93834 , n16642 );
or ( n93836 , n93833 , n93835 );
not ( n93837 , n93836 );
or ( n93838 , n93832 , n93837 );
nand ( n93839 , n93838 , n13570 );
xor ( n93840 , n93831 , n93839 );
not ( n93841 , n12638 );
not ( n93842 , n93760 );
or ( n93843 , n93841 , n93842 );
not ( n93844 , n491 );
not ( n93845 , n13370 );
or ( n93846 , n93844 , n93845 );
nand ( n93847 , n12610 , n13369 );
nand ( n93848 , n93846 , n93847 );
nand ( n93849 , n93848 , n12595 );
nand ( n93850 , n93843 , n93849 );
not ( n93851 , n12580 );
not ( n93852 , n93772 );
or ( n93853 , n93851 , n93852 );
and ( n93854 , n489 , n12674 );
not ( n93855 , n489 );
and ( n93856 , n93855 , n13357 );
nor ( n93857 , n93854 , n93856 );
nand ( n93858 , n93857 , n12542 );
nand ( n93859 , n93853 , n93858 );
xor ( n93860 , n93850 , n93859 );
not ( n93861 , n13032 );
not ( n93862 , n93780 );
or ( n93863 , n93861 , n93862 );
not ( n93864 , n495 );
not ( n93865 , n13255 );
or ( n93866 , n93864 , n93865 );
not ( n93867 , n495 );
nand ( n93868 , n93867 , n13258 );
nand ( n93869 , n93866 , n93868 );
nand ( n93870 , n93869 , n12969 );
nand ( n93871 , n93863 , n93870 );
and ( n93872 , n93860 , n93871 );
and ( n93873 , n93850 , n93859 );
or ( n93874 , n93872 , n93873 );
and ( n93875 , n93840 , n93874 );
and ( n93876 , n93831 , n93839 );
or ( n93877 , n93875 , n93876 );
xor ( n93878 , n93744 , n93753 );
xor ( n93879 , n93878 , n93787 );
xor ( n93880 , n93877 , n93879 );
xor ( n93881 , n93764 , n93774 );
xor ( n93882 , n93881 , n93784 );
not ( n93883 , n12758 );
not ( n93884 , n93804 );
or ( n93885 , n93883 , n93884 );
not ( n93886 , n493 );
not ( n93887 , n15563 );
or ( n93888 , n93886 , n93887 );
nand ( n93889 , n15566 , n12775 );
nand ( n93890 , n93888 , n93889 );
nand ( n93891 , n93890 , n15344 );
nand ( n93892 , n93885 , n93891 );
not ( n93893 , n12470 );
not ( n93894 , n93810 );
or ( n93895 , n93893 , n93894 );
xor ( n93896 , n497 , n16253 );
nand ( n93897 , n93896 , n12517 );
nand ( n93898 , n93895 , n93897 );
xor ( n93899 , n93892 , n93898 );
not ( n93900 , n12650 );
not ( n93901 , n93836 );
or ( n93902 , n93900 , n93901 );
not ( n93903 , n499 );
not ( n93904 , n16318 );
or ( n93905 , n93903 , n93904 );
nand ( n93906 , n12467 , n16321 );
nand ( n93907 , n93905 , n93906 );
nand ( n93908 , n93907 , n12702 );
nand ( n93909 , n93902 , n93908 );
and ( n93910 , n93899 , n93909 );
and ( n93911 , n93892 , n93898 );
or ( n93912 , n93910 , n93911 );
xor ( n93913 , n93882 , n93912 );
xor ( n93914 , n93806 , n93807 );
xor ( n93915 , n93914 , n93814 );
and ( n93916 , n93913 , n93915 );
and ( n93917 , n93882 , n93912 );
or ( n93918 , n93916 , n93917 );
and ( n93919 , n93880 , n93918 );
and ( n93920 , n93877 , n93879 );
or ( n93921 , n93919 , n93920 );
xor ( n93922 , n93822 , n93921 );
not ( n93923 , n93922 );
xor ( n93924 , n93793 , n93795 );
xor ( n93925 , n93924 , n93817 );
xor ( n93926 , n93877 , n93879 );
xor ( n93927 , n93926 , n93918 );
xor ( n93928 , n93925 , n93927 );
not ( n93929 , n12542 );
not ( n93930 , n489 );
not ( n93931 , n12694 );
or ( n93932 , n93930 , n93931 );
not ( n93933 , n489 );
nand ( n93934 , n93933 , n12693 );
nand ( n93935 , n93932 , n93934 );
not ( n93936 , n93935 );
or ( n93937 , n93929 , n93936 );
nand ( n93938 , n93857 , n12580 );
nand ( n93939 , n93937 , n93938 );
xor ( n93940 , n93939 , n93827 );
nand ( n93941 , n12509 , n489 );
not ( n93942 , n12462 );
nand ( n93943 , n93942 , n70376 );
nand ( n93944 , n93941 , n93943 );
and ( n93945 , n93940 , n93944 );
and ( n93946 , n93939 , n93827 );
or ( n93947 , n93945 , n93946 );
xor ( n93948 , n93824 , n93825 );
xor ( n93949 , n93948 , n93828 );
xor ( n93950 , n93947 , n93949 );
not ( n93951 , n93890 );
not ( n93952 , n12758 );
or ( n93953 , n93951 , n93952 );
not ( n93954 , n12885 );
not ( n93955 , n12775 );
or ( n93956 , n93954 , n93955 );
nand ( n93957 , n12886 , n493 );
nand ( n93958 , n93956 , n93957 );
nand ( n93959 , n93958 , n15344 );
nand ( n93960 , n93953 , n93959 );
not ( n93961 , n12638 );
not ( n93962 , n93848 );
or ( n93963 , n93961 , n93962 );
not ( n93964 , n12824 );
not ( n93965 , n12829 );
or ( n93966 , n93964 , n93965 );
nand ( n93967 , n93966 , n12834 );
and ( n93968 , n93967 , n12610 );
not ( n93969 , n93967 );
and ( n93970 , n93969 , n491 );
or ( n93971 , n93968 , n93970 );
nand ( n93972 , n93971 , n12595 );
nand ( n93973 , n93963 , n93972 );
xor ( n93974 , n93960 , n93973 );
not ( n93975 , n12470 );
not ( n93976 , n93896 );
or ( n93977 , n93975 , n93976 );
and ( n93978 , n15538 , n497 );
not ( n93979 , n15538 );
and ( n93980 , n93979 , n70541 );
nor ( n93981 , n93978 , n93980 );
nand ( n93982 , n93981 , n12517 );
nand ( n93983 , n93977 , n93982 );
and ( n93984 , n93974 , n93983 );
and ( n93985 , n93960 , n93973 );
or ( n93986 , n93984 , n93985 );
and ( n93987 , n93950 , n93986 );
and ( n93988 , n93947 , n93949 );
or ( n93989 , n93987 , n93988 );
xor ( n93990 , n93831 , n93839 );
xor ( n93991 , n93990 , n93874 );
xor ( n93992 , n93989 , n93991 );
xor ( n93993 , n93850 , n93859 );
xor ( n93994 , n93993 , n93871 );
xor ( n93995 , n93892 , n93898 );
xor ( n93996 , n93995 , n93909 );
xor ( n93997 , n93994 , n93996 );
not ( n93998 , n13032 );
not ( n93999 , n93869 );
or ( n94000 , n93998 , n93999 );
not ( n94001 , n3325 );
not ( n94002 , n12418 );
or ( n94003 , n94001 , n94002 );
nand ( n94004 , n495 , n15438 );
nand ( n94005 , n94003 , n94004 );
nand ( n94006 , n94005 , n12969 );
nand ( n94007 , n94000 , n94006 );
not ( n94008 , n12650 );
not ( n94009 , n93907 );
or ( n94010 , n94008 , n94009 );
not ( n94011 , n499 );
not ( n94012 , n93711 );
or ( n94013 , n94011 , n94012 );
nand ( n94014 , n15928 , n12467 );
nand ( n94015 , n94013 , n94014 );
nand ( n94016 , n94015 , n12702 );
nand ( n94017 , n94010 , n94016 );
xor ( n94018 , n94007 , n94017 );
not ( n94019 , n12822 );
not ( n94020 , n501 );
not ( n94021 , n16643 );
or ( n94022 , n94020 , n94021 );
nand ( n94023 , n71522 , n16642 );
nand ( n94024 , n94022 , n94023 );
not ( n94025 , n94024 );
or ( n94026 , n94019 , n94025 );
nand ( n94027 , n94026 , n16254 );
and ( n94028 , n94018 , n94027 );
and ( n94029 , n94007 , n94017 );
or ( n94030 , n94028 , n94029 );
and ( n94031 , n93997 , n94030 );
and ( n94032 , n93994 , n93996 );
or ( n94033 , n94031 , n94032 );
and ( n94034 , n93992 , n94033 );
and ( n94035 , n93989 , n93991 );
or ( n94036 , n94034 , n94035 );
and ( n94037 , n93928 , n94036 );
and ( n94038 , n93925 , n93927 );
or ( n94039 , n94037 , n94038 );
not ( n94040 , n94039 );
nand ( n94041 , n93923 , n94040 );
not ( n94042 , n94041 );
xor ( n94043 , n93882 , n93912 );
xor ( n94044 , n94043 , n93915 );
xor ( n94045 , n93989 , n93991 );
xor ( n94046 , n94045 , n94033 );
xor ( n94047 , n94044 , n94046 );
xor ( n94048 , n93947 , n93949 );
xor ( n94049 , n94048 , n93986 );
not ( n94050 , n12580 );
not ( n94051 , n93935 );
or ( n94052 , n94050 , n94051 );
nand ( n94053 , n87483 , n12542 );
nand ( n94054 , n94052 , n94053 );
not ( n94055 , n87476 );
and ( n94056 , n87487 , n94055 );
xor ( n94057 , n94054 , n94056 );
or ( n94058 , n93941 , n93943 );
nand ( n94059 , n94058 , n93944 );
and ( n94060 , n94057 , n94059 );
and ( n94061 , n94054 , n94056 );
or ( n94062 , n94060 , n94061 );
xor ( n94063 , n93939 , n93827 );
xor ( n94064 , n94063 , n93944 );
xor ( n94065 , n94062 , n94064 );
xor ( n94066 , n93960 , n93973 );
xor ( n94067 , n94066 , n93983 );
and ( n94068 , n94065 , n94067 );
and ( n94069 , n94062 , n94064 );
or ( n94070 , n94068 , n94069 );
xor ( n94071 , n94049 , n94070 );
not ( n94072 , n12758 );
not ( n94073 , n93958 );
or ( n94074 , n94072 , n94073 );
nand ( n94075 , n17776 , n15344 );
nand ( n94076 , n94074 , n94075 );
not ( n94077 , n12638 );
not ( n94078 , n93971 );
or ( n94079 , n94077 , n94078 );
nand ( n94080 , n12595 , n87471 );
nand ( n94081 , n94079 , n94080 );
xor ( n94082 , n94076 , n94081 );
not ( n94083 , n12470 );
not ( n94084 , n93981 );
or ( n94085 , n94083 , n94084 );
not ( n94086 , n497 );
not ( n94087 , n13255 );
or ( n94088 , n94086 , n94087 );
nand ( n94089 , n13258 , n12486 );
nand ( n94090 , n94088 , n94089 );
nand ( n94091 , n94090 , n12517 );
nand ( n94092 , n94085 , n94091 );
and ( n94093 , n94082 , n94092 );
and ( n94094 , n94076 , n94081 );
or ( n94095 , n94093 , n94094 );
not ( n94096 , n13032 );
not ( n94097 , n94005 );
or ( n94098 , n94096 , n94097 );
nand ( n94099 , n17766 , n12969 );
nand ( n94100 , n94098 , n94099 );
not ( n94101 , n12702 );
not ( n94102 , n87416 );
or ( n94103 , n94101 , n94102 );
nand ( n94104 , n94015 , n12650 );
nand ( n94105 , n94103 , n94104 );
xor ( n94106 , n94100 , n94105 );
not ( n94107 , n12843 );
not ( n94108 , n94024 );
or ( n94109 , n94107 , n94108 );
not ( n94110 , n501 );
not ( n94111 , n16318 );
or ( n94112 , n94110 , n94111 );
nand ( n94113 , n16321 , n12856 );
nand ( n94114 , n94112 , n94113 );
nand ( n94115 , n94114 , n12822 );
nand ( n94116 , n94109 , n94115 );
and ( n94117 , n94106 , n94116 );
and ( n94118 , n94100 , n94105 );
or ( n94119 , n94117 , n94118 );
xor ( n94120 , n94095 , n94119 );
xor ( n94121 , n94007 , n94017 );
xor ( n94122 , n94121 , n94027 );
and ( n94123 , n94120 , n94122 );
and ( n94124 , n94095 , n94119 );
or ( n94125 , n94123 , n94124 );
and ( n94126 , n94071 , n94125 );
and ( n94127 , n94049 , n94070 );
or ( n94128 , n94126 , n94127 );
xor ( n94129 , n94047 , n94128 );
xor ( n94130 , n93994 , n93996 );
xor ( n94131 , n94130 , n94030 );
xor ( n94132 , n87473 , n87474 );
and ( n94133 , n94132 , n87491 );
and ( n94134 , n87473 , n87474 );
or ( n94135 , n94133 , n94134 );
xor ( n94136 , n94054 , n94056 );
xor ( n94137 , n94136 , n94059 );
xor ( n94138 , n94135 , n94137 );
xor ( n94139 , n17768 , n17781 );
and ( n94140 , n94139 , n87418 );
and ( n94141 , n17768 , n17781 );
or ( n94142 , n94140 , n94141 );
and ( n94143 , n94138 , n94142 );
and ( n94144 , n94135 , n94137 );
or ( n94145 , n94143 , n94144 );
xor ( n94146 , n94062 , n94064 );
xor ( n94147 , n94146 , n94067 );
xor ( n94148 , n94145 , n94147 );
xor ( n94149 , n94076 , n94081 );
xor ( n94150 , n94149 , n94092 );
xor ( n94151 , n87444 , n87453 );
and ( n94152 , n94151 , n87458 );
and ( n94153 , n87444 , n87453 );
or ( n94154 , n94152 , n94153 );
xor ( n94155 , n94150 , n94154 );
xor ( n94156 , n94100 , n94105 );
xor ( n94157 , n94156 , n94116 );
and ( n94158 , n94155 , n94157 );
and ( n94159 , n94150 , n94154 );
or ( n94160 , n94158 , n94159 );
and ( n94161 , n94148 , n94160 );
and ( n94162 , n94145 , n94147 );
or ( n94163 , n94161 , n94162 );
xor ( n94164 , n94131 , n94163 );
xor ( n94165 , n94049 , n94070 );
xor ( n94166 , n94165 , n94125 );
and ( n94167 , n94164 , n94166 );
and ( n94168 , n94131 , n94163 );
or ( n94169 , n94167 , n94168 );
nor ( n94170 , n94129 , n94169 );
xor ( n94171 , n93925 , n93927 );
xor ( n94172 , n94171 , n94036 );
xor ( n94173 , n94044 , n94046 );
and ( n94174 , n94173 , n94128 );
and ( n94175 , n94044 , n94046 );
or ( n94176 , n94174 , n94175 );
nor ( n94177 , n94172 , n94176 );
nor ( n94178 , n94170 , n94177 );
not ( n94179 , n94178 );
xor ( n94180 , n87429 , n87504 );
and ( n94181 , n94180 , n87509 );
and ( n94182 , n87429 , n87504 );
or ( n94183 , n94181 , n94182 );
xor ( n94184 , n87419 , n87423 );
and ( n94185 , n94184 , n87428 );
and ( n94186 , n87419 , n87423 );
or ( n94187 , n94185 , n94186 );
xor ( n94188 , n87459 , n87498 );
and ( n94189 , n94188 , n87503 );
and ( n94190 , n87459 , n87498 );
or ( n94191 , n94189 , n94190 );
xor ( n94192 , n94187 , n94191 );
xor ( n94193 , n87463 , n87492 );
and ( n94194 , n94193 , n87497 );
and ( n94195 , n87463 , n87492 );
or ( n94196 , n94194 , n94195 );
xor ( n94197 , n94135 , n94137 );
xor ( n94198 , n94197 , n94142 );
xor ( n94199 , n94196 , n94198 );
xor ( n94200 , n94150 , n94154 );
xor ( n94201 , n94200 , n94157 );
xor ( n94202 , n94199 , n94201 );
xor ( n94203 , n94192 , n94202 );
nor ( n94204 , n94183 , n94203 );
not ( n94205 , n94204 );
xor ( n94206 , n94095 , n94119 );
xor ( n94207 , n94206 , n94122 );
xor ( n94208 , n94145 , n94147 );
xor ( n94209 , n94208 , n94160 );
xor ( n94210 , n94207 , n94209 );
xor ( n94211 , n94196 , n94198 );
and ( n94212 , n94211 , n94201 );
and ( n94213 , n94196 , n94198 );
or ( n94214 , n94212 , n94213 );
xor ( n94215 , n94210 , n94214 );
xor ( n94216 , n94187 , n94191 );
and ( n94217 , n94216 , n94202 );
and ( n94218 , n94187 , n94191 );
or ( n94219 , n94217 , n94218 );
nor ( n94220 , n94215 , n94219 );
not ( n94221 , n94220 );
xor ( n94222 , n94207 , n94209 );
and ( n94223 , n94222 , n94214 );
and ( n94224 , n94207 , n94209 );
or ( n94225 , n94223 , n94224 );
not ( n94226 , n94225 );
xor ( n94227 , n94131 , n94163 );
xor ( n94228 , n94227 , n94166 );
not ( n94229 , n94228 );
nand ( n94230 , n94226 , n94229 );
nand ( n94231 , n94205 , n87520 , n94221 , n94230 );
nor ( n94232 , n17754 , n94231 );
not ( n94233 , n94203 );
not ( n94234 , n94183 );
or ( n94235 , n94233 , n94234 );
nand ( n94236 , n94228 , n94225 );
nand ( n94237 , n94235 , n94236 );
and ( n94238 , n94215 , n94219 );
nor ( n94239 , n94237 , n94238 );
not ( n94240 , n94204 );
nand ( n94241 , n94240 , n87517 );
and ( n94242 , n94239 , n94241 );
not ( n94243 , n94215 );
not ( n94244 , n94219 );
nand ( n94245 , n94243 , n94244 );
nand ( n94246 , n94230 , n94245 );
nand ( n94247 , n94225 , n94228 );
and ( n94248 , n94246 , n94247 );
nor ( n94249 , n94242 , n94248 );
nor ( n94250 , n94232 , n94249 );
not ( n94251 , n15777 );
not ( n94252 , n15771 );
or ( n94253 , n94251 , n94252 );
nor ( n94254 , n94231 , n87381 );
nand ( n94255 , n94253 , n94254 );
nand ( n94256 , n94250 , n94255 );
not ( n94257 , n94256 );
or ( n94258 , n94179 , n94257 );
nor ( n94259 , n94172 , n94176 );
nand ( n94260 , n94129 , n94169 );
or ( n94261 , n94259 , n94260 );
nand ( n94262 , n94172 , n94176 );
nand ( n94263 , n94261 , n94262 );
not ( n94264 , n94263 );
nand ( n94265 , n94258 , n94264 );
not ( n94266 , n94265 );
or ( n94267 , n94042 , n94266 );
nand ( n94268 , n93922 , n94039 );
nand ( n94269 , n94267 , n94268 );
xor ( n94270 , n93702 , n93821 );
and ( n94271 , n94270 , n93921 );
and ( n94272 , n93702 , n93821 );
or ( n94273 , n94271 , n94272 );
xor ( n94274 , n93642 , n93677 );
and ( n94275 , n94274 , n93701 );
and ( n94276 , n93642 , n93677 );
or ( n94277 , n94275 , n94276 );
xor ( n94278 , n93718 , n93728 );
and ( n94279 , n94278 , n93736 );
and ( n94280 , n93718 , n93728 );
or ( n94281 , n94279 , n94280 );
not ( n94282 , n12580 );
not ( n94283 , n489 );
not ( n94284 , n12419 );
or ( n94285 , n94283 , n94284 );
nand ( n94286 , n12422 , n12560 );
nand ( n94287 , n94285 , n94286 );
not ( n94288 , n94287 );
or ( n94289 , n94282 , n94288 );
nand ( n94290 , n93733 , n12542 );
nand ( n94291 , n94289 , n94290 );
not ( n94292 , n15344 );
not ( n94293 , n93685 );
or ( n94294 , n94292 , n94293 );
not ( n94295 , n493 );
not ( n94296 , n93711 );
or ( n94297 , n94295 , n94296 );
nand ( n94298 , n93714 , n12775 );
nand ( n94299 , n94297 , n94298 );
nand ( n94300 , n94299 , n12758 );
nand ( n94301 , n94294 , n94300 );
xor ( n94302 , n94291 , n94301 );
not ( n94303 , n13032 );
and ( n94304 , n495 , n93723 );
not ( n94305 , n495 );
and ( n94306 , n94305 , n93720 );
or ( n94307 , n94304 , n94306 );
not ( n94308 , n94307 );
or ( n94309 , n94303 , n94308 );
nand ( n94310 , n93708 , n12969 );
nand ( n94311 , n94309 , n94310 );
xor ( n94312 , n94302 , n94311 );
xor ( n94313 , n94281 , n94312 );
xor ( n94314 , n93679 , n93689 );
and ( n94315 , n94314 , n93700 );
and ( n94316 , n93679 , n93689 );
or ( n94317 , n94315 , n94316 );
xor ( n94318 , n93735 , n94317 );
or ( n94319 , n12517 , n12470 );
nand ( n94320 , n94319 , n497 );
and ( n94321 , n489 , n13046 );
xor ( n94322 , n94320 , n94321 );
not ( n94323 , n12638 );
not ( n94324 , n491 );
not ( n94325 , n15543 );
or ( n94326 , n94324 , n94325 );
nand ( n94327 , n15544 , n12610 );
nand ( n94328 , n94326 , n94327 );
not ( n94329 , n94328 );
or ( n94330 , n94323 , n94329 );
nand ( n94331 , n93698 , n12595 );
nand ( n94332 , n94330 , n94331 );
xor ( n94333 , n94322 , n94332 );
xor ( n94334 , n94318 , n94333 );
xor ( n94335 , n94313 , n94334 );
xor ( n94336 , n94277 , n94335 );
xor ( n94337 , n93737 , n93790 );
and ( n94338 , n94337 , n93820 );
and ( n94339 , n93737 , n93790 );
or ( n94340 , n94338 , n94339 );
xor ( n94341 , n94336 , n94340 );
or ( n94342 , n94273 , n94341 );
nand ( n94343 , n94341 , n94273 );
nand ( n94344 , n94342 , n94343 );
not ( n94345 , n94344 );
and ( n94346 , n94269 , n94345 );
not ( n94347 , n94269 );
xnor ( n94348 , n94273 , n94341 );
and ( n94349 , n94347 , n94348 );
nor ( n94350 , n94346 , n94349 );
not ( n94351 , n94350 );
or ( n94352 , n93628 , n94351 );
nand ( n94353 , n16505 , n16402 );
and ( n94354 , n16396 , n94353 );
not ( n94355 , n87651 );
not ( n94356 , n16501 );
not ( n94357 , n16402 );
nand ( n94358 , n94356 , n94357 );
nand ( n94359 , n94355 , n94358 );
nor ( n94360 , n94354 , n94359 );
not ( n94361 , n87654 );
nor ( n94362 , n94360 , n94361 );
not ( n94363 , n16391 );
not ( n94364 , n87651 );
nand ( n94365 , n94364 , n94358 );
nor ( n94366 , n94363 , n94365 );
nand ( n94367 , n94366 , n9922 );
nand ( n94368 , n94362 , n94367 );
or ( n94369 , n6955 , n6811 );
nand ( n94370 , n94369 , n547 );
not ( n94371 , n537 );
nor ( n94372 , n94371 , n7378 );
xor ( n94373 , n94370 , n94372 );
nor ( n94374 , n6885 , n5123 );
and ( n94375 , n94373 , n94374 );
and ( n94376 , n94370 , n94372 );
or ( n94377 , n94375 , n94376 );
not ( n94378 , n75018 );
and ( n94379 , n9553 , n4440 );
not ( n94380 , n9553 );
and ( n94381 , n94380 , n545 );
or ( n94382 , n94379 , n94381 );
not ( n94383 , n94382 );
or ( n94384 , n94378 , n94383 );
not ( n94385 , n70470 );
not ( n94386 , n9845 );
or ( n94387 , n94385 , n94386 );
nand ( n94388 , n9794 , n455 );
nand ( n94389 , n94387 , n94388 );
and ( n94390 , n94389 , n545 );
not ( n94391 , n94389 );
and ( n94392 , n94391 , n5268 );
nor ( n94393 , n94390 , n94392 );
nand ( n94394 , n94393 , n5399 );
nand ( n94395 , n94384 , n94394 );
not ( n94396 , n5590 );
not ( n94397 , n541 );
not ( n94398 , n9735 );
or ( n94399 , n94397 , n94398 );
nand ( n94400 , n9734 , n5538 );
nand ( n94401 , n94399 , n94400 );
not ( n94402 , n94401 );
or ( n94403 , n94396 , n94402 );
not ( n94404 , n541 );
not ( n94405 , n9945 );
or ( n94406 , n94404 , n94405 );
nand ( n94407 , n76644 , n5538 );
nand ( n94408 , n94406 , n94407 );
nand ( n94409 , n94408 , n9938 );
nand ( n94410 , n94403 , n94409 );
xor ( n94411 , n94395 , n94410 );
not ( n94412 , n4434 );
not ( n94413 , n539 );
not ( n94414 , n6867 );
or ( n94415 , n94413 , n94414 );
not ( n94416 , n6867 );
nand ( n94417 , n94416 , n4251 );
nand ( n94418 , n94415 , n94417 );
not ( n94419 , n94418 );
or ( n94420 , n94412 , n94419 );
not ( n94421 , n4251 );
not ( n94422 , n7175 );
not ( n94423 , n94422 );
or ( n94424 , n94421 , n94423 );
nand ( n94425 , n7175 , n539 );
nand ( n94426 , n94424 , n94425 );
nand ( n94427 , n94426 , n4224 );
nand ( n94428 , n94420 , n94427 );
and ( n94429 , n94411 , n94428 );
and ( n94430 , n94395 , n94410 );
or ( n94431 , n94429 , n94430 );
xor ( n94432 , n94377 , n94431 );
not ( n94433 , n5590 );
not ( n94434 , n541 );
not ( n94435 , n9382 );
or ( n94436 , n94434 , n94435 );
nand ( n94437 , n7160 , n5538 );
nand ( n94438 , n94436 , n94437 );
not ( n94439 , n94438 );
or ( n94440 , n94433 , n94439 );
nand ( n94441 , n94401 , n9938 );
nand ( n94442 , n94440 , n94441 );
nand ( n94443 , n7304 , n537 );
xor ( n94444 , n94442 , n94443 );
not ( n94445 , n75018 );
and ( n94446 , n94389 , n545 );
not ( n94447 , n94389 );
and ( n94448 , n94447 , n4440 );
nor ( n94449 , n94446 , n94448 );
not ( n94450 , n94449 );
or ( n94451 , n94445 , n94450 );
nand ( n94452 , n5399 , n545 );
nand ( n94453 , n94451 , n94452 );
xor ( n94454 , n94444 , n94453 );
and ( n94455 , n94432 , n94454 );
and ( n94456 , n94377 , n94431 );
or ( n94457 , n94455 , n94456 );
not ( n94458 , n5501 );
not ( n94459 , n537 );
not ( n94460 , n6867 );
or ( n94461 , n94459 , n94460 );
nand ( n94462 , n94416 , n5409 );
nand ( n94463 , n94461 , n94462 );
not ( n94464 , n94463 );
or ( n94465 , n94458 , n94464 );
not ( n94466 , n537 );
not ( n94467 , n7175 );
or ( n94468 , n94466 , n94467 );
nand ( n94469 , n94422 , n5409 );
nand ( n94470 , n94468 , n94469 );
nand ( n94471 , n94470 , n16155 );
nand ( n94472 , n94465 , n94471 );
not ( n94473 , n5590 );
not ( n94474 , n541 );
not ( n94475 , n9557 );
or ( n94476 , n94474 , n94475 );
not ( n94477 , n9557 );
nand ( n94478 , n94477 , n5538 );
nand ( n94479 , n94476 , n94478 );
not ( n94480 , n94479 );
or ( n94481 , n94473 , n94480 );
nand ( n94482 , n94438 , n9938 );
nand ( n94483 , n94481 , n94482 );
xor ( n94484 , n94472 , n94483 );
and ( n94485 , n537 , n6848 );
xor ( n94486 , n94484 , n94485 );
or ( n94487 , n75018 , n5399 );
nand ( n94488 , n94487 , n545 );
not ( n94489 , n4445 );
not ( n94490 , n543 );
not ( n94491 , n9554 );
or ( n94492 , n94490 , n94491 );
nand ( n94493 , n9757 , n4938 );
nand ( n94494 , n94492 , n94493 );
not ( n94495 , n94494 );
or ( n94496 , n94489 , n94495 );
not ( n94497 , n543 );
not ( n94498 , n9848 );
or ( n94499 , n94497 , n94498 );
buf ( n94500 , n79653 );
nand ( n94501 , n94500 , n4938 );
nand ( n94502 , n94499 , n94501 );
nand ( n94503 , n94502 , n9595 );
nand ( n94504 , n94496 , n94503 );
xor ( n94505 , n94488 , n94504 );
not ( n94506 , n4434 );
not ( n94507 , n539 );
not ( n94508 , n9735 );
or ( n94509 , n94507 , n94508 );
not ( n94510 , n9735 );
nand ( n94511 , n94510 , n4251 );
nand ( n94512 , n94509 , n94511 );
not ( n94513 , n94512 );
or ( n94514 , n94506 , n94513 );
not ( n94515 , n539 );
buf ( n94516 , n76644 );
not ( n94517 , n94516 );
not ( n94518 , n94517 );
or ( n94519 , n94515 , n94518 );
nand ( n94520 , n94516 , n4251 );
nand ( n94521 , n94519 , n94520 );
nand ( n94522 , n4224 , n94521 );
nand ( n94523 , n94514 , n94522 );
xor ( n94524 , n94505 , n94523 );
xor ( n94525 , n94486 , n94524 );
not ( n94526 , n94443 );
not ( n94527 , n4445 );
not ( n94528 , n543 );
not ( n94529 , n9557 );
or ( n94530 , n94528 , n94529 );
nand ( n94531 , n94477 , n4938 );
nand ( n94532 , n94530 , n94531 );
not ( n94533 , n94532 );
or ( n94534 , n94527 , n94533 );
nand ( n94535 , n94494 , n9595 );
nand ( n94536 , n94534 , n94535 );
not ( n94537 , n4433 );
not ( n94538 , n94521 );
or ( n94539 , n94537 , n94538 );
nand ( n94540 , n94418 , n4224 );
nand ( n94541 , n94539 , n94540 );
xor ( n94542 , n94536 , n94541 );
not ( n94543 , n94470 );
not ( n94544 , n5501 );
or ( n94545 , n94543 , n94544 );
xor ( n94546 , n537 , n6848 );
not ( n94547 , n94546 );
not ( n94548 , n16155 );
or ( n94549 , n94547 , n94548 );
nand ( n94550 , n94545 , n94549 );
and ( n94551 , n94542 , n94550 );
and ( n94552 , n94536 , n94541 );
or ( n94553 , n94551 , n94552 );
xor ( n94554 , n94526 , n94553 );
xor ( n94555 , n94442 , n94443 );
and ( n94556 , n94555 , n94453 );
and ( n94557 , n94442 , n94443 );
or ( n94558 , n94556 , n94557 );
xor ( n94559 , n94554 , n94558 );
xor ( n94560 , n94525 , n94559 );
xor ( n94561 , n94457 , n94560 );
xor ( n94562 , n94536 , n94541 );
xor ( n94563 , n94562 , n94550 );
not ( n94564 , n5501 );
not ( n94565 , n94546 );
or ( n94566 , n94564 , n94565 );
not ( n94567 , n537 );
not ( n94568 , n7303 );
or ( n94569 , n94567 , n94568 );
nand ( n94570 , n5392 , n5409 );
nand ( n94571 , n94569 , n94570 );
nand ( n94572 , n94571 , n16155 );
nand ( n94573 , n94566 , n94572 );
not ( n94574 , n9595 );
not ( n94575 , n94532 );
or ( n94576 , n94574 , n94575 );
not ( n94577 , n543 );
not ( n94578 , n9382 );
or ( n94579 , n94577 , n94578 );
not ( n94580 , n9382 );
nand ( n94581 , n94580 , n4938 );
nand ( n94582 , n94579 , n94581 );
nand ( n94583 , n94582 , n4445 );
nand ( n94584 , n94576 , n94583 );
xor ( n94585 , n94573 , n94584 );
xor ( n94586 , n94370 , n94372 );
xor ( n94587 , n94586 , n94374 );
and ( n94588 , n94585 , n94587 );
and ( n94589 , n94573 , n94584 );
or ( n94590 , n94588 , n94589 );
xor ( n94591 , n94563 , n94590 );
not ( n94592 , n5501 );
not ( n94593 , n94571 );
or ( n94594 , n94592 , n94593 );
nand ( n94595 , n87587 , n16155 );
nand ( n94596 , n94594 , n94595 );
not ( n94597 , n94374 );
xor ( n94598 , n94596 , n94597 );
not ( n94599 , n87575 );
or ( n94600 , n94599 , n75017 );
not ( n94601 , n94382 );
or ( n94602 , n94601 , n7649 );
nand ( n94603 , n94600 , n94602 );
and ( n94604 , n94598 , n94603 );
and ( n94605 , n94596 , n94597 );
or ( n94606 , n94604 , n94605 );
not ( n94607 , n5590 );
not ( n94608 , n94408 );
or ( n94609 , n94607 , n94608 );
nand ( n94610 , n87551 , n9938 );
nand ( n94611 , n94609 , n94610 );
xor ( n94612 , n87616 , n87617 );
and ( n94613 , n94612 , n87619 );
and ( n94614 , n87616 , n87617 );
or ( n94615 , n94613 , n94614 );
xor ( n94616 , n94611 , n94615 );
not ( n94617 , n94426 );
or ( n94618 , n94617 , n5780 );
not ( n94619 , n87560 );
or ( n94620 , n94619 , n5771 );
nand ( n94621 , n94618 , n94620 );
and ( n94622 , n94616 , n94621 );
and ( n94623 , n94611 , n94615 );
or ( n94624 , n94622 , n94623 );
xor ( n94625 , n94606 , n94624 );
xor ( n94626 , n94395 , n94410 );
xor ( n94627 , n94626 , n94428 );
and ( n94628 , n94625 , n94627 );
and ( n94629 , n94606 , n94624 );
or ( n94630 , n94628 , n94629 );
and ( n94631 , n94591 , n94630 );
and ( n94632 , n94563 , n94590 );
or ( n94633 , n94631 , n94632 );
xor ( n94634 , n94561 , n94633 );
not ( n94635 , n94634 );
xor ( n94636 , n94377 , n94431 );
xor ( n94637 , n94636 , n94454 );
xor ( n94638 , n94563 , n94590 );
xor ( n94639 , n94638 , n94630 );
xor ( n94640 , n94637 , n94639 );
xor ( n94641 , n94573 , n94584 );
xor ( n94642 , n94641 , n94587 );
not ( n94643 , n6854 );
not ( n94644 , n87608 );
or ( n94645 , n94643 , n94644 );
nand ( n94646 , n94645 , n7637 );
not ( n94647 , n4445 );
not ( n94648 , n87597 );
or ( n94649 , n94647 , n94648 );
nand ( n94650 , n94582 , n9595 );
nand ( n94651 , n94649 , n94650 );
xor ( n94652 , n94646 , n94651 );
xor ( n94653 , n87555 , n87568 );
and ( n94654 , n94653 , n87579 );
and ( n94655 , n87555 , n87568 );
or ( n94656 , n94654 , n94655 );
and ( n94657 , n94652 , n94656 );
and ( n94658 , n94646 , n94651 );
or ( n94659 , n94657 , n94658 );
xor ( n94660 , n94642 , n94659 );
xor ( n94661 , n94606 , n94624 );
xor ( n94662 , n94661 , n94627 );
and ( n94663 , n94660 , n94662 );
and ( n94664 , n94642 , n94659 );
or ( n94665 , n94663 , n94664 );
and ( n94666 , n94640 , n94665 );
and ( n94667 , n94637 , n94639 );
or ( n94668 , n94666 , n94667 );
not ( n94669 , n94668 );
nand ( n94670 , n94635 , n94669 );
xor ( n94671 , n87591 , n87601 );
and ( n94672 , n94671 , n87612 );
and ( n94673 , n87591 , n87601 );
or ( n94674 , n94672 , n94673 );
xor ( n94675 , n94596 , n94597 );
xor ( n94676 , n94675 , n94603 );
xor ( n94677 , n94674 , n94676 );
xor ( n94678 , n94611 , n94615 );
xor ( n94679 , n94678 , n94621 );
and ( n94680 , n94677 , n94679 );
and ( n94681 , n94674 , n94676 );
or ( n94682 , n94680 , n94681 );
xor ( n94683 , n94642 , n94659 );
xor ( n94684 , n94683 , n94662 );
xor ( n94685 , n94682 , n94684 );
xor ( n94686 , n94646 , n94651 );
xor ( n94687 , n94686 , n94656 );
xor ( n94688 , n87620 , n87624 );
and ( n94689 , n94688 , n87629 );
and ( n94690 , n87620 , n87624 );
or ( n94691 , n94689 , n94690 );
xor ( n94692 , n94687 , n94691 );
xor ( n94693 , n87545 , n87580 );
and ( n94694 , n94693 , n87613 );
and ( n94695 , n87545 , n87580 );
or ( n94696 , n94694 , n94695 );
and ( n94697 , n94692 , n94696 );
and ( n94698 , n94687 , n94691 );
or ( n94699 , n94697 , n94698 );
xor ( n94700 , n94685 , n94699 );
xor ( n94701 , n94674 , n94676 );
xor ( n94702 , n94701 , n94679 );
xor ( n94703 , n94687 , n94691 );
xor ( n94704 , n94703 , n94696 );
xor ( n94705 , n94702 , n94704 );
xor ( n94706 , n87630 , n87634 );
and ( n94707 , n94706 , n87639 );
and ( n94708 , n87630 , n87634 );
or ( n94709 , n94707 , n94708 );
and ( n94710 , n94705 , n94709 );
and ( n94711 , n94702 , n94704 );
or ( n94712 , n94710 , n94711 );
nor ( n94713 , n94700 , n94712 );
xor ( n94714 , n94637 , n94639 );
xor ( n94715 , n94714 , n94665 );
xor ( n94716 , n94682 , n94684 );
and ( n94717 , n94716 , n94699 );
and ( n94718 , n94682 , n94684 );
or ( n94719 , n94717 , n94718 );
nor ( n94720 , n94715 , n94719 );
xor ( n94721 , n94702 , n94704 );
xor ( n94722 , n94721 , n94709 );
xor ( n94723 , n87614 , n87640 );
and ( n94724 , n94723 , n87645 );
and ( n94725 , n87614 , n87640 );
or ( n94726 , n94724 , n94725 );
nor ( n94727 , n94722 , n94726 );
nor ( n94728 , n94713 , n94720 , n94727 );
nand ( n94729 , n94670 , n94728 );
xor ( n94730 , n94457 , n94560 );
and ( n94731 , n94730 , n94633 );
and ( n94732 , n94457 , n94560 );
or ( n94733 , n94731 , n94732 );
not ( n94734 , n94733 );
xor ( n94735 , n94526 , n94553 );
and ( n94736 , n94735 , n94558 );
and ( n94737 , n94526 , n94553 );
or ( n94738 , n94736 , n94737 );
xor ( n94739 , n94488 , n94504 );
and ( n94740 , n94739 , n94523 );
and ( n94741 , n94488 , n94504 );
or ( n94742 , n94740 , n94741 );
not ( n94743 , n5501 );
not ( n94744 , n537 );
not ( n94745 , n94517 );
or ( n94746 , n94744 , n94745 );
nand ( n94747 , n94516 , n5409 );
nand ( n94748 , n94746 , n94747 );
not ( n94749 , n94748 );
or ( n94750 , n94743 , n94749 );
nand ( n94751 , n94463 , n16155 );
nand ( n94752 , n94750 , n94751 );
not ( n94753 , n94422 );
nor ( n94754 , n94753 , n5409 );
xor ( n94755 , n94752 , n94754 );
not ( n94756 , n4445 );
not ( n94757 , n94502 );
or ( n94758 , n94756 , n94757 );
nand ( n94759 , n94758 , n7444 );
xor ( n94760 , n94755 , n94759 );
xor ( n94761 , n94742 , n94760 );
not ( n94762 , n4434 );
and ( n94763 , n94580 , n4251 );
not ( n94764 , n94580 );
and ( n94765 , n94764 , n539 );
or ( n94766 , n94763 , n94765 );
not ( n94767 , n94766 );
or ( n94768 , n94762 , n94767 );
nand ( n94769 , n94512 , n4224 );
nand ( n94770 , n94768 , n94769 );
not ( n94771 , n5590 );
nand ( n94772 , n541 , n9758 );
nand ( n94773 , n9757 , n5538 );
nand ( n94774 , n94772 , n94773 );
not ( n94775 , n94774 );
or ( n94776 , n94771 , n94775 );
nand ( n94777 , n9938 , n94479 );
nand ( n94778 , n94776 , n94777 );
not ( n94779 , n94778 );
xor ( n94780 , n94770 , n94779 );
xor ( n94781 , n94472 , n94483 );
and ( n94782 , n94781 , n94485 );
and ( n94783 , n94472 , n94483 );
or ( n94784 , n94782 , n94783 );
xor ( n94785 , n94780 , n94784 );
xor ( n94786 , n94761 , n94785 );
xor ( n94787 , n94738 , n94786 );
xor ( n94788 , n94486 , n94524 );
and ( n94789 , n94788 , n94559 );
and ( n94790 , n94486 , n94524 );
or ( n94791 , n94789 , n94790 );
xor ( n94792 , n94787 , n94791 );
not ( n94793 , n94792 );
nand ( n94794 , n94734 , n94793 );
xor ( n94795 , n94738 , n94786 );
and ( n94796 , n94795 , n94791 );
and ( n94797 , n94738 , n94786 );
or ( n94798 , n94796 , n94797 );
xor ( n94799 , n94770 , n94779 );
and ( n94800 , n94799 , n94784 );
and ( n94801 , n94770 , n94779 );
or ( n94802 , n94800 , n94801 );
xor ( n94803 , n94752 , n94754 );
and ( n94804 , n94803 , n94759 );
and ( n94805 , n94752 , n94754 );
or ( n94806 , n94804 , n94805 );
or ( n94807 , n4445 , n9595 );
nand ( n94808 , n94807 , n543 );
not ( n94809 , n9938 );
not ( n94810 , n94774 );
or ( n94811 , n94809 , n94810 );
not ( n94812 , n541 );
not ( n94813 , n9848 );
or ( n94814 , n94812 , n94813 );
nand ( n94815 , n94500 , n5538 );
nand ( n94816 , n94814 , n94815 );
nand ( n94817 , n94816 , n5590 );
nand ( n94818 , n94811 , n94817 );
xor ( n94819 , n94808 , n94818 );
not ( n94820 , n5501 );
not ( n94821 , n537 );
not ( n94822 , n9735 );
or ( n94823 , n94821 , n94822 );
nand ( n94824 , n94510 , n5409 );
nand ( n94825 , n94823 , n94824 );
not ( n94826 , n94825 );
or ( n94827 , n94820 , n94826 );
nand ( n94828 , n94748 , n16155 );
nand ( n94829 , n94827 , n94828 );
xor ( n94830 , n94819 , n94829 );
xor ( n94831 , n94806 , n94830 );
and ( n94832 , n94416 , n537 );
not ( n94833 , n4434 );
not ( n94834 , n539 );
not ( n94835 , n9557 );
or ( n94836 , n94834 , n94835 );
nand ( n94837 , n4251 , n94477 );
nand ( n94838 , n94836 , n94837 );
not ( n94839 , n94838 );
or ( n94840 , n94833 , n94839 );
nand ( n94841 , n94766 , n4224 );
nand ( n94842 , n94840 , n94841 );
xor ( n94843 , n94832 , n94842 );
xor ( n94844 , n94843 , n94778 );
xor ( n94845 , n94831 , n94844 );
xor ( n94846 , n94802 , n94845 );
xor ( n94847 , n94742 , n94760 );
and ( n94848 , n94847 , n94785 );
and ( n94849 , n94742 , n94760 );
or ( n94850 , n94848 , n94849 );
xor ( n94851 , n94846 , n94850 );
nor ( n94852 , n94798 , n94851 );
not ( n94853 , n94852 );
nand ( n94854 , n94794 , n94853 );
nor ( n94855 , n94729 , n94854 );
nand ( n94856 , n94368 , n94855 );
nand ( n94857 , n94634 , n94668 );
not ( n94858 , n94857 );
nand ( n94859 , n94719 , n94715 );
not ( n94860 , n94859 );
nand ( n94861 , n94722 , n94726 );
nor ( n94862 , n94700 , n94712 );
or ( n94863 , n94861 , n94862 );
nand ( n94864 , n94700 , n94712 );
nand ( n94865 , n94863 , n94864 );
not ( n94866 , n94719 );
not ( n94867 , n94715 );
nand ( n94868 , n94866 , n94867 );
nand ( n94869 , n94865 , n94868 );
not ( n94870 , n94869 );
or ( n94871 , n94860 , n94870 );
nand ( n94872 , n94635 , n94669 );
nand ( n94873 , n94871 , n94872 );
not ( n94874 , n94873 );
or ( n94875 , n94858 , n94874 );
not ( n94876 , n94854 );
nand ( n94877 , n94875 , n94876 );
nand ( n94878 , n94733 , n94792 );
nor ( n94879 , n94798 , n94851 );
or ( n94880 , n94878 , n94879 );
nand ( n94881 , n94798 , n94851 );
nand ( n94882 , n94880 , n94881 );
not ( n94883 , n94882 );
nand ( n94884 , n94856 , n94877 , n94883 );
xor ( n94885 , n94832 , n94842 );
and ( n94886 , n94885 , n94778 );
and ( n94887 , n94832 , n94842 );
or ( n94888 , n94886 , n94887 );
not ( n94889 , n7440 );
not ( n94890 , n5538 );
and ( n94891 , n94889 , n94890 );
and ( n94892 , n94816 , n9938 );
nor ( n94893 , n94891 , n94892 );
xor ( n94894 , n94808 , n94818 );
and ( n94895 , n94894 , n94829 );
and ( n94896 , n94808 , n94818 );
or ( n94897 , n94895 , n94896 );
xor ( n94898 , n94893 , n94897 );
and ( n94899 , n94516 , n537 );
not ( n94900 , n4434 );
not ( n94901 , n539 );
not ( n94902 , n9758 );
or ( n94903 , n94901 , n94902 );
nand ( n94904 , n4251 , n9757 );
nand ( n94905 , n94903 , n94904 );
not ( n94906 , n94905 );
or ( n94907 , n94900 , n94906 );
nand ( n94908 , n94838 , n4224 );
nand ( n94909 , n94907 , n94908 );
xor ( n94910 , n94899 , n94909 );
not ( n94911 , n16155 );
not ( n94912 , n94825 );
or ( n94913 , n94911 , n94912 );
xor ( n94914 , n537 , n94580 );
nand ( n94915 , n94914 , n5501 );
nand ( n94916 , n94913 , n94915 );
xor ( n94917 , n94910 , n94916 );
xor ( n94918 , n94898 , n94917 );
xor ( n94919 , n94888 , n94918 );
xor ( n94920 , n94806 , n94830 );
and ( n94921 , n94920 , n94844 );
and ( n94922 , n94806 , n94830 );
or ( n94923 , n94921 , n94922 );
xor ( n94924 , n94919 , n94923 );
xor ( n94925 , n94802 , n94845 );
and ( n94926 , n94925 , n94850 );
and ( n94927 , n94802 , n94845 );
or ( n94928 , n94926 , n94927 );
or ( n94929 , n94924 , n94928 );
nand ( n94930 , n94928 , n94924 );
nand ( n94931 , n94929 , n94930 );
not ( n94932 , n94931 );
and ( n94933 , n94884 , n94932 );
not ( n94934 , n94884 );
and ( n94935 , n94934 , n94931 );
nor ( n94936 , n94933 , n94935 );
nand ( n94937 , n94936 , n454 );
nand ( n94938 , n94352 , n94937 );
and ( n94939 , n94938 , n472 );
not ( n94940 , n10061 );
buf ( n94941 , n94256 );
nand ( n94942 , n94129 , n94169 );
not ( n94943 , n94942 );
nor ( n94944 , n94943 , n94170 );
and ( n94945 , n94941 , n94944 );
not ( n94946 , n94941 );
not ( n94947 , n94944 );
and ( n94948 , n94946 , n94947 );
nor ( n94949 , n94945 , n94948 );
not ( n94950 , n94949 );
or ( n94951 , n94940 , n94950 );
and ( n94952 , n94872 , n94857 );
not ( n94953 , n94952 );
buf ( n94954 , n94728 );
not ( n94955 , n94954 );
not ( n94956 , n94360 );
nand ( n94957 , n94956 , n94367 );
not ( n94958 , n94957 );
or ( n94959 , n94955 , n94958 );
nand ( n94960 , n94954 , n94361 );
buf ( n94961 , n94869 );
nand ( n94962 , n94960 , n94961 , n94859 );
not ( n94963 , n94962 );
nand ( n94964 , n94959 , n94963 );
not ( n94965 , n94964 );
or ( n94966 , n94953 , n94965 );
nand ( n94967 , n94957 , n94954 );
nor ( n94968 , n94962 , n94952 );
and ( n94969 , n94967 , n94968 );
not ( n94970 , n454 );
nor ( n94971 , n94969 , n94970 );
nand ( n94972 , n94966 , n94971 );
nand ( n94973 , n94951 , n94972 );
and ( n94974 , n94973 , n470 );
nor ( n94975 , n94360 , n94361 );
not ( n94976 , n94975 );
not ( n94977 , n94367 );
or ( n94978 , n94976 , n94977 );
buf ( n94979 , n94727 );
not ( n94980 , n94979 );
nand ( n94981 , n94978 , n94980 );
buf ( n94982 , n94862 );
or ( n94983 , n94981 , n94982 );
buf ( n94984 , n94865 );
not ( n94985 , n94984 );
and ( n94986 , n94719 , n94867 );
not ( n94987 , n94719 );
and ( n94988 , n94987 , n94715 );
nor ( n94989 , n94986 , n94988 );
not ( n94990 , n94989 );
and ( n94991 , n94985 , n94990 );
nand ( n94992 , n94983 , n94991 );
not ( n94993 , n94992 );
not ( n94994 , n94981 );
not ( n94995 , n94982 );
nand ( n94996 , n94995 , n94989 );
not ( n94997 , n94996 );
and ( n94998 , n94994 , n94997 );
nor ( n94999 , n94985 , n94990 );
nor ( n95000 , n94998 , n94999 );
not ( n95001 , n95000 );
or ( n95002 , n94993 , n95001 );
nand ( n95003 , n95002 , n454 );
not ( n95004 , n94238 );
or ( n95005 , n94183 , n94203 );
nand ( n95006 , n95005 , n87517 );
buf ( n95007 , n94183 );
nand ( n95008 , n95007 , n94203 );
and ( n95009 , n95006 , n95008 );
nand ( n95010 , n95004 , n95009 );
not ( n95011 , n95010 );
and ( n95012 , n94230 , n94247 );
not ( n95013 , n95012 );
nand ( n95014 , n17751 , n17755 );
nor ( n95015 , n95013 , n95014 );
nand ( n95016 , n95011 , n95015 );
buf ( n95017 , n94245 );
not ( n95018 , n95017 );
nor ( n95019 , n95018 , n95009 );
not ( n95020 , n95004 );
or ( n95021 , n95019 , n95020 );
nand ( n95022 , n95021 , n95013 );
not ( n95023 , n87520 );
not ( n95024 , n95005 );
nor ( n95025 , n95023 , n95024 );
nor ( n95026 , n95025 , n95010 );
not ( n95027 , n95004 );
nor ( n95028 , n95027 , n95017 );
or ( n95029 , n95026 , n95028 );
nand ( n95030 , n95029 , n95012 );
nand ( n95031 , n95016 , n95022 , n95030 );
nand ( n95032 , n17751 , n17755 );
and ( n95033 , n95013 , n95032 , n95025 , n95017 );
or ( n95034 , n95031 , n95033 );
nand ( n95035 , n95034 , n10061 );
and ( n95036 , n95003 , n95035 );
nor ( n95037 , n95036 , n16056 );
xor ( n95038 , n94974 , n95037 );
not ( n95039 , n10061 );
nand ( n95040 , n94041 , n94268 );
xnor ( n95041 , n94265 , n95040 );
not ( n95042 , n95041 );
or ( n95043 , n95039 , n95042 );
not ( n95044 , n94975 );
not ( n95045 , n94367 );
or ( n95046 , n95044 , n95045 );
not ( n95047 , n94733 );
nand ( n95048 , n95047 , n94793 );
buf ( n95049 , n95048 );
not ( n95050 , n95049 );
nor ( n95051 , n95050 , n94729 );
nand ( n95052 , n95046 , n95051 );
xnor ( n95053 , n94798 , n94851 );
and ( n95054 , n95053 , n454 );
or ( n95055 , n95052 , n95054 );
not ( n95056 , n94857 );
not ( n95057 , n94873 );
or ( n95058 , n95056 , n95057 );
nand ( n95059 , n95058 , n95049 );
not ( n95060 , n95059 );
not ( n95061 , n95054 );
and ( n95062 , n95060 , n95061 );
not ( n95063 , n95054 );
not ( n95064 , n94878 );
and ( n95065 , n95063 , n95064 );
nor ( n95066 , n95062 , n95065 );
not ( n95067 , n95053 );
and ( n95068 , n95067 , n454 );
nor ( n95069 , n95068 , n95064 );
nand ( n95070 , n95052 , n95059 , n95069 );
nand ( n95071 , n95055 , n95066 , n95070 );
nand ( n95072 , n95043 , n95071 );
and ( n95073 , n95072 , n472 );
and ( n95074 , n95038 , n95073 );
and ( n95075 , n94974 , n95037 );
or ( n95076 , n95074 , n95075 );
xor ( n95077 , n94939 , n95076 );
not ( n95078 , n10061 );
not ( n95079 , n94949 );
or ( n95080 , n95078 , n95079 );
nand ( n95081 , n95080 , n94972 );
and ( n95082 , n95081 , n469 );
and ( n95083 , n95072 , n471 );
xor ( n95084 , n95082 , n95083 );
not ( n95085 , n454 );
not ( n95086 , n94729 );
not ( n95087 , n95086 );
not ( n95088 , n94368 );
or ( n95089 , n95087 , n95088 );
and ( n95090 , n94873 , n94857 );
nand ( n95091 , n95089 , n95090 );
nand ( n95092 , n95049 , n94878 );
not ( n95093 , n95092 );
and ( n95094 , n95091 , n95093 );
not ( n95095 , n95091 );
and ( n95096 , n95095 , n95092 );
nor ( n95097 , n95094 , n95096 );
not ( n95098 , n95097 );
or ( n95099 , n95085 , n95098 );
not ( n95100 , n94170 );
not ( n95101 , n95100 );
not ( n95102 , n94941 );
or ( n95103 , n95101 , n95102 );
nand ( n95104 , n95103 , n94942 );
not ( n95105 , n94177 );
nand ( n95106 , n95105 , n94262 );
not ( n95107 , n95106 );
and ( n95108 , n95104 , n95107 );
not ( n95109 , n95104 );
and ( n95110 , n95109 , n95106 );
nor ( n95111 , n95108 , n95110 );
nand ( n95112 , n95111 , n10061 );
nand ( n95113 , n95099 , n95112 );
and ( n95114 , n95113 , n470 );
xor ( n95115 , n95084 , n95114 );
xor ( n95116 , n95077 , n95115 );
not ( n95117 , n95116 );
buf ( n95118 , n95113 );
and ( n95119 , n95118 , n471 );
and ( n95120 , n95081 , n471 );
not ( n95121 , n10061 );
not ( n95122 , n95025 );
not ( n95123 , n95032 );
or ( n95124 , n95122 , n95123 );
buf ( n95125 , n95009 );
nand ( n95126 , n95124 , n95125 );
and ( n95127 , n95017 , n95004 );
xor ( n95128 , n95126 , n95127 );
not ( n95129 , n95128 );
or ( n95130 , n95121 , n95129 );
buf ( n95131 , n94861 );
and ( n95132 , n94981 , n95131 );
not ( n95133 , n94982 );
buf ( n95134 , n94864 );
nand ( n95135 , n95133 , n95134 );
and ( n95136 , n95135 , n454 );
or ( n95137 , n95132 , n95136 );
not ( n95138 , n95135 );
nand ( n95139 , n95138 , n454 );
nand ( n95140 , n95139 , n94981 , n95131 );
nand ( n95141 , n95137 , n95140 );
nand ( n95142 , n95130 , n95141 );
not ( n95143 , n95142 );
nor ( n95144 , n95143 , n16056 );
xor ( n95145 , n95120 , n95144 );
nand ( n95146 , n95035 , n95003 );
not ( n95147 , n95146 );
nor ( n95148 , n95147 , n2359 );
and ( n95149 , n95145 , n95148 );
and ( n95150 , n95120 , n95144 );
or ( n95151 , n95149 , n95150 );
xor ( n95152 , n95119 , n95151 );
xor ( n95153 , n94974 , n95037 );
xor ( n95154 , n95153 , n95073 );
and ( n95155 , n95152 , n95154 );
and ( n95156 , n95119 , n95151 );
or ( n95157 , n95155 , n95156 );
not ( n95158 , n95157 );
and ( n95159 , n95117 , n95158 );
and ( n95160 , n95118 , n472 );
and ( n95161 , n94973 , n472 );
not ( n95162 , n10061 );
not ( n95163 , n87521 );
not ( n95164 , n95032 );
or ( n95165 , n95163 , n95164 );
nand ( n95166 , n95165 , n87518 );
not ( n95167 , n95008 );
nor ( n95168 , n95167 , n95024 );
xor ( n95169 , n95166 , n95168 );
not ( n95170 , n95169 );
or ( n95171 , n95162 , n95170 );
nand ( n95172 , n94980 , n94861 );
xnor ( n95173 , n94368 , n95172 );
nand ( n95174 , n95173 , n454 );
nand ( n95175 , n95171 , n95174 );
and ( n95176 , n95175 , n469 );
xor ( n95177 , n95161 , n95176 );
and ( n95178 , n95142 , n470 );
and ( n95179 , n95177 , n95178 );
and ( n95180 , n95161 , n95176 );
or ( n95181 , n95179 , n95180 );
xor ( n95182 , n95160 , n95181 );
xor ( n95183 , n95120 , n95144 );
xor ( n95184 , n95183 , n95148 );
and ( n95185 , n95182 , n95184 );
and ( n95186 , n95160 , n95181 );
or ( n95187 , n95185 , n95186 );
not ( n95188 , n95187 );
xor ( n95189 , n95119 , n95151 );
xor ( n95190 , n95189 , n95154 );
not ( n95191 , n95190 );
and ( n95192 , n95188 , n95191 );
nor ( n95193 , n95159 , n95192 );
buf ( n95194 , n95193 );
not ( n95195 , n95194 );
xor ( n95196 , n95160 , n95181 );
xor ( n95197 , n95196 , n95184 );
not ( n95198 , n95197 );
not ( n95199 , n95147 );
and ( n95200 , n95199 , n471 );
not ( n95201 , n454 );
not ( n95202 , n87660 );
or ( n95203 , n95201 , n95202 );
and ( n95204 , n95014 , n87523 );
not ( n95205 , n95014 );
and ( n95206 , n95205 , n87522 );
nor ( n95207 , n95204 , n95206 );
nand ( n95208 , n95207 , n10061 );
nand ( n95209 , n95203 , n95208 );
and ( n95210 , n95209 , n469 );
nor ( n95211 , n95143 , n17275 );
xor ( n95212 , n95210 , n95211 );
and ( n95213 , n95175 , n470 );
and ( n95214 , n95212 , n95213 );
and ( n95215 , n95210 , n95211 );
or ( n95216 , n95214 , n95215 );
xor ( n95217 , n95200 , n95216 );
xor ( n95218 , n95161 , n95176 );
xor ( n95219 , n95218 , n95178 );
and ( n95220 , n95217 , n95219 );
and ( n95221 , n95200 , n95216 );
or ( n95222 , n95220 , n95221 );
not ( n95223 , n95222 );
nand ( n95224 , n95198 , n95223 );
not ( n95225 , n95224 );
xor ( n95226 , n95200 , n95216 );
xor ( n95227 , n95226 , n95219 );
and ( n95228 , n95199 , n472 );
and ( n95229 , n95209 , n470 );
and ( n95230 , n16704 , n469 );
xor ( n95231 , n95229 , n95230 );
and ( n95232 , n95142 , n472 );
and ( n95233 , n95231 , n95232 );
and ( n95234 , n95229 , n95230 );
or ( n95235 , n95233 , n95234 );
xor ( n95236 , n95228 , n95235 );
xor ( n95237 , n95210 , n95211 );
xor ( n95238 , n95237 , n95213 );
and ( n95239 , n95236 , n95238 );
and ( n95240 , n95228 , n95235 );
or ( n95241 , n95239 , n95240 );
nor ( n95242 , n95227 , n95241 );
xor ( n95243 , n95228 , n95235 );
xor ( n95244 , n95243 , n95238 );
and ( n95245 , n95175 , n471 );
and ( n95246 , n87661 , n87528 );
not ( n95247 , n471 );
nor ( n95248 , n95246 , n95247 );
and ( n95249 , n16381 , n469 );
xor ( n95250 , n95248 , n95249 );
and ( n95251 , n16704 , n470 );
and ( n95252 , n95250 , n95251 );
and ( n95253 , n95248 , n95249 );
or ( n95254 , n95252 , n95253 );
xor ( n95255 , n95245 , n95254 );
xor ( n95256 , n95229 , n95230 );
xor ( n95257 , n95256 , n95232 );
and ( n95258 , n95255 , n95257 );
and ( n95259 , n95245 , n95254 );
or ( n95260 , n95258 , n95259 );
nand ( n95261 , n95244 , n95260 );
or ( n95262 , n95242 , n95261 );
nand ( n95263 , n95227 , n95241 );
nand ( n95264 , n95262 , n95263 );
not ( n95265 , n95264 );
or ( n95266 , n95225 , n95265 );
buf ( n95267 , n95197 );
nand ( n95268 , n95267 , n95222 );
nand ( n95269 , n95266 , n95268 );
not ( n95270 , n95269 );
not ( n95271 , n17736 );
not ( n95272 , n87358 );
nand ( n95273 , n17508 , n17525 );
nand ( n95274 , n17664 , n17629 , n95273 );
nand ( n95275 , n17628 , n95274 , n17631 , n17633 );
nand ( n95276 , n95275 , n17712 , n17689 );
not ( n95277 , n95276 );
or ( n95278 , n95272 , n95277 );
nand ( n95279 , n95278 , n16772 );
not ( n95280 , n95279 );
or ( n95281 , n95271 , n95280 );
and ( n95282 , n95175 , n472 );
xor ( n95283 , n87663 , n87664 );
and ( n95284 , n95283 , n87666 );
and ( n95285 , n87663 , n87664 );
or ( n95286 , n95284 , n95285 );
xor ( n95287 , n95282 , n95286 );
xor ( n95288 , n95248 , n95249 );
xor ( n95289 , n95288 , n95251 );
and ( n95290 , n95287 , n95289 );
and ( n95291 , n95282 , n95286 );
or ( n95292 , n95290 , n95291 );
not ( n95293 , n95292 );
not ( n95294 , n95293 );
xor ( n95295 , n95245 , n95254 );
xor ( n95296 , n95295 , n95257 );
not ( n95297 , n95296 );
not ( n95298 , n95297 );
or ( n95299 , n95294 , n95298 );
xor ( n95300 , n95282 , n95286 );
xor ( n95301 , n95300 , n95289 );
not ( n95302 , n95301 );
xor ( n95303 , n17738 , n17742 );
and ( n95304 , n95303 , n87667 );
and ( n95305 , n17738 , n17742 );
or ( n95306 , n95304 , n95305 );
not ( n95307 , n95306 );
and ( n95308 , n95302 , n95307 );
nor ( n95309 , n95308 , n87673 );
nand ( n95310 , n95299 , n95309 );
not ( n95311 , n95310 );
nand ( n95312 , n95281 , n95311 );
not ( n95313 , n95312 );
nor ( n95314 , n95301 , n95306 );
or ( n95315 , n95314 , n87676 );
nand ( n95316 , n95301 , n95306 );
nand ( n95317 , n95315 , n95316 );
nand ( n95318 , n95293 , n95297 );
and ( n95319 , n95317 , n95318 );
nand ( n95320 , n95296 , n95292 );
not ( n95321 , n95320 );
nor ( n95322 , n95319 , n95321 );
not ( n95323 , n95322 );
or ( n95324 , n95313 , n95323 );
not ( n95325 , n95227 );
not ( n95326 , n95241 );
nand ( n95327 , n95325 , n95326 );
not ( n95328 , n95244 );
not ( n95329 , n95260 );
nand ( n95330 , n95328 , n95329 );
and ( n95331 , n95327 , n95330 , n95224 );
nand ( n95332 , n95324 , n95331 );
nand ( n95333 , n95270 , n95332 );
not ( n95334 , n95333 );
or ( n95335 , n95195 , n95334 );
not ( n95336 , n95116 );
nand ( n95337 , n95336 , n95158 );
not ( n95338 , n95337 );
nand ( n95339 , n95187 , n95190 );
not ( n95340 , n95339 );
not ( n95341 , n95340 );
or ( n95342 , n95338 , n95341 );
nand ( n95343 , n95116 , n95157 );
nand ( n95344 , n95342 , n95343 );
buf ( n95345 , n95344 );
not ( n95346 , n95345 );
nand ( n95347 , n95335 , n95346 );
and ( n95348 , n94938 , n471 );
xor ( n95349 , n95082 , n95083 );
and ( n95350 , n95349 , n95114 );
and ( n95351 , n95082 , n95083 );
or ( n95352 , n95350 , n95351 );
xor ( n95353 , n95348 , n95352 );
nand ( n95354 , n93923 , n94040 );
and ( n95355 , n94178 , n95354 , n94342 );
not ( n95356 , n95355 );
not ( n95357 , n94256 );
or ( n95358 , n95356 , n95357 );
not ( n95359 , n94342 );
not ( n95360 , n95354 );
not ( n95361 , n94263 );
or ( n95362 , n95360 , n95361 );
nand ( n95363 , n95362 , n94268 );
not ( n95364 , n95363 );
or ( n95365 , n95359 , n95364 );
nand ( n95366 , n95365 , n94343 );
not ( n95367 , n95366 );
nand ( n95368 , n95358 , n95367 );
and ( n95369 , n489 , n15566 );
not ( n95370 , n95369 );
not ( n95371 , n12969 );
not ( n95372 , n94307 );
or ( n95373 , n95371 , n95372 );
nand ( n95374 , n13032 , n495 );
nand ( n95375 , n95373 , n95374 );
xor ( n95376 , n95370 , n95375 );
xor ( n95377 , n94320 , n94321 );
and ( n95378 , n95377 , n94332 );
and ( n95379 , n94320 , n94321 );
or ( n95380 , n95378 , n95379 );
xor ( n95381 , n95376 , n95380 );
xor ( n95382 , n94291 , n94301 );
and ( n95383 , n95382 , n94311 );
and ( n95384 , n94291 , n94301 );
or ( n95385 , n95383 , n95384 );
not ( n95386 , n12638 );
and ( n95387 , n15696 , n12610 );
not ( n95388 , n15696 );
and ( n95389 , n95388 , n491 );
or ( n95390 , n95387 , n95389 );
not ( n95391 , n95390 );
or ( n95392 , n95386 , n95391 );
nand ( n95393 , n12595 , n94328 );
nand ( n95394 , n95392 , n95393 );
not ( n95395 , n12542 );
not ( n95396 , n94287 );
or ( n95397 , n95395 , n95396 );
xor ( n95398 , n489 , n87441 );
nand ( n95399 , n95398 , n12795 );
nand ( n95400 , n95397 , n95399 );
xor ( n95401 , n95394 , n95400 );
not ( n95402 , n12758 );
not ( n95403 , n493 );
not ( n95404 , n16321 );
not ( n95405 , n95404 );
or ( n95406 , n95403 , n95405 );
nand ( n95407 , n16321 , n12775 );
nand ( n95408 , n95406 , n95407 );
not ( n95409 , n95408 );
or ( n95410 , n95402 , n95409 );
nand ( n95411 , n94299 , n15344 );
nand ( n95412 , n95410 , n95411 );
xor ( n95413 , n95401 , n95412 );
xor ( n95414 , n95385 , n95413 );
xor ( n95415 , n93735 , n94317 );
and ( n95416 , n95415 , n94333 );
and ( n95417 , n93735 , n94317 );
or ( n95418 , n95416 , n95417 );
xor ( n95419 , n95414 , n95418 );
xor ( n95420 , n95381 , n95419 );
xor ( n95421 , n94281 , n94312 );
and ( n95422 , n95421 , n94334 );
and ( n95423 , n94281 , n94312 );
or ( n95424 , n95422 , n95423 );
xor ( n95425 , n95420 , n95424 );
not ( n95426 , n95425 );
xor ( n95427 , n94277 , n94335 );
and ( n95428 , n95427 , n94340 );
and ( n95429 , n94277 , n94335 );
or ( n95430 , n95428 , n95429 );
not ( n95431 , n95430 );
nand ( n95432 , n95426 , n95431 );
buf ( n95433 , n95432 );
and ( n95434 , n95430 , n95425 );
not ( n95435 , n95434 );
nand ( n95436 , n95433 , n95435 );
not ( n95437 , n95436 );
and ( n95438 , n95368 , n95437 );
not ( n95439 , n95368 );
and ( n95440 , n95439 , n95436 );
nor ( n95441 , n95438 , n95440 );
nand ( n95442 , n95441 , n10061 );
not ( n95443 , n95442 );
not ( n95444 , n94929 );
not ( n95445 , n94882 );
or ( n95446 , n95444 , n95445 );
nand ( n95447 , n95446 , n94930 );
not ( n95448 , n95447 );
not ( n95449 , n95448 );
or ( n95450 , n94957 , n94361 );
or ( n95451 , n94924 , n94928 );
nand ( n95452 , n95048 , n94853 , n95451 );
nor ( n95453 , n95452 , n94729 );
nand ( n95454 , n95450 , n95453 );
not ( n95455 , n95454 );
or ( n95456 , n95449 , n95455 );
or ( n95457 , n9938 , n5590 );
nand ( n95458 , n95457 , n541 );
not ( n95459 , n4224 );
not ( n95460 , n94905 );
or ( n95461 , n95459 , n95460 );
not ( n95462 , n539 );
not ( n95463 , n9848 );
or ( n95464 , n95462 , n95463 );
not ( n95465 , n9848 );
nand ( n95466 , n95465 , n4251 );
nand ( n95467 , n95464 , n95466 );
nand ( n95468 , n95467 , n4434 );
nand ( n95469 , n95461 , n95468 );
xor ( n95470 , n95458 , n95469 );
nor ( n95471 , n9735 , n5409 );
xor ( n95472 , n95470 , n95471 );
not ( n95473 , n5501 );
xor ( n95474 , n94477 , n537 );
not ( n95475 , n95474 );
or ( n95476 , n95473 , n95475 );
nand ( n95477 , n94914 , n16155 );
nand ( n95478 , n95476 , n95477 );
not ( n95479 , n94893 );
xor ( n95480 , n95478 , n95479 );
xor ( n95481 , n94899 , n94909 );
and ( n95482 , n95481 , n94916 );
and ( n95483 , n94899 , n94909 );
or ( n95484 , n95482 , n95483 );
xor ( n95485 , n95480 , n95484 );
xor ( n95486 , n95472 , n95485 );
xor ( n95487 , n94893 , n94897 );
and ( n95488 , n95487 , n94917 );
and ( n95489 , n94893 , n94897 );
or ( n95490 , n95488 , n95489 );
xor ( n95491 , n95486 , n95490 );
xor ( n95492 , n94888 , n94918 );
and ( n95493 , n95492 , n94923 );
and ( n95494 , n94888 , n94918 );
or ( n95495 , n95493 , n95494 );
and ( n95496 , n95491 , n95495 );
not ( n95497 , n95496 );
nor ( n95498 , n95495 , n95491 );
not ( n95499 , n95498 );
and ( n95500 , n95497 , n95499 );
nand ( n95501 , n95456 , n95500 );
not ( n95502 , n94857 );
not ( n95503 , n94873 );
or ( n95504 , n95502 , n95503 );
not ( n95505 , n95452 );
nand ( n95506 , n95504 , n95505 );
not ( n95507 , n95500 );
or ( n95508 , n95506 , n95507 );
nand ( n95509 , n95508 , n454 );
not ( n95510 , n95509 );
nor ( n95511 , n95447 , n95500 );
nand ( n95512 , n95454 , n95506 , n95511 );
nand ( n95513 , n95501 , n95510 , n95512 );
not ( n95514 , n95513 );
or ( n95515 , n95443 , n95514 );
nand ( n95516 , n95515 , n472 );
not ( n95517 , n95516 );
and ( n95518 , n95113 , n469 );
xor ( n95519 , n95517 , n95518 );
and ( n95520 , n95072 , n470 );
xor ( n95521 , n95519 , n95520 );
xor ( n95522 , n95353 , n95521 );
xor ( n95523 , n94939 , n95076 );
and ( n95524 , n95523 , n95115 );
and ( n95525 , n94939 , n95076 );
or ( n95526 , n95524 , n95525 );
or ( n95527 , n95522 , n95526 );
nand ( n95528 , n95522 , n95526 );
nand ( n95529 , n95527 , n95528 );
and ( n95530 , n95347 , n95529 );
nand ( n95531 , n95333 , n95194 );
nor ( n95532 , n95529 , n95345 );
and ( n95533 , n95531 , n95532 );
nor ( n95534 , n95530 , n95533 );
or ( n95535 , n95534 , n87684 );
not ( n95536 , n90370 );
not ( n95537 , n90555 );
or ( n95538 , n95536 , n95537 );
nand ( n95539 , n90690 , n90722 );
nand ( n95540 , n95538 , n95539 );
not ( n95541 , n95540 );
not ( n95542 , n90324 );
not ( n95543 , n90305 );
not ( n95544 , n90815 );
or ( n95545 , n95543 , n95544 );
nand ( n95546 , n90814 , n90321 );
nand ( n95547 , n95545 , n95546 );
not ( n95548 , n95547 );
or ( n95549 , n95542 , n95548 );
not ( n95550 , n90305 );
not ( n95551 , n90873 );
or ( n95552 , n95550 , n95551 );
nand ( n95553 , n90870 , n90321 );
nand ( n95554 , n95552 , n95553 );
nand ( n95555 , n95554 , n90279 );
nand ( n95556 , n95549 , n95555 );
xor ( n95557 , n95541 , n95556 );
not ( n95558 , n90405 );
not ( n95559 , n90407 );
not ( n95560 , n90858 );
or ( n95561 , n95559 , n95560 );
nand ( n95562 , n90855 , n90422 );
nand ( n95563 , n95561 , n95562 );
not ( n95564 , n95563 );
or ( n95565 , n95558 , n95564 );
not ( n95566 , n90407 );
not ( n95567 , n90577 );
or ( n95568 , n95566 , n95567 );
nand ( n95569 , n90576 , n90422 );
nand ( n95570 , n95568 , n95569 );
nand ( n95571 , n95570 , n90442 );
nand ( n95572 , n95565 , n95571 );
xor ( n95573 , n95557 , n95572 );
not ( n95574 , n90840 );
not ( n95575 , n90844 );
not ( n95576 , n90135 );
or ( n95577 , n87716 , n87826 );
nand ( n95578 , n95577 , n87718 );
or ( n95579 , n90128 , n87918 );
and ( n95580 , n87857 , n87922 );
and ( n95581 , n88115 , n87921 );
nor ( n95582 , n95580 , n95581 );
or ( n95583 , n95582 , n87966 );
nand ( n95584 , n95579 , n95583 );
xor ( n95585 , n95578 , n95584 );
nor ( n95586 , n87998 , n87921 );
xor ( n95587 , n95585 , n95586 );
xor ( n95588 , n95576 , n95587 );
xor ( n95589 , n90130 , n90131 );
and ( n95590 , n95589 , n90135 );
and ( n95591 , n90130 , n90131 );
or ( n95592 , n95590 , n95591 );
and ( n95593 , n95588 , n95592 );
and ( n95594 , n95576 , n95587 );
or ( n95595 , n95593 , n95594 );
nor ( n95596 , n88094 , n87921 );
not ( n95597 , n95582 );
and ( n95598 , n95597 , n87919 );
and ( n95599 , n87967 , n87922 );
nor ( n95600 , n95598 , n95599 );
xor ( n95601 , n95596 , n95600 );
xor ( n95602 , n95578 , n95584 );
and ( n95603 , n95602 , n95586 );
and ( n95604 , n95578 , n95584 );
or ( n95605 , n95603 , n95604 );
xor ( n95606 , n95601 , n95605 );
or ( n95607 , n95595 , n95606 );
nand ( n95608 , n95595 , n95606 );
nand ( n95609 , n95607 , n95608 );
not ( n95610 , n95609 );
not ( n95611 , n95610 );
nand ( n95612 , n90143 , n90092 );
nor ( n95613 , n88321 , n95612 );
nand ( n95614 , n88276 , n95613 );
nor ( n95615 , n90035 , n95614 );
not ( n95616 , n95615 );
not ( n95617 , n90008 );
or ( n95618 , n95616 , n95617 );
or ( n95619 , n90044 , n88277 );
nand ( n95620 , n95619 , n90048 );
buf ( n95621 , n95613 );
and ( n95622 , n95620 , n95621 );
not ( n95623 , n90143 );
not ( n95624 , n90092 );
or ( n95625 , n90050 , n95624 );
nand ( n95626 , n95625 , n90093 );
not ( n95627 , n95626 );
or ( n95628 , n95623 , n95627 );
nand ( n95629 , n95628 , n90144 );
nor ( n95630 , n95622 , n95629 );
nand ( n95631 , n95618 , n95630 );
xor ( n95632 , n90122 , n90136 );
and ( n95633 , n95632 , n90141 );
and ( n95634 , n90122 , n90136 );
or ( n95635 , n95633 , n95634 );
xor ( n95636 , n95576 , n95587 );
xor ( n95637 , n95636 , n95592 );
or ( n95638 , n95635 , n95637 );
and ( n95639 , n95631 , n95638 );
and ( n95640 , n95635 , n95637 );
nor ( n95641 , n95639 , n95640 );
not ( n95642 , n95641 );
or ( n95643 , n95611 , n95642 );
not ( n95644 , n95641 );
nand ( n95645 , n95644 , n95609 );
nand ( n95646 , n95643 , n95645 );
not ( n95647 , n95646 );
not ( n95648 , n95647 );
or ( n95649 , n95575 , n95648 );
not ( n95650 , n95610 );
not ( n95651 , n95641 );
or ( n95652 , n95650 , n95651 );
nand ( n95653 , n95652 , n95645 );
nand ( n95654 , n95653 , n90843 );
nand ( n95655 , n95649 , n95654 );
not ( n95656 , n95655 );
or ( n95657 , n95574 , n95656 );
and ( n95658 , n95638 , n95607 );
not ( n95659 , n95658 );
not ( n95660 , n95631 );
or ( n95661 , n95659 , n95660 );
and ( n95662 , n95607 , n95640 );
not ( n95663 , n95608 );
nor ( n95664 , n95662 , n95663 );
nand ( n95665 , n95661 , n95664 );
xor ( n95666 , n95596 , n95600 );
and ( n95667 , n95666 , n95605 );
and ( n95668 , n95596 , n95600 );
or ( n95669 , n95667 , n95668 );
or ( n95670 , n87919 , n87967 );
nand ( n95671 , n95670 , n87922 );
nor ( n95672 , n87857 , n87921 );
xor ( n95673 , n95671 , n95672 );
not ( n95674 , n95600 );
xor ( n95675 , n95673 , n95674 );
xor ( n95676 , n95669 , n95675 );
xor ( n95677 , n95665 , n95676 );
buf ( n95678 , n95677 );
and ( n95679 , n90844 , n95678 );
not ( n95680 , n90844 );
not ( n95681 , n95677 );
and ( n95682 , n95680 , n95681 );
nor ( n95683 , n95679 , n95682 );
nand ( n95684 , n95683 , n90876 );
nand ( n95685 , n95657 , n95684 );
not ( n95686 , n90680 );
and ( n95687 , n90660 , n91071 );
not ( n95688 , n90660 );
and ( n95689 , n95688 , n91068 );
nor ( n95690 , n95687 , n95689 );
not ( n95691 , n95690 );
or ( n95692 , n95686 , n95691 );
and ( n95693 , n90660 , n90099 );
not ( n95694 , n90660 );
and ( n95695 , n95694 , n90102 );
nor ( n95696 , n95693 , n95695 );
nand ( n95697 , n95696 , n91011 );
nand ( n95698 , n95692 , n95697 );
xor ( n95699 , n95685 , n95698 );
not ( n95700 , n90582 );
not ( n95701 , n90540 );
not ( n95702 , n95640 );
nand ( n95703 , n95702 , n95638 );
and ( n95704 , n95631 , n95703 );
not ( n95705 , n95631 );
not ( n95706 , n95703 );
and ( n95707 , n95705 , n95706 );
or ( n95708 , n95704 , n95707 );
not ( n95709 , n95708 );
not ( n95710 , n95709 );
or ( n95711 , n95701 , n95710 );
nand ( n95712 , n95708 , n90539 );
nand ( n95713 , n95711 , n95712 );
not ( n95714 , n95713 );
or ( n95715 , n95700 , n95714 );
and ( n95716 , n90890 , n90151 );
not ( n95717 , n90890 );
and ( n95718 , n95717 , n90154 );
nor ( n95719 , n95716 , n95718 );
nand ( n95720 , n95719 , n90537 );
nand ( n95721 , n95715 , n95720 );
and ( n95722 , n95699 , n95721 );
and ( n95723 , n95685 , n95698 );
or ( n95724 , n95722 , n95723 );
xor ( n95725 , n95573 , n95724 );
not ( n95726 , n90844 );
not ( n95727 , n90876 );
or ( n95728 , n95726 , n95727 );
nand ( n95729 , n95683 , n90840 );
nand ( n95730 , n95728 , n95729 );
not ( n95731 , n90722 );
not ( n95732 , n90669 );
or ( n95733 , n95731 , n95732 );
nand ( n95734 , n90690 , n90370 );
nand ( n95735 , n95733 , n95734 );
or ( n95736 , n90825 , n90782 );
nand ( n95737 , n95736 , n90788 );
or ( n95738 , n95735 , n95737 );
not ( n95739 , n95738 );
not ( n95740 , n90405 );
not ( n95741 , n95570 );
or ( n95742 , n95740 , n95741 );
not ( n95743 , n90407 );
not ( n95744 , n90552 );
or ( n95745 , n95743 , n95744 );
nand ( n95746 , n90555 , n90422 );
nand ( n95747 , n95745 , n95746 );
nand ( n95748 , n95747 , n90442 );
nand ( n95749 , n95742 , n95748 );
not ( n95750 , n95749 );
or ( n95751 , n95739 , n95750 );
nand ( n95752 , n95735 , n95737 );
nand ( n95753 , n95751 , n95752 );
xor ( n95754 , n95730 , n95753 );
not ( n95755 , n90657 );
not ( n95756 , n90612 );
not ( n95757 , n90796 );
or ( n95758 , n95756 , n95757 );
nand ( n95759 , n90795 , n90630 );
nand ( n95760 , n95758 , n95759 );
not ( n95761 , n95760 );
or ( n95762 , n95755 , n95761 );
and ( n95763 , n90612 , n91071 );
not ( n95764 , n90612 );
and ( n95765 , n95764 , n91068 );
nor ( n95766 , n95763 , n95765 );
nand ( n95767 , n95766 , n90610 );
nand ( n95768 , n95762 , n95767 );
xor ( n95769 , n95754 , n95768 );
xor ( n95770 , n95725 , n95769 );
not ( n95771 , n91011 );
and ( n95772 , n90660 , n90151 );
not ( n95773 , n90660 );
and ( n95774 , n95773 , n90154 );
nor ( n95775 , n95772 , n95774 );
not ( n95776 , n95775 );
or ( n95777 , n95771 , n95776 );
nand ( n95778 , n95696 , n90680 );
nand ( n95779 , n95777 , n95778 );
not ( n95780 , n90582 );
and ( n95781 , n90890 , n95646 );
not ( n95782 , n90890 );
and ( n95783 , n95782 , n95647 );
nor ( n95784 , n95781 , n95783 );
not ( n95785 , n95784 );
or ( n95786 , n95780 , n95785 );
nand ( n95787 , n95713 , n90537 );
nand ( n95788 , n95786 , n95787 );
xor ( n95789 , n95779 , n95788 );
and ( n95790 , n90669 , n90370 );
and ( n95791 , n90622 , n90722 );
nor ( n95792 , n95790 , n95791 );
not ( n95793 , n95792 );
not ( n95794 , n90610 );
not ( n95795 , n95760 );
or ( n95796 , n95794 , n95795 );
not ( n95797 , n90612 );
not ( n95798 , n90815 );
or ( n95799 , n95797 , n95798 );
nand ( n95800 , n90814 , n90630 );
nand ( n95801 , n95799 , n95800 );
nand ( n95802 , n95801 , n90656 );
nand ( n95803 , n95796 , n95802 );
xor ( n95804 , n95793 , n95803 );
not ( n95805 , n90324 );
not ( n95806 , n95554 );
or ( n95807 , n95805 , n95806 );
not ( n95808 , n90305 );
not ( n95809 , n90858 );
or ( n95810 , n95808 , n95809 );
nand ( n95811 , n90855 , n90321 );
nand ( n95812 , n95810 , n95811 );
nand ( n95813 , n95812 , n90279 );
nand ( n95814 , n95807 , n95813 );
and ( n95815 , n95804 , n95814 );
and ( n95816 , n95793 , n95803 );
or ( n95817 , n95815 , n95816 );
xor ( n95818 , n95789 , n95817 );
and ( n95819 , n90622 , n90370 );
and ( n95820 , n90646 , n90722 );
nor ( n95821 , n95819 , n95820 );
and ( n95822 , n87701 , n92472 );
nor ( n95823 , n95822 , n87705 );
nand ( n95824 , n95821 , n95823 );
xor ( n95825 , n95824 , n95792 );
not ( n95826 , n90405 );
not ( n95827 , n95747 );
or ( n95828 , n95826 , n95827 );
not ( n95829 , n90683 );
not ( n95830 , n90422 );
and ( n95831 , n95829 , n95830 );
not ( n95832 , n95829 );
not ( n95833 , n90407 );
and ( n95834 , n95832 , n95833 );
or ( n95835 , n95831 , n95834 );
and ( n95836 , n90685 , n95835 );
not ( n95837 , n90685 );
not ( n95838 , n90422 );
and ( n95839 , n90683 , n95838 );
not ( n95840 , n90683 );
not ( n95841 , n90407 );
and ( n95842 , n95840 , n95841 );
or ( n95843 , n95839 , n95842 );
and ( n95844 , n95837 , n95843 );
or ( n95845 , n95836 , n95844 );
nand ( n95846 , n95845 , n90442 );
nand ( n95847 , n95828 , n95846 );
and ( n95848 , n95825 , n95847 );
and ( n95849 , n95824 , n95792 );
or ( n95850 , n95848 , n95849 );
xor ( n95851 , n95735 , n95737 );
xor ( n95852 , n95749 , n95851 );
xor ( n95853 , n95850 , n95852 );
xor ( n95854 , n95793 , n95803 );
xor ( n95855 , n95854 , n95814 );
and ( n95856 , n95853 , n95855 );
and ( n95857 , n95850 , n95852 );
or ( n95858 , n95856 , n95857 );
xor ( n95859 , n95818 , n95858 );
not ( n95860 , n90610 );
not ( n95861 , n95801 );
or ( n95862 , n95860 , n95861 );
and ( n95863 , n90869 , n90612 );
not ( n95864 , n90869 );
and ( n95865 , n95864 , n90630 );
nor ( n95866 , n95863 , n95865 );
nand ( n95867 , n95866 , n90657 );
nand ( n95868 , n95862 , n95867 );
not ( n95869 , n90324 );
not ( n95870 , n95812 );
or ( n95871 , n95869 , n95870 );
not ( n95872 , n90305 );
not ( n95873 , n90577 );
or ( n95874 , n95872 , n95873 );
nand ( n95875 , n90576 , n90321 );
nand ( n95876 , n95874 , n95875 );
nand ( n95877 , n95876 , n90279 );
nand ( n95878 , n95871 , n95877 );
xor ( n95879 , n95868 , n95878 );
not ( n95880 , n90680 );
not ( n95881 , n90660 );
not ( n95882 , n90796 );
or ( n95883 , n95881 , n95882 );
nand ( n95884 , n90795 , n91164 );
nand ( n95885 , n95883 , n95884 );
not ( n95886 , n95885 );
or ( n95887 , n95880 , n95886 );
nand ( n95888 , n95690 , n91011 );
nand ( n95889 , n95887 , n95888 );
and ( n95890 , n95879 , n95889 );
and ( n95891 , n95868 , n95878 );
or ( n95892 , n95890 , n95891 );
or ( n95893 , n95821 , n95823 );
nand ( n95894 , n95893 , n95824 );
not ( n95895 , n90442 );
not ( n95896 , n90407 );
not ( n95897 , n90672 );
or ( n95898 , n95896 , n95897 );
nand ( n95899 , n90669 , n90422 );
nand ( n95900 , n95898 , n95899 );
not ( n95901 , n95900 );
or ( n95902 , n95895 , n95901 );
nand ( n95903 , n95845 , n90405 );
nand ( n95904 , n95902 , n95903 );
xor ( n95905 , n95894 , n95904 );
not ( n95906 , n90279 );
not ( n95907 , n90286 );
not ( n95908 , n90552 );
or ( n95909 , n95907 , n95908 );
or ( n95910 , n90552 , n90286 );
nand ( n95911 , n95909 , n95910 );
not ( n95912 , n95911 );
or ( n95913 , n95906 , n95912 );
nand ( n95914 , n95876 , n90324 );
nand ( n95915 , n95913 , n95914 );
and ( n95916 , n95905 , n95915 );
and ( n95917 , n95894 , n95904 );
or ( n95918 , n95916 , n95917 );
not ( n95919 , n90825 );
not ( n95920 , n90788 );
not ( n95921 , n95681 );
or ( n95922 , n95920 , n95921 );
nand ( n95923 , n95678 , n90801 );
nand ( n95924 , n95922 , n95923 );
not ( n95925 , n95924 );
or ( n95926 , n95919 , n95925 );
nand ( n95927 , n90782 , n90788 );
nand ( n95928 , n95926 , n95927 );
xor ( n95929 , n95918 , n95928 );
and ( n95930 , n90844 , n95708 );
not ( n95931 , n90844 );
and ( n95932 , n95931 , n95709 );
nor ( n95933 , n95930 , n95932 );
not ( n95934 , n95933 );
not ( n95935 , n90840 );
or ( n95936 , n95934 , n95935 );
not ( n95937 , n95655 );
or ( n95938 , n95937 , n90838 );
nand ( n95939 , n95936 , n95938 );
and ( n95940 , n95929 , n95939 );
and ( n95941 , n95918 , n95928 );
or ( n95942 , n95940 , n95941 );
xor ( n95943 , n95892 , n95942 );
xor ( n95944 , n95685 , n95698 );
xor ( n95945 , n95944 , n95721 );
and ( n95946 , n95943 , n95945 );
and ( n95947 , n95892 , n95942 );
or ( n95948 , n95946 , n95947 );
xor ( n95949 , n95859 , n95948 );
xor ( n95950 , n95770 , n95949 );
xor ( n95951 , n95850 , n95852 );
xor ( n95952 , n95951 , n95855 );
not ( n95953 , n90582 );
not ( n95954 , n95719 );
or ( n95955 , n95953 , n95954 );
and ( n95956 , n90890 , n90099 );
not ( n95957 , n90890 );
and ( n95958 , n95957 , n90102 );
nor ( n95959 , n95956 , n95958 );
nand ( n95960 , n95959 , n90537 );
nand ( n95961 , n95955 , n95960 );
not ( n95962 , n95961 );
not ( n95963 , n90370 );
not ( n95964 , n90646 );
or ( n95965 , n95963 , n95964 );
or ( n95966 , n90318 , n90387 );
nand ( n95967 , n95965 , n95966 );
not ( n95968 , n90405 );
not ( n95969 , n95900 );
or ( n95970 , n95968 , n95969 );
not ( n95971 , n90407 );
not ( n95972 , n90623 );
or ( n95973 , n95971 , n95972 );
nand ( n95974 , n90629 , n90422 );
nand ( n95975 , n95973 , n95974 );
nand ( n95976 , n95975 , n90442 );
nand ( n95977 , n95970 , n95976 );
and ( n95978 , n95967 , n95977 );
not ( n95979 , n90656 );
not ( n95980 , n90612 );
not ( n95981 , n90858 );
or ( n95982 , n95980 , n95981 );
nand ( n95983 , n90855 , n90630 );
nand ( n95984 , n95982 , n95983 );
not ( n95985 , n95984 );
or ( n95986 , n95979 , n95985 );
nand ( n95987 , n95866 , n90610 );
nand ( n95988 , n95986 , n95987 );
xor ( n95989 , n95978 , n95988 );
not ( n95990 , n91011 );
not ( n95991 , n95885 );
or ( n95992 , n95990 , n95991 );
not ( n95993 , n90660 );
not ( n95994 , n90815 );
or ( n95995 , n95993 , n95994 );
nand ( n95996 , n90814 , n91164 );
nand ( n95997 , n95995 , n95996 );
nand ( n95998 , n95997 , n90680 );
nand ( n95999 , n95992 , n95998 );
and ( n96000 , n95989 , n95999 );
and ( n96001 , n95978 , n95988 );
or ( n96002 , n96000 , n96001 );
not ( n96003 , n96002 );
or ( n96004 , n95962 , n96003 );
or ( n96005 , n96002 , n95961 );
xor ( n96006 , n95824 , n95792 );
xor ( n96007 , n96006 , n95847 );
nand ( n96008 , n96005 , n96007 );
nand ( n96009 , n96004 , n96008 );
xor ( n96010 , n95952 , n96009 );
xor ( n96011 , n95892 , n95942 );
xor ( n96012 , n96011 , n95945 );
and ( n96013 , n96010 , n96012 );
and ( n96014 , n95952 , n96009 );
or ( n96015 , n96013 , n96014 );
xor ( n96016 , n95950 , n96015 );
xor ( n96017 , n95952 , n96009 );
xor ( n96018 , n96017 , n96012 );
xor ( n96019 , n95868 , n95878 );
xor ( n96020 , n96019 , n95889 );
not ( n96021 , n90825 );
not ( n96022 , n90788 );
not ( n96023 , n95647 );
or ( n96024 , n96022 , n96023 );
nand ( n96025 , n95653 , n90801 );
nand ( n96026 , n96024 , n96025 );
not ( n96027 , n96026 );
or ( n96028 , n96021 , n96027 );
nand ( n96029 , n95924 , n90782 );
nand ( n96030 , n96028 , n96029 );
not ( n96031 , n90876 );
not ( n96032 , n95933 );
or ( n96033 , n96031 , n96032 );
not ( n96034 , n90844 );
not ( n96035 , n90154 );
or ( n96036 , n96034 , n96035 );
nand ( n96037 , n90151 , n90843 );
nand ( n96038 , n96036 , n96037 );
nand ( n96039 , n96038 , n90840 );
nand ( n96040 , n96033 , n96039 );
xor ( n96041 , n96030 , n96040 );
not ( n96042 , n90537 );
and ( n96043 , n90890 , n91071 );
not ( n96044 , n90890 );
and ( n96045 , n96044 , n91068 );
nor ( n96046 , n96043 , n96045 );
not ( n96047 , n96046 );
or ( n96048 , n96042 , n96047 );
nand ( n96049 , n95959 , n90582 );
nand ( n96050 , n96048 , n96049 );
and ( n96051 , n96041 , n96050 );
and ( n96052 , n96030 , n96040 );
or ( n96053 , n96051 , n96052 );
xor ( n96054 , n96020 , n96053 );
xor ( n96055 , n95918 , n95928 );
xor ( n96056 , n96055 , n95939 );
and ( n96057 , n96054 , n96056 );
and ( n96058 , n96020 , n96053 );
or ( n96059 , n96057 , n96058 );
or ( n96060 , n96018 , n96059 );
and ( n96061 , n95961 , n96007 );
not ( n96062 , n95961 );
not ( n96063 , n96007 );
and ( n96064 , n96062 , n96063 );
or ( n96065 , n96061 , n96064 );
xor ( n96066 , n96002 , n96065 );
not ( n96067 , n96066 );
not ( n96068 , n96067 );
xor ( n96069 , n96020 , n96053 );
xor ( n96070 , n96069 , n96056 );
not ( n96071 , n96070 );
or ( n96072 , n96068 , n96071 );
or ( n96073 , n96070 , n96067 );
xor ( n96074 , n95894 , n95904 );
xor ( n96075 , n96074 , n95915 );
xor ( n96076 , n95967 , n95977 );
buf ( n96077 , n96076 );
not ( n96078 , n96077 );
not ( n96079 , n90370 );
not ( n96080 , n90765 );
or ( n96081 , n96079 , n96080 );
or ( n96082 , n90300 , n90387 );
nand ( n96083 , n96081 , n96082 );
not ( n96084 , n90405 );
not ( n96085 , n95975 );
or ( n96086 , n96084 , n96085 );
and ( n96087 , n90407 , n90646 );
not ( n96088 , n90407 );
and ( n96089 , n96088 , n90649 );
nor ( n96090 , n96087 , n96089 );
nand ( n96091 , n96090 , n90442 );
nand ( n96092 , n96086 , n96091 );
and ( n96093 , n96083 , n96092 );
buf ( n96094 , n96093 );
not ( n96095 , n96094 );
or ( n96096 , n96078 , n96095 );
not ( n96097 , n96094 );
not ( n96098 , n96097 );
not ( n96099 , n96077 );
not ( n96100 , n96099 );
or ( n96101 , n96098 , n96100 );
and ( n96102 , n90305 , n90690 );
not ( n96103 , n90305 );
and ( n96104 , n96103 , n90693 );
nor ( n96105 , n96102 , n96104 );
and ( n96106 , n96105 , n90279 );
and ( n96107 , n95911 , n90248 );
nor ( n96108 , n96106 , n96107 );
not ( n96109 , n96108 );
nand ( n96110 , n96101 , n96109 );
nand ( n96111 , n96096 , n96110 );
xor ( n96112 , n96075 , n96111 );
not ( n96113 , n90680 );
and ( n96114 , n90660 , n90870 );
not ( n96115 , n90660 );
and ( n96116 , n96115 , n90873 );
nor ( n96117 , n96114 , n96116 );
not ( n96118 , n96117 );
or ( n96119 , n96113 , n96118 );
nand ( n96120 , n95997 , n91011 );
nand ( n96121 , n96119 , n96120 );
not ( n96122 , n95984 );
or ( n96123 , n96122 , n90609 );
not ( n96124 , n90612 );
not ( n96125 , n90577 );
or ( n96126 , n96124 , n96125 );
nand ( n96127 , n90576 , n90630 );
nand ( n96128 , n96126 , n96127 );
nand ( n96129 , n96128 , n90656 );
nand ( n96130 , n96123 , n96129 );
xor ( n96131 , n96121 , n96130 );
xor ( n96132 , n96083 , n96092 );
not ( n96133 , n90370 );
not ( n96134 , n90297 );
or ( n96135 , n96133 , n96134 );
or ( n96136 , n90464 , n90387 );
nand ( n96137 , n96135 , n96136 );
not ( n96138 , n90405 );
not ( n96139 , n96090 );
or ( n96140 , n96138 , n96139 );
not ( n96141 , n90407 );
not ( n96142 , n90318 );
or ( n96143 , n96141 , n96142 );
nand ( n96144 , n90765 , n90422 );
nand ( n96145 , n96143 , n96144 );
nand ( n96146 , n96145 , n90442 );
nand ( n96147 , n96140 , n96146 );
and ( n96148 , n96137 , n96147 );
xor ( n96149 , n96132 , n96148 );
not ( n96150 , n90279 );
not ( n96151 , n90305 );
not ( n96152 , n90672 );
or ( n96153 , n96151 , n96152 );
nand ( n96154 , n90669 , n90321 );
nand ( n96155 , n96153 , n96154 );
not ( n96156 , n96155 );
or ( n96157 , n96150 , n96156 );
nand ( n96158 , n96105 , n90324 );
nand ( n96159 , n96157 , n96158 );
and ( n96160 , n96149 , n96159 );
and ( n96161 , n96132 , n96148 );
or ( n96162 , n96160 , n96161 );
and ( n96163 , n96131 , n96162 );
and ( n96164 , n96121 , n96130 );
or ( n96165 , n96163 , n96164 );
and ( n96166 , n96112 , n96165 );
and ( n96167 , n96075 , n96111 );
or ( n96168 , n96166 , n96167 );
nand ( n96169 , n96073 , n96168 );
nand ( n96170 , n96072 , n96169 );
nand ( n96171 , n96060 , n96170 );
nand ( n96172 , n96018 , n96059 );
nand ( n96173 , n96171 , n96172 );
or ( n96174 , n96016 , n96173 );
nand ( n96175 , n96016 , n96173 );
nand ( n96176 , n96174 , n96175 );
not ( n96177 , n90582 );
not ( n96178 , n90540 );
not ( n96179 , n90796 );
or ( n96180 , n96178 , n96179 );
nand ( n96181 , n90795 , n90539 );
nand ( n96182 , n96180 , n96181 );
not ( n96183 , n96182 );
or ( n96184 , n96177 , n96183 );
not ( n96185 , n90540 );
not ( n96186 , n90815 );
or ( n96187 , n96185 , n96186 );
nand ( n96188 , n90814 , n90539 );
nand ( n96189 , n96187 , n96188 );
nand ( n96190 , n96189 , n90537 );
nand ( n96191 , n96184 , n96190 );
not ( n96192 , n87689 );
not ( n96193 , n87706 );
not ( n96194 , n95681 );
or ( n96195 , n96193 , n96194 );
nand ( n96196 , n95678 , n87705 );
nand ( n96197 , n96195 , n96196 );
not ( n96198 , n96197 );
or ( n96199 , n96192 , n96198 );
not ( n96200 , n87706 );
not ( n96201 , n95647 );
or ( n96202 , n96200 , n96201 );
nand ( n96203 , n95653 , n87705 );
nand ( n96204 , n96202 , n96203 );
nand ( n96205 , n96204 , n87702 );
nand ( n96206 , n96199 , n96205 );
xor ( n96207 , n96191 , n96206 );
not ( n96208 , n90825 );
and ( n96209 , n90801 , n90154 );
not ( n96210 , n90801 );
and ( n96211 , n96210 , n90151 );
or ( n96212 , n96209 , n96211 );
not ( n96213 , n96212 );
not ( n96214 , n96213 );
or ( n96215 , n96208 , n96214 );
not ( n96216 , n90788 );
not ( n96217 , n95709 );
or ( n96218 , n96216 , n96217 );
nand ( n96219 , n95708 , n90801 );
nand ( n96220 , n96218 , n96219 );
nand ( n96221 , n96220 , n90782 );
nand ( n96222 , n96215 , n96221 );
and ( n96223 , n96207 , n96222 );
and ( n96224 , n96191 , n96206 );
or ( n96225 , n96223 , n96224 );
xor ( n96226 , n96121 , n96130 );
xor ( n96227 , n96226 , n96162 );
xor ( n96228 , n96225 , n96227 );
not ( n96229 , n90582 );
not ( n96230 , n96046 );
or ( n96231 , n96229 , n96230 );
nand ( n96232 , n96182 , n90537 );
nand ( n96233 , n96231 , n96232 );
not ( n96234 , n90825 );
not ( n96235 , n96220 );
or ( n96236 , n96234 , n96235 );
nand ( n96237 , n96026 , n90782 );
nand ( n96238 , n96236 , n96237 );
xor ( n96239 , n96233 , n96238 );
not ( n96240 , n87706 );
not ( n96241 , n87689 );
or ( n96242 , n96240 , n96241 );
not ( n96243 , n96197 );
or ( n96244 , n96243 , n87701 );
nand ( n96245 , n96242 , n96244 );
xor ( n96246 , n96239 , n96245 );
xor ( n96247 , n96228 , n96246 );
xor ( n96248 , n96132 , n96148 );
xor ( n96249 , n96248 , n96159 );
not ( n96250 , n90840 );
not ( n96251 , n90844 );
not ( n96252 , n91068 );
or ( n96253 , n96251 , n96252 );
nand ( n96254 , n91071 , n90843 );
nand ( n96255 , n96253 , n96254 );
not ( n96256 , n96255 );
or ( n96257 , n96250 , n96256 );
not ( n96258 , n90844 );
not ( n96259 , n90102 );
or ( n96260 , n96258 , n96259 );
nand ( n96261 , n90099 , n90843 );
nand ( n96262 , n96260 , n96261 );
nand ( n96263 , n96262 , n90876 );
nand ( n96264 , n96257 , n96263 );
xor ( n96265 , n96249 , n96264 );
not ( n96266 , n91110 );
nor ( n96267 , n96266 , n91115 );
not ( n96268 , n90324 );
not ( n96269 , n90321 );
not ( n96270 , n90622 );
or ( n96271 , n96269 , n96270 );
nand ( n96272 , n90623 , n90305 );
nand ( n96273 , n96271 , n96272 );
not ( n96274 , n96273 );
or ( n96275 , n96268 , n96274 );
nand ( n96276 , n91094 , n90279 );
nand ( n96277 , n96275 , n96276 );
xor ( n96278 , n96267 , n96277 );
not ( n96279 , n90370 );
not ( n96280 , n90471 );
or ( n96281 , n96279 , n96280 );
nand ( n96282 , n90418 , n90722 );
nand ( n96283 , n96281 , n96282 );
not ( n96284 , n90442 );
not ( n96285 , n91108 );
or ( n96286 , n96284 , n96285 );
nand ( n96287 , n96145 , n90405 );
nand ( n96288 , n96286 , n96287 );
xor ( n96289 , n96283 , n96288 );
and ( n96290 , n96278 , n96289 );
and ( n96291 , n96267 , n96277 );
or ( n96292 , n96290 , n96291 );
not ( n96293 , n90612 );
not ( n96294 , n90552 );
or ( n96295 , n96293 , n96294 );
nand ( n96296 , n90555 , n90630 );
nand ( n96297 , n96295 , n96296 );
not ( n96298 , n96297 );
or ( n96299 , n96298 , n90609 );
not ( n96300 , n90612 );
not ( n96301 , n90693 );
or ( n96302 , n96300 , n96301 );
nand ( n96303 , n90690 , n90630 );
nand ( n96304 , n96302 , n96303 );
nand ( n96305 , n96304 , n90657 );
nand ( n96306 , n96299 , n96305 );
xor ( n96307 , n96292 , n96306 );
not ( n96308 , n90680 );
not ( n96309 , n90660 );
not ( n96310 , n90577 );
or ( n96311 , n96309 , n96310 );
nand ( n96312 , n90576 , n91164 );
nand ( n96313 , n96311 , n96312 );
not ( n96314 , n96313 );
or ( n96315 , n96308 , n96314 );
and ( n96316 , n90660 , n90855 );
not ( n96317 , n90660 );
and ( n96318 , n96317 , n90858 );
nor ( n96319 , n96316 , n96318 );
nand ( n96320 , n96319 , n91011 );
nand ( n96321 , n96315 , n96320 );
and ( n96322 , n96307 , n96321 );
and ( n96323 , n96292 , n96306 );
or ( n96324 , n96322 , n96323 );
and ( n96325 , n96265 , n96324 );
and ( n96326 , n96249 , n96264 );
or ( n96327 , n96325 , n96326 );
not ( n96328 , n90840 );
not ( n96329 , n96262 );
or ( n96330 , n96328 , n96329 );
nand ( n96331 , n96038 , n90876 );
nand ( n96332 , n96330 , n96331 );
xor ( n96333 , n96108 , n96094 );
and ( n96334 , n96333 , n96099 );
not ( n96335 , n96333 );
and ( n96336 , n96335 , n96077 );
nor ( n96337 , n96334 , n96336 );
xor ( n96338 , n96332 , n96337 );
not ( n96339 , n90656 );
not ( n96340 , n96297 );
or ( n96341 , n96339 , n96340 );
nand ( n96342 , n96128 , n90610 );
nand ( n96343 , n96341 , n96342 );
not ( n96344 , n91011 );
not ( n96345 , n96117 );
or ( n96346 , n96344 , n96345 );
nand ( n96347 , n96319 , n90680 );
nand ( n96348 , n96346 , n96347 );
xor ( n96349 , n96343 , n96348 );
and ( n96350 , n96283 , n96288 );
not ( n96351 , n90324 );
not ( n96352 , n96155 );
or ( n96353 , n96351 , n96352 );
nand ( n96354 , n96273 , n90279 );
nand ( n96355 , n96353 , n96354 );
xor ( n96356 , n96350 , n96355 );
xor ( n96357 , n96137 , n96147 );
and ( n96358 , n96356 , n96357 );
and ( n96359 , n96350 , n96355 );
or ( n96360 , n96358 , n96359 );
and ( n96361 , n96349 , n96360 );
and ( n96362 , n96343 , n96348 );
or ( n96363 , n96361 , n96362 );
xor ( n96364 , n96338 , n96363 );
xor ( n96365 , n96327 , n96364 );
xor ( n96366 , n96343 , n96348 );
xor ( n96367 , n96366 , n96360 );
not ( n96368 , n90582 );
not ( n96369 , n96189 );
or ( n96370 , n96368 , n96369 );
not ( n96371 , n90890 );
not ( n96372 , n90873 );
or ( n96373 , n96371 , n96372 );
nand ( n96374 , n90870 , n90539 );
nand ( n96375 , n96373 , n96374 );
nand ( n96376 , n96375 , n90537 );
nand ( n96377 , n96370 , n96376 );
not ( n96378 , n87689 );
not ( n96379 , n96204 );
or ( n96380 , n96378 , n96379 );
not ( n96381 , n87706 );
not ( n96382 , n95709 );
or ( n96383 , n96381 , n96382 );
nand ( n96384 , n95708 , n87705 );
nand ( n96385 , n96383 , n96384 );
nand ( n96386 , n96385 , n87702 );
nand ( n96387 , n96380 , n96386 );
xor ( n96388 , n96377 , n96387 );
not ( n96389 , n90788 );
not ( n96390 , n90102 );
or ( n96391 , n96389 , n96390 );
nand ( n96392 , n90801 , n90099 );
nand ( n96393 , n96391 , n96392 );
not ( n96394 , n96393 );
not ( n96395 , n90825 );
or ( n96396 , n96394 , n96395 );
not ( n96397 , n90782 );
or ( n96398 , n96212 , n96397 );
nand ( n96399 , n96396 , n96398 );
and ( n96400 , n96388 , n96399 );
and ( n96401 , n96377 , n96387 );
or ( n96402 , n96400 , n96401 );
xor ( n96403 , n96367 , n96402 );
xor ( n96404 , n96350 , n96355 );
xor ( n96405 , n96404 , n96357 );
not ( n96406 , n90610 );
not ( n96407 , n96304 );
or ( n96408 , n96406 , n96407 );
nand ( n96409 , n91152 , n90656 );
nand ( n96410 , n96408 , n96409 );
not ( n96411 , n91011 );
not ( n96412 , n96313 );
or ( n96413 , n96411 , n96412 );
nand ( n96414 , n91166 , n90680 );
nand ( n96415 , n96413 , n96414 );
xor ( n96416 , n96410 , n96415 );
xor ( n96417 , n91089 , n91098 );
and ( n96418 , n96417 , n91116 );
and ( n96419 , n91089 , n91098 );
or ( n96420 , n96418 , n96419 );
and ( n96421 , n96416 , n96420 );
and ( n96422 , n96410 , n96415 );
or ( n96423 , n96421 , n96422 );
xor ( n96424 , n96405 , n96423 );
not ( n96425 , n96255 );
or ( n96426 , n96425 , n90838 );
not ( n96427 , n90844 );
not ( n96428 , n90796 );
or ( n96429 , n96427 , n96428 );
nand ( n96430 , n90795 , n90843 );
nand ( n96431 , n96429 , n96430 );
nand ( n96432 , n96431 , n90840 );
nand ( n96433 , n96426 , n96432 );
and ( n96434 , n96424 , n96433 );
and ( n96435 , n96405 , n96423 );
or ( n96436 , n96434 , n96435 );
and ( n96437 , n96403 , n96436 );
and ( n96438 , n96367 , n96402 );
or ( n96439 , n96437 , n96438 );
xor ( n96440 , n96365 , n96439 );
xor ( n96441 , n96247 , n96440 );
xor ( n96442 , n96191 , n96206 );
xor ( n96443 , n96442 , n96222 );
xor ( n96444 , n96249 , n96264 );
xor ( n96445 , n96444 , n96324 );
xor ( n96446 , n96443 , n96445 );
xor ( n96447 , n96292 , n96306 );
xor ( n96448 , n96447 , n96321 );
not ( n96449 , n96448 );
not ( n96450 , n90825 );
not ( n96451 , n91178 );
or ( n96452 , n96450 , n96451 );
nand ( n96453 , n96393 , n90782 );
nand ( n96454 , n96452 , n96453 );
not ( n96455 , n87702 );
not ( n96456 , n90156 );
or ( n96457 , n96455 , n96456 );
nand ( n96458 , n96385 , n87689 );
nand ( n96459 , n96457 , n96458 );
xor ( n96460 , n96454 , n96459 );
xor ( n96461 , n91146 , n91156 );
and ( n96462 , n96461 , n91168 );
and ( n96463 , n91146 , n91156 );
or ( n96464 , n96462 , n96463 );
and ( n96465 , n96460 , n96464 );
and ( n96466 , n96454 , n96459 );
or ( n96467 , n96465 , n96466 );
not ( n96468 , n96467 );
or ( n96469 , n96449 , n96468 );
or ( n96470 , n96467 , n96448 );
xor ( n96471 , n96267 , n96277 );
xor ( n96472 , n96471 , n96289 );
not ( n96473 , n90537 );
not ( n96474 , n91133 );
or ( n96475 , n96473 , n96474 );
nand ( n96476 , n96375 , n90582 );
nand ( n96477 , n96475 , n96476 );
xor ( n96478 , n96472 , n96477 );
not ( n96479 , n90876 );
not ( n96480 , n96431 );
or ( n96481 , n96479 , n96480 );
nand ( n96482 , n91125 , n90840 );
nand ( n96483 , n96481 , n96482 );
and ( n96484 , n96478 , n96483 );
and ( n96485 , n96472 , n96477 );
or ( n96486 , n96484 , n96485 );
nand ( n96487 , n96470 , n96486 );
nand ( n96488 , n96469 , n96487 );
and ( n96489 , n96446 , n96488 );
and ( n96490 , n96443 , n96445 );
or ( n96491 , n96489 , n96490 );
xor ( n96492 , n96441 , n96491 );
xor ( n96493 , n96367 , n96402 );
xor ( n96494 , n96493 , n96436 );
buf ( n96495 , n96494 );
not ( n96496 , n96495 );
xor ( n96497 , n96443 , n96445 );
xor ( n96498 , n96497 , n96488 );
not ( n96499 , n96498 );
or ( n96500 , n96496 , n96499 );
or ( n96501 , n96498 , n96495 );
xor ( n96502 , n96377 , n96387 );
xor ( n96503 , n96502 , n96399 );
xor ( n96504 , n96405 , n96423 );
xor ( n96505 , n96504 , n96433 );
xor ( n96506 , n96503 , n96505 );
xor ( n96507 , n96410 , n96415 );
xor ( n96508 , n96507 , n96420 );
xor ( n96509 , n91117 , n91127 );
and ( n96510 , n96509 , n91137 );
and ( n96511 , n91117 , n91127 );
or ( n96512 , n96510 , n96511 );
xor ( n96513 , n96508 , n96512 );
xor ( n96514 , n91142 , n91169 );
and ( n96515 , n96514 , n91180 );
and ( n96516 , n91142 , n91169 );
or ( n96517 , n96515 , n96516 );
and ( n96518 , n96513 , n96517 );
and ( n96519 , n96508 , n96512 );
or ( n96520 , n96518 , n96519 );
and ( n96521 , n96506 , n96520 );
and ( n96522 , n96503 , n96505 );
or ( n96523 , n96521 , n96522 );
nand ( n96524 , n96501 , n96523 );
nand ( n96525 , n96500 , n96524 );
nor ( n96526 , n96492 , n96525 );
xor ( n96527 , n96332 , n96337 );
and ( n96528 , n96527 , n96363 );
and ( n96529 , n96332 , n96337 );
or ( n96530 , n96528 , n96529 );
xor ( n96531 , n96075 , n96111 );
xor ( n96532 , n96531 , n96165 );
xor ( n96533 , n96530 , n96532 );
xor ( n96534 , n95978 , n95988 );
xor ( n96535 , n96534 , n95999 );
xor ( n96536 , n96233 , n96238 );
and ( n96537 , n96536 , n96245 );
and ( n96538 , n96233 , n96238 );
or ( n96539 , n96537 , n96538 );
xor ( n96540 , n96535 , n96539 );
xor ( n96541 , n96030 , n96040 );
xor ( n96542 , n96541 , n96050 );
xor ( n96543 , n96540 , n96542 );
xor ( n96544 , n96533 , n96543 );
not ( n96545 , n96544 );
xor ( n96546 , n96327 , n96364 );
and ( n96547 , n96546 , n96439 );
and ( n96548 , n96327 , n96364 );
or ( n96549 , n96547 , n96548 );
not ( n96550 , n96549 );
xor ( n96551 , n96225 , n96227 );
and ( n96552 , n96551 , n96246 );
and ( n96553 , n96225 , n96227 );
or ( n96554 , n96552 , n96553 );
not ( n96555 , n96554 );
not ( n96556 , n96555 );
and ( n96557 , n96550 , n96556 );
and ( n96558 , n96549 , n96555 );
nor ( n96559 , n96557 , n96558 );
not ( n96560 , n96559 );
or ( n96561 , n96545 , n96560 );
or ( n96562 , n96544 , n96559 );
nand ( n96563 , n96561 , n96562 );
xor ( n96564 , n96247 , n96440 );
and ( n96565 , n96564 , n96491 );
and ( n96566 , n96247 , n96440 );
or ( n96567 , n96565 , n96566 );
nor ( n96568 , n96563 , n96567 );
nor ( n96569 , n96526 , n96568 );
xor ( n96570 , n96535 , n96539 );
and ( n96571 , n96570 , n96542 );
and ( n96572 , n96535 , n96539 );
or ( n96573 , n96571 , n96572 );
not ( n96574 , n96573 );
not ( n96575 , n96574 );
not ( n96576 , n96070 );
xor ( n96577 , n96168 , n96066 );
not ( n96578 , n96577 );
and ( n96579 , n96576 , n96578 );
and ( n96580 , n96070 , n96577 );
nor ( n96581 , n96579 , n96580 );
not ( n96582 , n96581 );
not ( n96583 , n96582 );
or ( n96584 , n96575 , n96583 );
nand ( n96585 , n96581 , n96573 );
nand ( n96586 , n96584 , n96585 );
xor ( n96587 , n96530 , n96532 );
and ( n96588 , n96587 , n96543 );
and ( n96589 , n96530 , n96532 );
or ( n96590 , n96588 , n96589 );
not ( n96591 , n96590 );
and ( n96592 , n96586 , n96591 );
not ( n96593 , n96586 );
and ( n96594 , n96593 , n96590 );
nor ( n96595 , n96592 , n96594 );
not ( n96596 , n96549 );
not ( n96597 , n96596 );
not ( n96598 , n96555 );
and ( n96599 , n96597 , n96598 );
nand ( n96600 , n96596 , n96555 );
and ( n96601 , n96544 , n96600 );
nor ( n96602 , n96599 , n96601 );
nand ( n96603 , n96595 , n96602 );
not ( n96604 , n96574 );
not ( n96605 , n96581 );
or ( n96606 , n96604 , n96605 );
nand ( n96607 , n96606 , n96590 );
nand ( n96608 , n96582 , n96573 );
and ( n96609 , n96607 , n96608 );
xor ( n96610 , n96059 , n96018 );
xnor ( n96611 , n96610 , n96170 );
nand ( n96612 , n96609 , n96611 );
and ( n96613 , n96569 , n96603 , n96612 );
not ( n96614 , n96613 );
xor ( n96615 , n96494 , n96523 );
xnor ( n96616 , n96615 , n96498 );
xor ( n96617 , n96503 , n96505 );
xor ( n96618 , n96617 , n96520 );
xor ( n96619 , n96448 , n96486 );
xnor ( n96620 , n96619 , n96467 );
not ( n96621 , n96620 );
or ( n96622 , n96618 , n96621 );
xor ( n96623 , n96472 , n96477 );
xor ( n96624 , n96623 , n96483 );
xor ( n96625 , n96454 , n96459 );
xor ( n96626 , n96625 , n96464 );
xor ( n96627 , n96624 , n96626 );
xor ( n96628 , n90158 , n90745 );
and ( n96629 , n96628 , n90881 );
and ( n96630 , n90158 , n90745 );
or ( n96631 , n96629 , n96630 );
and ( n96632 , n96627 , n96631 );
and ( n96633 , n96624 , n96626 );
or ( n96634 , n96632 , n96633 );
nand ( n96635 , n96622 , n96634 );
nand ( n96636 , n96618 , n96621 );
and ( n96637 , n96635 , n96636 );
nand ( n96638 , n96616 , n96637 );
xor ( n96639 , n96634 , n96620 );
xor ( n96640 , n96639 , n96618 );
xor ( n96641 , n96624 , n96626 );
xor ( n96642 , n96641 , n96631 );
xor ( n96643 , n96508 , n96512 );
xor ( n96644 , n96643 , n96517 );
or ( n96645 , n96642 , n96644 );
xor ( n96646 , n91138 , n91181 );
and ( n96647 , n96646 , n91227 );
and ( n96648 , n91138 , n91181 );
or ( n96649 , n96647 , n96648 );
and ( n96650 , n96645 , n96649 );
and ( n96651 , n96644 , n96642 );
nor ( n96652 , n96650 , n96651 );
nand ( n96653 , n96640 , n96652 );
and ( n96654 , n96638 , n96653 );
not ( n96655 , n96654 );
xor ( n96656 , n96644 , n96642 );
xor ( n96657 , n96656 , n96649 );
not ( n96658 , n96657 );
or ( n96659 , n91228 , n90882 );
nand ( n96660 , n96659 , n91087 );
nand ( n96661 , n91228 , n90882 );
nand ( n96662 , n96660 , n96661 );
not ( n96663 , n96662 );
nand ( n96664 , n96658 , n96663 );
and ( n96665 , n96664 , n91468 );
not ( n96666 , n96665 );
not ( n96667 , n93512 );
or ( n96668 , n96666 , n96667 );
and ( n96669 , n96664 , n91466 );
and ( n96670 , n96657 , n96662 );
nor ( n96671 , n96669 , n96670 );
nand ( n96672 , n96668 , n96671 );
not ( n96673 , n96672 );
or ( n96674 , n96655 , n96673 );
nor ( n96675 , n96640 , n96652 );
and ( n96676 , n96638 , n96675 );
nor ( n96677 , n96616 , n96637 );
nor ( n96678 , n96676 , n96677 );
nand ( n96679 , n96674 , n96678 );
not ( n96680 , n96679 );
or ( n96681 , n96614 , n96680 );
not ( n96682 , n96603 );
nand ( n96683 , n96492 , n96525 );
or ( n96684 , n96683 , n96568 );
nand ( n96685 , n96563 , n96567 );
nand ( n96686 , n96684 , n96685 );
not ( n96687 , n96686 );
or ( n96688 , n96682 , n96687 );
not ( n96689 , n96595 );
not ( n96690 , n96602 );
nand ( n96691 , n96689 , n96690 );
nand ( n96692 , n96688 , n96691 );
and ( n96693 , n96692 , n96612 );
nor ( n96694 , n96609 , n96611 );
nor ( n96695 , n96693 , n96694 );
nand ( n96696 , n96681 , n96695 );
xor ( n96697 , n96176 , n96696 );
or ( n96698 , n96697 , n93514 );
nand ( n96699 , n95535 , n96698 );
not ( n96700 , n17569 );
not ( n96701 , n96700 );
not ( n96702 , n93590 );
or ( n96703 , n96701 , n96702 );
not ( n96704 , n17651 );
nand ( n96705 , n96703 , n96704 );
not ( n96706 , n17650 );
nor ( n96707 , n96706 , n17654 );
and ( n96708 , n96705 , n96707 );
not ( n96709 , n96705 );
not ( n96710 , n96707 );
and ( n96711 , n96709 , n96710 );
or ( n96712 , n96708 , n96711 );
or ( n96713 , n96712 , n93521 );
nor ( n96714 , n93620 , n93479 );
xor ( n96715 , n96714 , n93619 );
or ( n96716 , n96715 , n93522 );
nand ( n96717 , n96713 , n96716 );
nand ( n96718 , n96700 , n96704 );
xor ( n96719 , n93590 , n96718 );
or ( n96720 , n96719 , n93521 );
nand ( n96721 , n93428 , n92736 );
xor ( n96722 , n96721 , n93424 );
or ( n96723 , n96722 , n93625 );
nand ( n96724 , n96720 , n96723 );
not ( n96725 , n17643 );
nor ( n96726 , n96725 , n16912 );
not ( n96727 , n96726 );
not ( n96728 , n16956 );
not ( n96729 , n96728 );
buf ( n96730 , n17381 );
not ( n96731 , n96730 );
or ( n96732 , n96729 , n96731 );
nand ( n96733 , n96732 , n17641 );
not ( n96734 , n96733 );
or ( n96735 , n96727 , n96734 );
or ( n96736 , n96726 , n96733 );
nand ( n96737 , n96735 , n96736 );
or ( n96738 , n96737 , n93521 );
xor ( n96739 , n92881 , n92883 );
xor ( n96740 , n96739 , n93421 );
not ( n96741 , n96740 );
or ( n96742 , n96741 , n93625 );
nand ( n96743 , n96738 , n96742 );
nor ( n96744 , n95187 , n95190 );
not ( n96745 , n96744 );
not ( n96746 , n95340 );
nand ( n96747 , n96745 , n96746 );
not ( n96748 , n95333 );
and ( n96749 , n96747 , n96748 );
not ( n96750 , n96747 );
and ( n96751 , n96750 , n95333 );
or ( n96752 , n96749 , n96751 );
or ( n96753 , n96752 , n87684 );
and ( n96754 , n96691 , n96603 );
and ( n96755 , n96679 , n96569 );
buf ( n96756 , n96686 );
nor ( n96757 , n96755 , n96756 );
xor ( n96758 , n96754 , n96757 );
or ( n96759 , n96758 , n93514 );
nand ( n96760 , n96753 , n96759 );
and ( n96761 , n96728 , n17641 );
not ( n96762 , n96761 );
not ( n96763 , n96730 );
or ( n96764 , n96762 , n96763 );
or ( n96765 , n96761 , n96730 );
nand ( n96766 , n96764 , n96765 );
or ( n96767 , n96766 , n93521 );
xor ( n96768 , n92910 , n92912 );
xor ( n96769 , n96768 , n93418 );
not ( n96770 , n96769 );
or ( n96771 , n96770 , n93625 );
nand ( n96772 , n96767 , n96771 );
nand ( n96773 , n17039 , n17376 );
xor ( n96774 , n96773 , n17372 );
or ( n96775 , n96774 , n93521 );
not ( n96776 , n93402 );
nand ( n96777 , n96776 , n93405 );
not ( n96778 , n96777 );
nand ( n96779 , n93374 , n93091 );
not ( n96780 , n96779 );
or ( n96781 , n96778 , n96780 );
or ( n96782 , n96779 , n96777 );
nand ( n96783 , n96781 , n96782 );
not ( n96784 , n96783 );
or ( n96785 , n96784 , n93625 );
nand ( n96786 , n96775 , n96785 );
not ( n96787 , n17360 );
and ( n96788 , n17150 , n17363 );
not ( n96789 , n96788 );
or ( n96790 , n96787 , n96789 );
or ( n96791 , n96788 , n17360 );
nand ( n96792 , n96790 , n96791 );
or ( n96793 , n96792 , n93521 );
xor ( n96794 , n93152 , n93154 );
xor ( n96795 , n96794 , n93365 );
not ( n96796 , n96795 );
or ( n96797 , n96796 , n93522 );
nand ( n96798 , n96793 , n96797 );
not ( n96799 , n17356 );
and ( n96800 , n17188 , n17359 );
not ( n96801 , n96800 );
or ( n96802 , n96799 , n96801 );
or ( n96803 , n96800 , n17356 );
nand ( n96804 , n96802 , n96803 );
or ( n96805 , n96804 , n93521 );
nand ( n96806 , n93364 , n93250 );
xor ( n96807 , n93360 , n96806 );
or ( n96808 , n96807 , n93625 );
nand ( n96809 , n96805 , n96808 );
not ( n96810 , n17736 );
not ( n96811 , n95279 );
or ( n96812 , n96810 , n96811 );
nand ( n96813 , n96812 , n95311 );
nand ( n96814 , n95322 , n96813 );
nand ( n96815 , n95330 , n95261 );
xor ( n96816 , n96814 , n96815 );
or ( n96817 , n96816 , n87684 );
not ( n96818 , n96677 );
nand ( n96819 , n96818 , n96638 );
not ( n96820 , n96653 );
not ( n96821 , n96672 );
or ( n96822 , n96820 , n96821 );
not ( n96823 , n96675 );
nand ( n96824 , n96822 , n96823 );
xor ( n96825 , n96819 , n96824 );
or ( n96826 , n96825 , n93514 );
nand ( n96827 , n96817 , n96826 );
and ( n96828 , n17355 , n17226 );
xnor ( n96829 , n17352 , n96828 );
or ( n96830 , n96829 , n93521 );
nand ( n96831 , n93359 , n93265 );
xor ( n96832 , n93355 , n96831 );
or ( n96833 , n96832 , n93625 );
nand ( n96834 , n96830 , n96833 );
not ( n96835 , n93514 );
not ( n96836 , n95314 );
nand ( n96837 , n96836 , n95316 );
not ( n96838 , n96837 );
nand ( n96839 , n17737 , n87675 );
nand ( n96840 , n96839 , n87676 );
not ( n96841 , n96840 );
or ( n96842 , n96838 , n96841 );
or ( n96843 , n96837 , n96840 );
nand ( n96844 , n96842 , n96843 );
not ( n96845 , n96844 );
or ( n96846 , n96835 , n96845 );
not ( n96847 , n96670 );
nand ( n96848 , n96847 , n96664 );
not ( n96849 , n96848 );
not ( n96850 , n91468 );
not ( n96851 , n93512 );
or ( n96852 , n96850 , n96851 );
nand ( n96853 , n96852 , n91467 );
not ( n96854 , n96853 );
or ( n96855 , n96849 , n96854 );
or ( n96856 , n96853 , n96848 );
nand ( n96857 , n96855 , n96856 );
nand ( n96858 , n96857 , n87684 );
nand ( n96859 , n96846 , n96858 );
and ( n96860 , n90555 , n90722 );
and ( n96861 , n90576 , n90370 );
nor ( n96862 , n96860 , n96861 );
not ( n96863 , n96862 );
or ( n96864 , n90839 , n90876 );
nand ( n96865 , n96864 , n90844 );
not ( n96866 , n96865 );
and ( n96867 , n96863 , n96866 );
and ( n96868 , n96862 , n96865 );
nor ( n96869 , n96867 , n96868 );
not ( n96870 , n96869 );
not ( n96871 , n90324 );
not ( n96872 , n90305 );
not ( n96873 , n90796 );
or ( n96874 , n96872 , n96873 );
nand ( n96875 , n90795 , n90321 );
nand ( n96876 , n96874 , n96875 );
not ( n96877 , n96876 );
or ( n96878 , n96871 , n96877 );
nand ( n96879 , n95547 , n90279 );
nand ( n96880 , n96878 , n96879 );
not ( n96881 , n96880 );
or ( n96882 , n96870 , n96881 );
or ( n96883 , n96880 , n96869 );
nand ( n96884 , n96882 , n96883 );
not ( n96885 , n90442 );
not ( n96886 , n95563 );
or ( n96887 , n96885 , n96886 );
and ( n96888 , n90407 , n90870 );
not ( n96889 , n90407 );
and ( n96890 , n96889 , n90873 );
nor ( n96891 , n96888 , n96890 );
nand ( n96892 , n96891 , n90405 );
nand ( n96893 , n96887 , n96892 );
xor ( n96894 , n95540 , n96893 );
not ( n96895 , n90610 );
not ( n96896 , n90612 );
not ( n96897 , n90102 );
or ( n96898 , n96896 , n96897 );
nand ( n96899 , n90630 , n90099 );
nand ( n96900 , n96898 , n96899 );
not ( n96901 , n96900 );
or ( n96902 , n96895 , n96901 );
nand ( n96903 , n95766 , n90656 );
nand ( n96904 , n96902 , n96903 );
xor ( n96905 , n96894 , n96904 );
xor ( n96906 , n96884 , n96905 );
xor ( n96907 , n95730 , n95753 );
and ( n96908 , n96907 , n95768 );
and ( n96909 , n95730 , n95753 );
or ( n96910 , n96908 , n96909 );
xor ( n96911 , n96906 , n96910 );
not ( n96912 , n90680 );
not ( n96913 , n95775 );
or ( n96914 , n96912 , n96913 );
not ( n96915 , n90660 );
not ( n96916 , n95709 );
or ( n96917 , n96915 , n96916 );
nand ( n96918 , n95708 , n91164 );
nand ( n96919 , n96917 , n96918 );
nand ( n96920 , n96919 , n91011 );
nand ( n96921 , n96914 , n96920 );
not ( n96922 , n90537 );
not ( n96923 , n95784 );
or ( n96924 , n96922 , n96923 );
not ( n96925 , n90540 );
not ( n96926 , n95681 );
or ( n96927 , n96925 , n96926 );
nand ( n96928 , n95678 , n90539 );
nand ( n96929 , n96927 , n96928 );
nand ( n96930 , n96929 , n90582 );
nand ( n96931 , n96924 , n96930 );
xor ( n96932 , n96921 , n96931 );
xor ( n96933 , n95541 , n95556 );
and ( n96934 , n96933 , n95572 );
and ( n96935 , n95541 , n95556 );
or ( n96936 , n96934 , n96935 );
xor ( n96937 , n96932 , n96936 );
xor ( n96938 , n95779 , n95788 );
and ( n96939 , n96938 , n95817 );
and ( n96940 , n95779 , n95788 );
or ( n96941 , n96939 , n96940 );
not ( n96942 , n96941 );
xor ( n96943 , n96937 , n96942 );
xor ( n96944 , n95573 , n95724 );
and ( n96945 , n96944 , n95769 );
and ( n96946 , n95573 , n95724 );
or ( n96947 , n96945 , n96946 );
xnor ( n96948 , n96943 , n96947 );
xor ( n96949 , n96911 , n96948 );
xor ( n96950 , n95818 , n95858 );
and ( n96951 , n96950 , n95948 );
and ( n96952 , n95818 , n95858 );
or ( n96953 , n96951 , n96952 );
xor ( n96954 , n96949 , n96953 );
xor ( n96955 , n95770 , n95949 );
and ( n96956 , n96955 , n96015 );
and ( n96957 , n95770 , n95949 );
or ( n96958 , n96956 , n96957 );
nand ( n96959 , n96954 , n96958 );
nor ( n96960 , n96954 , n96958 );
not ( n96961 , n96960 );
nand ( n96962 , n96959 , n96961 );
not ( n96963 , n96962 );
not ( n96964 , n96613 );
not ( n96965 , n96679 );
or ( n96966 , n96964 , n96965 );
nand ( n96967 , n96966 , n96695 );
nand ( n96968 , n96967 , n96174 );
nand ( n96969 , n96968 , n96175 );
not ( n96970 , n96969 );
or ( n96971 , n96963 , n96970 );
or ( n96972 , n96969 , n96962 );
nand ( n96973 , n96971 , n96972 );
nand ( n96974 , n96973 , n87684 );
not ( n96975 , n93371 );
nand ( n96976 , n93091 , n93373 );
not ( n96977 , n96976 );
or ( n96978 , n96975 , n96977 );
or ( n96979 , n96976 , n93371 );
nand ( n96980 , n96978 , n96979 );
and ( n96981 , n96980 , n93521 );
not ( n96982 , n454 );
not ( n96983 , n9091 );
or ( n96984 , n96982 , n96983 );
or ( n96985 , n14998 , n454 );
nand ( n96986 , n96984 , n96985 );
not ( n96987 , n96986 );
not ( n96988 , n93284 );
nand ( n96989 , n96988 , n93340 );
xor ( n96990 , n93338 , n96989 );
and ( n96991 , n93521 , n96990 );
not ( n96992 , n93521 );
not ( n96993 , n17342 );
not ( n96994 , n96993 );
not ( n96995 , n17306 );
nand ( n96996 , n96995 , n17344 );
not ( n96997 , n96996 );
or ( n96998 , n96994 , n96997 );
or ( n96999 , n96993 , n96996 );
nand ( n97000 , n96998 , n96999 );
and ( n97001 , n96992 , n97000 );
or ( n97002 , n96991 , n97001 );
not ( n97003 , n454 );
nand ( n97004 , n94853 , n94794 , n95451 );
xor ( n97005 , n95458 , n95469 );
and ( n97006 , n97005 , n95471 );
and ( n97007 , n95458 , n95469 );
or ( n97008 , n97006 , n97007 );
not ( n97009 , n16155 );
not ( n97010 , n95474 );
or ( n97011 , n97009 , n97010 );
and ( n97012 , n537 , n9757 );
not ( n97013 , n537 );
and ( n97014 , n97013 , n9758 );
nor ( n97015 , n97012 , n97014 );
nand ( n97016 , n97015 , n5501 );
nand ( n97017 , n97011 , n97016 );
and ( n97018 , n537 , n94580 );
xor ( n97019 , n97017 , n97018 );
and ( n97020 , n95467 , n4224 );
nor ( n97021 , n97020 , n5781 );
xor ( n97022 , n97019 , n97021 );
xor ( n97023 , n97008 , n97022 );
xor ( n97024 , n95478 , n95479 );
and ( n97025 , n97024 , n95484 );
and ( n97026 , n95478 , n95479 );
or ( n97027 , n97025 , n97026 );
xor ( n97028 , n97023 , n97027 );
not ( n97029 , n97028 );
xor ( n97030 , n95472 , n95485 );
and ( n97031 , n97030 , n95490 );
and ( n97032 , n95472 , n95485 );
or ( n97033 , n97031 , n97032 );
not ( n97034 , n97033 );
nand ( n97035 , n97029 , n97034 );
not ( n97036 , n97035 );
nor ( n97037 , n97036 , n95498 );
not ( n97038 , n97021 );
or ( n97039 , n4224 , n4433 );
nand ( n97040 , n97039 , n539 );
not ( n97041 , n16155 );
not ( n97042 , n97015 );
or ( n97043 , n97041 , n97042 );
xor ( n97044 , n537 , n95465 );
nand ( n97045 , n97044 , n5501 );
nand ( n97046 , n97043 , n97045 );
xor ( n97047 , n97040 , n97046 );
and ( n97048 , n94477 , n537 );
xor ( n97049 , n97047 , n97048 );
xor ( n97050 , n97038 , n97049 );
xor ( n97051 , n97017 , n97018 );
and ( n97052 , n97051 , n97021 );
and ( n97053 , n97017 , n97018 );
or ( n97054 , n97052 , n97053 );
xor ( n97055 , n97050 , n97054 );
xor ( n97056 , n97008 , n97022 );
and ( n97057 , n97056 , n97027 );
and ( n97058 , n97008 , n97022 );
or ( n97059 , n97057 , n97058 );
or ( n97060 , n97055 , n97059 );
nand ( n97061 , n97037 , n97060 );
nor ( n97062 , n97004 , n97061 );
not ( n97063 , n97062 );
not ( n97064 , n95091 );
or ( n97065 , n97063 , n97064 );
and ( n97066 , n95496 , n97035 );
and ( n97067 , n97033 , n97028 );
nor ( n97068 , n97066 , n97067 );
not ( n97069 , n97068 );
and ( n97070 , n97055 , n97059 );
nor ( n97071 , n97069 , n97070 );
not ( n97072 , n97071 );
not ( n97073 , n95448 );
or ( n97074 , n97072 , n97073 );
not ( n97075 , n97060 );
not ( n97076 , n97070 );
and ( n97077 , n97075 , n97076 );
nor ( n97078 , n97070 , n97037 );
and ( n97079 , n97068 , n97078 );
nor ( n97080 , n97077 , n97079 );
nand ( n97081 , n97074 , n97080 );
nand ( n97082 , n97065 , n97081 );
not ( n97083 , n97044 );
or ( n97084 , n97083 , n94548 );
or ( n97085 , n5408 , n5409 );
nand ( n97086 , n97084 , n97085 );
nand ( n97087 , n9757 , n537 );
xor ( n97088 , n97086 , n97087 );
xor ( n97089 , n97040 , n97046 );
and ( n97090 , n97089 , n97048 );
and ( n97091 , n97040 , n97046 );
or ( n97092 , n97090 , n97091 );
xor ( n97093 , n97088 , n97092 );
not ( n97094 , n97093 );
not ( n97095 , n97094 );
xor ( n97096 , n97038 , n97049 );
and ( n97097 , n97096 , n97054 );
and ( n97098 , n97038 , n97049 );
or ( n97099 , n97097 , n97098 );
not ( n97100 , n97099 );
not ( n97101 , n97100 );
or ( n97102 , n97095 , n97101 );
or ( n97103 , n97100 , n97094 );
nand ( n97104 , n97102 , n97103 );
not ( n97105 , n97104 );
and ( n97106 , n97082 , n97105 );
not ( n97107 , n97082 );
and ( n97108 , n97107 , n97104 );
nor ( n97109 , n97106 , n97108 );
not ( n97110 , n97109 );
or ( n97111 , n97003 , n97110 );
xor ( n97112 , n95381 , n95419 );
and ( n97113 , n97112 , n95424 );
and ( n97114 , n95381 , n95419 );
or ( n97115 , n97113 , n97114 );
not ( n97116 , n97115 );
xor ( n97117 , n95370 , n95375 );
and ( n97118 , n97117 , n95380 );
and ( n97119 , n95370 , n95375 );
or ( n97120 , n97118 , n97119 );
or ( n97121 , n12969 , n13032 );
nand ( n97122 , n97121 , n495 );
not ( n97123 , n12542 );
not ( n97124 , n95398 );
or ( n97125 , n97123 , n97124 );
xor ( n97126 , n489 , n15544 );
nand ( n97127 , n12795 , n97126 );
nand ( n97128 , n97125 , n97127 );
xor ( n97129 , n97122 , n97128 );
and ( n97130 , n12422 , n489 );
xor ( n97131 , n97129 , n97130 );
xor ( n97132 , n95394 , n95400 );
and ( n97133 , n97132 , n95412 );
and ( n97134 , n95394 , n95400 );
or ( n97135 , n97133 , n97134 );
xor ( n97136 , n97131 , n97135 );
not ( n97137 , n12595 );
not ( n97138 , n95390 );
or ( n97139 , n97137 , n97138 );
not ( n97140 , n491 );
not ( n97141 , n93711 );
or ( n97142 , n97140 , n97141 );
nand ( n97143 , n93714 , n12610 );
nand ( n97144 , n97142 , n97143 );
nand ( n97145 , n97144 , n12638 );
nand ( n97146 , n97139 , n97145 );
not ( n97147 , n12758 );
and ( n97148 , n493 , n93720 );
not ( n97149 , n493 );
and ( n97150 , n97149 , n93723 );
nor ( n97151 , n97148 , n97150 );
not ( n97152 , n97151 );
or ( n97153 , n97147 , n97152 );
nand ( n97154 , n95408 , n15344 );
nand ( n97155 , n97153 , n97154 );
xor ( n97156 , n97146 , n97155 );
xor ( n97157 , n97156 , n95369 );
xor ( n97158 , n97136 , n97157 );
xor ( n97159 , n97120 , n97158 );
xor ( n97160 , n95385 , n95413 );
and ( n97161 , n97160 , n95418 );
and ( n97162 , n95385 , n95413 );
or ( n97163 , n97161 , n97162 );
xor ( n97164 , n97159 , n97163 );
not ( n97165 , n97164 );
nand ( n97166 , n97116 , n97165 );
nand ( n97167 , n97166 , n95432 );
xor ( n97168 , n97120 , n97158 );
and ( n97169 , n97168 , n97163 );
and ( n97170 , n97120 , n97158 );
or ( n97171 , n97169 , n97170 );
and ( n97172 , n489 , n87441 );
not ( n97173 , n12638 );
not ( n97174 , n491 );
not ( n97175 , n95404 );
or ( n97176 , n97174 , n97175 );
not ( n97177 , n95404 );
nand ( n97178 , n97177 , n12610 );
nand ( n97179 , n97176 , n97178 );
not ( n97180 , n97179 );
or ( n97181 , n97173 , n97180 );
nand ( n97182 , n97144 , n12595 );
nand ( n97183 , n97181 , n97182 );
xor ( n97184 , n97172 , n97183 );
not ( n97185 , n15344 );
not ( n97186 , n97151 );
or ( n97187 , n97185 , n97186 );
nand ( n97188 , n12758 , n493 );
nand ( n97189 , n97187 , n97188 );
xor ( n97190 , n97184 , n97189 );
buf ( n97191 , n93681 );
and ( n97192 , n97191 , n12560 );
not ( n97193 , n97191 );
and ( n97194 , n97193 , n489 );
or ( n97195 , n97192 , n97194 );
not ( n97196 , n97195 );
nor ( n97197 , n97196 , n12539 );
not ( n97198 , n97126 );
nor ( n97199 , n97198 , n12541 );
nor ( n97200 , n97197 , n97199 );
xor ( n97201 , n97122 , n97128 );
and ( n97202 , n97201 , n97130 );
and ( n97203 , n97122 , n97128 );
or ( n97204 , n97202 , n97203 );
xor ( n97205 , n97200 , n97204 );
xor ( n97206 , n97146 , n97155 );
and ( n97207 , n97206 , n95369 );
and ( n97208 , n97146 , n97155 );
or ( n97209 , n97207 , n97208 );
xor ( n97210 , n97205 , n97209 );
xor ( n97211 , n97190 , n97210 );
xor ( n97212 , n97131 , n97135 );
and ( n97213 , n97212 , n97157 );
and ( n97214 , n97131 , n97135 );
or ( n97215 , n97213 , n97214 );
xor ( n97216 , n97211 , n97215 );
nor ( n97217 , n97171 , n97216 );
nor ( n97218 , n97167 , n97217 );
buf ( n97219 , n97218 );
not ( n97220 , n97219 );
not ( n97221 , n95368 );
or ( n97222 , n97220 , n97221 );
not ( n97223 , n97217 );
not ( n97224 , n97223 );
not ( n97225 , n97166 );
not ( n97226 , n95434 );
or ( n97227 , n97225 , n97226 );
nand ( n97228 , n97115 , n97164 );
nand ( n97229 , n97227 , n97228 );
not ( n97230 , n97229 );
or ( n97231 , n97224 , n97230 );
nand ( n97232 , n97171 , n97216 );
nand ( n97233 , n97231 , n97232 );
not ( n97234 , n97233 );
nand ( n97235 , n97222 , n97234 );
xor ( n97236 , n97190 , n97210 );
and ( n97237 , n97236 , n97215 );
and ( n97238 , n97190 , n97210 );
or ( n97239 , n97237 , n97238 );
not ( n97240 , n97239 );
xor ( n97241 , n97172 , n97183 );
and ( n97242 , n97241 , n97189 );
and ( n97243 , n97172 , n97183 );
or ( n97244 , n97242 , n97243 );
not ( n97245 , n12638 );
and ( n97246 , n491 , n93723 );
not ( n97247 , n491 );
and ( n97248 , n97247 , n93720 );
or ( n97249 , n97246 , n97248 );
not ( n97250 , n97249 );
or ( n97251 , n97245 , n97250 );
nand ( n97252 , n97179 , n12595 );
nand ( n97253 , n97251 , n97252 );
not ( n97254 , n97200 );
xor ( n97255 , n97253 , n97254 );
or ( n97256 , n15344 , n12758 );
nand ( n97257 , n97256 , n493 );
and ( n97258 , n489 , n15544 );
xor ( n97259 , n97257 , n97258 );
not ( n97260 , n12580 );
xor ( n97261 , n489 , n93714 );
not ( n97262 , n97261 );
or ( n97263 , n97260 , n97262 );
nand ( n97264 , n97195 , n12542 );
nand ( n97265 , n97263 , n97264 );
xor ( n97266 , n97259 , n97265 );
xor ( n97267 , n97255 , n97266 );
xor ( n97268 , n97244 , n97267 );
xor ( n97269 , n97200 , n97204 );
and ( n97270 , n97269 , n97209 );
and ( n97271 , n97200 , n97204 );
or ( n97272 , n97270 , n97271 );
xor ( n97273 , n97268 , n97272 );
not ( n97274 , n97273 );
nand ( n97275 , n97240 , n97274 );
buf ( n97276 , n97275 );
not ( n97277 , n97274 );
nand ( n97278 , n97277 , n97239 );
nand ( n97279 , n97276 , n97278 );
not ( n97280 , n97279 );
and ( n97281 , n97235 , n97280 );
not ( n97282 , n97235 );
and ( n97283 , n97282 , n97279 );
nor ( n97284 , n97281 , n97283 );
nand ( n97285 , n97284 , n10061 );
nand ( n97286 , n97111 , n97285 );
xor ( n97287 , n97086 , n97087 );
and ( n97288 , n97287 , n97092 );
and ( n97289 , n97086 , n97087 );
or ( n97290 , n97288 , n97289 );
or ( n97291 , n97100 , n97094 );
nand ( n97292 , n97100 , n97094 );
not ( n97293 , n9107 );
not ( n97294 , n78927 );
nand ( n97295 , n97294 , n9071 );
not ( n97296 , n97295 );
or ( n97297 , n97293 , n97296 );
or ( n97298 , n9107 , n97295 );
nand ( n97299 , n97297 , n97298 );
not ( n97300 , n9102 );
nand ( n97301 , n9080 , n9106 );
not ( n97302 , n97301 );
or ( n97303 , n97300 , n97302 );
or ( n97304 , n9102 , n97301 );
nand ( n97305 , n97303 , n97304 );
xor ( n97306 , n9082 , n9093 );
xor ( n97307 , n97306 , n9099 );
and ( n97308 , n9090 , n9092 );
nor ( n97309 , n97308 , n9093 );
or ( n97310 , n16155 , n5501 );
nand ( n97311 , n97310 , n537 );
not ( n97312 , n97087 );
and ( n97313 , n537 , n95465 );
xor ( n97314 , n97311 , n97313 );
xor ( n97315 , n97314 , n97312 );
not ( n97316 , n90407 );
not ( n97317 , n95681 );
or ( n97318 , n97316 , n97317 );
buf ( n97319 , n95677 );
nand ( n97320 , n97319 , n90422 );
nand ( n97321 , n97318 , n97320 );
not ( n97322 , n97321 );
or ( n97323 , n97322 , n90441 );
or ( n97324 , n90995 , n90422 );
nand ( n97325 , n97323 , n97324 );
not ( n97326 , n95709 );
not ( n97327 , n90387 );
and ( n97328 , n97326 , n97327 );
and ( n97329 , n95646 , n90370 );
nor ( n97330 , n97328 , n97329 );
xor ( n97331 , n97325 , n97330 );
or ( n97332 , n90279 , n90324 );
nand ( n97333 , n97332 , n90305 );
not ( n97334 , n97333 );
not ( n97335 , n90722 );
not ( n97336 , n90151 );
or ( n97337 , n97335 , n97336 );
nand ( n97338 , n95708 , n90370 );
nand ( n97339 , n97337 , n97338 );
not ( n97340 , n97339 );
or ( n97341 , n97334 , n97340 );
or ( n97342 , n97339 , n97333 );
not ( n97343 , n90405 );
not ( n97344 , n97321 );
or ( n97345 , n97343 , n97344 );
not ( n97346 , n90407 );
not ( n97347 , n95647 );
or ( n97348 , n97346 , n97347 );
nand ( n97349 , n95653 , n90422 );
nand ( n97350 , n97348 , n97349 );
nand ( n97351 , n97350 , n90442 );
nand ( n97352 , n97345 , n97351 );
nand ( n97353 , n97342 , n97352 );
nand ( n97354 , n97341 , n97353 );
and ( n97355 , n97331 , n97354 );
and ( n97356 , n97325 , n97330 );
nor ( n97357 , n97355 , n97356 );
and ( n97358 , n90441 , n90995 );
nor ( n97359 , n97358 , n90422 );
xor ( n97360 , n97330 , n97359 );
and ( n97361 , n95646 , n90722 );
and ( n97362 , n97319 , n90370 );
nor ( n97363 , n97361 , n97362 );
xor ( n97364 , n97360 , n97363 );
nand ( n97365 , n97357 , n97364 );
or ( n97366 , n97357 , n97364 );
nand ( n97367 , n97365 , n97366 );
not ( n97368 , n97367 );
not ( n97369 , n90370 );
not ( n97370 , n91071 );
or ( n97371 , n97369 , n97370 );
nand ( n97372 , n90795 , n90722 );
nand ( n97373 , n97371 , n97372 );
not ( n97374 , n90405 );
not ( n97375 , n90407 );
not ( n97376 , n90154 );
or ( n97377 , n97375 , n97376 );
nand ( n97378 , n90151 , n90422 );
nand ( n97379 , n97377 , n97378 );
not ( n97380 , n97379 );
or ( n97381 , n97374 , n97380 );
buf ( n97382 , n90099 );
and ( n97383 , n90407 , n97382 );
not ( n97384 , n90407 );
and ( n97385 , n97384 , n90102 );
nor ( n97386 , n97383 , n97385 );
nand ( n97387 , n97386 , n90442 );
nand ( n97388 , n97381 , n97387 );
xor ( n97389 , n97373 , n97388 );
not ( n97390 , n90324 );
and ( n97391 , n90305 , n95646 );
not ( n97392 , n90305 );
and ( n97393 , n97392 , n95647 );
nor ( n97394 , n97391 , n97393 );
not ( n97395 , n97394 );
or ( n97396 , n97390 , n97395 );
not ( n97397 , n90305 );
not ( n97398 , n95709 );
or ( n97399 , n97397 , n97398 );
nand ( n97400 , n95708 , n90321 );
nand ( n97401 , n97399 , n97400 );
nand ( n97402 , n97401 , n90279 );
nand ( n97403 , n97396 , n97402 );
xor ( n97404 , n97389 , n97403 );
not ( n97405 , n90609 );
not ( n97406 , n90630 );
and ( n97407 , n97405 , n97406 );
not ( n97408 , n90612 );
not ( n97409 , n95681 );
or ( n97410 , n97408 , n97409 );
nand ( n97411 , n97319 , n90630 );
nand ( n97412 , n97410 , n97411 );
and ( n97413 , n97412 , n90657 );
nor ( n97414 , n97407 , n97413 );
or ( n97415 , n90680 , n91011 );
nand ( n97416 , n97415 , n90660 );
not ( n97417 , n90370 );
not ( n97418 , n90795 );
or ( n97419 , n97417 , n97418 );
nand ( n97420 , n90814 , n90722 );
nand ( n97421 , n97419 , n97420 );
xor ( n97422 , n97416 , n97421 );
not ( n97423 , n90442 );
not ( n97424 , n90407 );
not ( n97425 , n91068 );
or ( n97426 , n97424 , n97425 );
nand ( n97427 , n91071 , n90422 );
nand ( n97428 , n97426 , n97427 );
not ( n97429 , n97428 );
or ( n97430 , n97423 , n97429 );
nand ( n97431 , n97386 , n90405 );
nand ( n97432 , n97430 , n97431 );
and ( n97433 , n97422 , n97432 );
and ( n97434 , n97416 , n97421 );
or ( n97435 , n97433 , n97434 );
xor ( n97436 , n97414 , n97435 );
not ( n97437 , n90873 );
not ( n97438 , n90387 );
and ( n97439 , n97437 , n97438 );
and ( n97440 , n90814 , n90370 );
nor ( n97441 , n97439 , n97440 );
not ( n97442 , n97441 );
not ( n97443 , n90610 );
not ( n97444 , n97412 );
or ( n97445 , n97443 , n97444 );
and ( n97446 , n90612 , n95646 );
not ( n97447 , n90612 );
and ( n97448 , n97447 , n95647 );
nor ( n97449 , n97446 , n97448 );
nand ( n97450 , n97449 , n90656 );
nand ( n97451 , n97445 , n97450 );
xor ( n97452 , n97442 , n97451 );
not ( n97453 , n90279 );
not ( n97454 , n90305 );
not ( n97455 , n90154 );
or ( n97456 , n97454 , n97455 );
nand ( n97457 , n90151 , n90321 );
nand ( n97458 , n97456 , n97457 );
not ( n97459 , n97458 );
or ( n97460 , n97453 , n97459 );
nand ( n97461 , n97401 , n90324 );
nand ( n97462 , n97460 , n97461 );
and ( n97463 , n97452 , n97462 );
and ( n97464 , n97442 , n97451 );
or ( n97465 , n97463 , n97464 );
xor ( n97466 , n97436 , n97465 );
xor ( n97467 , n97404 , n97466 );
xor ( n97468 , n97416 , n97421 );
xor ( n97469 , n97468 , n97432 );
xor ( n97470 , n97442 , n97451 );
xor ( n97471 , n97470 , n97462 );
xor ( n97472 , n97469 , n97471 );
not ( n97473 , n90680 );
not ( n97474 , n90660 );
not ( n97475 , n95681 );
or ( n97476 , n97474 , n97475 );
nand ( n97477 , n97319 , n91164 );
nand ( n97478 , n97476 , n97477 );
not ( n97479 , n97478 );
or ( n97480 , n97473 , n97479 );
nand ( n97481 , n91011 , n90660 );
nand ( n97482 , n97480 , n97481 );
not ( n97483 , n90656 );
not ( n97484 , n90612 );
not ( n97485 , n95709 );
or ( n97486 , n97484 , n97485 );
nand ( n97487 , n90630 , n95708 );
nand ( n97488 , n97486 , n97487 );
not ( n97489 , n97488 );
or ( n97490 , n97483 , n97489 );
nand ( n97491 , n97449 , n90610 );
nand ( n97492 , n97490 , n97491 );
xor ( n97493 , n97482 , n97492 );
not ( n97494 , n90405 );
not ( n97495 , n97428 );
or ( n97496 , n97494 , n97495 );
and ( n97497 , n90407 , n90795 );
not ( n97498 , n90407 );
and ( n97499 , n97498 , n90796 );
nor ( n97500 , n97497 , n97499 );
nand ( n97501 , n97500 , n90442 );
nand ( n97502 , n97496 , n97501 );
and ( n97503 , n97493 , n97502 );
and ( n97504 , n97482 , n97492 );
or ( n97505 , n97503 , n97504 );
and ( n97506 , n97472 , n97505 );
and ( n97507 , n97469 , n97471 );
or ( n97508 , n97506 , n97507 );
and ( n97509 , n97467 , n97508 );
and ( n97510 , n97404 , n97466 );
or ( n97511 , n97509 , n97510 );
or ( n97512 , n90657 , n90610 );
nand ( n97513 , n97512 , n90612 );
not ( n97514 , n90722 );
not ( n97515 , n91071 );
or ( n97516 , n97514 , n97515 );
nand ( n97517 , n97382 , n90370 );
nand ( n97518 , n97516 , n97517 );
xor ( n97519 , n97513 , n97518 );
not ( n97520 , n90324 );
and ( n97521 , n90305 , n97319 );
not ( n97522 , n90305 );
and ( n97523 , n97522 , n95681 );
nor ( n97524 , n97521 , n97523 );
not ( n97525 , n97524 );
or ( n97526 , n97520 , n97525 );
nand ( n97527 , n97394 , n90279 );
nand ( n97528 , n97526 , n97527 );
xor ( n97529 , n97519 , n97528 );
xor ( n97530 , n97414 , n97435 );
and ( n97531 , n97530 , n97465 );
and ( n97532 , n97414 , n97435 );
or ( n97533 , n97531 , n97532 );
xor ( n97534 , n97529 , n97533 );
not ( n97535 , n97414 );
and ( n97536 , n90422 , n95708 );
not ( n97537 , n90422 );
and ( n97538 , n97537 , n95709 );
nor ( n97539 , n97536 , n97538 );
nor ( n97540 , n97539 , n90995 );
not ( n97541 , n97379 );
nor ( n97542 , n97541 , n90441 );
or ( n97543 , n97540 , n97542 );
xor ( n97544 , n97535 , n97543 );
xor ( n97545 , n97373 , n97388 );
and ( n97546 , n97545 , n97403 );
and ( n97547 , n97373 , n97388 );
or ( n97548 , n97546 , n97547 );
xor ( n97549 , n97544 , n97548 );
xor ( n97550 , n97534 , n97549 );
nor ( n97551 , n97511 , n97550 );
not ( n97552 , n97551 );
not ( n97553 , n90324 );
not ( n97554 , n97458 );
or ( n97555 , n97553 , n97554 );
not ( n97556 , n90305 );
not ( n97557 , n90102 );
or ( n97558 , n97556 , n97557 );
nand ( n97559 , n97382 , n90321 );
nand ( n97560 , n97558 , n97559 );
nand ( n97561 , n97560 , n90279 );
nand ( n97562 , n97555 , n97561 );
xor ( n97563 , n97441 , n97562 );
or ( n97564 , n90537 , n90582 );
nand ( n97565 , n97564 , n90890 );
not ( n97566 , n90722 );
not ( n97567 , n90855 );
or ( n97568 , n97566 , n97567 );
nand ( n97569 , n90370 , n90870 );
nand ( n97570 , n97568 , n97569 );
xor ( n97571 , n97565 , n97570 );
not ( n97572 , n90405 );
not ( n97573 , n97500 );
or ( n97574 , n97572 , n97573 );
and ( n97575 , n90407 , n90814 );
not ( n97576 , n90407 );
and ( n97577 , n97576 , n90815 );
nor ( n97578 , n97575 , n97577 );
nand ( n97579 , n97578 , n90442 );
nand ( n97580 , n97574 , n97579 );
and ( n97581 , n97571 , n97580 );
and ( n97582 , n97565 , n97570 );
or ( n97583 , n97581 , n97582 );
and ( n97584 , n97563 , n97583 );
and ( n97585 , n97441 , n97562 );
or ( n97586 , n97584 , n97585 );
xor ( n97587 , n97469 , n97471 );
xor ( n97588 , n97587 , n97505 );
xor ( n97589 , n97586 , n97588 );
not ( n97590 , n91011 );
not ( n97591 , n97478 );
or ( n97592 , n97590 , n97591 );
not ( n97593 , n90660 );
not ( n97594 , n95647 );
or ( n97595 , n97593 , n97594 );
nand ( n97596 , n95653 , n91164 );
nand ( n97597 , n97595 , n97596 );
nand ( n97598 , n97597 , n90680 );
nand ( n97599 , n97592 , n97598 );
not ( n97600 , n90657 );
not ( n97601 , n90612 );
not ( n97602 , n90154 );
or ( n97603 , n97601 , n97602 );
nand ( n97604 , n90151 , n90630 );
nand ( n97605 , n97603 , n97604 );
not ( n97606 , n97605 );
or ( n97607 , n97600 , n97606 );
nand ( n97608 , n97488 , n90610 );
nand ( n97609 , n97607 , n97608 );
xor ( n97610 , n97599 , n97609 );
not ( n97611 , n90279 );
not ( n97612 , n90305 );
not ( n97613 , n91068 );
or ( n97614 , n97612 , n97613 );
nand ( n97615 , n91071 , n90321 );
nand ( n97616 , n97614 , n97615 );
not ( n97617 , n97616 );
or ( n97618 , n97611 , n97617 );
nand ( n97619 , n97560 , n90324 );
nand ( n97620 , n97618 , n97619 );
and ( n97621 , n97610 , n97620 );
and ( n97622 , n97599 , n97609 );
or ( n97623 , n97621 , n97622 );
xor ( n97624 , n97482 , n97492 );
xor ( n97625 , n97624 , n97502 );
xor ( n97626 , n97623 , n97625 );
xor ( n97627 , n97441 , n97562 );
xor ( n97628 , n97627 , n97583 );
and ( n97629 , n97626 , n97628 );
and ( n97630 , n97623 , n97625 );
or ( n97631 , n97629 , n97630 );
and ( n97632 , n97589 , n97631 );
and ( n97633 , n97586 , n97588 );
or ( n97634 , n97632 , n97633 );
xor ( n97635 , n97404 , n97466 );
xor ( n97636 , n97635 , n97508 );
or ( n97637 , n97634 , n97636 );
nand ( n97638 , n97552 , n97637 );
xor ( n97639 , n97513 , n97518 );
and ( n97640 , n97639 , n97528 );
and ( n97641 , n97513 , n97518 );
or ( n97642 , n97640 , n97641 );
not ( n97643 , n90442 );
not ( n97644 , n97539 );
not ( n97645 , n97644 );
or ( n97646 , n97643 , n97645 );
nand ( n97647 , n97350 , n90405 );
nand ( n97648 , n97646 , n97647 );
not ( n97649 , n97648 );
not ( n97650 , n90102 );
not ( n97651 , n90387 );
and ( n97652 , n97650 , n97651 );
and ( n97653 , n90151 , n90370 );
nor ( n97654 , n97652 , n97653 );
not ( n97655 , n97654 );
and ( n97656 , n97649 , n97655 );
and ( n97657 , n97648 , n97654 );
nor ( n97658 , n97656 , n97657 );
not ( n97659 , n97524 );
not ( n97660 , n90279 );
or ( n97661 , n97659 , n97660 );
nand ( n97662 , n90324 , n90305 );
nand ( n97663 , n97661 , n97662 );
and ( n97664 , n97658 , n97663 );
not ( n97665 , n97658 );
not ( n97666 , n97663 );
and ( n97667 , n97665 , n97666 );
nor ( n97668 , n97664 , n97667 );
xor ( n97669 , n97642 , n97668 );
xor ( n97670 , n97535 , n97543 );
and ( n97671 , n97670 , n97548 );
and ( n97672 , n97535 , n97543 );
or ( n97673 , n97671 , n97672 );
xor ( n97674 , n97669 , n97673 );
xor ( n97675 , n97529 , n97533 );
and ( n97676 , n97675 , n97549 );
and ( n97677 , n97529 , n97533 );
or ( n97678 , n97676 , n97677 );
or ( n97679 , n97674 , n97678 );
xor ( n97680 , n97333 , n97339 );
xnor ( n97681 , n97680 , n97352 );
and ( n97682 , n97681 , n97663 );
not ( n97683 , n97681 );
and ( n97684 , n97683 , n97666 );
or ( n97685 , n97682 , n97684 );
not ( n97686 , n97654 );
not ( n97687 , n97663 );
or ( n97688 , n97686 , n97687 );
nand ( n97689 , n97688 , n97648 );
not ( n97690 , n97654 );
nand ( n97691 , n97690 , n97666 );
and ( n97692 , n97689 , n97691 );
xnor ( n97693 , n97685 , n97692 );
xor ( n97694 , n97642 , n97668 );
and ( n97695 , n97694 , n97673 );
and ( n97696 , n97642 , n97668 );
or ( n97697 , n97695 , n97696 );
or ( n97698 , n97693 , n97697 );
xor ( n97699 , n97325 , n97330 );
xor ( n97700 , n97699 , n97354 );
not ( n97701 , n97700 );
not ( n97702 , n97681 );
not ( n97703 , n97666 );
and ( n97704 , n97702 , n97703 );
and ( n97705 , n97681 , n97666 );
nor ( n97706 , n97705 , n97692 );
nor ( n97707 , n97704 , n97706 );
nand ( n97708 , n97701 , n97707 );
nand ( n97709 , n97679 , n97698 , n97708 );
nor ( n97710 , n97638 , n97709 );
not ( n97711 , n97710 );
not ( n97712 , n90442 );
not ( n97713 , n96891 );
or ( n97714 , n97712 , n97713 );
nand ( n97715 , n97578 , n90405 );
nand ( n97716 , n97714 , n97715 );
xor ( n97717 , n97565 , n97570 );
xor ( n97718 , n97717 , n97580 );
xor ( n97719 , n97716 , n97718 );
not ( n97720 , n90324 );
not ( n97721 , n97616 );
or ( n97722 , n97720 , n97721 );
nand ( n97723 , n96876 , n90279 );
nand ( n97724 , n97722 , n97723 );
not ( n97725 , n90577 );
not ( n97726 , n90387 );
and ( n97727 , n97725 , n97726 );
and ( n97728 , n90855 , n90370 );
nor ( n97729 , n97727 , n97728 );
not ( n97730 , n97729 );
nor ( n97731 , n97724 , n97730 );
not ( n97732 , n90537 );
not ( n97733 , n96929 );
or ( n97734 , n97732 , n97733 );
nand ( n97735 , n90582 , n90890 );
nand ( n97736 , n97734 , n97735 );
not ( n97737 , n97736 );
or ( n97738 , n97731 , n97737 );
nand ( n97739 , n97724 , n97730 );
nand ( n97740 , n97738 , n97739 );
and ( n97741 , n97719 , n97740 );
and ( n97742 , n97716 , n97718 );
or ( n97743 , n97741 , n97742 );
xor ( n97744 , n97623 , n97625 );
xor ( n97745 , n97744 , n97628 );
xor ( n97746 , n97743 , n97745 );
xor ( n97747 , n97599 , n97609 );
xor ( n97748 , n97747 , n97620 );
not ( n97749 , n97748 );
and ( n97750 , n97597 , n91011 );
and ( n97751 , n96919 , n90680 );
nor ( n97752 , n97750 , n97751 );
xor ( n97753 , n97716 , n97752 );
and ( n97754 , n96900 , n90656 );
and ( n97755 , n97605 , n90610 );
nor ( n97756 , n97754 , n97755 );
and ( n97757 , n97753 , n97756 );
and ( n97758 , n97716 , n97752 );
or ( n97759 , n97757 , n97758 );
nand ( n97760 , n97749 , n97759 );
not ( n97761 , n97760 );
xor ( n97762 , n97716 , n97718 );
xor ( n97763 , n97762 , n97740 );
not ( n97764 , n97763 );
or ( n97765 , n97761 , n97764 );
not ( n97766 , n97759 );
nand ( n97767 , n97766 , n97748 );
nand ( n97768 , n97765 , n97767 );
xor ( n97769 , n97746 , n97768 );
xor ( n97770 , n97759 , n97748 );
xor ( n97771 , n97770 , n97763 );
not ( n97772 , n97771 );
not ( n97773 , n97772 );
not ( n97774 , n96862 );
not ( n97775 , n96880 );
not ( n97776 , n97775 );
or ( n97777 , n97774 , n97776 );
nand ( n97778 , n97777 , n96865 );
not ( n97779 , n96862 );
nand ( n97780 , n97779 , n96880 );
and ( n97781 , n97778 , n97780 );
not ( n97782 , n97781 );
not ( n97783 , n97782 );
xor ( n97784 , n97716 , n97752 );
xor ( n97785 , n97784 , n97756 );
not ( n97786 , n97785 );
not ( n97787 , n97786 );
or ( n97788 , n97783 , n97787 );
not ( n97789 , n97781 );
not ( n97790 , n97785 );
or ( n97791 , n97789 , n97790 );
xor ( n97792 , n95540 , n96893 );
and ( n97793 , n97792 , n96904 );
and ( n97794 , n95540 , n96893 );
or ( n97795 , n97793 , n97794 );
nand ( n97796 , n97791 , n97795 );
nand ( n97797 , n97788 , n97796 );
not ( n97798 , n97797 );
or ( n97799 , n97773 , n97798 );
not ( n97800 , n97797 );
not ( n97801 , n97800 );
not ( n97802 , n97771 );
or ( n97803 , n97801 , n97802 );
xor ( n97804 , n96921 , n96931 );
and ( n97805 , n97804 , n96936 );
and ( n97806 , n96921 , n96931 );
or ( n97807 , n97805 , n97806 );
not ( n97808 , n97807 );
xor ( n97809 , n97736 , n97729 );
xor ( n97810 , n97809 , n97724 );
nand ( n97811 , n97808 , n97810 );
not ( n97812 , n97811 );
xor ( n97813 , n96884 , n96905 );
and ( n97814 , n97813 , n96910 );
and ( n97815 , n96884 , n96905 );
or ( n97816 , n97814 , n97815 );
not ( n97817 , n97816 );
or ( n97818 , n97812 , n97817 );
not ( n97819 , n97810 );
nand ( n97820 , n97819 , n97807 );
nand ( n97821 , n97818 , n97820 );
nand ( n97822 , n97803 , n97821 );
nand ( n97823 , n97799 , n97822 );
or ( n97824 , n97769 , n97823 );
xor ( n97825 , n97743 , n97745 );
and ( n97826 , n97825 , n97768 );
and ( n97827 , n97743 , n97745 );
or ( n97828 , n97826 , n97827 );
xor ( n97829 , n97586 , n97588 );
xor ( n97830 , n97829 , n97631 );
nor ( n97831 , n97828 , n97830 );
not ( n97832 , n97831 );
and ( n97833 , n97824 , n97832 );
not ( n97834 , n97833 );
and ( n97835 , n97795 , n97781 );
not ( n97836 , n97795 );
and ( n97837 , n97836 , n97782 );
nor ( n97838 , n97835 , n97837 );
and ( n97839 , n97838 , n97786 );
not ( n97840 , n97838 );
and ( n97841 , n97840 , n97785 );
nor ( n97842 , n97839 , n97841 );
not ( n97843 , n97807 );
not ( n97844 , n97810 );
and ( n97845 , n97843 , n97844 );
and ( n97846 , n97807 , n97810 );
nor ( n97847 , n97845 , n97846 );
xor ( n97848 , n97816 , n97847 );
xor ( n97849 , n97842 , n97848 );
not ( n97850 , n96937 );
nand ( n97851 , n97850 , n96942 );
and ( n97852 , n96947 , n97851 );
nor ( n97853 , n97850 , n96942 );
nor ( n97854 , n97852 , n97853 );
xor ( n97855 , n97849 , n97854 );
or ( n97856 , n96911 , n96948 );
and ( n97857 , n97856 , n96953 );
and ( n97858 , n96911 , n96948 );
nor ( n97859 , n97857 , n97858 );
nand ( n97860 , n97855 , n97859 );
and ( n97861 , n97821 , n97797 );
not ( n97862 , n97821 );
and ( n97863 , n97862 , n97800 );
nor ( n97864 , n97861 , n97863 );
and ( n97865 , n97864 , n97771 );
not ( n97866 , n97864 );
and ( n97867 , n97866 , n97772 );
nor ( n97868 , n97865 , n97867 );
xor ( n97869 , n97842 , n97848 );
and ( n97870 , n97869 , n97854 );
and ( n97871 , n97842 , n97848 );
or ( n97872 , n97870 , n97871 );
nand ( n97873 , n97868 , n97872 );
nand ( n97874 , n96174 , n96961 , n97860 , n97873 );
not ( n97875 , n97874 );
not ( n97876 , n97875 );
not ( n97877 , n96967 );
or ( n97878 , n97876 , n97877 );
not ( n97879 , n97873 );
not ( n97880 , n97860 );
or ( n97881 , n96175 , n96960 );
nand ( n97882 , n97881 , n96959 );
not ( n97883 , n97882 );
or ( n97884 , n97880 , n97883 );
or ( n97885 , n97855 , n97859 );
nand ( n97886 , n97884 , n97885 );
not ( n97887 , n97886 );
or ( n97888 , n97879 , n97887 );
or ( n97889 , n97868 , n97872 );
nand ( n97890 , n97888 , n97889 );
not ( n97891 , n97890 );
nand ( n97892 , n97878 , n97891 );
not ( n97893 , n97892 );
or ( n97894 , n97834 , n97893 );
nand ( n97895 , n97769 , n97823 );
or ( n97896 , n97895 , n97831 );
nand ( n97897 , n97828 , n97830 );
nand ( n97898 , n97896 , n97897 );
not ( n97899 , n97898 );
nand ( n97900 , n97894 , n97899 );
not ( n97901 , n97900 );
or ( n97902 , n97711 , n97901 );
nand ( n97903 , n97634 , n97636 );
not ( n97904 , n97903 );
not ( n97905 , n97551 );
and ( n97906 , n97904 , n97905 );
and ( n97907 , n97511 , n97550 );
nor ( n97908 , n97906 , n97907 );
or ( n97909 , n97908 , n97709 );
nand ( n97910 , n97674 , n97678 );
nor ( n97911 , n97693 , n97697 );
or ( n97912 , n97910 , n97911 );
nand ( n97913 , n97693 , n97697 );
nand ( n97914 , n97912 , n97913 );
and ( n97915 , n97914 , n97708 );
not ( n97916 , n97700 );
nor ( n97917 , n97916 , n97707 );
nor ( n97918 , n97915 , n97917 );
nand ( n97919 , n97909 , n97918 );
not ( n97920 , n97919 );
nand ( n97921 , n97902 , n97920 );
not ( n97922 , n97921 );
or ( n97923 , n97368 , n97922 );
or ( n97924 , n97921 , n97367 );
nand ( n97925 , n97923 , n97924 );
nor ( n97926 , n96968 , n96960 );
nor ( n97927 , n97926 , n97882 );
not ( n97928 , n97927 );
nand ( n97929 , n97928 , n97860 );
nand ( n97930 , n97929 , n97885 );
not ( n97931 , n96603 );
or ( n97932 , n96757 , n97931 );
nand ( n97933 , n97932 , n96691 );
not ( n97934 , n96679 );
or ( n97935 , n97934 , n96526 );
nand ( n97936 , n97935 , n96683 );
not ( n97937 , n93510 );
nand ( n97938 , n97937 , n91518 );
not ( n97939 , n97938 );
not ( n97940 , n93505 );
not ( n97941 , n91790 );
or ( n97942 , n97940 , n97941 );
not ( n97943 , n93508 );
nand ( n97944 , n97942 , n97943 );
not ( n97945 , n97944 );
or ( n97946 , n97939 , n97945 );
or ( n97947 , n97944 , n97938 );
nand ( n97948 , n97946 , n97947 );
nor ( n97949 , n93508 , n97941 );
and ( n97950 , n97949 , n93505 );
not ( n97951 , n97949 );
and ( n97952 , n97951 , n97940 );
nor ( n97953 , n97950 , n97952 );
and ( n97954 , n93486 , n93606 );
nor ( n97955 , n97954 , n93490 );
xor ( n97956 , n92493 , n92495 );
xor ( n97957 , n97956 , n93483 );
not ( n97958 , n93489 );
nor ( n97959 , n97958 , n93492 );
not ( n97960 , n96683 );
nor ( n97961 , n97960 , n96526 );
not ( n97962 , n96568 );
nand ( n97963 , n97962 , n96685 );
nand ( n97964 , n96653 , n96823 );
xor ( n97965 , n93109 , n93111 );
xor ( n97966 , n97965 , n93368 );
not ( n97967 , n96694 );
nand ( n97968 , n97967 , n96612 );
nand ( n97969 , n97833 , n97710 , n97365 );
nor ( n97970 , n97969 , n97874 );
and ( n97971 , n97710 , n97898 );
nor ( n97972 , n97971 , n97919 );
not ( n97973 , n97365 );
or ( n97974 , n97972 , n97973 );
nand ( n97975 , n97974 , n97366 );
nand ( n97976 , n97889 , n97873 );
and ( n97977 , n97885 , n97860 );
nor ( n97978 , n97907 , n97551 );
not ( n97979 , n97903 );
not ( n97980 , n97637 );
nor ( n97981 , n97979 , n97980 );
not ( n97982 , n93341 );
nand ( n97983 , n93351 , n93354 );
not ( n97984 , n97983 );
or ( n97985 , n97982 , n97984 );
or ( n97986 , n97983 , n93341 );
nand ( n97987 , n97985 , n97986 );
nand ( n97988 , n97679 , n97910 );
nand ( n97989 , n97698 , n97913 );
xor ( n97990 , n93301 , n93308 );
xor ( n97991 , n97990 , n93331 );
nor ( n97992 , n95681 , n90387 );
not ( n97993 , n97992 );
xor ( n97994 , n97330 , n97359 );
and ( n97995 , n97994 , n97363 );
and ( n97996 , n97330 , n97359 );
or ( n97997 , n97995 , n97996 );
not ( n97998 , n97997 );
or ( n97999 , n97993 , n97998 );
or ( n98000 , n97997 , n97992 );
nand ( n98001 , n97999 , n98000 );
xor ( n98002 , n93310 , n93323 );
xor ( n98003 , n98002 , n93329 );
not ( n98004 , n97679 );
not ( n98005 , n97638 );
nand ( n98006 , n98005 , n97900 );
nand ( n98007 , n98006 , n97908 );
not ( n98008 , n98007 );
or ( n98009 , n98004 , n98008 );
nand ( n98010 , n98009 , n97910 );
xnor ( n98011 , n98010 , n97989 );
xor ( n98012 , n97257 , n97258 );
and ( n98013 , n98012 , n97265 );
and ( n98014 , n97257 , n97258 );
or ( n98015 , n98013 , n98014 );
xor ( n98016 , n97253 , n97254 );
and ( n98017 , n98016 , n97266 );
and ( n98018 , n97253 , n97254 );
or ( n98019 , n98017 , n98018 );
xor ( n98020 , n97244 , n97267 );
and ( n98021 , n98020 , n97272 );
and ( n98022 , n97244 , n97267 );
or ( n98023 , n98021 , n98022 );
not ( n98024 , n12580 );
not ( n98025 , n489 );
not ( n98026 , n95404 );
or ( n98027 , n98025 , n98026 );
nand ( n98028 , n97177 , n12560 );
nand ( n98029 , n98027 , n98028 );
not ( n98030 , n98029 );
or ( n98031 , n98024 , n98030 );
nand ( n98032 , n97261 , n12542 );
nand ( n98033 , n98031 , n98032 );
not ( n98034 , n12595 );
not ( n98035 , n97249 );
or ( n98036 , n98034 , n98035 );
nand ( n98037 , n12638 , n491 );
nand ( n98038 , n98036 , n98037 );
xor ( n98039 , n98033 , n98038 );
nand ( n98040 , n97191 , n489 );
xor ( n98041 , n98039 , n98040 );
xor ( n98042 , n98033 , n98038 );
and ( n98043 , n98042 , n98040 );
and ( n98044 , n98033 , n98038 );
or ( n98045 , n98043 , n98044 );
xor ( n98046 , n98015 , n98041 );
xor ( n98047 , n98046 , n98019 );
xor ( n98048 , n98015 , n98041 );
and ( n98049 , n98048 , n98019 );
and ( n98050 , n98015 , n98041 );
or ( n98051 , n98049 , n98050 );
or ( n98052 , n12595 , n12638 );
nand ( n98053 , n98052 , n491 );
and ( n98054 , n489 , n93714 );
xor ( n98055 , n98053 , n98054 );
not ( n98056 , n12580 );
xor ( n98057 , n489 , n93720 );
not ( n98058 , n98057 );
or ( n98059 , n98056 , n98058 );
nand ( n98060 , n98029 , n12542 );
nand ( n98061 , n98059 , n98060 );
xor ( n98062 , n98055 , n98061 );
xor ( n98063 , n98053 , n98054 );
and ( n98064 , n98063 , n98061 );
and ( n98065 , n98053 , n98054 );
or ( n98066 , n98064 , n98065 );
not ( n98067 , n98040 );
xor ( n98068 , n98067 , n98062 );
xor ( n98069 , n98068 , n98045 );
xor ( n98070 , n98067 , n98062 );
and ( n98071 , n98070 , n98045 );
and ( n98072 , n98067 , n98062 );
or ( n98073 , n98071 , n98072 );
not ( n98074 , n98057 );
or ( n98075 , n98074 , n12541 );
or ( n98076 , n12539 , n12560 );
nand ( n98077 , n98075 , n98076 );
nand ( n98078 , n97177 , n489 );
xor ( n98079 , n98077 , n98078 );
xor ( n98080 , n98079 , n98066 );
xor ( n98081 , n98077 , n98078 );
and ( n98082 , n98081 , n98066 );
and ( n98083 , n98077 , n98078 );
or ( n98084 , n98082 , n98083 );
not ( n98085 , n98023 );
not ( n98086 , n98047 );
nand ( n98087 , n98085 , n98086 );
nand ( n98088 , n97275 , n98087 );
nor ( n98089 , n98051 , n98069 );
nor ( n98090 , n98088 , n98089 );
and ( n98091 , n98090 , n97218 );
nand ( n98092 , n98091 , n95366 );
nand ( n98093 , n97166 , n97228 );
not ( n98094 , n98089 );
not ( n98095 , n98094 );
not ( n98096 , n98087 );
or ( n98097 , n98096 , n97278 );
not ( n98098 , n98086 );
nand ( n98099 , n98098 , n98023 );
nand ( n98100 , n98097 , n98099 );
not ( n98101 , n98100 );
or ( n98102 , n98095 , n98101 );
nand ( n98103 , n98051 , n98069 );
nand ( n98104 , n98102 , n98103 );
not ( n98105 , n98104 );
nand ( n98106 , n98087 , n98099 );
not ( n98107 , n15020 );
not ( n98108 , n14972 );
nand ( n98109 , n98108 , n15023 );
not ( n98110 , n98109 );
or ( n98111 , n98107 , n98110 );
or ( n98112 , n98109 , n15020 );
nand ( n98113 , n98111 , n98112 );
nand ( n98114 , n98073 , n98080 );
xor ( n98115 , n14978 , n14988 );
xor ( n98116 , n98115 , n15017 );
or ( n98117 , n14996 , n14999 );
nand ( n98118 , n98117 , n15000 );
not ( n98119 , n98118 );
or ( n98120 , n12542 , n12795 );
nand ( n98121 , n98120 , n489 );
not ( n98122 , n98078 );
and ( n98123 , n489 , n93720 );
xor ( n98124 , n98121 , n98123 );
xor ( n98125 , n98124 , n98122 );
xor ( n98126 , n95517 , n95518 );
and ( n98127 , n98126 , n95520 );
and ( n98128 , n95517 , n95518 );
or ( n98129 , n98127 , n98128 );
xor ( n98130 , n95348 , n95352 );
and ( n98131 , n98130 , n95521 );
and ( n98132 , n95348 , n95352 );
or ( n98133 , n98131 , n98132 );
nand ( n98134 , n95513 , n95442 );
and ( n98135 , n98134 , n471 );
and ( n98136 , n95072 , n469 );
xor ( n98137 , n98135 , n98136 );
and ( n98138 , n94938 , n470 );
xor ( n98139 , n98137 , n98138 );
xor ( n98140 , n98135 , n98136 );
and ( n98141 , n98140 , n98138 );
and ( n98142 , n98135 , n98136 );
or ( n98143 , n98141 , n98142 );
not ( n98144 , n10061 );
not ( n98145 , n95433 );
not ( n98146 , n95368 );
or ( n98147 , n98145 , n98146 );
nand ( n98148 , n98147 , n95435 );
xnor ( n98149 , n98148 , n98093 );
not ( n98150 , n98149 );
or ( n98151 , n98144 , n98150 );
not ( n98152 , n97067 );
nand ( n98153 , n98152 , n97035 );
nand ( n98154 , n98153 , n454 );
not ( n98155 , n98154 );
nor ( n98156 , n97004 , n95498 );
not ( n98157 , n98156 );
not ( n98158 , n95086 );
not ( n98159 , n94368 );
or ( n98160 , n98158 , n98159 );
nand ( n98161 , n98160 , n95090 );
not ( n98162 , n98161 );
or ( n98163 , n98157 , n98162 );
and ( n98164 , n95447 , n95499 );
nor ( n98165 , n98164 , n95496 );
nand ( n98166 , n98163 , n98165 );
not ( n98167 , n98166 );
or ( n98168 , n98155 , n98167 );
not ( n98169 , n454 );
nor ( n98170 , n98169 , n98153 );
or ( n98171 , n98166 , n98170 );
nand ( n98172 , n98168 , n98171 );
nand ( n98173 , n98151 , n98172 );
and ( n98174 , n98173 , n472 );
xor ( n98175 , n98174 , n98129 );
xor ( n98176 , n98175 , n98139 );
xor ( n98177 , n98174 , n98129 );
and ( n98178 , n98177 , n98139 );
and ( n98179 , n98174 , n98129 );
or ( n98180 , n98178 , n98179 );
nand ( n98181 , n95513 , n95442 );
and ( n98182 , n98181 , n470 );
not ( n98183 , n94938 );
nor ( n98184 , n98183 , n16056 );
xor ( n98185 , n98182 , n98184 );
not ( n98186 , n97167 );
not ( n98187 , n98186 );
not ( n98188 , n95355 );
not ( n98189 , n94256 );
or ( n98190 , n98188 , n98189 );
nand ( n98191 , n98190 , n95367 );
not ( n98192 , n98191 );
or ( n98193 , n98187 , n98192 );
not ( n98194 , n97229 );
buf ( n98195 , n98194 );
nand ( n98196 , n98193 , n98195 );
nand ( n98197 , n97223 , n97232 );
nand ( n98198 , n98197 , n10061 );
and ( n98199 , n98196 , n98198 );
not ( n98200 , n98196 );
not ( n98201 , n98197 );
nand ( n98202 , n98201 , n10061 );
and ( n98203 , n98200 , n98202 );
or ( n98204 , n98199 , n98203 );
not ( n98205 , n94930 );
nand ( n98206 , n98205 , n97037 );
nand ( n98207 , n97068 , n98206 );
and ( n98208 , n97037 , n94929 );
or ( n98209 , n98207 , n98208 );
not ( n98210 , n98209 );
nor ( n98211 , n98207 , n94882 );
nand ( n98212 , n94877 , n94856 , n98211 );
not ( n98213 , n98212 );
or ( n98214 , n98210 , n98213 );
nand ( n98215 , n97055 , n97059 );
nand ( n98216 , n97060 , n98215 );
not ( n98217 , n98216 );
nand ( n98218 , n98214 , n98217 );
not ( n98219 , n98218 );
nand ( n98220 , n98219 , n454 );
not ( n98221 , n98212 );
and ( n98222 , n98216 , n454 );
nand ( n98223 , n98209 , n98222 );
nor ( n98224 , n98221 , n98223 );
not ( n98225 , n98224 );
nand ( n98226 , n98204 , n98220 , n98225 );
and ( n98227 , n98226 , n472 );
xor ( n98228 , n98185 , n98227 );
xor ( n98229 , n98182 , n98184 );
and ( n98230 , n98229 , n98227 );
and ( n98231 , n98182 , n98184 );
or ( n98232 , n98230 , n98231 );
and ( n98233 , n98173 , n471 );
xor ( n98234 , n98233 , n98143 );
xor ( n98235 , n98234 , n98228 );
xor ( n98236 , n98233 , n98143 );
and ( n98237 , n98236 , n98228 );
and ( n98238 , n98233 , n98143 );
or ( n98239 , n98237 , n98238 );
and ( n98240 , n98181 , n469 );
and ( n98241 , n98209 , n98212 );
nand ( n98242 , n98217 , n454 );
nor ( n98243 , n98241 , n98242 );
nor ( n98244 , n98243 , n98224 );
nand ( n98245 , n98244 , n98204 );
and ( n98246 , n98245 , n471 );
xor ( n98247 , n98240 , n98246 );
and ( n98248 , n98173 , n470 );
xor ( n98249 , n98247 , n98248 );
xor ( n98250 , n98240 , n98246 );
and ( n98251 , n98250 , n98248 );
and ( n98252 , n98240 , n98246 );
or ( n98253 , n98251 , n98252 );
and ( n98254 , n97286 , n472 );
xor ( n98255 , n98254 , n98232 );
xor ( n98256 , n98255 , n98249 );
xor ( n98257 , n98254 , n98232 );
and ( n98258 , n98257 , n98249 );
and ( n98259 , n98254 , n98232 );
or ( n98260 , n98258 , n98259 );
not ( n98261 , n10061 );
not ( n98262 , n98191 );
not ( n98263 , n97278 );
nor ( n98264 , n98263 , n98106 );
nand ( n98265 , n98262 , n97234 , n98264 );
and ( n98266 , n98106 , n97276 );
and ( n98267 , n98266 , n97218 );
and ( n98268 , n98191 , n98267 );
or ( n98269 , n98106 , n97276 );
and ( n98270 , n97278 , n98269 );
not ( n98271 , n97278 );
not ( n98272 , n98106 );
and ( n98273 , n98271 , n98272 );
nor ( n98274 , n98270 , n98273 );
nor ( n98275 , n98268 , n98274 );
nand ( n98276 , n98272 , n97278 );
nor ( n98277 , n98276 , n97219 );
and ( n98278 , n97234 , n98277 );
not ( n98279 , n97234 );
and ( n98280 , n98279 , n98266 );
nor ( n98281 , n98278 , n98280 );
nand ( n98282 , n98265 , n98275 , n98281 );
not ( n98283 , n98282 );
or ( n98284 , n98261 , n98283 );
xnor ( n98285 , n97290 , n97315 );
not ( n98286 , n98285 );
nand ( n98287 , n98286 , n454 );
nor ( n98288 , n97292 , n98287 );
and ( n98289 , n97291 , n98288 );
not ( n98290 , n97291 );
nand ( n98291 , n98285 , n454 );
not ( n98292 , n98291 );
and ( n98293 , n98290 , n98292 );
nor ( n98294 , n98289 , n98293 );
not ( n98295 , n98294 );
not ( n98296 , n97292 );
nor ( n98297 , n98296 , n98291 );
nor ( n98298 , n98295 , n98297 );
not ( n98299 , n98298 );
not ( n98300 , n97082 );
or ( n98301 , n98299 , n98300 );
nand ( n98302 , n97062 , n98161 );
not ( n98303 , n98287 );
nand ( n98304 , n98303 , n97291 );
and ( n98305 , n98294 , n98304 );
nand ( n98306 , n98302 , n97081 , n98305 );
nand ( n98307 , n98301 , n98306 );
nand ( n98308 , n98284 , n98307 );
and ( n98309 , n98308 , n472 );
and ( n98310 , n98173 , n469 );
xor ( n98311 , n98309 , n98310 );
and ( n98312 , n98226 , n470 );
xor ( n98313 , n98311 , n98312 );
xor ( n98314 , n98309 , n98310 );
and ( n98315 , n98314 , n98312 );
and ( n98316 , n98309 , n98310 );
or ( n98317 , n98315 , n98316 );
and ( n98318 , n97286 , n471 );
xor ( n98319 , n98318 , n98253 );
xor ( n98320 , n98319 , n98313 );
xor ( n98321 , n98318 , n98253 );
and ( n98322 , n98321 , n98313 );
and ( n98323 , n98318 , n98253 );
or ( n98324 , n98322 , n98323 );
nor ( n98325 , n98088 , n97217 );
not ( n98326 , n98325 );
not ( n98327 , n98196 );
or ( n98328 , n98326 , n98327 );
and ( n98329 , n98094 , n98103 );
not ( n98330 , n98329 );
not ( n98331 , n98088 );
not ( n98332 , n98331 );
not ( n98333 , n97232 );
not ( n98334 , n98333 );
or ( n98335 , n98332 , n98334 );
not ( n98336 , n98100 );
nand ( n98337 , n98335 , n98336 );
nor ( n98338 , n98330 , n98337 );
nand ( n98339 , n98328 , n98338 );
not ( n98340 , n98186 );
not ( n98341 , n98191 );
or ( n98342 , n98340 , n98341 );
nand ( n98343 , n98342 , n98194 );
not ( n98344 , n98325 );
nor ( n98345 , n98344 , n98329 );
and ( n98346 , n98343 , n98345 );
not ( n98347 , n98337 );
nor ( n98348 , n98347 , n98329 );
nor ( n98349 , n98346 , n98348 );
nand ( n98350 , n98339 , n98349 );
and ( n98351 , n98350 , n472 , n10061 );
and ( n98352 , n469 , n98245 );
xor ( n98353 , n98351 , n98352 );
and ( n98354 , n97286 , n470 );
xor ( n98355 , n98353 , n98354 );
xor ( n98356 , n98351 , n98352 );
and ( n98357 , n98356 , n98354 );
and ( n98358 , n98351 , n98352 );
or ( n98359 , n98357 , n98358 );
buf ( n98360 , n98308 );
and ( n98361 , n98360 , n471 );
xor ( n98362 , n98361 , n98317 );
xor ( n98363 , n98362 , n98355 );
xor ( n98364 , n98361 , n98317 );
and ( n98365 , n98364 , n98355 );
and ( n98366 , n98361 , n98317 );
or ( n98367 , n98365 , n98366 );
and ( n98368 , n98350 , n471 , n10061 );
not ( n98369 , n98090 );
not ( n98370 , n97233 );
or ( n98371 , n98369 , n98370 );
nand ( n98372 , n98371 , n98105 );
not ( n98373 , n98372 );
and ( n98374 , n98091 , n95355 );
not ( n98375 , n98374 );
not ( n98376 , n94232 );
nand ( n98377 , n98376 , n94255 );
not ( n98378 , n98377 );
buf ( n98379 , n94249 );
not ( n98380 , n98379 );
nand ( n98381 , n98378 , n98380 );
not ( n98382 , n98381 );
or ( n98383 , n98375 , n98382 );
nand ( n98384 , n98383 , n98092 );
not ( n98385 , n98384 );
nand ( n98386 , n98373 , n98385 );
or ( n98387 , n98073 , n98080 );
not ( n98388 , n98387 );
not ( n98389 , n98388 );
nand ( n98390 , n98389 , n98114 );
and ( n98391 , n10061 , n472 );
and ( n98392 , n98390 , n98391 );
and ( n98393 , n98386 , n98392 );
not ( n98394 , n98386 );
not ( n98395 , n98391 );
nor ( n98396 , n98395 , n98390 );
and ( n98397 , n98394 , n98396 );
or ( n98398 , n98393 , n98397 );
xor ( n98399 , n98368 , n98398 );
and ( n98400 , n98308 , n470 );
xor ( n98401 , n98399 , n98400 );
xor ( n98402 , n98368 , n98398 );
and ( n98403 , n98402 , n98400 );
and ( n98404 , n98368 , n98398 );
or ( n98405 , n98403 , n98404 );
and ( n98406 , n97286 , n469 );
xor ( n98407 , n98406 , n98401 );
xor ( n98408 , n98407 , n98359 );
xor ( n98409 , n98406 , n98401 );
and ( n98410 , n98409 , n98359 );
and ( n98411 , n98406 , n98401 );
or ( n98412 , n98410 , n98411 );
not ( n98413 , n98125 );
not ( n98414 , n98084 );
or ( n98415 , n98413 , n98414 );
or ( n98416 , n98125 , n98084 );
nand ( n98417 , n98415 , n98416 );
nand ( n98418 , n98417 , n10061 );
nor ( n98419 , n98418 , n98388 );
not ( n98420 , n98419 );
not ( n98421 , n98420 );
not ( n98422 , n98374 );
not ( n98423 , n98381 );
or ( n98424 , n98422 , n98423 );
nand ( n98425 , n98424 , n98092 );
not ( n98426 , n98425 );
or ( n98427 , n98421 , n98426 );
not ( n98428 , n10061 );
nor ( n98429 , n98428 , n98417 );
nand ( n98430 , n98429 , n98114 );
nor ( n98431 , n98372 , n98430 );
nand ( n98432 , n98427 , n98431 );
and ( n98433 , n98372 , n98419 );
or ( n98434 , n98418 , n98114 );
nand ( n98435 , n98429 , n98114 , n98388 );
nand ( n98436 , n98434 , n98435 );
nor ( n98437 , n98433 , n98436 );
nand ( n98438 , n98425 , n98419 );
nand ( n98439 , n98432 , n98437 , n98438 );
and ( n98440 , n98439 , n472 );
and ( n98441 , n98350 , n10061 );
and ( n98442 , n98441 , n470 );
xor ( n98443 , n98440 , n98442 );
not ( n98444 , n98385 );
nor ( n98445 , n98372 , n98390 , n454 );
not ( n98446 , n98445 );
or ( n98447 , n98444 , n98446 );
or ( n98448 , n98384 , n98372 );
and ( n98449 , n98390 , n10061 );
nand ( n98450 , n98448 , n98449 );
nand ( n98451 , n98447 , n98450 );
and ( n98452 , n98451 , n471 );
xor ( n98453 , n98443 , n98452 );
xor ( n98454 , n98440 , n98442 );
and ( n98455 , n98454 , n98452 );
and ( n98456 , n98440 , n98442 );
or ( n98457 , n98455 , n98456 );
and ( n98458 , n98360 , n469 );
xor ( n98459 , n98458 , n98453 );
xor ( n98460 , n98459 , n98405 );
xor ( n98461 , n98458 , n98453 );
and ( n98462 , n98461 , n98405 );
and ( n98463 , n98458 , n98453 );
or ( n98464 , n98462 , n98463 );
buf ( n98465 , n98451 );
and ( n98466 , n98465 , n470 );
not ( n98467 , n98387 );
not ( n98468 , n98384 );
or ( n98469 , n98467 , n98468 );
and ( n98470 , n98372 , n98387 );
not ( n98471 , n98114 );
nor ( n98472 , n98470 , n98471 );
nand ( n98473 , n98469 , n98472 );
and ( n98474 , n98473 , n98418 );
not ( n98475 , n98473 );
not ( n98476 , n98417 );
nand ( n98477 , n98476 , n10061 );
and ( n98478 , n98475 , n98477 );
nor ( n98479 , n98474 , n98478 );
and ( n98480 , n98479 , n471 );
and ( n98481 , n98441 , n469 );
xor ( n98482 , n98480 , n98481 );
xor ( n98483 , n98466 , n98482 );
xor ( n98484 , n98483 , n98457 );
not ( n98485 , n16771 );
not ( n98486 , n98485 );
nor ( n98487 , n17690 , n93531 );
not ( n98488 , n98487 );
not ( n98489 , n93539 );
or ( n98490 , n98488 , n98489 );
not ( n98491 , n17690 );
not ( n98492 , n93542 );
and ( n98493 , n98491 , n98492 );
nor ( n98494 , n98493 , n17722 );
nand ( n98495 , n98490 , n98494 );
not ( n98496 , n98495 );
or ( n98497 , n98486 , n98496 );
nand ( n98498 , n98497 , n17729 );
not ( n98499 , n98320 );
not ( n98500 , n98260 );
nand ( n98501 , n98499 , n98500 );
nor ( n98502 , n98256 , n98239 );
nor ( n98503 , n98235 , n98180 );
nor ( n98504 , n98502 , n98503 );
nand ( n98505 , n98501 , n98504 );
nor ( n98506 , n98363 , n98324 );
nor ( n98507 , n98505 , n98506 );
not ( n98508 , n98507 );
not ( n98509 , n98408 );
not ( n98510 , n98367 );
nand ( n98511 , n98509 , n98510 );
not ( n98512 , n98460 );
not ( n98513 , n98412 );
nand ( n98514 , n98512 , n98513 );
nand ( n98515 , n98511 , n98514 );
nor ( n98516 , n98508 , n98515 );
nand ( n98517 , n98464 , n98484 );
not ( n98518 , n95264 );
nand ( n98519 , n17116 , n17367 );
not ( n98520 , n98176 );
not ( n98521 , n98133 );
nand ( n98522 , n98520 , n98521 );
nand ( n98523 , n98176 , n98133 );
nand ( n98524 , n98522 , n98523 );
or ( n98525 , n98180 , n98235 );
nand ( n98526 , n98235 , n98180 );
and ( n98527 , n98525 , n98526 );
and ( n98528 , n95318 , n95320 );
not ( n98529 , n98528 );
xor ( n98530 , n17307 , n17309 );
xor ( n98531 , n98530 , n17329 );
nor ( n98532 , n98510 , n98509 );
not ( n98533 , n96839 );
and ( n98534 , n17300 , n17351 );
not ( n98535 , n17341 );
nand ( n98536 , n98535 , n17339 );
xnor ( n98537 , n17364 , n98519 );
and ( n98538 , n17072 , n17371 );
not ( n98539 , n98513 );
nand ( n98540 , n98539 , n98460 );
xor ( n98541 , n97968 , n97933 );
nor ( n98542 , n98176 , n98133 );
nor ( n98543 , n95522 , n95526 );
nor ( n98544 , n98542 , n98543 );
not ( n98545 , n98544 );
not ( n98546 , n95344 );
or ( n98547 , n98545 , n98546 );
not ( n98548 , n95528 );
and ( n98549 , n98522 , n98548 );
not ( n98550 , n98523 );
nor ( n98551 , n98549 , n98550 );
nand ( n98552 , n98547 , n98551 );
not ( n98553 , n98552 );
not ( n98554 , n95322 );
not ( n98555 , n96813 );
or ( n98556 , n98554 , n98555 );
nand ( n98557 , n98544 , n95193 );
nand ( n98558 , n95327 , n95330 , n95224 );
nor ( n98559 , n98557 , n98558 );
nand ( n98560 , n98556 , n98559 );
not ( n98561 , n98557 );
nand ( n98562 , n95269 , n98561 );
nand ( n98563 , n98553 , n98560 , n98562 );
buf ( n98564 , n98563 );
not ( n98565 , n98564 );
nand ( n98566 , n98514 , n98540 );
not ( n98567 , n98500 );
not ( n98568 , n98320 );
not ( n98569 , n98568 );
or ( n98570 , n98567 , n98569 );
nor ( n98571 , n98239 , n98256 );
or ( n98572 , n98571 , n98526 );
nand ( n98573 , n98256 , n98239 );
nand ( n98574 , n98572 , n98573 );
nand ( n98575 , n98570 , n98574 );
buf ( n98576 , n98320 );
nand ( n98577 , n98260 , n98576 );
nand ( n98578 , n98324 , n98363 );
nand ( n98579 , n98575 , n98577 , n98578 );
not ( n98580 , n98579 );
not ( n98581 , n98363 );
not ( n98582 , n98324 );
nand ( n98583 , n98581 , n98582 );
not ( n98584 , n98583 );
nor ( n98585 , n98580 , n98584 );
nand ( n98586 , n98509 , n98510 );
and ( n98587 , n98585 , n98586 );
nor ( n98588 , n98587 , n98532 );
nand ( n98589 , n98576 , n98260 );
nand ( n98590 , n98501 , n98589 );
not ( n98591 , n97917 );
nand ( n98592 , n98591 , n97708 );
buf ( n98593 , n98504 );
not ( n98594 , n97970 );
not ( n98595 , n96696 );
or ( n98596 , n98594 , n98595 );
not ( n98597 , n97969 );
and ( n98598 , n98597 , n97890 );
nor ( n98599 , n98598 , n97975 );
nand ( n98600 , n98596 , n98599 );
or ( n98601 , n98590 , n87684 );
not ( n98602 , n98593 );
not ( n98603 , n98564 );
or ( n98604 , n98602 , n98603 );
not ( n98605 , n98574 );
nand ( n98606 , n98604 , n98605 );
not ( n98607 , n98590 );
nor ( n98608 , n98607 , n87684 );
nand ( n98609 , n98606 , n98608 );
and ( n98610 , n97895 , n97824 );
xnor ( n98611 , n97892 , n98610 );
or ( n98612 , n98611 , n93514 );
not ( n98613 , n98502 );
nand ( n98614 , n98613 , n98573 );
not ( n98615 , n98614 );
nor ( n98616 , n98615 , n87684 );
or ( n98617 , n98363 , n98324 );
nand ( n98618 , n98617 , n98578 );
and ( n98619 , n98618 , n93514 );
not ( n98620 , n95527 );
nand ( n98621 , n95522 , n95526 );
nand ( n98622 , n98620 , n98621 );
not ( n98623 , n98508 );
or ( n98624 , n98529 , n87684 );
not ( n98625 , n96836 );
not ( n98626 , n98533 );
or ( n98627 , n98625 , n98626 );
not ( n98628 , n95317 );
nand ( n98629 , n98627 , n98628 );
or ( n98630 , n98624 , n98629 );
not ( n98631 , n98629 );
or ( n98632 , n98528 , n87684 );
or ( n98633 , n98631 , n98632 );
xor ( n98634 , n97964 , n96672 );
or ( n98635 , n98634 , n93514 );
nand ( n98636 , n98630 , n98633 , n98635 );
buf ( n98637 , n95327 );
nand ( n98638 , n98637 , n95263 );
or ( n98639 , n98638 , n87684 );
not ( n98640 , n95330 );
not ( n98641 , n96814 );
or ( n98642 , n98640 , n98641 );
nand ( n98643 , n98642 , n95261 );
or ( n98644 , n98639 , n98643 );
not ( n98645 , n98638 );
nor ( n98646 , n98645 , n87684 );
nand ( n98647 , n98643 , n98646 );
and ( n98648 , n97961 , n96679 );
not ( n98649 , n97961 );
and ( n98650 , n98649 , n97934 );
or ( n98651 , n98648 , n98650 );
or ( n98652 , n98651 , n93514 );
nand ( n98653 , n98644 , n98647 , n98652 );
nand ( n98654 , n95337 , n95343 );
or ( n98655 , n98654 , n87684 );
or ( n98656 , n96748 , n96744 );
nand ( n98657 , n98656 , n96746 );
or ( n98658 , n98655 , n98657 );
not ( n98659 , n98654 );
nor ( n98660 , n98659 , n87684 );
nand ( n98661 , n98657 , n98660 );
or ( n98662 , n98541 , n93514 );
nand ( n98663 , n98658 , n98661 , n98662 );
nand ( n98664 , n95268 , n95224 );
not ( n98665 , n98664 );
nand ( n98666 , n98665 , n93514 );
nand ( n98667 , n95330 , n98637 );
not ( n98668 , n98667 );
not ( n98669 , n98668 );
not ( n98670 , n96814 );
or ( n98671 , n98669 , n98670 );
nand ( n98672 , n98671 , n98518 );
or ( n98673 , n98666 , n98672 );
not ( n98674 , n98664 );
not ( n98675 , n93514 );
nor ( n98676 , n98674 , n98675 );
nand ( n98677 , n98672 , n98676 );
xnor ( n98678 , n97963 , n97936 );
nand ( n98679 , n98678 , n98675 );
nand ( n98680 , n98673 , n98677 , n98679 );
and ( n98681 , n98589 , n98578 );
or ( n98682 , n98320 , n98260 );
nand ( n98683 , n98682 , n98574 );
and ( n98684 , n98683 , n98589 );
not ( n98685 , n17315 );
or ( n98686 , n17328 , n98685 );
or ( n98687 , n98685 , n17324 );
and ( n98688 , n98685 , n17323 , n86977 );
nor ( n98689 , n86977 , n17315 , n17323 );
nor ( n98690 , n98688 , n98689 );
nand ( n98691 , n98686 , n98687 , n98690 );
and ( n98692 , n17265 , n472 );
not ( n98693 , n98527 );
nand ( n98694 , n98693 , n93514 );
or ( n98695 , n98565 , n98694 );
and ( n98696 , n98527 , n93514 );
nand ( n98697 , n98565 , n98696 );
buf ( n98698 , n97927 );
not ( n98699 , n98698 );
not ( n98700 , n97977 );
or ( n98701 , n98699 , n98700 );
or ( n98702 , n98698 , n97977 );
nand ( n98703 , n98701 , n98702 );
nand ( n98704 , n98703 , n87684 );
nand ( n98705 , n98695 , n98697 , n98704 );
nand ( n98706 , n98553 , n98560 , n98562 );
not ( n98707 , n98588 );
not ( n98708 , n98586 );
nor ( n98709 , n98708 , n98508 );
nand ( n98710 , n98564 , n98709 );
not ( n98711 , n98710 );
or ( n98712 , n98707 , n98711 );
and ( n98713 , n98566 , n93514 );
nand ( n98714 , n98712 , n98713 );
nor ( n98715 , n98566 , n87684 );
nand ( n98716 , n98588 , n98710 , n98715 );
not ( n98717 , n97637 );
not ( n98718 , n97833 );
not ( n98719 , n97892 );
or ( n98720 , n98718 , n98719 );
nand ( n98721 , n98720 , n97899 );
not ( n98722 , n98721 );
or ( n98723 , n98717 , n98722 );
nand ( n98724 , n98723 , n97903 );
xor ( n98725 , n98724 , n97978 );
nand ( n98726 , n98725 , n87684 );
nand ( n98727 , n98714 , n98716 , n98726 );
not ( n98728 , n98532 );
not ( n98729 , n98514 );
or ( n98730 , n98728 , n98729 );
nand ( n98731 , n98730 , n98540 );
not ( n98732 , n97913 );
and ( n98733 , n98006 , n97910 , n97908 );
nand ( n98734 , n97679 , n97698 );
nor ( n98735 , n98733 , n98734 );
nor ( n98736 , n98732 , n98735 );
xor ( n98737 , n98592 , n98736 );
nand ( n98738 , n98737 , n93521 );
nand ( n98739 , C1 , n98738 );
nor ( n98740 , n98515 , n98584 );
and ( n98741 , n98579 , n98740 );
nor ( n98742 , n98741 , n98731 );
and ( n98743 , n98683 , n98681 );
nor ( n98744 , n98743 , n98584 );
not ( n98745 , n98744 );
and ( n98746 , n97925 , n87684 );
nor ( n98747 , C0 , n98746 );
nand ( n98748 , n98747 , C1 , C1 , C1 );
and ( n98749 , n93375 , n93403 );
nor ( n98750 , n98749 , n93406 );
not ( n98751 , n98750 );
and ( n98752 , n98751 , n93415 );
nor ( n98753 , n98750 , n93417 );
nor ( n98754 , n98752 , n98753 );
not ( n98755 , n93414 );
nand ( n98756 , n98755 , n98750 , n93409 );
not ( n98757 , n93409 );
nand ( n98758 , n98757 , n98750 , n93414 );
nand ( n98759 , n98754 , n98756 , n98758 );
not ( n98760 , n98623 );
not ( n98761 , n98564 );
or ( n98762 , n98760 , n98761 );
nand ( n98763 , n98762 , n98745 );
or ( n98764 , n98601 , n98606 );
nand ( n98765 , n98764 , n98609 , n98612 );
not ( n98766 , n98684 );
not ( n98767 , n98505 );
nand ( n98768 , n98564 , n98767 );
not ( n98769 , n98768 );
or ( n98770 , n98766 , n98769 );
nand ( n98771 , n98770 , n98619 );
not ( n98772 , n93514 );
nor ( n98773 , n98772 , n98618 );
and ( n98774 , n98768 , n98684 , n98773 );
not ( n98775 , n97897 );
nor ( n98776 , n98775 , n97831 );
not ( n98777 , n98776 );
not ( n98778 , n97875 );
not ( n98779 , n96967 );
or ( n98780 , n98778 , n98779 );
nand ( n98781 , n98780 , n97891 );
and ( n98782 , n98781 , n97824 );
not ( n98783 , n97895 );
nor ( n98784 , n98782 , n98783 );
not ( n98785 , n98784 );
or ( n98786 , n98777 , n98785 );
or ( n98787 , n98784 , n98776 );
nand ( n98788 , n98786 , n98787 );
and ( n98789 , n98788 , n87684 );
nor ( n98790 , n98774 , n98789 );
nand ( n98791 , n98771 , n98790 );
not ( n98792 , n93514 );
nand ( n98793 , n98792 , n98011 );
nand ( n98794 , C1 , C1 , n98793 , C1 );
nand ( n98795 , n98525 , n98706 , n98616 );
not ( n98796 , n97930 );
nor ( n98797 , n97976 , n93514 );
nand ( n98798 , n98796 , n98797 );
and ( n98799 , n97976 , n87684 );
nand ( n98800 , n97930 , n98799 );
not ( n98801 , n98525 );
not ( n98802 , n98614 );
nand ( n98803 , n98801 , n98802 , n98526 , n93514 );
and ( n98804 , n98798 , n98800 , n98803 );
not ( n98805 , n98526 );
nand ( n98806 , n98805 , n98616 );
not ( n98807 , n98706 );
and ( n98808 , n98802 , n98526 , n93514 );
nand ( n98809 , n98807 , n98808 );
nand ( n98810 , n98795 , n98804 , n98806 , n98809 );
not ( n98811 , n98621 );
buf ( n98812 , n98524 );
not ( n98813 , n98812 );
or ( n98814 , n98811 , n98813 );
not ( n98815 , n98622 );
or ( n98816 , n98815 , n98812 );
nand ( n98817 , n98814 , n98816 );
not ( n98818 , n98817 );
not ( n98819 , n98524 );
nand ( n98820 , n98819 , n95346 , n98621 );
not ( n98821 , n98820 );
nand ( n98822 , n98821 , n95531 );
not ( n98823 , n98822 );
or ( n98824 , n98818 , n98823 );
nand ( n98825 , n98824 , n93514 );
and ( n98826 , n98524 , n95527 , n93514 );
nand ( n98827 , n95347 , n98826 );
nand ( n98828 , n98825 , n98827 , n96974 );
not ( n98829 , n98532 );
and ( n98830 , n98586 , n98829 );
nor ( n98831 , n98830 , n87684 );
nand ( n98832 , n98763 , n98831 );
nand ( n98833 , n98623 , n98564 );
not ( n98834 , n87684 );
nand ( n98835 , n98834 , n98829 , n98586 );
nor ( n98836 , n98744 , n98835 );
and ( n98837 , n98833 , n98836 );
xnor ( n98838 , n97981 , n98721 );
nor ( n98839 , n98838 , n93514 );
nor ( n98840 , n98837 , n98839 );
nand ( n98841 , n98832 , n98840 );
nand ( n98842 , n15014 , n15003 );
or ( n98843 , n15001 , n98842 );
not ( n98844 , n15003 );
and ( n98845 , n15001 , n15014 , n98844 );
not ( n98846 , n15014 );
and ( n98847 , n15004 , n98846 );
nor ( n98848 , n98845 , n98847 );
nand ( n98849 , n98843 , C1 , n98848 );
not ( n98850 , n17634 );
not ( n98851 , n93596 );
or ( n98852 , n98850 , n98851 );
nand ( n98853 , n98852 , n93598 );
not ( n98854 , n96981 );
xor ( n98855 , n17368 , n98538 );
nand ( n98856 , n93522 , n98855 );
nand ( n98857 , n98854 , n98856 );
xor ( n98858 , n98534 , n17345 );
not ( n98859 , n454 );
and ( n98860 , n97299 , n454 );
and ( n98861 , n98113 , n98859 );
nor ( n98862 , n98860 , n98861 );
not ( n98863 , n98862 );
not ( n98864 , n93522 );
not ( n98865 , n98692 );
or ( n98866 , n98864 , n98865 );
not ( n98867 , n93321 );
nand ( n98868 , n98867 , n93521 );
nand ( n98869 , n98866 , n98868 );
and ( n98870 , n97305 , n454 );
and ( n98871 , n98116 , n98859 );
nor ( n98872 , n98870 , n98871 );
not ( n98873 , n98872 );
and ( n98874 , n97309 , n454 );
and ( n98875 , n98119 , n98859 );
nor ( n98876 , n98874 , n98875 );
not ( n98877 , n98876 );
not ( n98878 , n93522 );
not ( n98879 , n98531 );
or ( n98880 , n98878 , n98879 );
nand ( n98881 , n97991 , n93521 );
nand ( n98882 , n98880 , n98881 );
and ( n98883 , n97307 , n454 );
and ( n98884 , n98849 , n98859 );
nor ( n98885 , n98883 , n98884 );
not ( n98886 , n17622 );
not ( n98887 , n93593 );
or ( n98888 , n98886 , n98887 );
not ( n98889 , n17660 );
nand ( n98890 , n98888 , n98889 );
not ( n98891 , n17662 );
and ( n98892 , n17659 , n98891 );
nand ( n98893 , n98892 , n93514 );
or ( n98894 , n98890 , n98893 );
not ( n98895 , n97957 );
or ( n98896 , n98895 , n93514 );
not ( n98897 , n98890 );
not ( n98898 , n98892 );
nand ( n98899 , n98898 , n93514 );
or ( n98900 , n98897 , n98899 );
nand ( n98901 , n98894 , n98896 , n98900 );
nand ( n98902 , n17633 , n17629 );
not ( n98903 , n98902 );
nand ( n98904 , n98903 , n93514 );
or ( n98905 , n98853 , n98904 );
xor ( n98906 , n97959 , n97955 );
or ( n98907 , n98906 , n93514 );
not ( n98908 , n98853 );
nand ( n98909 , n98902 , n93514 );
or ( n98910 , n98908 , n98909 );
nand ( n98911 , n98905 , n98907 , n98910 );
nand ( n98912 , n98001 , n93521 );
and ( n98913 , n98600 , n98912 );
not ( n98914 , n98600 );
not ( n98915 , n98001 );
nand ( n98916 , n98915 , n93521 );
and ( n98917 , n98914 , n98916 );
nor ( n98918 , n98913 , n98917 );
not ( n98919 , n93522 );
not ( n98920 , n98537 );
or ( n98921 , n98919 , n98920 );
nand ( n98922 , n97966 , n93521 );
nand ( n98923 , n98921 , n98922 );
not ( n98924 , n93522 );
not ( n98925 , n98858 );
or ( n98926 , n98924 , n98925 );
nand ( n98927 , n97987 , n93521 );
nand ( n98928 , n98926 , n98927 );
nand ( n98929 , n98759 , n93521 );
not ( n98930 , n16961 );
nand ( n98931 , n98930 , n16996 );
buf ( n98932 , n17377 );
or ( n98933 , n98931 , n98932 );
not ( n98934 , n16996 );
nand ( n98935 , n98934 , n16961 );
or ( n98936 , n98935 , n98932 );
not ( n98937 , n17380 );
not ( n98938 , n16997 );
or ( n98939 , n98937 , n98938 );
nand ( n98940 , n98939 , n98932 );
nand ( n98941 , n98933 , n98936 , n98940 );
nand ( n98942 , n93522 , n98941 );
nand ( n98943 , n98929 , n98942 );
not ( n98944 , n93625 );
not ( n98945 , n98691 );
or ( n98946 , n98944 , n98945 );
nand ( n98947 , n98003 , n93521 );
nand ( n98948 , n98946 , n98947 );
or ( n98949 , n98464 , n98484 );
nand ( n98950 , n98949 , n98517 );
not ( n98951 , n98516 );
not ( n98952 , n98564 );
or ( n98953 , n98951 , n98952 );
nand ( n98954 , n98953 , n98742 );
not ( n98955 , n98950 );
nor ( n98956 , n98955 , n87684 );
nand ( n98957 , n98954 , n98956 );
xor ( n98958 , n98007 , n97988 );
or ( n98959 , n98958 , n93514 );
nand ( n98960 , C1 , n98957 , n98959 );
not ( n98961 , n17735 );
nand ( n98962 , n98961 , n17733 );
not ( n98963 , n98962 );
nand ( n98964 , n98963 , n93514 );
or ( n98965 , n98498 , n98964 );
and ( n98966 , n98962 , n93514 );
nand ( n98967 , n98498 , n98966 );
nand ( n98968 , n97948 , n87684 );
nand ( n98969 , n98965 , n98967 , n98968 );
nand ( n98970 , n98485 , n17729 );
not ( n98971 , n98970 );
nand ( n98972 , n98971 , n93514 );
nand ( n98973 , n97953 , n87684 );
not ( n98974 , n93527 );
not ( n98975 , n98885 );
xor ( n98976 , n93286 , n93295 );
xor ( n98977 , n98976 , n93334 );
not ( n98978 , n17332 );
not ( n98979 , n98536 );
or ( n98980 , n98978 , n98979 );
or ( n98981 , n17332 , n98536 );
nand ( n98982 , n98980 , n98981 );
and ( n98983 , n93522 , n98982 );
and ( n98984 , n98977 , n93521 );
nor ( n98985 , n98983 , n98984 );
not ( n98986 , n98985 );
or ( n98987 , n98972 , n98495 );
and ( n98988 , n98970 , n93514 );
nand ( n98989 , n98495 , n98988 );
nand ( n98990 , n98987 , n98989 , n98973 );
nand ( n98991 , n87528 , n87661 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
not ( C1n , n0 );
or ( C1 , C1n , n0 );
endmodule
