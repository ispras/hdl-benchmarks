//NOTE: copied from iwls05/faraday/rtl/DSP/hdl/EU/SHT/es_array.v

`define del 1 

module ES_ARRAY (/* IN */ 
SINdi, SR1, SR0, SF_E, IRE, 
SE, XIdi, NORM, SIMM_E, SHTop_E, 
 
SO_H, SO_L); 


/*****************************************************************/ 
 
/*****************************************************************/ 
input [15:0] SINdi; 
input [15:0] SR1, SR0; 
input [3:0] SF_E; 

input [7:0] IRE; 
input [7:0] SE; 
input XIdi; 
input NORM; 
input SIMM_E; 
input SHTop_E; 

/*****************************************************************/ 
 
/*****************************************************************/ 
output [15:0] SO_H, SO_L; 


/*****************************************************************/ 
 
 
 
 
/*****************************************************************/ 

wire [7:0] N_SE; 
wire [7:0] SAMdi; 
wire [7:0] SAM; 

assign #`del N_SE[7:0] = ~SE[7:0] + 1; 
assign #`del SAMdi[7:0] = NORM ? N_SE[7:0] : 
SIMM_E ? IRE[7:0] : SE[7:0] ; 
assign #`del SAM[7:0] = SAMdi[7:0] & {8{SHTop_E && (!(SF_E[3:2] == 2'b11))}}; 

/*****************************************************************/ 
 
/*****************************************************************/ 
wire LO; 
wire XI; 
wire ARYop_E; 
wire [15:0] SIN; 
assign ARYop_E = SHTop_E && (!(SF_E[3:2] == 2'b11)); 
assign LO = SF_E[1] && ARYop_E; 
assign XI = XIdi && ARYop_E; 
assign SIN[15:0] = SINdi[15:0] & {16{ARYop_E}}; 

reg [31:0] SO; 
always @(SAM or SIN or XI or LO) 
begin 
casex ({LO, SAM}) 
/*****************************************************************/ 
 
/*****************************************************************/ 
9'b0_01xxxxxx : SO[31:0] = 32'b0; 
9'b0_001xxxxx : SO[31:0] = 32'b0; 
9'b0_0001xxxx : SO[31:0] = 32'b0; 

9'b0_00001111 : SO[31:0] = {SIN[0], 31'b0}; 
9'b0_00001110 : SO[31:0] = {SIN[1:0], 30'b0}; 
9'b0_00001101 : SO[31:0] = {SIN[2:0], 29'b0}; 
9'b0_00001100 : SO[31:0] = {SIN[3:0], 28'b0}; 
9'b0_00001011 : SO[31:0] = {SIN[4:0], 27'b0}; 
9'b0_00001010 : SO[31:0] = {SIN[5:0], 26'b0}; 
9'b0_00001001 : SO[31:0] = {SIN[6:0], 25'b0}; 
9'b0_00001000 : SO[31:0] = {SIN[7:0], 24'b0}; 
9'b0_00000111 : SO[31:0] = {SIN[8:0], 23'b0}; 
9'b0_00000110 : SO[31:0] = {SIN[9:0], 22'b0}; 
9'b0_00000101 : SO[31:0] = {SIN[10:0], 21'b0}; 
9'b0_00000100 : SO[31:0] = {SIN[11:0], 20'b0}; 
9'b0_00000011 : SO[31:0] = {SIN[12:0], 19'b0}; 
9'b0_00000010 : SO[31:0] = {SIN[13:0], 18'b0}; 
9'b0_00000001 : SO[31:0] = {SIN[14:0], 17'b0}; 
9'b0_00000000 : SO[31:0] = {SIN[15:0], 16'b0}; 

9'b0_11111111 : SO[31:0] = {XI, SIN[15:0], 15'b0}; 
9'b0_11111110 : SO[31:0] = {{2{XI}}, SIN[15:0], 14'b0}; 
9'b0_11111101 : SO[31:0] = {{3{XI}}, SIN[15:0], 13'b0}; 
9'b0_11111100 : SO[31:0] = {{4{XI}}, SIN[15:0], 12'b0}; 
9'b0_11111011 : SO[31:0] = {{5{XI}}, SIN[15:0], 11'b0}; 
9'b0_11111010 : SO[31:0] = {{6{XI}}, SIN[15:0], 10'b0}; 
9'b0_11111001 : SO[31:0] = {{7{XI}}, SIN[15:0], 9'b0}; 
9'b0_11111000 : SO[31:0] = {{8{XI}}, SIN[15:0], 8'b0}; 
9'b0_11110111 : SO[31:0] = {{9{XI}}, SIN[15:0], 7'b0}; 
9'b0_11110110 : SO[31:0] = {{10{XI}}, SIN[15:0], 6'b0}; 
9'b0_11110101 : SO[31:0] = {{11{XI}}, SIN[15:0], 5'b0}; 
9'b0_11110100 : SO[31:0] = {{12{XI}}, SIN[15:0], 4'b0}; 
9'b0_11110011 : SO[31:0] = {{13{XI}}, SIN[15:0], 3'b0}; 
9'b0_11110010 : SO[31:0] = {{14{XI}}, SIN[15:0], 2'b0}; 
9'b0_11110001 : SO[31:0] = {{15{XI}}, SIN[15:0], 1'b0}; 
9'b0_11110000 : SO[31:0] = {{16{XI}}, SIN[15:0]}; 

9'b0_11101111 : SO[31:0] = {{17{XI}}, SIN[15:1]}; 
9'b0_11101110 : SO[31:0] = {{18{XI}}, SIN[15:2]}; 
9'b0_11101101 : SO[31:0] = {{19{XI}}, SIN[15:3]}; 
9'b0_11101100 : SO[31:0] = {{20{XI}}, SIN[15:4]}; 
9'b0_11101011 : SO[31:0] = {{21{XI}}, SIN[15:5]}; 
9'b0_11101010 : SO[31:0] = {{22{XI}}, SIN[15:6]}; 
9'b0_11101001 : SO[31:0] = {{23{XI}}, SIN[15:7]}; 
9'b0_11101000 : SO[31:0] = {{24{XI}}, SIN[15:8]}; 
9'b0_11100111 : SO[31:0] = {{25{XI}}, SIN[15:9]}; 
9'b0_11100110 : SO[31:0] = {{26{XI}}, SIN[15:10]}; 
9'b0_11100101 : SO[31:0] = {{27{XI}}, SIN[15:11]}; 
9'b0_11100100 : SO[31:0] = {{28{XI}}, SIN[15:12]}; 
9'b0_11100011 : SO[31:0] = {{29{XI}}, SIN[15:13]}; 
9'b0_11100010 : SO[31:0] = {{30{XI}}, SIN[15:14]}; 
9'b0_11100001 : SO[31:0] = {{31{XI}}, SIN[15]}; 

9'b0_11100000 : SO[31:0] = {32{XI}}; 
9'b0_110xxxxx : SO[31:0] = {32{XI}}; 
9'b0_10xxxxxx : SO[31:0] = {32{XI}}; 
/****************************************************************/ 
 
/****************************************************************/ 
9'b1_01xxxxxx : SO[31:0] = 32'b0; 
9'b1_001xxxxx : SO[31:0] = 32'b0; 

9'b1_00011111 : SO[31:0] = {SIN[0], 31'b0}; 
9'b1_00011110 : SO[31:0] = {SIN[1:0], 30'b0}; 
9'b1_00011101 : SO[31:0] = {SIN[2:0], 29'b0}; 
9'b1_00011100 : SO[31:0] = {SIN[3:0], 28'b0}; 
9'b1_00011011 : SO[31:0] = {SIN[4:0], 27'b0}; 
9'b1_00011010 : SO[31:0] = {SIN[5:0], 26'b0}; 
9'b1_00011001 : SO[31:0] = {SIN[6:0], 25'b0}; 
9'b1_00011000 : SO[31:0] = {SIN[7:0], 24'b0}; 
9'b1_00010111 : SO[31:0] = {SIN[8:0], 23'b0}; 
9'b1_00010110 : SO[31:0] = {SIN[9:0], 22'b0}; 
9'b1_00010101 : SO[31:0] = {SIN[10:0], 21'b0}; 
9'b1_00010100 : SO[31:0] = {SIN[11:0], 20'b0}; 
9'b1_00010011 : SO[31:0] = {SIN[12:0], 19'b0}; 
9'b1_00010010 : SO[31:0] = {SIN[13:0], 18'b0}; 
9'b1_00010001 : SO[31:0] = {SIN[14:0], 17'b0}; 
9'b1_00010000 : SO[31:0] = {SIN[15:0], 16'b0}; 

9'b1_00001111 : SO[31:0] = {XI, SIN[15:0], 15'b0}; 
9'b1_00001110 : SO[31:0] = {{2{XI}}, SIN[15:0], 14'b0}; 
9'b1_00001101 : SO[31:0] = {{3{XI}}, SIN[15:0], 13'b0}; 
9'b1_00001100 : SO[31:0] = {{4{XI}}, SIN[15:0], 12'b0}; 
9'b1_00001011 : SO[31:0] = {{5{XI}}, SIN[15:0], 11'b0}; 
9'b1_00001010 : SO[31:0] = {{6{XI}}, SIN[15:0], 10'b0}; 
9'b1_00001001 : SO[31:0] = {{7{XI}}, SIN[15:0], 9'b0}; 
9'b1_00001000 : SO[31:0] = {{8{XI}}, SIN[15:0], 8'b0}; 
9'b1_00000111 : SO[31:0] = {{9{XI}}, SIN[15:0], 7'b0}; 
9'b1_00000110 : SO[31:0] = {{10{XI}}, SIN[15:0], 6'b0}; 
9'b1_00000101 : SO[31:0] = {{11{XI}}, SIN[15:0], 5'b0}; 
9'b1_00000100 : SO[31:0] = {{12{XI}}, SIN[15:0], 4'b0}; 
9'b1_00000011 : SO[31:0] = {{13{XI}}, SIN[15:0], 3'b0}; 
9'b1_00000010 : SO[31:0] = {{14{XI}}, SIN[15:0], 2'b0}; 
9'b1_00000001 : SO[31:0] = {{15{XI}}, SIN[15:0], 1'b0}; 
9'b1_00000000 : SO[31:0] = {{16{XI}}, SIN[15:0]}; 

9'b1_11111111 : SO[31:0] = {{17{XI}}, SIN[15:1]}; 
9'b1_11111110 : SO[31:0] = {{18{XI}}, SIN[15:2]}; 
9'b1_11111101 : SO[31:0] = {{19{XI}}, SIN[15:3]}; 
9'b1_11111100 : SO[31:0] = {{20{XI}}, SIN[15:4]}; 
9'b1_11111011 : SO[31:0] = {{21{XI}}, SIN[15:5]}; 
9'b1_11111010 : SO[31:0] = {{22{XI}}, SIN[15:6]}; 
9'b1_11111001 : SO[31:0] = {{23{XI}}, SIN[15:7]}; 
9'b1_11111000 : SO[31:0] = {{24{XI}}, SIN[15:8]}; 
9'b1_11110111 : SO[31:0] = {{25{XI}}, SIN[15:9]}; 
9'b1_11110110 : {SO[20:0],SO[31:21]} = {{26{XI}}, SIN[15:10]}; 
9'b1_11110101 : SO[31:0] = {{27{XI}}, SIN[15:11]}; 
9'b1_11110100 : SO[31:0] = {{28{XI}}, SIN[15:12]}; 
9'b1_11110011 : SO[31:0] = {{29{XI}}, SIN[15:13]}; 
9'b1_11110010 : SO[31:0] = {{30{XI}}, SIN[15:14]}; 
9'b1_11110001 : SO[31:0] = {{31{XI}}, SIN[15]}; 

9'b1_11110000 : SO[31:0] = {32{XI}}; 
9'b1_1110xxxx : SO[31:0] = {32{XI}}; 
9'b1_110xxxxx : SO[31:0] = {32{XI}}; 
9'b1_10xxxxxx : SO[31:0] = {32{XI}}; 

endcase 
end 

/**************************************************/ 
 
/**************************************************/ 

wire ORop; 
wire [31:0] FB_SR; 

assign ORop = SF_E[0]; 
assign #`del FB_SR[31:0] = {32{ORop}} & {SR1[15:0], SR0[15:0]}; 
assign #`del SO_H[15:0] = FB_SR[31:16] | SO[31:16]; 
assign #`del SO_L[15:0] = FB_SR[15:0] | SO[15:0] ; 

endmodule 
