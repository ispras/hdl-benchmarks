module neg_2(a, b);
  input [1:0] a;
  output [2:0] b;
  assign b = -a;
endmodule
