module bitwise_or_4_6_1(a, b, c);
  input [3:0] a;
  input [5:0] b;
  output c;
  assign c = a | b;
endmodule
