//NOTE: no-implementation module stub

module REG12LC (
    input OSC,
    input OSCNTR_enb,
    input OSCNTR_ena,
    input OSCNTR_nx,
    output [11:0] OSCNTR,
    input OSCNTR_clr,
    input SCAN_TEST
);

endmodule
