module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 ;
output n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , 
 n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , 
 n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , 
 n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , 
 n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , 
 n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , 
 n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , 
 n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , 
 n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , 
 n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , 
 n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , 
 n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , 
 n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 ;
wire n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , 
 n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , 
 n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , 
 n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , 
 n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , 
 n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , 
 n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , 
 n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , 
 n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , 
 n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , 
 n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , 
 n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , 
 n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , 
 n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , 
 n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , 
 n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , 
 n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , 
 n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , 
 n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , 
 n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , 
 n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , 
 n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , 
 n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , 
 n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , 
 n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , 
 n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , 
 n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , 
 n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , 
 n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , 
 n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , 
 n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , 
 n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , 
 n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , 
 n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , 
 n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , 
 n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , 
 n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , 
 n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , 
 n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , 
 n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , 
 n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , 
 n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , 
 n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , 
 n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , 
 n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , 
 n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , 
 n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , 
 n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , 
 n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , 
 n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , 
 n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , 
 n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , 
 n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , 
 n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , 
 n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , 
 n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , 
 n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , 
 n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , 
 n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , 
 n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , 
 n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , 
 n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , 
 n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , 
 n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , 
 n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , 
 n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , 
 n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , 
 n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , 
 n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , 
 n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , 
 n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , 
 n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , 
 n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , 
 n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , 
 n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , 
 n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , 
 n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , 
 n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , 
 n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , 
 n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , 
 n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , 
 n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , 
 n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , 
 n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , 
 n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , 
 n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , 
 n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , 
 n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , 
 n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , 
 n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , 
 n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , 
 n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , 
 n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , 
 n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , 
 n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , 
 n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , 
 n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , 
 n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , 
 n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , 
 n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , 
 n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , 
 n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , 
 n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , 
 n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , 
 n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , 
 n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , 
 n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , 
 n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , 
 n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , 
 n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , 
 n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , 
 n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , 
 n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , 
 n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , 
 n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , 
 n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , 
 n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , 
 n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , 
 n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , 
 n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , 
 n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , 
 n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , 
 n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , 
 n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , 
 n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , 
 n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , 
 n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , 
 n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , 
 n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , 
 n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , 
 n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , 
 n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , 
 n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , 
 n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , 
 n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , 
 n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , 
 n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , 
 n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , 
 n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , 
 n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , 
 n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , 
 n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , 
 n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , 
 n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , 
 n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , 
 n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , 
 n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , 
 n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , 
 n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , 
 n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , 
 n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , 
 n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , 
 n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , 
 n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , 
 n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , 
 n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , 
 n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , 
 n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , 
 n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , 
 n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , 
 n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , 
 n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , 
 n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , 
 n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , 
 n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , 
 n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , 
 n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , 
 n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , 
 n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , 
 n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , 
 n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , 
 n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , 
 n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , 
 n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , 
 n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , 
 n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , 
 n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , 
 n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , 
 n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , 
 n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , 
 n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , 
 n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , 
 n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , 
 n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , 
 n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , 
 n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , 
 n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , 
 n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , 
 n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , 
 n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , 
 n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , 
 n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , 
 n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , 
 n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , 
 n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , 
 n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , 
 n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
 n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
 n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , 
 n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
 n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
 n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
 n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
 n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , 
 n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , 
 n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , 
 n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , 
 n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , 
 n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , 
 n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , 
 n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , 
 n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , 
 n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , 
 n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , 
 n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , 
 n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , 
 n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , 
 n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , 
 n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , 
 n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , 
 n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , 
 n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , 
 n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , 
 n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , 
 n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , 
 n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , 
 n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , 
 n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , 
 n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , 
 n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , 
 n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , 
 n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , 
 n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , 
 n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , 
 n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , 
 n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , 
 n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , 
 n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , 
 n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , 
 n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , 
 n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , 
 n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , 
 n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , 
 n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , 
 n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , 
 n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , 
 n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , 
 n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , 
 n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , 
 n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , 
 n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , 
 n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , 
 n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , 
 n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , 
 n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , 
 n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , 
 n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , 
 n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , 
 n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , 
 n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , 
 n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , 
 n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , 
 n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , 
 n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , 
 n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , 
 n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , 
 n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , 
 n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , 
 n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , 
 n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , 
 n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , 
 n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , 
 n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , 
 n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , 
 n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , 
 n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , 
 n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , 
 n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , 
 n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , 
 n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , 
 n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , 
 n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , 
 n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , 
 n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , 
 n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , 
 n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , 
 n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , 
 n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , 
 n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , 
 n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , 
 n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , 
 n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , 
 n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , 
 n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , 
 n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , 
 n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , 
 n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , 
 n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , 
 n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , 
 n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , 
 n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , 
 n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , 
 n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , 
 n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , 
 n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , 
 n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , 
 n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , 
 n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , 
 n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , 
 n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , 
 n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , 
 n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , 
 n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , 
 n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , 
 n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , 
 n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , 
 n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , 
 n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , 
 n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , 
 n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , 
 n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , 
 n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , 
 n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , 
 n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , 
 n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , 
 n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , 
 n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , 
 n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , 
 n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , 
 n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , 
 n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , 
 n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , 
 n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , 
 n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , 
 n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , 
 n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , 
 n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , 
 n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , 
 n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , 
 n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , 
 n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , 
 n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , 
 n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , 
 n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , 
 n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , 
 n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , 
 n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , 
 n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , 
 n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , 
 n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , 
 n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , 
 n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , 
 n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , 
 n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , 
 n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , 
 n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , 
 n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , 
 n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , 
 n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , 
 n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , 
 n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , 
 n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , 
 n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , 
 n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , 
 n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , 
 n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , 
 n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , 
 n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , 
 n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , 
 n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , 
 n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , 
 n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , 
 n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , 
 n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , 
 n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , 
 n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , 
 n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , 
 n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , 
 n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , 
 n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , 
 n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , 
 n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , 
 n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , 
 n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , 
 n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , 
 n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , 
 n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , 
 n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , 
 n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , 
 n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , 
 n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , 
 n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , 
 n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , 
 n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , 
 n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , 
 n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , 
 n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , 
 n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , 
 n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , 
 n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , 
 n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , 
 n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , 
 n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , 
 n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , 
 n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , 
 n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , 
 n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , 
 n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , 
 n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , 
 n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , 
 n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , 
 n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , 
 n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , 
 n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , 
 n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , 
 n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , 
 n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , 
 n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , 
 n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , 
 n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , 
 n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , 
 n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , 
 n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , 
 n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , 
 n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , 
 n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , 
 n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , 
 n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , 
 n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , 
 n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , 
 n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , 
 n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , 
 n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , 
 n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , 
 n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , 
 n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , 
 n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , 
 n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , 
 n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , 
 n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , 
 n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , 
 n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , 
 n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , 
 n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , 
 n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , 
 n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , 
 n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , 
 n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , 
 n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , 
 n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , 
 n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , 
 n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , 
 n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , 
 n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , 
 n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , 
 n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , 
 n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , 
 n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , 
 n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , 
 n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , 
 n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , 
 n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , 
 n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , 
 n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , 
 n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , 
 n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , 
 n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , 
 n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , 
 n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , 
 n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , 
 n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , 
 n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , 
 n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , 
 n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , 
 n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , 
 n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , 
 n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , 
 n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , 
 n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , 
 n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , 
 n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , 
 n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , 
 n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , 
 n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , 
 n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , 
 n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , 
 n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , 
 n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , 
 n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , 
 n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , 
 n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , 
 n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , 
 n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , 
 n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , 
 n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , 
 n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , 
 n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , 
 n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , 
 n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , 
 n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , 
 n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , 
 n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , 
 n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , 
 n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , 
 n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , 
 n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , 
 n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , 
 n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , 
 n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , 
 n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , 
 n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , 
 n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , 
 n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , 
 n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , 
 n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , 
 n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , 
 n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , 
 n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , 
 n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , 
 n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , 
 n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , 
 n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , 
 n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , 
 n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , 
 n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , 
 n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , 
 n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , 
 n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , 
 n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , 
 n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , 
 n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , 
 n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , 
 n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , 
 n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , 
 n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , 
 n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , 
 n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , 
 n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , 
 n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , 
 n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , 
 n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , 
 n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , 
 n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , 
 n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , 
 n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , 
 n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , 
 n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , 
 n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , 
 n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , 
 n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , 
 n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , 
 n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , 
 n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , 
 n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , 
 n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , 
 n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , 
 n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , 
 n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , 
 n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , 
 n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , 
 n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , 
 n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , 
 n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , 
 n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , 
 n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , 
 n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , 
 n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , 
 n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , 
 n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , 
 n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , 
 n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , 
 n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , 
 n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , 
 n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , 
 n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , 
 n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , 
 n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , 
 n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , 
 n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , 
 n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , 
 n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , 
 n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , 
 n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , 
 n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , 
 n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , 
 n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , 
 n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , 
 n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , 
 n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , 
 n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , 
 n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , 
 n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , 
 n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , 
 n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , 
 n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , 
 n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , 
 n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , 
 n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , 
 n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , 
 n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , 
 n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , 
 n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , 
 n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , 
 n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , 
 n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , 
 n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , 
 n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , 
 n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , 
 n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , 
 n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , 
 n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , 
 n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , 
 n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , 
 n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , 
 n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , 
 n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , 
 n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , 
 n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , 
 n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , 
 n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , 
 n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , 
 n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , 
 n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , 
 n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , 
 n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , 
 n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , 
 n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , 
 n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , 
 n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , 
 n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , 
 n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , 
 n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , 
 n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , 
 n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , 
 n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , 
 n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , 
 n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , 
 n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , 
 n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , 
 n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , 
 n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , 
 n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , 
 n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , 
 n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , 
 n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , 
 n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , 
 n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , 
 n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , 
 n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , 
 n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , 
 n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , 
 n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , 
 n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , 
 n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , 
 n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , 
 n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , 
 n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , 
 n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , 
 n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , 
 n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , 
 n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , 
 n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , 
 n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , 
 n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , 
 n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , 
 n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , 
 n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , 
 n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , 
 n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , 
 n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , 
 n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , 
 n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , 
 n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , 
 n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , 
 n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , 
 n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , 
 n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , 
 n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , 
 n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , 
 n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , 
 n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , 
 n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , 
 n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , 
 n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , 
 n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , 
 n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , 
 n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , 
 n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , 
 n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , 
 n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , 
 n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , 
 n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , 
 n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , 
 n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , 
 n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , 
 n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , 
 n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , 
 n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , 
 n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , 
 n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , 
 n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , 
 n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , 
 n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , 
 n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , 
 n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , 
 n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , 
 n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , 
 n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , 
 n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , 
 n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , 
 n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , 
 n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , 
 n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , 
 n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , 
 n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , 
 n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , 
 n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , 
 n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , 
 n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , 
 n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , 
 n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , 
 n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , 
 n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , 
 n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , 
 n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , 
 n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , 
 n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , 
 n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , 
 n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , 
 n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , 
 n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , 
 n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , 
 n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , 
 n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , 
 n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , 
 n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , 
 n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , 
 n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , 
 n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , 
 n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , 
 n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , 
 n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , 
 n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , 
 n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , 
 n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , 
 n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , 
 n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , 
 n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , 
 n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , 
 n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , 
 n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , 
 n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , 
 n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , 
 n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , 
 n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , 
 n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , 
 n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , 
 n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , 
 n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , 
 n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , 
 n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , 
 n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , 
 n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , 
 n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , 
 n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , 
 n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , 
 n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , 
 n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , 
 n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , 
 n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , 
 n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , 
 n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , 
 n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , 
 n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , 
 n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , 
 n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , 
 n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , 
 n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , 
 n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , 
 n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , 
 n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , 
 n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , 
 n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , 
 n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , 
 n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , 
 n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , 
 n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , 
 n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , 
 n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , 
 n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , 
 n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , 
 n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , 
 n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , 
 n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , 
 n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , 
 n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , 
 n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , 
 n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , 
 n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , 
 n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , 
 n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , 
 n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , 
 n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , 
 n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , 
 n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , 
 n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , 
 n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , 
 n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , 
 n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , 
 n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , 
 n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , 
 n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , 
 n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , 
 n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , 
 n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , 
 n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , 
 n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , 
 n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , 
 n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , 
 n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , 
 n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , 
 n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , 
 n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , 
 n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , 
 n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , 
 n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , 
 n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , 
 n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , 
 n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , 
 n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , 
 n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , 
 n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , 
 n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , 
 n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , 
 n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , 
 n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , 
 n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , 
 n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , 
 n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , 
 n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , 
 n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , 
 n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , 
 n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , 
 n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , 
 n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , 
 n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , 
 n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , 
 n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , 
 n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , 
 n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , 
 n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , 
 n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , 
 n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , 
 n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , 
 n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , 
 n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , 
 n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , 
 n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , 
 n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , 
 n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , 
 n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , 
 n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , 
 n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , 
 n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , 
 n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , 
 n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , 
 n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , 
 n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , 
 n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , 
 n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , 
 n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , 
 n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , 
 n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , 
 n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , 
 n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , 
 n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , 
 n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , 
 n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , 
 n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , 
 n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , 
 n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , 
 n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , 
 n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , 
 n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , 
 n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , 
 n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , 
 n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , 
 n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , 
 n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , 
 n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , 
 n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , 
 n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , 
 n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , 
 n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , 
 n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , 
 n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , 
 n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , 
 n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , 
 n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , 
 n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , 
 n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , 
 n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , 
 n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , 
 n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , 
 n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , 
 n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , 
 n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , 
 n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , 
 n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , 
 n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , 
 n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , 
 n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , 
 n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , 
 n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , 
 n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , 
 n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , 
 n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , 
 n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , 
 n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , 
 n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , 
 n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , 
 n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , 
 n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , 
 n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , 
 n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , 
 n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , 
 n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , 
 n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , 
 n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , 
 n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , 
 n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , 
 n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , 
 n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , 
 n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , 
 n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , 
 n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , 
 n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , 
 n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , 
 n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , 
 n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , 
 n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , 
 n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , 
 n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , 
 n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , 
 n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , 
 n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , 
 n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , 
 n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , 
 n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , 
 n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , 
 n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , 
 n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , 
 n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , 
 n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , 
 n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , 
 n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , 
 n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , 
 n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , 
 n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , 
 n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , 
 n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , 
 n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , 
 n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , 
 n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , 
 n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , 
 n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , 
 n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , 
 n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , 
 n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , 
 n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , 
 n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , 
 n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , 
 n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , 
 n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , 
 n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , 
 n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , 
 n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , 
 n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , 
 n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , 
 n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , 
 n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , 
 n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , 
 n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , 
 n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , 
 n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , 
 n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , 
 n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , 
 n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , 
 n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , 
 n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , 
 n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , 
 n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , 
 n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , 
 n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , 
 n10321 , C0n , C0 ;
buf ( n370 , n0 );
buf ( n371 , n1 );
buf ( n372 , n2 );
buf ( n373 , n3 );
buf ( n374 , n4 );
buf ( n375 , n5 );
buf ( n376 , n6 );
buf ( n377 , n7 );
buf ( n378 , n8 );
buf ( n379 , n9 );
buf ( n380 , n10 );
buf ( n381 , n11 );
buf ( n382 , n12 );
buf ( n383 , n13 );
buf ( n384 , n14 );
buf ( n385 , n15 );
buf ( n386 , n16 );
buf ( n387 , n17 );
buf ( n388 , n18 );
buf ( n389 , n19 );
buf ( n390 , n20 );
buf ( n391 , n21 );
buf ( n392 , n22 );
buf ( n393 , n23 );
buf ( n394 , n24 );
buf ( n395 , n25 );
buf ( n396 , n26 );
buf ( n397 , n27 );
buf ( n398 , n28 );
buf ( n399 , n29 );
buf ( n400 , n30 );
buf ( n401 , n31 );
buf ( n402 , n32 );
buf ( n403 , n33 );
buf ( n404 , n34 );
buf ( n405 , n35 );
buf ( n406 , n36 );
buf ( n407 , n37 );
buf ( n408 , n38 );
buf ( n409 , n39 );
buf ( n410 , n40 );
buf ( n411 , n41 );
buf ( n412 , n42 );
buf ( n413 , n43 );
buf ( n414 , n44 );
buf ( n415 , n45 );
buf ( n416 , n46 );
buf ( n417 , n47 );
buf ( n418 , n48 );
buf ( n419 , n49 );
buf ( n420 , n50 );
buf ( n421 , n51 );
buf ( n422 , n52 );
buf ( n423 , n53 );
buf ( n424 , n54 );
buf ( n425 , n55 );
buf ( n56 , n426 );
buf ( n57 , n427 );
buf ( n58 , n428 );
buf ( n59 , n429 );
buf ( n60 , n430 );
buf ( n61 , n431 );
buf ( n62 , n432 );
buf ( n63 , n433 );
buf ( n64 , n434 );
buf ( n65 , n435 );
buf ( n66 , n436 );
buf ( n67 , n437 );
buf ( n68 , n438 );
buf ( n69 , n439 );
buf ( n70 , n440 );
buf ( n71 , n441 );
buf ( n72 , n442 );
buf ( n73 , n443 );
buf ( n74 , n444 );
buf ( n75 , n445 );
buf ( n76 , n446 );
buf ( n77 , n447 );
buf ( n78 , n448 );
buf ( n79 , n449 );
buf ( n80 , n450 );
buf ( n81 , n451 );
buf ( n82 , n452 );
buf ( n83 , n453 );
buf ( n84 , n454 );
buf ( n85 , n455 );
buf ( n86 , n456 );
buf ( n87 , n457 );
buf ( n88 , n458 );
buf ( n89 , n459 );
buf ( n90 , n460 );
buf ( n91 , n461 );
buf ( n92 , n462 );
buf ( n93 , n463 );
buf ( n94 , n464 );
buf ( n95 , n465 );
buf ( n96 , n466 );
buf ( n97 , n467 );
buf ( n98 , n468 );
buf ( n99 , n469 );
buf ( n100 , n470 );
buf ( n101 , n471 );
buf ( n102 , n472 );
buf ( n103 , n473 );
buf ( n104 , n474 );
buf ( n105 , n475 );
buf ( n106 , n476 );
buf ( n107 , n477 );
buf ( n108 , n478 );
buf ( n109 , n479 );
buf ( n110 , n480 );
buf ( n111 , n481 );
buf ( n112 , n482 );
buf ( n113 , n483 );
buf ( n114 , n484 );
buf ( n115 , n485 );
buf ( n116 , n486 );
buf ( n117 , n487 );
buf ( n118 , n488 );
buf ( n119 , n489 );
buf ( n120 , n490 );
buf ( n121 , n491 );
buf ( n122 , n492 );
buf ( n123 , n493 );
buf ( n124 , n494 );
buf ( n125 , n495 );
buf ( n126 , n496 );
buf ( n127 , n497 );
buf ( n128 , n498 );
buf ( n129 , n499 );
buf ( n130 , n500 );
buf ( n131 , n501 );
buf ( n132 , n502 );
buf ( n133 , n503 );
buf ( n134 , n504 );
buf ( n135 , n505 );
buf ( n136 , n506 );
buf ( n137 , n507 );
buf ( n138 , n508 );
buf ( n139 , n509 );
buf ( n140 , n510 );
buf ( n141 , n511 );
buf ( n142 , n512 );
buf ( n143 , n513 );
buf ( n144 , n514 );
buf ( n145 , n515 );
buf ( n146 , n516 );
buf ( n147 , n517 );
buf ( n148 , n518 );
buf ( n149 , n519 );
buf ( n150 , n520 );
buf ( n151 , n521 );
buf ( n152 , n522 );
buf ( n153 , n523 );
buf ( n154 , n524 );
buf ( n155 , n525 );
buf ( n156 , n526 );
buf ( n157 , n527 );
buf ( n158 , n528 );
buf ( n159 , n529 );
buf ( n160 , n530 );
buf ( n161 , n531 );
buf ( n162 , n532 );
buf ( n163 , n533 );
buf ( n164 , n534 );
buf ( n165 , n535 );
buf ( n166 , n536 );
buf ( n167 , n537 );
buf ( n168 , n538 );
buf ( n169 , n539 );
buf ( n170 , n540 );
buf ( n171 , n541 );
buf ( n172 , n542 );
buf ( n173 , n543 );
buf ( n174 , n544 );
buf ( n175 , n545 );
buf ( n176 , n546 );
buf ( n177 , n547 );
buf ( n178 , n548 );
buf ( n179 , n549 );
buf ( n180 , n550 );
buf ( n181 , n551 );
buf ( n182 , n552 );
buf ( n183 , n553 );
buf ( n184 , n554 );
buf ( n426 , C0 );
buf ( n427 , C0 );
buf ( n428 , C0 );
buf ( n429 , C0 );
buf ( n430 , C0 );
buf ( n431 , C0 );
buf ( n432 , C0 );
buf ( n433 , C0 );
buf ( n434 , C0 );
buf ( n435 , C0 );
buf ( n436 , C0 );
buf ( n437 , C0 );
buf ( n438 , C0 );
buf ( n439 , C0 );
buf ( n440 , C0 );
buf ( n441 , C0 );
buf ( n442 , C0 );
buf ( n443 , C0 );
buf ( n444 , C0 );
buf ( n445 , C0 );
buf ( n446 , C0 );
buf ( n447 , C0 );
buf ( n448 , C0 );
buf ( n449 , C0 );
buf ( n450 , C0 );
buf ( n451 , C0 );
buf ( n452 , C0 );
buf ( n453 , C0 );
buf ( n454 , C0 );
buf ( n455 , C0 );
buf ( n456 , C0 );
buf ( n457 , C0 );
buf ( n458 , C0 );
buf ( n459 , C0 );
buf ( n460 , C0 );
buf ( n461 , C0 );
buf ( n462 , C0 );
buf ( n463 , C0 );
buf ( n464 , C0 );
buf ( n465 , C0 );
buf ( n466 , C0 );
buf ( n467 , C0 );
buf ( n468 , C0 );
buf ( n469 , C0 );
buf ( n470 , C0 );
buf ( n471 , C0 );
buf ( n472 , C0 );
buf ( n473 , C0 );
buf ( n474 , C0 );
buf ( n475 , C0 );
buf ( n476 , C0 );
buf ( n477 , C0 );
buf ( n478 , C0 );
buf ( n479 , C0 );
buf ( n480 , C0 );
buf ( n481 , C0 );
buf ( n482 , C0 );
buf ( n483 , C0 );
buf ( n484 , C0 );
buf ( n485 , C0 );
buf ( n486 , C0 );
buf ( n487 , C0 );
buf ( n488 , C0 );
buf ( n489 , C0 );
buf ( n490 , n10187 );
buf ( n491 , n10189 );
buf ( n492 , n10191 );
buf ( n493 , n10193 );
buf ( n494 , n10195 );
buf ( n495 , n10197 );
buf ( n496 , n10199 );
buf ( n497 , n10201 );
buf ( n498 , n10203 );
buf ( n499 , n10205 );
buf ( n500 , n10207 );
buf ( n501 , n10209 );
buf ( n502 , n10211 );
buf ( n503 , n10213 );
buf ( n504 , n10215 );
buf ( n505 , n10217 );
buf ( n506 , n10219 );
buf ( n507 , n10221 );
buf ( n508 , n10223 );
buf ( n509 , n10225 );
buf ( n510 , n10227 );
buf ( n511 , n10229 );
buf ( n512 , n10231 );
buf ( n513 , n10233 );
buf ( n514 , n10235 );
buf ( n515 , n10237 );
buf ( n516 , n10239 );
buf ( n517 , n10241 );
buf ( n518 , n10243 );
buf ( n519 , n10245 );
buf ( n520 , n10247 );
buf ( n521 , n10249 );
buf ( n522 , n10251 );
buf ( n523 , n10253 );
buf ( n524 , n10255 );
buf ( n525 , n10257 );
buf ( n526 , n10259 );
buf ( n527 , n10261 );
buf ( n528 , n10263 );
buf ( n529 , n10265 );
buf ( n530 , n10267 );
buf ( n531 , n10269 );
buf ( n532 , n10271 );
buf ( n533 , n10273 );
buf ( n534 , n10275 );
buf ( n535 , n10277 );
buf ( n536 , n10279 );
buf ( n537 , n10281 );
buf ( n538 , n10283 );
buf ( n539 , n10285 );
buf ( n540 , n10287 );
buf ( n541 , n10289 );
buf ( n542 , n10291 );
buf ( n543 , n10293 );
buf ( n544 , n10295 );
buf ( n545 , n10297 );
buf ( n546 , n10299 );
buf ( n547 , n10301 );
buf ( n548 , n10303 );
buf ( n549 , n10305 );
buf ( n550 , n10307 );
buf ( n551 , n10310 );
buf ( n552 , n10313 );
buf ( n553 , n10317 );
buf ( n554 , n10321 );
buf ( n555 , n418 );
buf ( n556 , n555 );
buf ( n557 , n556 );
buf ( n558 , n419 );
buf ( n559 , n558 );
buf ( n560 , n418 );
buf ( n561 , n560 );
and ( n562 , n559 , n561 );
buf ( n563 , n419 );
buf ( n564 , n563 );
and ( n565 , n556 , n564 );
and ( n566 , n562 , n565 );
and ( n567 , n557 , n566 );
xor ( n568 , n557 , n566 );
buf ( n569 , n420 );
buf ( n570 , n569 );
and ( n571 , n556 , n570 );
buf ( n572 , n559 );
or ( n573 , n571 , n572 );
xor ( n574 , n562 , n565 );
and ( n575 , n573 , n574 );
buf ( n576 , n420 );
buf ( n577 , n576 );
and ( n578 , n577 , n561 );
xnor ( n579 , n571 , n572 );
and ( n580 , n578 , n579 );
and ( n581 , n574 , n580 );
and ( n582 , n573 , n580 );
or ( n583 , n575 , n581 , n582 );
and ( n584 , n568 , n583 );
buf ( n585 , n421 );
buf ( n586 , n585 );
and ( n587 , n556 , n586 );
buf ( n588 , n421 );
buf ( n589 , n588 );
and ( n590 , n589 , n561 );
and ( n591 , n587 , n590 );
and ( n592 , n577 , n564 );
and ( n593 , n559 , n570 );
and ( n594 , n592 , n593 );
and ( n595 , n591 , n594 );
xor ( n596 , n587 , n590 );
buf ( n597 , n422 );
buf ( n598 , n597 );
and ( n599 , n556 , n598 );
buf ( n600 , n422 );
buf ( n601 , n600 );
and ( n602 , n601 , n561 );
and ( n603 , n599 , n602 );
and ( n604 , n596 , n603 );
and ( n605 , n559 , n586 );
and ( n606 , n589 , n564 );
and ( n607 , n605 , n606 );
and ( n608 , n603 , n607 );
and ( n609 , n596 , n607 );
or ( n610 , n604 , n608 , n609 );
and ( n611 , n594 , n610 );
and ( n612 , n591 , n610 );
or ( n613 , n595 , n611 , n612 );
xor ( n614 , n573 , n574 );
xor ( n615 , n614 , n580 );
and ( n616 , n613 , n615 );
xor ( n617 , n578 , n579 );
xor ( n618 , n592 , n593 );
buf ( n619 , n577 );
xor ( n620 , n599 , n602 );
and ( n621 , n619 , n620 );
and ( n622 , n618 , n621 );
xor ( n623 , n605 , n606 );
buf ( n624 , n423 );
buf ( n625 , n624 );
and ( n626 , n556 , n625 );
buf ( n627 , n423 );
buf ( n628 , n627 );
and ( n629 , n628 , n561 );
and ( n630 , n626 , n629 );
and ( n631 , n623 , n630 );
and ( n632 , n559 , n598 );
and ( n633 , n601 , n564 );
and ( n634 , n632 , n633 );
and ( n635 , n630 , n634 );
and ( n636 , n623 , n634 );
or ( n637 , n631 , n635 , n636 );
and ( n638 , n621 , n637 );
and ( n639 , n618 , n637 );
or ( n640 , n622 , n638 , n639 );
and ( n641 , n617 , n640 );
xor ( n642 , n591 , n594 );
xor ( n643 , n642 , n610 );
and ( n644 , n640 , n643 );
and ( n645 , n617 , n643 );
or ( n646 , n641 , n644 , n645 );
and ( n647 , n615 , n646 );
and ( n648 , n613 , n646 );
or ( n649 , n616 , n647 , n648 );
and ( n650 , n583 , n649 );
and ( n651 , n568 , n649 );
or ( n652 , n584 , n650 , n651 );
and ( n653 , n567 , n652 );
xor ( n654 , n567 , n652 );
xor ( n655 , n568 , n583 );
xor ( n656 , n655 , n649 );
xor ( n657 , n613 , n615 );
xor ( n658 , n657 , n646 );
xor ( n659 , n596 , n603 );
xor ( n660 , n659 , n607 );
and ( n661 , n577 , n586 );
and ( n662 , n589 , n570 );
and ( n663 , n661 , n662 );
and ( n664 , n628 , n564 );
and ( n665 , n601 , n570 );
or ( n666 , n664 , n665 );
and ( n667 , n559 , n625 );
and ( n668 , n577 , n598 );
or ( n669 , n667 , n668 );
and ( n670 , n666 , n669 );
and ( n671 , n663 , n670 );
xor ( n672 , n626 , n629 );
xor ( n673 , n632 , n633 );
and ( n674 , n672 , n673 );
and ( n675 , n670 , n674 );
and ( n676 , n663 , n674 );
or ( n677 , n671 , n675 , n676 );
and ( n678 , n660 , n677 );
xor ( n679 , n661 , n662 );
buf ( n680 , n589 );
buf ( n681 , n418 );
buf ( n682 , n681 );
or ( n683 , n680 , n682 );
and ( n684 , n679 , n683 );
buf ( n685 , n424 );
buf ( n686 , n685 );
and ( n687 , n556 , n686 );
buf ( n688 , n424 );
buf ( n689 , n688 );
and ( n690 , n689 , n561 );
and ( n691 , n687 , n690 );
and ( n692 , n683 , n691 );
and ( n693 , n679 , n691 );
or ( n694 , n684 , n692 , n693 );
xor ( n695 , n619 , n620 );
and ( n696 , n694 , n695 );
xor ( n697 , n623 , n630 );
xor ( n698 , n697 , n634 );
and ( n699 , n695 , n698 );
and ( n700 , n694 , n698 );
or ( n701 , n696 , n699 , n700 );
and ( n702 , n677 , n701 );
and ( n703 , n660 , n701 );
or ( n704 , n678 , n702 , n703 );
xor ( n705 , n617 , n640 );
xor ( n706 , n705 , n643 );
and ( n707 , n704 , n706 );
xor ( n708 , n618 , n621 );
xor ( n709 , n708 , n637 );
xor ( n710 , n666 , n669 );
buf ( n711 , n425 );
buf ( n712 , n711 );
and ( n713 , n556 , n712 );
buf ( n714 , n425 );
buf ( n715 , n714 );
and ( n716 , n715 , n561 );
and ( n717 , n713 , n716 );
xnor ( n718 , n680 , n682 );
and ( n719 , n717 , n718 );
and ( n720 , n710 , n719 );
and ( n721 , n628 , n570 );
and ( n722 , n601 , n586 );
or ( n723 , n721 , n722 );
and ( n724 , n577 , n625 );
and ( n725 , n589 , n598 );
or ( n726 , n724 , n725 );
and ( n727 , n723 , n726 );
and ( n728 , n719 , n727 );
and ( n729 , n710 , n727 );
or ( n730 , n720 , n728 , n729 );
xnor ( n731 , n664 , n665 );
xnor ( n732 , n667 , n668 );
and ( n733 , n731 , n732 );
xor ( n734 , n672 , n673 );
and ( n735 , n733 , n734 );
xor ( n736 , n679 , n683 );
xor ( n737 , n736 , n691 );
and ( n738 , n734 , n737 );
and ( n739 , n733 , n737 );
or ( n740 , n735 , n738 , n739 );
and ( n741 , n730 , n740 );
xor ( n742 , n663 , n670 );
xor ( n743 , n742 , n674 );
and ( n744 , n740 , n743 );
and ( n745 , n730 , n743 );
or ( n746 , n741 , n744 , n745 );
and ( n747 , n709 , n746 );
xor ( n748 , n660 , n677 );
xor ( n749 , n748 , n701 );
and ( n750 , n746 , n749 );
and ( n751 , n709 , n749 );
or ( n752 , n747 , n750 , n751 );
and ( n753 , n706 , n752 );
and ( n754 , n704 , n752 );
or ( n755 , n707 , n753 , n754 );
or ( n756 , n658 , n755 );
or ( n757 , n656 , n756 );
or ( n758 , n654 , n757 );
and ( n759 , n653 , n758 );
not ( n760 , n759 );
xor ( n761 , n653 , n758 );
not ( n762 , n761 );
xnor ( n763 , n654 , n757 );
xnor ( n764 , n656 , n756 );
xnor ( n765 , n658 , n755 );
xor ( n766 , n704 , n706 );
xor ( n767 , n766 , n752 );
xor ( n768 , n694 , n695 );
xor ( n769 , n768 , n698 );
xor ( n770 , n687 , n690 );
and ( n771 , n559 , n686 );
and ( n772 , n689 , n564 );
and ( n773 , n771 , n772 );
and ( n774 , n770 , n773 );
xor ( n775 , n717 , n718 );
and ( n776 , n773 , n775 );
and ( n777 , n770 , n775 );
or ( n778 , n774 , n776 , n777 );
xor ( n779 , n723 , n726 );
xor ( n780 , n731 , n732 );
and ( n781 , n779 , n780 );
and ( n782 , n689 , n570 );
and ( n783 , n628 , n586 );
and ( n784 , n782 , n783 );
and ( n785 , n577 , n686 );
and ( n786 , n589 , n625 );
and ( n787 , n785 , n786 );
and ( n788 , n784 , n787 );
and ( n789 , n780 , n788 );
and ( n790 , n779 , n788 );
or ( n791 , n781 , n789 , n790 );
and ( n792 , n778 , n791 );
xor ( n793 , n710 , n719 );
xor ( n794 , n793 , n727 );
and ( n795 , n791 , n794 );
and ( n796 , n778 , n794 );
or ( n797 , n792 , n795 , n796 );
and ( n798 , n769 , n797 );
xor ( n799 , n730 , n740 );
xor ( n800 , n799 , n743 );
and ( n801 , n797 , n800 );
and ( n802 , n769 , n800 );
or ( n803 , n798 , n801 , n802 );
xor ( n804 , n709 , n746 );
xor ( n805 , n804 , n749 );
and ( n806 , n803 , n805 );
xor ( n807 , n733 , n734 );
xor ( n808 , n807 , n737 );
xnor ( n809 , n721 , n722 );
xnor ( n810 , n724 , n725 );
and ( n811 , n809 , n810 );
buf ( n812 , n419 );
buf ( n813 , n812 );
buf ( n814 , n370 );
buf ( n815 , n814 );
not ( n816 , n815 );
and ( n817 , n813 , n816 );
xor ( n818 , n713 , n716 );
and ( n819 , n816 , n818 );
and ( n820 , n813 , n818 );
or ( n821 , n817 , n819 , n820 );
and ( n822 , n811 , n821 );
buf ( n823 , n601 );
buf ( n824 , n420 );
buf ( n825 , n824 );
and ( n826 , n823 , n825 );
buf ( n827 , n371 );
buf ( n828 , n827 );
not ( n829 , n828 );
and ( n830 , n825 , n829 );
and ( n831 , n823 , n829 );
or ( n832 , n826 , n830 , n831 );
xor ( n833 , n782 , n783 );
xor ( n834 , n785 , n786 );
and ( n835 , n833 , n834 );
and ( n836 , n832 , n835 );
and ( n837 , n821 , n836 );
and ( n838 , n811 , n836 );
or ( n839 , n822 , n837 , n838 );
and ( n840 , n808 , n839 );
xor ( n841 , n771 , n772 );
and ( n842 , n559 , n712 );
and ( n843 , n715 , n564 );
and ( n844 , n842 , n843 );
and ( n845 , n841 , n844 );
xor ( n846 , n784 , n787 );
and ( n847 , n844 , n846 );
and ( n848 , n841 , n846 );
or ( n849 , n845 , n847 , n848 );
xor ( n850 , n809 , n810 );
and ( n851 , n715 , n570 );
and ( n852 , n689 , n586 );
and ( n853 , n851 , n852 );
and ( n854 , n628 , n598 );
and ( n855 , n852 , n854 );
and ( n856 , n851 , n854 );
or ( n857 , n853 , n855 , n856 );
and ( n858 , n577 , n712 );
and ( n859 , n589 , n686 );
and ( n860 , n858 , n859 );
and ( n861 , n601 , n625 );
and ( n862 , n859 , n861 );
and ( n863 , n858 , n861 );
or ( n864 , n860 , n862 , n863 );
and ( n865 , n857 , n864 );
and ( n866 , n850 , n865 );
xor ( n867 , n813 , n816 );
xor ( n868 , n867 , n818 );
and ( n869 , n865 , n868 );
and ( n870 , n850 , n868 );
or ( n871 , n866 , n869 , n870 );
and ( n872 , n849 , n871 );
xor ( n873 , n770 , n773 );
xor ( n874 , n873 , n775 );
and ( n875 , n871 , n874 );
and ( n876 , n849 , n874 );
or ( n877 , n872 , n875 , n876 );
and ( n878 , n839 , n877 );
and ( n879 , n808 , n877 );
or ( n880 , n840 , n878 , n879 );
xor ( n881 , n769 , n797 );
xor ( n882 , n881 , n800 );
and ( n883 , n880 , n882 );
xor ( n884 , n778 , n791 );
xor ( n885 , n884 , n794 );
xor ( n886 , n779 , n780 );
xor ( n887 , n886 , n788 );
xor ( n888 , n832 , n835 );
and ( n889 , n601 , n686 );
and ( n890 , n689 , n598 );
and ( n891 , n889 , n890 );
buf ( n892 , n421 );
buf ( n893 , n892 );
and ( n894 , n891 , n893 );
buf ( n895 , n372 );
buf ( n896 , n895 );
not ( n897 , n896 );
and ( n898 , n893 , n897 );
and ( n899 , n891 , n897 );
or ( n900 , n894 , n898 , n899 );
xor ( n901 , n851 , n852 );
xor ( n902 , n901 , n854 );
xor ( n903 , n858 , n859 );
xor ( n904 , n903 , n861 );
and ( n905 , n902 , n904 );
and ( n906 , n900 , n905 );
xor ( n907 , n823 , n825 );
xor ( n908 , n907 , n829 );
and ( n909 , n905 , n908 );
and ( n910 , n900 , n908 );
or ( n911 , n906 , n909 , n910 );
and ( n912 , n888 , n911 );
xor ( n913 , n842 , n843 );
xor ( n914 , n857 , n864 );
and ( n915 , n913 , n914 );
xor ( n916 , n833 , n834 );
and ( n917 , n914 , n916 );
and ( n918 , n913 , n916 );
or ( n919 , n915 , n917 , n918 );
and ( n920 , n911 , n919 );
and ( n921 , n888 , n919 );
or ( n922 , n912 , n920 , n921 );
and ( n923 , n887 , n922 );
xor ( n924 , n811 , n821 );
xor ( n925 , n924 , n836 );
and ( n926 , n922 , n925 );
and ( n927 , n887 , n925 );
or ( n928 , n923 , n926 , n927 );
and ( n929 , n885 , n928 );
xor ( n930 , n808 , n839 );
xor ( n931 , n930 , n877 );
and ( n932 , n928 , n931 );
and ( n933 , n885 , n931 );
or ( n934 , n929 , n932 , n933 );
and ( n935 , n882 , n934 );
and ( n936 , n880 , n934 );
or ( n937 , n883 , n935 , n936 );
and ( n938 , n805 , n937 );
and ( n939 , n803 , n937 );
or ( n940 , n806 , n938 , n939 );
and ( n941 , n767 , n940 );
xor ( n942 , n767 , n940 );
xor ( n943 , n803 , n805 );
xor ( n944 , n943 , n937 );
not ( n945 , n944 );
xor ( n946 , n880 , n882 );
xor ( n947 , n946 , n934 );
xor ( n948 , n849 , n871 );
xor ( n949 , n948 , n874 );
xor ( n950 , n841 , n844 );
xor ( n951 , n950 , n846 );
xor ( n952 , n850 , n865 );
xor ( n953 , n952 , n868 );
and ( n954 , n951 , n953 );
buf ( n955 , n628 );
buf ( n956 , n422 );
buf ( n957 , n956 );
and ( n958 , n955 , n957 );
buf ( n959 , n373 );
buf ( n960 , n959 );
not ( n961 , n960 );
and ( n962 , n957 , n961 );
and ( n963 , n955 , n961 );
or ( n964 , n958 , n962 , n963 );
and ( n965 , n589 , n712 );
and ( n966 , n715 , n586 );
and ( n967 , n965 , n966 );
and ( n968 , n964 , n967 );
xor ( n969 , n891 , n893 );
xor ( n970 , n969 , n897 );
and ( n971 , n967 , n970 );
and ( n972 , n964 , n970 );
or ( n973 , n968 , n971 , n972 );
xor ( n974 , n900 , n905 );
xor ( n975 , n974 , n908 );
or ( n976 , n973 , n975 );
and ( n977 , n953 , n976 );
and ( n978 , n951 , n976 );
or ( n979 , n954 , n977 , n978 );
and ( n980 , n949 , n979 );
xor ( n981 , n887 , n922 );
xor ( n982 , n981 , n925 );
and ( n983 , n979 , n982 );
and ( n984 , n949 , n982 );
or ( n985 , n980 , n983 , n984 );
xor ( n986 , n885 , n928 );
xor ( n987 , n986 , n931 );
and ( n988 , n985 , n987 );
xor ( n989 , n888 , n911 );
xor ( n990 , n989 , n919 );
xor ( n991 , n902 , n904 );
and ( n992 , n715 , n598 );
and ( n993 , n689 , n625 );
or ( n994 , n992 , n993 );
and ( n995 , n601 , n712 );
and ( n996 , n628 , n686 );
or ( n997 , n995 , n996 );
and ( n998 , n994 , n997 );
and ( n999 , n991 , n998 );
xor ( n1000 , n955 , n957 );
xor ( n1001 , n1000 , n961 );
xor ( n1002 , n965 , n966 );
and ( n1003 , n1001 , n1002 );
xor ( n1004 , n889 , n890 );
and ( n1005 , n1002 , n1004 );
and ( n1006 , n1001 , n1004 );
or ( n1007 , n1003 , n1005 , n1006 );
and ( n1008 , n998 , n1007 );
and ( n1009 , n991 , n1007 );
or ( n1010 , n999 , n1008 , n1009 );
xor ( n1011 , n913 , n914 );
xor ( n1012 , n1011 , n916 );
and ( n1013 , n1010 , n1012 );
xnor ( n1014 , n973 , n975 );
and ( n1015 , n1012 , n1014 );
and ( n1016 , n1010 , n1014 );
or ( n1017 , n1013 , n1015 , n1016 );
and ( n1018 , n990 , n1017 );
xor ( n1019 , n951 , n953 );
xor ( n1020 , n1019 , n976 );
and ( n1021 , n1017 , n1020 );
and ( n1022 , n990 , n1020 );
or ( n1023 , n1018 , n1021 , n1022 );
xor ( n1024 , n949 , n979 );
xor ( n1025 , n1024 , n982 );
and ( n1026 , n1023 , n1025 );
xor ( n1027 , n990 , n1017 );
xor ( n1028 , n1027 , n1020 );
xor ( n1029 , n964 , n967 );
xor ( n1030 , n1029 , n970 );
xor ( n1031 , n994 , n997 );
buf ( n1032 , n424 );
buf ( n1033 , n1032 );
buf ( n1034 , n1033 );
buf ( n1035 , n423 );
buf ( n1036 , n1035 );
and ( n1037 , n1034 , n1036 );
buf ( n1038 , n374 );
buf ( n1039 , n1038 );
not ( n1040 , n1039 );
and ( n1041 , n1036 , n1040 );
and ( n1042 , n1034 , n1040 );
or ( n1043 , n1037 , n1041 , n1042 );
and ( n1044 , n1031 , n1043 );
xnor ( n1045 , n992 , n993 );
xnor ( n1046 , n995 , n996 );
and ( n1047 , n1045 , n1046 );
and ( n1048 , n1043 , n1047 );
and ( n1049 , n1031 , n1047 );
or ( n1050 , n1044 , n1048 , n1049 );
and ( n1051 , n1030 , n1050 );
xor ( n1052 , n991 , n998 );
xor ( n1053 , n1052 , n1007 );
and ( n1054 , n1050 , n1053 );
and ( n1055 , n1030 , n1053 );
or ( n1056 , n1051 , n1054 , n1055 );
xor ( n1057 , n1010 , n1012 );
xor ( n1058 , n1057 , n1014 );
and ( n1059 , n1056 , n1058 );
xor ( n1060 , n1001 , n1002 );
xor ( n1061 , n1060 , n1004 );
and ( n1062 , n628 , n712 );
and ( n1063 , n715 , n625 );
and ( n1064 , n1062 , n1063 );
xor ( n1065 , n1034 , n1036 );
xor ( n1066 , n1065 , n1040 );
and ( n1067 , n1064 , n1066 );
xor ( n1068 , n1045 , n1046 );
and ( n1069 , n1066 , n1068 );
and ( n1070 , n1064 , n1068 );
or ( n1071 , n1067 , n1069 , n1070 );
and ( n1072 , n1061 , n1071 );
xor ( n1073 , n1031 , n1043 );
xor ( n1074 , n1073 , n1047 );
and ( n1075 , n1071 , n1074 );
and ( n1076 , n1061 , n1074 );
or ( n1077 , n1072 , n1075 , n1076 );
xor ( n1078 , n1030 , n1050 );
xor ( n1079 , n1078 , n1053 );
and ( n1080 , n1077 , n1079 );
buf ( n1081 , n375 );
buf ( n1082 , n1081 );
not ( n1083 , n1082 );
xor ( n1084 , n1062 , n1063 );
and ( n1085 , n1083 , n1084 );
buf ( n1086 , n1085 );
and ( n1087 , n689 , n712 );
and ( n1088 , n715 , n686 );
and ( n1089 , n1087 , n1088 );
buf ( n1090 , n425 );
buf ( n1091 , n1090 );
buf ( n1092 , n376 );
buf ( n1093 , n1092 );
not ( n1094 , n1093 );
and ( n1095 , n1091 , n1094 );
xor ( n1096 , n1087 , n1088 );
and ( n1097 , n1094 , n1096 );
and ( n1098 , n1091 , n1096 );
or ( n1099 , n1095 , n1097 , n1098 );
and ( n1100 , n1089 , n1099 );
xor ( n1101 , n1083 , n1084 );
buf ( n1102 , n1101 );
and ( n1103 , n1099 , n1102 );
and ( n1104 , n1089 , n1102 );
or ( n1105 , n1100 , n1103 , n1104 );
and ( n1106 , n1086 , n1105 );
xor ( n1107 , n1064 , n1066 );
xor ( n1108 , n1107 , n1068 );
and ( n1109 , n1105 , n1108 );
and ( n1110 , n1086 , n1108 );
or ( n1111 , n1106 , n1109 , n1110 );
xor ( n1112 , n1061 , n1071 );
xor ( n1113 , n1112 , n1074 );
or ( n1114 , n1111 , n1113 );
and ( n1115 , n1079 , n1114 );
and ( n1116 , n1077 , n1114 );
or ( n1117 , n1080 , n1115 , n1116 );
and ( n1118 , n1058 , n1117 );
and ( n1119 , n1056 , n1117 );
or ( n1120 , n1059 , n1118 , n1119 );
or ( n1121 , n1028 , n1120 );
and ( n1122 , n1025 , n1121 );
and ( n1123 , n1023 , n1121 );
or ( n1124 , n1026 , n1122 , n1123 );
and ( n1125 , n987 , n1124 );
and ( n1126 , n985 , n1124 );
or ( n1127 , n988 , n1125 , n1126 );
and ( n1128 , n947 , n1127 );
xor ( n1129 , n947 , n1127 );
xor ( n1130 , n985 , n987 );
xor ( n1131 , n1130 , n1124 );
not ( n1132 , n1131 );
xor ( n1133 , n1023 , n1025 );
xor ( n1134 , n1133 , n1121 );
xnor ( n1135 , n1028 , n1120 );
xor ( n1136 , n1056 , n1058 );
xor ( n1137 , n1136 , n1117 );
xor ( n1138 , n1077 , n1079 );
xor ( n1139 , n1138 , n1114 );
not ( n1140 , n1139 );
xnor ( n1141 , n1111 , n1113 );
xor ( n1142 , n1086 , n1105 );
xor ( n1143 , n1142 , n1108 );
xor ( n1144 , n1089 , n1099 );
xor ( n1145 , n1144 , n1102 );
buf ( n1146 , n715 );
buf ( n1147 , n377 );
buf ( n1148 , n1147 );
not ( n1149 , n1148 );
and ( n1150 , n1146 , n1149 );
xor ( n1151 , n1091 , n1094 );
xor ( n1152 , n1151 , n1096 );
and ( n1153 , n1150 , n1152 );
xor ( n1154 , n1150 , n1152 );
xor ( n1155 , n1146 , n1149 );
and ( n1156 , n1154 , n1155 );
or ( n1157 , n1153 , n1156 );
and ( n1158 , n1145 , n1157 );
and ( n1159 , n1143 , n1158 );
and ( n1160 , n1141 , n1159 );
and ( n1161 , n1140 , n1160 );
or ( n1162 , n1139 , n1161 );
and ( n1163 , n1137 , n1162 );
and ( n1164 , n1135 , n1163 );
and ( n1165 , n1134 , n1164 );
and ( n1166 , n1132 , n1165 );
or ( n1167 , n1131 , n1166 );
and ( n1168 , n1129 , n1167 );
or ( n1169 , n1128 , n1168 );
and ( n1170 , n945 , n1169 );
or ( n1171 , n944 , n1170 );
and ( n1172 , n942 , n1171 );
or ( n1173 , n941 , n1172 );
and ( n1174 , n765 , n1173 );
and ( n1175 , n764 , n1174 );
and ( n1176 , n763 , n1175 );
and ( n1177 , n762 , n1176 );
or ( n1178 , n761 , n1177 );
and ( n1179 , n760 , n1178 );
or ( n1180 , n759 , n1179 );
not ( n1181 , n1180 );
buf ( n1182 , n1181 );
buf ( n1183 , n1182 );
buf ( n1184 , n1183 );
buf ( n1185 , n1184 );
buf ( n1186 , n410 );
buf ( n1187 , n1186 );
buf ( n1188 , n411 );
buf ( n1189 , n1188 );
xor ( n1190 , n1187 , n1189 );
not ( n1191 , n1190 );
and ( n1192 , n1187 , n1191 );
and ( n1193 , n1185 , n1192 );
buf ( n1194 , n413 );
buf ( n1195 , n1194 );
buf ( n1196 , n414 );
buf ( n1197 , n1196 );
buf ( n1198 , n415 );
buf ( n1199 , n1198 );
and ( n1200 , n1197 , n1199 );
not ( n1201 , n1200 );
and ( n1202 , n1195 , n1201 );
not ( n1203 , n1202 );
buf ( n1204 , n1181 );
buf ( n1205 , n1204 );
buf ( n1206 , n1205 );
buf ( n1207 , n1206 );
buf ( n1208 , n412 );
buf ( n1209 , n1208 );
xor ( n1210 , n1189 , n1209 );
xor ( n1211 , n1209 , n1195 );
not ( n1212 , n1211 );
and ( n1213 , n1210 , n1212 );
and ( n1214 , n1207 , n1213 );
and ( n1215 , n1185 , n1211 );
nor ( n1216 , n1214 , n1215 );
and ( n1217 , n1209 , n1195 );
not ( n1218 , n1217 );
and ( n1219 , n1189 , n1218 );
xnor ( n1220 , n1216 , n1219 );
and ( n1221 , n1203 , n1220 );
buf ( n1222 , n1181 );
buf ( n1223 , n1222 );
buf ( n1224 , n1223 );
buf ( n1225 , n1224 );
and ( n1226 , n1225 , n1192 );
buf ( n1227 , n1181 );
buf ( n1228 , n1227 );
buf ( n1229 , n1228 );
buf ( n1230 , n1229 );
and ( n1231 , n1230 , n1190 );
nor ( n1232 , n1226 , n1231 );
not ( n1233 , n1232 );
and ( n1234 , n1220 , n1233 );
and ( n1235 , n1203 , n1233 );
or ( n1236 , n1221 , n1234 , n1235 );
and ( n1237 , n1185 , n1213 );
not ( n1238 , n1237 );
xnor ( n1239 , n1238 , n1219 );
and ( n1240 , n1236 , n1239 );
and ( n1241 , n1230 , n1192 );
and ( n1242 , n1207 , n1190 );
nor ( n1243 , n1241 , n1242 );
and ( n1244 , n1239 , n1243 );
and ( n1245 , n1236 , n1243 );
or ( n1246 , n1240 , n1244 , n1245 );
not ( n1247 , n1219 );
or ( n1248 , n1246 , n1247 );
and ( n1249 , n1193 , n1248 );
and ( n1250 , n1207 , n1192 );
and ( n1251 , n1185 , n1190 );
nor ( n1252 , n1250 , n1251 );
not ( n1253 , n1252 );
not ( n1254 , n1243 );
buf ( n1255 , n1254 );
and ( n1256 , n1253 , n1255 );
and ( n1257 , n1248 , n1256 );
and ( n1258 , n1193 , n1256 );
or ( n1259 , n1249 , n1257 , n1258 );
not ( n1260 , n1259 );
xor ( n1261 , n1193 , n1248 );
xor ( n1262 , n1261 , n1256 );
xnor ( n1263 , n1246 , n1247 );
xor ( n1264 , n1253 , n1255 );
and ( n1265 , n1263 , n1264 );
xor ( n1266 , n1236 , n1239 );
xor ( n1267 , n1266 , n1243 );
xor ( n1268 , n1203 , n1220 );
xor ( n1269 , n1268 , n1233 );
xor ( n1270 , n1195 , n1197 );
xor ( n1271 , n1197 , n1199 );
not ( n1272 , n1271 );
and ( n1273 , n1270 , n1272 );
and ( n1274 , n1185 , n1273 );
not ( n1275 , n1274 );
xnor ( n1276 , n1275 , n1202 );
and ( n1277 , n1230 , n1213 );
and ( n1278 , n1207 , n1211 );
nor ( n1279 , n1277 , n1278 );
xnor ( n1280 , n1279 , n1219 );
and ( n1281 , n1276 , n1280 );
and ( n1282 , n1269 , n1281 );
and ( n1283 , n1230 , n1273 );
and ( n1284 , n1207 , n1271 );
nor ( n1285 , n1283 , n1284 );
xnor ( n1286 , n1285 , n1202 );
buf ( n1287 , n1181 );
buf ( n1288 , n1287 );
buf ( n1289 , n1288 );
buf ( n1290 , n1289 );
and ( n1291 , n1290 , n1192 );
buf ( n1292 , n1181 );
buf ( n1293 , n1292 );
buf ( n1294 , n1293 );
buf ( n1295 , n1294 );
and ( n1296 , n1295 , n1190 );
nor ( n1297 , n1291 , n1296 );
not ( n1298 , n1297 );
or ( n1299 , n1286 , n1298 );
buf ( n1300 , n416 );
buf ( n1301 , n1300 );
xor ( n1302 , n1199 , n1301 );
not ( n1303 , n1301 );
and ( n1304 , n1302 , n1303 );
and ( n1305 , n1185 , n1304 );
not ( n1306 , n1305 );
xnor ( n1307 , n1306 , n1199 );
buf ( n1308 , n1307 );
and ( n1309 , n1299 , n1308 );
and ( n1310 , n1225 , n1213 );
and ( n1311 , n1230 , n1211 );
nor ( n1312 , n1310 , n1311 );
xnor ( n1313 , n1312 , n1219 );
and ( n1314 , n1308 , n1313 );
and ( n1315 , n1299 , n1313 );
or ( n1316 , n1309 , n1314 , n1315 );
and ( n1317 , n1207 , n1273 );
and ( n1318 , n1185 , n1271 );
nor ( n1319 , n1317 , n1318 );
xnor ( n1320 , n1319 , n1202 );
and ( n1321 , n1295 , n1192 );
buf ( n1322 , n1181 );
buf ( n1323 , n1322 );
buf ( n1324 , n1323 );
buf ( n1325 , n1324 );
and ( n1326 , n1325 , n1190 );
nor ( n1327 , n1321 , n1326 );
not ( n1328 , n1327 );
or ( n1329 , n1320 , n1328 );
and ( n1330 , n1316 , n1329 );
and ( n1331 , n1281 , n1330 );
and ( n1332 , n1269 , n1330 );
or ( n1333 , n1282 , n1331 , n1332 );
and ( n1334 , n1267 , n1333 );
and ( n1335 , n1325 , n1192 );
and ( n1336 , n1225 , n1190 );
nor ( n1337 , n1335 , n1336 );
not ( n1338 , n1337 );
xor ( n1339 , n1276 , n1280 );
and ( n1340 , n1338 , n1339 );
xor ( n1341 , n1316 , n1329 );
and ( n1342 , n1339 , n1341 );
and ( n1343 , n1338 , n1341 );
or ( n1344 , n1340 , n1342 , n1343 );
xor ( n1345 , n1269 , n1281 );
xor ( n1346 , n1345 , n1330 );
and ( n1347 , n1344 , n1346 );
xor ( n1348 , n1299 , n1308 );
xor ( n1349 , n1348 , n1313 );
xnor ( n1350 , n1320 , n1328 );
or ( n1351 , n1349 , n1350 );
not ( n1352 , n1199 );
not ( n1353 , n1307 );
and ( n1354 , n1325 , n1213 );
and ( n1355 , n1225 , n1211 );
nor ( n1356 , n1354 , n1355 );
xnor ( n1357 , n1356 , n1219 );
and ( n1358 , n1353 , n1357 );
and ( n1359 , n1352 , n1358 );
xnor ( n1360 , n1286 , n1298 );
xor ( n1361 , n1353 , n1357 );
and ( n1362 , n1360 , n1361 );
and ( n1363 , n1207 , n1304 );
and ( n1364 , n1185 , n1301 );
nor ( n1365 , n1363 , n1364 );
xnor ( n1366 , n1365 , n1199 );
and ( n1367 , n1225 , n1273 );
and ( n1368 , n1230 , n1271 );
nor ( n1369 , n1367 , n1368 );
xnor ( n1370 , n1369 , n1202 );
and ( n1371 , n1366 , n1370 );
and ( n1372 , n1295 , n1213 );
and ( n1373 , n1325 , n1211 );
nor ( n1374 , n1372 , n1373 );
xnor ( n1375 , n1374 , n1219 );
and ( n1376 , n1370 , n1375 );
and ( n1377 , n1366 , n1375 );
or ( n1378 , n1371 , n1376 , n1377 );
and ( n1379 , n1361 , n1378 );
and ( n1380 , n1360 , n1378 );
or ( n1381 , n1362 , n1379 , n1380 );
and ( n1382 , n1358 , n1381 );
and ( n1383 , n1352 , n1381 );
or ( n1384 , n1359 , n1382 , n1383 );
and ( n1385 , n1351 , n1384 );
xor ( n1386 , n1338 , n1339 );
xor ( n1387 , n1386 , n1341 );
and ( n1388 , n1384 , n1387 );
and ( n1389 , n1351 , n1387 );
or ( n1390 , n1385 , n1388 , n1389 );
and ( n1391 , n1346 , n1390 );
and ( n1392 , n1344 , n1390 );
or ( n1393 , n1347 , n1391 , n1392 );
and ( n1394 , n1333 , n1393 );
and ( n1395 , n1267 , n1393 );
or ( n1396 , n1334 , n1394 , n1395 );
and ( n1397 , n1264 , n1396 );
and ( n1398 , n1263 , n1396 );
or ( n1399 , n1265 , n1397 , n1398 );
and ( n1400 , n1262 , n1399 );
xor ( n1401 , n1262 , n1399 );
xor ( n1402 , n1263 , n1264 );
xor ( n1403 , n1402 , n1396 );
xor ( n1404 , n1267 , n1333 );
xor ( n1405 , n1404 , n1393 );
xor ( n1406 , n1344 , n1346 );
xor ( n1407 , n1406 , n1390 );
xor ( n1408 , n1351 , n1384 );
xor ( n1409 , n1408 , n1387 );
xnor ( n1410 , n1349 , n1350 );
xor ( n1411 , n1352 , n1358 );
xor ( n1412 , n1411 , n1381 );
and ( n1413 , n1410 , n1412 );
buf ( n1414 , n1181 );
buf ( n1415 , n1414 );
buf ( n1416 , n1415 );
buf ( n1417 , n1416 );
and ( n1418 , n1417 , n1192 );
and ( n1419 , n1290 , n1190 );
nor ( n1420 , n1418 , n1419 );
not ( n1421 , n1420 );
xor ( n1422 , n1366 , n1370 );
xor ( n1423 , n1422 , n1375 );
and ( n1424 , n1421 , n1423 );
and ( n1425 , n1230 , n1304 );
and ( n1426 , n1207 , n1301 );
nor ( n1427 , n1425 , n1426 );
xnor ( n1428 , n1427 , n1199 );
and ( n1429 , n1325 , n1273 );
and ( n1430 , n1225 , n1271 );
nor ( n1431 , n1429 , n1430 );
xnor ( n1432 , n1431 , n1202 );
and ( n1433 , n1428 , n1432 );
and ( n1434 , n1290 , n1213 );
and ( n1435 , n1295 , n1211 );
nor ( n1436 , n1434 , n1435 );
xnor ( n1437 , n1436 , n1219 );
and ( n1438 , n1432 , n1437 );
and ( n1439 , n1428 , n1437 );
or ( n1440 , n1433 , n1438 , n1439 );
and ( n1441 , n1423 , n1440 );
and ( n1442 , n1421 , n1440 );
or ( n1443 , n1424 , n1441 , n1442 );
xor ( n1444 , n1360 , n1361 );
xor ( n1445 , n1444 , n1378 );
and ( n1446 , n1443 , n1445 );
buf ( n1447 , n1181 );
buf ( n1448 , n1447 );
buf ( n1449 , n1448 );
buf ( n1450 , n1449 );
and ( n1451 , n1450 , n1192 );
and ( n1452 , n1417 , n1190 );
nor ( n1453 , n1451 , n1452 );
not ( n1454 , n1453 );
xor ( n1455 , n1428 , n1432 );
xor ( n1456 , n1455 , n1437 );
and ( n1457 , n1454 , n1456 );
and ( n1458 , n1225 , n1304 );
and ( n1459 , n1230 , n1301 );
nor ( n1460 , n1458 , n1459 );
xnor ( n1461 , n1460 , n1199 );
and ( n1462 , n1295 , n1273 );
and ( n1463 , n1325 , n1271 );
nor ( n1464 , n1462 , n1463 );
xnor ( n1465 , n1464 , n1202 );
and ( n1466 , n1461 , n1465 );
and ( n1467 , n1417 , n1213 );
and ( n1468 , n1290 , n1211 );
nor ( n1469 , n1467 , n1468 );
xnor ( n1470 , n1469 , n1219 );
and ( n1471 , n1465 , n1470 );
and ( n1472 , n1461 , n1470 );
or ( n1473 , n1466 , n1471 , n1472 );
and ( n1474 , n1456 , n1473 );
and ( n1475 , n1454 , n1473 );
or ( n1476 , n1457 , n1474 , n1475 );
xor ( n1477 , n1421 , n1423 );
xor ( n1478 , n1477 , n1440 );
and ( n1479 , n1476 , n1478 );
buf ( n1480 , n1181 );
buf ( n1481 , n1480 );
buf ( n1482 , n1481 );
buf ( n1483 , n1482 );
and ( n1484 , n1483 , n1192 );
and ( n1485 , n1450 , n1190 );
nor ( n1486 , n1484 , n1485 );
not ( n1487 , n1486 );
xor ( n1488 , n1461 , n1465 );
xor ( n1489 , n1488 , n1470 );
and ( n1490 , n1487 , n1489 );
and ( n1491 , n1325 , n1304 );
and ( n1492 , n1225 , n1301 );
nor ( n1493 , n1491 , n1492 );
xnor ( n1494 , n1493 , n1199 );
and ( n1495 , n1290 , n1273 );
and ( n1496 , n1295 , n1271 );
nor ( n1497 , n1495 , n1496 );
xnor ( n1498 , n1497 , n1202 );
and ( n1499 , n1494 , n1498 );
and ( n1500 , n1450 , n1213 );
and ( n1501 , n1417 , n1211 );
nor ( n1502 , n1500 , n1501 );
xnor ( n1503 , n1502 , n1219 );
and ( n1504 , n1498 , n1503 );
and ( n1505 , n1494 , n1503 );
or ( n1506 , n1499 , n1504 , n1505 );
and ( n1507 , n1489 , n1506 );
and ( n1508 , n1487 , n1506 );
or ( n1509 , n1490 , n1507 , n1508 );
xor ( n1510 , n1454 , n1456 );
xor ( n1511 , n1510 , n1473 );
and ( n1512 , n1509 , n1511 );
buf ( n1513 , n1181 );
buf ( n1514 , n1513 );
buf ( n1515 , n1514 );
buf ( n1516 , n1515 );
and ( n1517 , n1516 , n1192 );
and ( n1518 , n1483 , n1190 );
nor ( n1519 , n1517 , n1518 );
not ( n1520 , n1519 );
xor ( n1521 , n1494 , n1498 );
xor ( n1522 , n1521 , n1503 );
and ( n1523 , n1520 , n1522 );
and ( n1524 , n1295 , n1304 );
and ( n1525 , n1325 , n1301 );
nor ( n1526 , n1524 , n1525 );
xnor ( n1527 , n1526 , n1199 );
and ( n1528 , n1417 , n1273 );
and ( n1529 , n1290 , n1271 );
nor ( n1530 , n1528 , n1529 );
xnor ( n1531 , n1530 , n1202 );
and ( n1532 , n1527 , n1531 );
and ( n1533 , n1483 , n1213 );
and ( n1534 , n1450 , n1211 );
nor ( n1535 , n1533 , n1534 );
xnor ( n1536 , n1535 , n1219 );
and ( n1537 , n1531 , n1536 );
and ( n1538 , n1527 , n1536 );
or ( n1539 , n1532 , n1537 , n1538 );
and ( n1540 , n1522 , n1539 );
and ( n1541 , n1520 , n1539 );
or ( n1542 , n1523 , n1540 , n1541 );
xor ( n1543 , n1487 , n1489 );
xor ( n1544 , n1543 , n1506 );
and ( n1545 , n1542 , n1544 );
buf ( n1546 , n1181 );
buf ( n1547 , n1546 );
buf ( n1548 , n1547 );
buf ( n1549 , n1548 );
and ( n1550 , n1549 , n1192 );
and ( n1551 , n1516 , n1190 );
nor ( n1552 , n1550 , n1551 );
not ( n1553 , n1552 );
xor ( n1554 , n1527 , n1531 );
xor ( n1555 , n1554 , n1536 );
and ( n1556 , n1553 , n1555 );
and ( n1557 , n1290 , n1304 );
and ( n1558 , n1295 , n1301 );
nor ( n1559 , n1557 , n1558 );
xnor ( n1560 , n1559 , n1199 );
and ( n1561 , n1450 , n1273 );
and ( n1562 , n1417 , n1271 );
nor ( n1563 , n1561 , n1562 );
xnor ( n1564 , n1563 , n1202 );
and ( n1565 , n1560 , n1564 );
and ( n1566 , n1516 , n1213 );
and ( n1567 , n1483 , n1211 );
nor ( n1568 , n1566 , n1567 );
xnor ( n1569 , n1568 , n1219 );
and ( n1570 , n1564 , n1569 );
and ( n1571 , n1560 , n1569 );
or ( n1572 , n1565 , n1570 , n1571 );
and ( n1573 , n1555 , n1572 );
and ( n1574 , n1553 , n1572 );
or ( n1575 , n1556 , n1573 , n1574 );
xor ( n1576 , n1520 , n1522 );
xor ( n1577 , n1576 , n1539 );
and ( n1578 , n1575 , n1577 );
buf ( n1579 , n1181 );
buf ( n1580 , n1579 );
buf ( n1581 , n1580 );
buf ( n1582 , n1581 );
and ( n1583 , n1582 , n1192 );
and ( n1584 , n1549 , n1190 );
nor ( n1585 , n1583 , n1584 );
not ( n1586 , n1585 );
xor ( n1587 , n1560 , n1564 );
xor ( n1588 , n1587 , n1569 );
and ( n1589 , n1586 , n1588 );
and ( n1590 , n1417 , n1304 );
and ( n1591 , n1290 , n1301 );
nor ( n1592 , n1590 , n1591 );
xnor ( n1593 , n1592 , n1199 );
and ( n1594 , n1483 , n1273 );
and ( n1595 , n1450 , n1271 );
nor ( n1596 , n1594 , n1595 );
xnor ( n1597 , n1596 , n1202 );
and ( n1598 , n1593 , n1597 );
and ( n1599 , n1549 , n1213 );
and ( n1600 , n1516 , n1211 );
nor ( n1601 , n1599 , n1600 );
xnor ( n1602 , n1601 , n1219 );
and ( n1603 , n1597 , n1602 );
and ( n1604 , n1593 , n1602 );
or ( n1605 , n1598 , n1603 , n1604 );
and ( n1606 , n1588 , n1605 );
and ( n1607 , n1586 , n1605 );
or ( n1608 , n1589 , n1606 , n1607 );
xor ( n1609 , n1553 , n1555 );
xor ( n1610 , n1609 , n1572 );
and ( n1611 , n1608 , n1610 );
buf ( n1612 , n1181 );
buf ( n1613 , n1612 );
buf ( n1614 , n1613 );
buf ( n1615 , n1614 );
and ( n1616 , n1615 , n1192 );
and ( n1617 , n1582 , n1190 );
nor ( n1618 , n1616 , n1617 );
not ( n1619 , n1618 );
xor ( n1620 , n1593 , n1597 );
xor ( n1621 , n1620 , n1602 );
and ( n1622 , n1619 , n1621 );
and ( n1623 , n1450 , n1304 );
and ( n1624 , n1417 , n1301 );
nor ( n1625 , n1623 , n1624 );
xnor ( n1626 , n1625 , n1199 );
and ( n1627 , n1516 , n1273 );
and ( n1628 , n1483 , n1271 );
nor ( n1629 , n1627 , n1628 );
xnor ( n1630 , n1629 , n1202 );
and ( n1631 , n1626 , n1630 );
and ( n1632 , n1582 , n1213 );
and ( n1633 , n1549 , n1211 );
nor ( n1634 , n1632 , n1633 );
xnor ( n1635 , n1634 , n1219 );
and ( n1636 , n1630 , n1635 );
and ( n1637 , n1626 , n1635 );
or ( n1638 , n1631 , n1636 , n1637 );
and ( n1639 , n1621 , n1638 );
and ( n1640 , n1619 , n1638 );
or ( n1641 , n1622 , n1639 , n1640 );
xor ( n1642 , n1586 , n1588 );
xor ( n1643 , n1642 , n1605 );
and ( n1644 , n1641 , n1643 );
buf ( n1645 , n1181 );
buf ( n1646 , n1645 );
buf ( n1647 , n1646 );
buf ( n1648 , n1647 );
and ( n1649 , n1648 , n1192 );
and ( n1650 , n1615 , n1190 );
nor ( n1651 , n1649 , n1650 );
not ( n1652 , n1651 );
xor ( n1653 , n1626 , n1630 );
xor ( n1654 , n1653 , n1635 );
and ( n1655 , n1652 , n1654 );
and ( n1656 , n1483 , n1304 );
and ( n1657 , n1450 , n1301 );
nor ( n1658 , n1656 , n1657 );
xnor ( n1659 , n1658 , n1199 );
and ( n1660 , n1549 , n1273 );
and ( n1661 , n1516 , n1271 );
nor ( n1662 , n1660 , n1661 );
xnor ( n1663 , n1662 , n1202 );
and ( n1664 , n1659 , n1663 );
and ( n1665 , n1615 , n1213 );
and ( n1666 , n1582 , n1211 );
nor ( n1667 , n1665 , n1666 );
xnor ( n1668 , n1667 , n1219 );
and ( n1669 , n1663 , n1668 );
and ( n1670 , n1659 , n1668 );
or ( n1671 , n1664 , n1669 , n1670 );
and ( n1672 , n1654 , n1671 );
and ( n1673 , n1652 , n1671 );
or ( n1674 , n1655 , n1672 , n1673 );
xor ( n1675 , n1619 , n1621 );
xor ( n1676 , n1675 , n1638 );
and ( n1677 , n1674 , n1676 );
buf ( n1678 , n1181 );
buf ( n1679 , n1678 );
buf ( n1680 , n1679 );
buf ( n1681 , n1680 );
and ( n1682 , n1681 , n1192 );
and ( n1683 , n1648 , n1190 );
nor ( n1684 , n1682 , n1683 );
not ( n1685 , n1684 );
xor ( n1686 , n1659 , n1663 );
xor ( n1687 , n1686 , n1668 );
and ( n1688 , n1685 , n1687 );
and ( n1689 , n1516 , n1304 );
and ( n1690 , n1483 , n1301 );
nor ( n1691 , n1689 , n1690 );
xnor ( n1692 , n1691 , n1199 );
and ( n1693 , n1582 , n1273 );
and ( n1694 , n1549 , n1271 );
nor ( n1695 , n1693 , n1694 );
xnor ( n1696 , n1695 , n1202 );
and ( n1697 , n1692 , n1696 );
and ( n1698 , n1648 , n1213 );
and ( n1699 , n1615 , n1211 );
nor ( n1700 , n1698 , n1699 );
xnor ( n1701 , n1700 , n1219 );
and ( n1702 , n1696 , n1701 );
and ( n1703 , n1692 , n1701 );
or ( n1704 , n1697 , n1702 , n1703 );
and ( n1705 , n1687 , n1704 );
and ( n1706 , n1685 , n1704 );
or ( n1707 , n1688 , n1705 , n1706 );
xor ( n1708 , n1652 , n1654 );
xor ( n1709 , n1708 , n1671 );
and ( n1710 , n1707 , n1709 );
buf ( n1711 , n1181 );
buf ( n1712 , n1711 );
buf ( n1713 , n1712 );
buf ( n1714 , n1713 );
and ( n1715 , n1714 , n1192 );
and ( n1716 , n1681 , n1190 );
nor ( n1717 , n1715 , n1716 );
not ( n1718 , n1717 );
xor ( n1719 , n1692 , n1696 );
xor ( n1720 , n1719 , n1701 );
and ( n1721 , n1718 , n1720 );
and ( n1722 , n1549 , n1304 );
and ( n1723 , n1516 , n1301 );
nor ( n1724 , n1722 , n1723 );
xnor ( n1725 , n1724 , n1199 );
and ( n1726 , n1615 , n1273 );
and ( n1727 , n1582 , n1271 );
nor ( n1728 , n1726 , n1727 );
xnor ( n1729 , n1728 , n1202 );
and ( n1730 , n1725 , n1729 );
and ( n1731 , n1681 , n1213 );
and ( n1732 , n1648 , n1211 );
nor ( n1733 , n1731 , n1732 );
xnor ( n1734 , n1733 , n1219 );
and ( n1735 , n1729 , n1734 );
and ( n1736 , n1725 , n1734 );
or ( n1737 , n1730 , n1735 , n1736 );
and ( n1738 , n1720 , n1737 );
and ( n1739 , n1718 , n1737 );
or ( n1740 , n1721 , n1738 , n1739 );
xor ( n1741 , n1685 , n1687 );
xor ( n1742 , n1741 , n1704 );
and ( n1743 , n1740 , n1742 );
buf ( n1744 , n1181 );
buf ( n1745 , n1744 );
buf ( n1746 , n1745 );
buf ( n1747 , n1746 );
and ( n1748 , n1747 , n1192 );
and ( n1749 , n1714 , n1190 );
nor ( n1750 , n1748 , n1749 );
not ( n1751 , n1750 );
xor ( n1752 , n1725 , n1729 );
xor ( n1753 , n1752 , n1734 );
and ( n1754 , n1751 , n1753 );
and ( n1755 , n1582 , n1304 );
and ( n1756 , n1549 , n1301 );
nor ( n1757 , n1755 , n1756 );
xnor ( n1758 , n1757 , n1199 );
and ( n1759 , n1648 , n1273 );
and ( n1760 , n1615 , n1271 );
nor ( n1761 , n1759 , n1760 );
xnor ( n1762 , n1761 , n1202 );
and ( n1763 , n1758 , n1762 );
and ( n1764 , n1714 , n1213 );
and ( n1765 , n1681 , n1211 );
nor ( n1766 , n1764 , n1765 );
xnor ( n1767 , n1766 , n1219 );
and ( n1768 , n1762 , n1767 );
and ( n1769 , n1758 , n1767 );
or ( n1770 , n1763 , n1768 , n1769 );
and ( n1771 , n1753 , n1770 );
and ( n1772 , n1751 , n1770 );
or ( n1773 , n1754 , n1771 , n1772 );
xor ( n1774 , n1718 , n1720 );
xor ( n1775 , n1774 , n1737 );
and ( n1776 , n1773 , n1775 );
buf ( n1777 , n1181 );
buf ( n1778 , n1777 );
buf ( n1779 , n1778 );
buf ( n1780 , n1779 );
and ( n1781 , n1780 , n1192 );
and ( n1782 , n1747 , n1190 );
nor ( n1783 , n1781 , n1782 );
not ( n1784 , n1783 );
xor ( n1785 , n1758 , n1762 );
xor ( n1786 , n1785 , n1767 );
and ( n1787 , n1784 , n1786 );
and ( n1788 , n1615 , n1304 );
and ( n1789 , n1582 , n1301 );
nor ( n1790 , n1788 , n1789 );
xnor ( n1791 , n1790 , n1199 );
and ( n1792 , n1681 , n1273 );
and ( n1793 , n1648 , n1271 );
nor ( n1794 , n1792 , n1793 );
xnor ( n1795 , n1794 , n1202 );
and ( n1796 , n1791 , n1795 );
and ( n1797 , n1747 , n1213 );
and ( n1798 , n1714 , n1211 );
nor ( n1799 , n1797 , n1798 );
xnor ( n1800 , n1799 , n1219 );
and ( n1801 , n1795 , n1800 );
and ( n1802 , n1791 , n1800 );
or ( n1803 , n1796 , n1801 , n1802 );
and ( n1804 , n1786 , n1803 );
and ( n1805 , n1784 , n1803 );
or ( n1806 , n1787 , n1804 , n1805 );
xor ( n1807 , n1751 , n1753 );
xor ( n1808 , n1807 , n1770 );
and ( n1809 , n1806 , n1808 );
buf ( n1810 , n1181 );
buf ( n1811 , n1810 );
buf ( n1812 , n1811 );
buf ( n1813 , n1812 );
and ( n1814 , n1813 , n1192 );
and ( n1815 , n1780 , n1190 );
nor ( n1816 , n1814 , n1815 );
not ( n1817 , n1816 );
xor ( n1818 , n1791 , n1795 );
xor ( n1819 , n1818 , n1800 );
and ( n1820 , n1817 , n1819 );
and ( n1821 , n1648 , n1304 );
and ( n1822 , n1615 , n1301 );
nor ( n1823 , n1821 , n1822 );
xnor ( n1824 , n1823 , n1199 );
and ( n1825 , n1714 , n1273 );
and ( n1826 , n1681 , n1271 );
nor ( n1827 , n1825 , n1826 );
xnor ( n1828 , n1827 , n1202 );
and ( n1829 , n1824 , n1828 );
and ( n1830 , n1780 , n1213 );
and ( n1831 , n1747 , n1211 );
nor ( n1832 , n1830 , n1831 );
xnor ( n1833 , n1832 , n1219 );
and ( n1834 , n1828 , n1833 );
and ( n1835 , n1824 , n1833 );
or ( n1836 , n1829 , n1834 , n1835 );
and ( n1837 , n1819 , n1836 );
and ( n1838 , n1817 , n1836 );
or ( n1839 , n1820 , n1837 , n1838 );
xor ( n1840 , n1784 , n1786 );
xor ( n1841 , n1840 , n1803 );
and ( n1842 , n1839 , n1841 );
buf ( n1843 , n1181 );
buf ( n1844 , n1843 );
buf ( n1845 , n1844 );
buf ( n1846 , n1845 );
and ( n1847 , n1846 , n1192 );
and ( n1848 , n1813 , n1190 );
nor ( n1849 , n1847 , n1848 );
not ( n1850 , n1849 );
xor ( n1851 , n1824 , n1828 );
xor ( n1852 , n1851 , n1833 );
and ( n1853 , n1850 , n1852 );
and ( n1854 , n1681 , n1304 );
and ( n1855 , n1648 , n1301 );
nor ( n1856 , n1854 , n1855 );
xnor ( n1857 , n1856 , n1199 );
and ( n1858 , n1747 , n1273 );
and ( n1859 , n1714 , n1271 );
nor ( n1860 , n1858 , n1859 );
xnor ( n1861 , n1860 , n1202 );
and ( n1862 , n1857 , n1861 );
and ( n1863 , n1813 , n1213 );
and ( n1864 , n1780 , n1211 );
nor ( n1865 , n1863 , n1864 );
xnor ( n1866 , n1865 , n1219 );
and ( n1867 , n1861 , n1866 );
and ( n1868 , n1857 , n1866 );
or ( n1869 , n1862 , n1867 , n1868 );
and ( n1870 , n1852 , n1869 );
and ( n1871 , n1850 , n1869 );
or ( n1872 , n1853 , n1870 , n1871 );
xor ( n1873 , n1817 , n1819 );
xor ( n1874 , n1873 , n1836 );
and ( n1875 , n1872 , n1874 );
buf ( n1876 , n1181 );
buf ( n1877 , n1876 );
buf ( n1878 , n1877 );
buf ( n1879 , n1878 );
and ( n1880 , n1879 , n1192 );
and ( n1881 , n1846 , n1190 );
nor ( n1882 , n1880 , n1881 );
not ( n1883 , n1882 );
xor ( n1884 , n1857 , n1861 );
xor ( n1885 , n1884 , n1866 );
and ( n1886 , n1883 , n1885 );
and ( n1887 , n1714 , n1304 );
and ( n1888 , n1681 , n1301 );
nor ( n1889 , n1887 , n1888 );
xnor ( n1890 , n1889 , n1199 );
and ( n1891 , n1780 , n1273 );
and ( n1892 , n1747 , n1271 );
nor ( n1893 , n1891 , n1892 );
xnor ( n1894 , n1893 , n1202 );
and ( n1895 , n1890 , n1894 );
and ( n1896 , n1846 , n1213 );
and ( n1897 , n1813 , n1211 );
nor ( n1898 , n1896 , n1897 );
xnor ( n1899 , n1898 , n1219 );
and ( n1900 , n1894 , n1899 );
and ( n1901 , n1890 , n1899 );
or ( n1902 , n1895 , n1900 , n1901 );
and ( n1903 , n1885 , n1902 );
and ( n1904 , n1883 , n1902 );
or ( n1905 , n1886 , n1903 , n1904 );
xor ( n1906 , n1850 , n1852 );
xor ( n1907 , n1906 , n1869 );
and ( n1908 , n1905 , n1907 );
buf ( n1909 , n1181 );
buf ( n1910 , n1909 );
buf ( n1911 , n1910 );
buf ( n1912 , n1911 );
and ( n1913 , n1912 , n1192 );
and ( n1914 , n1879 , n1190 );
nor ( n1915 , n1913 , n1914 );
not ( n1916 , n1915 );
xor ( n1917 , n1890 , n1894 );
xor ( n1918 , n1917 , n1899 );
and ( n1919 , n1916 , n1918 );
and ( n1920 , n1747 , n1304 );
and ( n1921 , n1714 , n1301 );
nor ( n1922 , n1920 , n1921 );
xnor ( n1923 , n1922 , n1199 );
and ( n1924 , n1813 , n1273 );
and ( n1925 , n1780 , n1271 );
nor ( n1926 , n1924 , n1925 );
xnor ( n1927 , n1926 , n1202 );
and ( n1928 , n1923 , n1927 );
and ( n1929 , n1879 , n1213 );
and ( n1930 , n1846 , n1211 );
nor ( n1931 , n1929 , n1930 );
xnor ( n1932 , n1931 , n1219 );
and ( n1933 , n1927 , n1932 );
and ( n1934 , n1923 , n1932 );
or ( n1935 , n1928 , n1933 , n1934 );
and ( n1936 , n1918 , n1935 );
and ( n1937 , n1916 , n1935 );
or ( n1938 , n1919 , n1936 , n1937 );
xor ( n1939 , n1883 , n1885 );
xor ( n1940 , n1939 , n1902 );
and ( n1941 , n1938 , n1940 );
buf ( n1942 , n1181 );
buf ( n1943 , n1942 );
buf ( n1944 , n1943 );
buf ( n1945 , n1944 );
and ( n1946 , n1945 , n1192 );
and ( n1947 , n1912 , n1190 );
nor ( n1948 , n1946 , n1947 );
not ( n1949 , n1948 );
xor ( n1950 , n1923 , n1927 );
xor ( n1951 , n1950 , n1932 );
and ( n1952 , n1949 , n1951 );
and ( n1953 , n1780 , n1304 );
and ( n1954 , n1747 , n1301 );
nor ( n1955 , n1953 , n1954 );
xnor ( n1956 , n1955 , n1199 );
and ( n1957 , n1846 , n1273 );
and ( n1958 , n1813 , n1271 );
nor ( n1959 , n1957 , n1958 );
xnor ( n1960 , n1959 , n1202 );
and ( n1961 , n1956 , n1960 );
and ( n1962 , n1912 , n1213 );
and ( n1963 , n1879 , n1211 );
nor ( n1964 , n1962 , n1963 );
xnor ( n1965 , n1964 , n1219 );
and ( n1966 , n1960 , n1965 );
and ( n1967 , n1956 , n1965 );
or ( n1968 , n1961 , n1966 , n1967 );
and ( n1969 , n1951 , n1968 );
and ( n1970 , n1949 , n1968 );
or ( n1971 , n1952 , n1969 , n1970 );
xor ( n1972 , n1916 , n1918 );
xor ( n1973 , n1972 , n1935 );
and ( n1974 , n1971 , n1973 );
buf ( n1975 , n1181 );
buf ( n1976 , n1975 );
buf ( n1977 , n1976 );
buf ( n1978 , n1977 );
and ( n1979 , n1978 , n1192 );
and ( n1980 , n1945 , n1190 );
nor ( n1981 , n1979 , n1980 );
not ( n1982 , n1981 );
xor ( n1983 , n1956 , n1960 );
xor ( n1984 , n1983 , n1965 );
and ( n1985 , n1982 , n1984 );
and ( n1986 , n1813 , n1304 );
and ( n1987 , n1780 , n1301 );
nor ( n1988 , n1986 , n1987 );
xnor ( n1989 , n1988 , n1199 );
and ( n1990 , n1879 , n1273 );
and ( n1991 , n1846 , n1271 );
nor ( n1992 , n1990 , n1991 );
xnor ( n1993 , n1992 , n1202 );
and ( n1994 , n1989 , n1993 );
and ( n1995 , n1945 , n1213 );
and ( n1996 , n1912 , n1211 );
nor ( n1997 , n1995 , n1996 );
xnor ( n1998 , n1997 , n1219 );
and ( n1999 , n1993 , n1998 );
and ( n2000 , n1989 , n1998 );
or ( n2001 , n1994 , n1999 , n2000 );
and ( n2002 , n1984 , n2001 );
and ( n2003 , n1982 , n2001 );
or ( n2004 , n1985 , n2002 , n2003 );
xor ( n2005 , n1949 , n1951 );
xor ( n2006 , n2005 , n1968 );
and ( n2007 , n2004 , n2006 );
buf ( n2008 , n1181 );
buf ( n2009 , n2008 );
buf ( n2010 , n2009 );
buf ( n2011 , n2010 );
and ( n2012 , n2011 , n1192 );
and ( n2013 , n1978 , n1190 );
nor ( n2014 , n2012 , n2013 );
not ( n2015 , n2014 );
xor ( n2016 , n1989 , n1993 );
xor ( n2017 , n2016 , n1998 );
and ( n2018 , n2015 , n2017 );
and ( n2019 , n1846 , n1304 );
and ( n2020 , n1813 , n1301 );
nor ( n2021 , n2019 , n2020 );
xnor ( n2022 , n2021 , n1199 );
and ( n2023 , n1912 , n1273 );
and ( n2024 , n1879 , n1271 );
nor ( n2025 , n2023 , n2024 );
xnor ( n2026 , n2025 , n1202 );
and ( n2027 , n2022 , n2026 );
and ( n2028 , n1978 , n1213 );
and ( n2029 , n1945 , n1211 );
nor ( n2030 , n2028 , n2029 );
xnor ( n2031 , n2030 , n1219 );
and ( n2032 , n2026 , n2031 );
and ( n2033 , n2022 , n2031 );
or ( n2034 , n2027 , n2032 , n2033 );
and ( n2035 , n2017 , n2034 );
and ( n2036 , n2015 , n2034 );
or ( n2037 , n2018 , n2035 , n2036 );
xor ( n2038 , n1982 , n1984 );
xor ( n2039 , n2038 , n2001 );
and ( n2040 , n2037 , n2039 );
buf ( n2041 , n1181 );
buf ( n2042 , n2041 );
buf ( n2043 , n2042 );
buf ( n2044 , n2043 );
and ( n2045 , n2044 , n1192 );
and ( n2046 , n2011 , n1190 );
nor ( n2047 , n2045 , n2046 );
not ( n2048 , n2047 );
xor ( n2049 , n2022 , n2026 );
xor ( n2050 , n2049 , n2031 );
and ( n2051 , n2048 , n2050 );
and ( n2052 , n1879 , n1304 );
and ( n2053 , n1846 , n1301 );
nor ( n2054 , n2052 , n2053 );
xnor ( n2055 , n2054 , n1199 );
and ( n2056 , n1945 , n1273 );
and ( n2057 , n1912 , n1271 );
nor ( n2058 , n2056 , n2057 );
xnor ( n2059 , n2058 , n1202 );
and ( n2060 , n2055 , n2059 );
and ( n2061 , n2011 , n1213 );
and ( n2062 , n1978 , n1211 );
nor ( n2063 , n2061 , n2062 );
xnor ( n2064 , n2063 , n1219 );
and ( n2065 , n2059 , n2064 );
and ( n2066 , n2055 , n2064 );
or ( n2067 , n2060 , n2065 , n2066 );
and ( n2068 , n2050 , n2067 );
and ( n2069 , n2048 , n2067 );
or ( n2070 , n2051 , n2068 , n2069 );
xor ( n2071 , n2015 , n2017 );
xor ( n2072 , n2071 , n2034 );
and ( n2073 , n2070 , n2072 );
buf ( n2074 , n1181 );
buf ( n2075 , n2074 );
buf ( n2076 , n2075 );
buf ( n2077 , n2076 );
and ( n2078 , n2077 , n1192 );
and ( n2079 , n2044 , n1190 );
nor ( n2080 , n2078 , n2079 );
not ( n2081 , n2080 );
xor ( n2082 , n2055 , n2059 );
xor ( n2083 , n2082 , n2064 );
and ( n2084 , n2081 , n2083 );
and ( n2085 , n1912 , n1304 );
and ( n2086 , n1879 , n1301 );
nor ( n2087 , n2085 , n2086 );
xnor ( n2088 , n2087 , n1199 );
and ( n2089 , n1978 , n1273 );
and ( n2090 , n1945 , n1271 );
nor ( n2091 , n2089 , n2090 );
xnor ( n2092 , n2091 , n1202 );
and ( n2093 , n2088 , n2092 );
and ( n2094 , n2044 , n1213 );
and ( n2095 , n2011 , n1211 );
nor ( n2096 , n2094 , n2095 );
xnor ( n2097 , n2096 , n1219 );
and ( n2098 , n2092 , n2097 );
and ( n2099 , n2088 , n2097 );
or ( n2100 , n2093 , n2098 , n2099 );
and ( n2101 , n2083 , n2100 );
and ( n2102 , n2081 , n2100 );
or ( n2103 , n2084 , n2101 , n2102 );
xor ( n2104 , n2048 , n2050 );
xor ( n2105 , n2104 , n2067 );
and ( n2106 , n2103 , n2105 );
buf ( n2107 , n1181 );
buf ( n2108 , n2107 );
buf ( n2109 , n2108 );
buf ( n2110 , n2109 );
and ( n2111 , n2110 , n1192 );
and ( n2112 , n2077 , n1190 );
nor ( n2113 , n2111 , n2112 );
not ( n2114 , n2113 );
xor ( n2115 , n2088 , n2092 );
xor ( n2116 , n2115 , n2097 );
and ( n2117 , n2114 , n2116 );
and ( n2118 , n1945 , n1304 );
and ( n2119 , n1912 , n1301 );
nor ( n2120 , n2118 , n2119 );
xnor ( n2121 , n2120 , n1199 );
and ( n2122 , n2011 , n1273 );
and ( n2123 , n1978 , n1271 );
nor ( n2124 , n2122 , n2123 );
xnor ( n2125 , n2124 , n1202 );
and ( n2126 , n2121 , n2125 );
and ( n2127 , n2077 , n1213 );
and ( n2128 , n2044 , n1211 );
nor ( n2129 , n2127 , n2128 );
xnor ( n2130 , n2129 , n1219 );
and ( n2131 , n2125 , n2130 );
and ( n2132 , n2121 , n2130 );
or ( n2133 , n2126 , n2131 , n2132 );
and ( n2134 , n2116 , n2133 );
and ( n2135 , n2114 , n2133 );
or ( n2136 , n2117 , n2134 , n2135 );
xor ( n2137 , n2081 , n2083 );
xor ( n2138 , n2137 , n2100 );
and ( n2139 , n2136 , n2138 );
buf ( n2140 , n1181 );
buf ( n2141 , n2140 );
buf ( n2142 , n2141 );
buf ( n2143 , n2142 );
and ( n2144 , n2143 , n1192 );
and ( n2145 , n2110 , n1190 );
nor ( n2146 , n2144 , n2145 );
not ( n2147 , n2146 );
xor ( n2148 , n2121 , n2125 );
xor ( n2149 , n2148 , n2130 );
and ( n2150 , n2147 , n2149 );
and ( n2151 , n1978 , n1304 );
and ( n2152 , n1945 , n1301 );
nor ( n2153 , n2151 , n2152 );
xnor ( n2154 , n2153 , n1199 );
and ( n2155 , n2044 , n1273 );
and ( n2156 , n2011 , n1271 );
nor ( n2157 , n2155 , n2156 );
xnor ( n2158 , n2157 , n1202 );
and ( n2159 , n2154 , n2158 );
and ( n2160 , n2110 , n1213 );
and ( n2161 , n2077 , n1211 );
nor ( n2162 , n2160 , n2161 );
xnor ( n2163 , n2162 , n1219 );
and ( n2164 , n2158 , n2163 );
and ( n2165 , n2154 , n2163 );
or ( n2166 , n2159 , n2164 , n2165 );
and ( n2167 , n2149 , n2166 );
and ( n2168 , n2147 , n2166 );
or ( n2169 , n2150 , n2167 , n2168 );
xor ( n2170 , n2114 , n2116 );
xor ( n2171 , n2170 , n2133 );
and ( n2172 , n2169 , n2171 );
buf ( n2173 , n1181 );
buf ( n2174 , n2173 );
buf ( n2175 , n2174 );
buf ( n2176 , n2175 );
and ( n2177 , n2176 , n1192 );
and ( n2178 , n2143 , n1190 );
nor ( n2179 , n2177 , n2178 );
not ( n2180 , n2179 );
xor ( n2181 , n2154 , n2158 );
xor ( n2182 , n2181 , n2163 );
and ( n2183 , n2180 , n2182 );
and ( n2184 , n2011 , n1304 );
and ( n2185 , n1978 , n1301 );
nor ( n2186 , n2184 , n2185 );
xnor ( n2187 , n2186 , n1199 );
and ( n2188 , n2077 , n1273 );
and ( n2189 , n2044 , n1271 );
nor ( n2190 , n2188 , n2189 );
xnor ( n2191 , n2190 , n1202 );
and ( n2192 , n2187 , n2191 );
and ( n2193 , n2143 , n1213 );
and ( n2194 , n2110 , n1211 );
nor ( n2195 , n2193 , n2194 );
xnor ( n2196 , n2195 , n1219 );
and ( n2197 , n2191 , n2196 );
and ( n2198 , n2187 , n2196 );
or ( n2199 , n2192 , n2197 , n2198 );
and ( n2200 , n2182 , n2199 );
and ( n2201 , n2180 , n2199 );
or ( n2202 , n2183 , n2200 , n2201 );
xor ( n2203 , n2147 , n2149 );
xor ( n2204 , n2203 , n2166 );
and ( n2205 , n2202 , n2204 );
buf ( n2206 , n1181 );
buf ( n2207 , n2206 );
buf ( n2208 , n2207 );
buf ( n2209 , n2208 );
and ( n2210 , n2209 , n1192 );
and ( n2211 , n2176 , n1190 );
nor ( n2212 , n2210 , n2211 );
not ( n2213 , n2212 );
xor ( n2214 , n2187 , n2191 );
xor ( n2215 , n2214 , n2196 );
and ( n2216 , n2213 , n2215 );
and ( n2217 , n2044 , n1304 );
and ( n2218 , n2011 , n1301 );
nor ( n2219 , n2217 , n2218 );
xnor ( n2220 , n2219 , n1199 );
and ( n2221 , n2110 , n1273 );
and ( n2222 , n2077 , n1271 );
nor ( n2223 , n2221 , n2222 );
xnor ( n2224 , n2223 , n1202 );
and ( n2225 , n2220 , n2224 );
and ( n2226 , n2176 , n1213 );
and ( n2227 , n2143 , n1211 );
nor ( n2228 , n2226 , n2227 );
xnor ( n2229 , n2228 , n1219 );
and ( n2230 , n2224 , n2229 );
and ( n2231 , n2220 , n2229 );
or ( n2232 , n2225 , n2230 , n2231 );
and ( n2233 , n2215 , n2232 );
and ( n2234 , n2213 , n2232 );
or ( n2235 , n2216 , n2233 , n2234 );
xor ( n2236 , n2180 , n2182 );
xor ( n2237 , n2236 , n2199 );
and ( n2238 , n2235 , n2237 );
buf ( n2239 , n1181 );
buf ( n2240 , n2239 );
buf ( n2241 , n2240 );
buf ( n2242 , n2241 );
and ( n2243 , n2242 , n1192 );
and ( n2244 , n2209 , n1190 );
nor ( n2245 , n2243 , n2244 );
not ( n2246 , n2245 );
xor ( n2247 , n2220 , n2224 );
xor ( n2248 , n2247 , n2229 );
and ( n2249 , n2246 , n2248 );
and ( n2250 , n2077 , n1304 );
and ( n2251 , n2044 , n1301 );
nor ( n2252 , n2250 , n2251 );
xnor ( n2253 , n2252 , n1199 );
and ( n2254 , n2143 , n1273 );
and ( n2255 , n2110 , n1271 );
nor ( n2256 , n2254 , n2255 );
xnor ( n2257 , n2256 , n1202 );
and ( n2258 , n2253 , n2257 );
and ( n2259 , n2209 , n1213 );
and ( n2260 , n2176 , n1211 );
nor ( n2261 , n2259 , n2260 );
xnor ( n2262 , n2261 , n1219 );
and ( n2263 , n2257 , n2262 );
and ( n2264 , n2253 , n2262 );
or ( n2265 , n2258 , n2263 , n2264 );
and ( n2266 , n2248 , n2265 );
and ( n2267 , n2246 , n2265 );
or ( n2268 , n2249 , n2266 , n2267 );
xor ( n2269 , n2213 , n2215 );
xor ( n2270 , n2269 , n2232 );
and ( n2271 , n2268 , n2270 );
buf ( n2272 , n1181 );
buf ( n2273 , n2272 );
buf ( n2274 , n2273 );
buf ( n2275 , n2274 );
and ( n2276 , n2275 , n1192 );
and ( n2277 , n2242 , n1190 );
nor ( n2278 , n2276 , n2277 );
not ( n2279 , n2278 );
xor ( n2280 , n2253 , n2257 );
xor ( n2281 , n2280 , n2262 );
and ( n2282 , n2279 , n2281 );
and ( n2283 , n2110 , n1304 );
and ( n2284 , n2077 , n1301 );
nor ( n2285 , n2283 , n2284 );
xnor ( n2286 , n2285 , n1199 );
and ( n2287 , n2176 , n1273 );
and ( n2288 , n2143 , n1271 );
nor ( n2289 , n2287 , n2288 );
xnor ( n2290 , n2289 , n1202 );
and ( n2291 , n2286 , n2290 );
and ( n2292 , n2242 , n1213 );
and ( n2293 , n2209 , n1211 );
nor ( n2294 , n2292 , n2293 );
xnor ( n2295 , n2294 , n1219 );
and ( n2296 , n2290 , n2295 );
and ( n2297 , n2286 , n2295 );
or ( n2298 , n2291 , n2296 , n2297 );
and ( n2299 , n2281 , n2298 );
and ( n2300 , n2279 , n2298 );
or ( n2301 , n2282 , n2299 , n2300 );
xor ( n2302 , n2246 , n2248 );
xor ( n2303 , n2302 , n2265 );
and ( n2304 , n2301 , n2303 );
buf ( n2305 , n1181 );
buf ( n2306 , n2305 );
buf ( n2307 , n2306 );
buf ( n2308 , n2307 );
and ( n2309 , n2308 , n1192 );
and ( n2310 , n2275 , n1190 );
nor ( n2311 , n2309 , n2310 );
not ( n2312 , n2311 );
xor ( n2313 , n2286 , n2290 );
xor ( n2314 , n2313 , n2295 );
and ( n2315 , n2312 , n2314 );
and ( n2316 , n2143 , n1304 );
and ( n2317 , n2110 , n1301 );
nor ( n2318 , n2316 , n2317 );
xnor ( n2319 , n2318 , n1199 );
and ( n2320 , n2209 , n1273 );
and ( n2321 , n2176 , n1271 );
nor ( n2322 , n2320 , n2321 );
xnor ( n2323 , n2322 , n1202 );
and ( n2324 , n2319 , n2323 );
and ( n2325 , n2275 , n1213 );
and ( n2326 , n2242 , n1211 );
nor ( n2327 , n2325 , n2326 );
xnor ( n2328 , n2327 , n1219 );
and ( n2329 , n2323 , n2328 );
and ( n2330 , n2319 , n2328 );
or ( n2331 , n2324 , n2329 , n2330 );
and ( n2332 , n2314 , n2331 );
and ( n2333 , n2312 , n2331 );
or ( n2334 , n2315 , n2332 , n2333 );
xor ( n2335 , n2279 , n2281 );
xor ( n2336 , n2335 , n2298 );
and ( n2337 , n2334 , n2336 );
buf ( n2338 , n1181 );
buf ( n2339 , n2338 );
buf ( n2340 , n2339 );
buf ( n2341 , n2340 );
and ( n2342 , n2341 , n1192 );
and ( n2343 , n2308 , n1190 );
nor ( n2344 , n2342 , n2343 );
not ( n2345 , n2344 );
xor ( n2346 , n2319 , n2323 );
xor ( n2347 , n2346 , n2328 );
and ( n2348 , n2345 , n2347 );
and ( n2349 , n2176 , n1304 );
and ( n2350 , n2143 , n1301 );
nor ( n2351 , n2349 , n2350 );
xnor ( n2352 , n2351 , n1199 );
and ( n2353 , n2242 , n1273 );
and ( n2354 , n2209 , n1271 );
nor ( n2355 , n2353 , n2354 );
xnor ( n2356 , n2355 , n1202 );
and ( n2357 , n2352 , n2356 );
and ( n2358 , n2308 , n1213 );
and ( n2359 , n2275 , n1211 );
nor ( n2360 , n2358 , n2359 );
xnor ( n2361 , n2360 , n1219 );
and ( n2362 , n2356 , n2361 );
and ( n2363 , n2352 , n2361 );
or ( n2364 , n2357 , n2362 , n2363 );
and ( n2365 , n2347 , n2364 );
and ( n2366 , n2345 , n2364 );
or ( n2367 , n2348 , n2365 , n2366 );
xor ( n2368 , n2312 , n2314 );
xor ( n2369 , n2368 , n2331 );
and ( n2370 , n2367 , n2369 );
buf ( n2371 , n1181 );
buf ( n2372 , n2371 );
buf ( n2373 , n2372 );
buf ( n2374 , n2373 );
and ( n2375 , n2374 , n1192 );
and ( n2376 , n2341 , n1190 );
nor ( n2377 , n2375 , n2376 );
not ( n2378 , n2377 );
xor ( n2379 , n2352 , n2356 );
xor ( n2380 , n2379 , n2361 );
and ( n2381 , n2378 , n2380 );
and ( n2382 , n2209 , n1304 );
and ( n2383 , n2176 , n1301 );
nor ( n2384 , n2382 , n2383 );
xnor ( n2385 , n2384 , n1199 );
and ( n2386 , n2275 , n1273 );
and ( n2387 , n2242 , n1271 );
nor ( n2388 , n2386 , n2387 );
xnor ( n2389 , n2388 , n1202 );
and ( n2390 , n2385 , n2389 );
and ( n2391 , n2341 , n1213 );
and ( n2392 , n2308 , n1211 );
nor ( n2393 , n2391 , n2392 );
xnor ( n2394 , n2393 , n1219 );
and ( n2395 , n2389 , n2394 );
and ( n2396 , n2385 , n2394 );
or ( n2397 , n2390 , n2395 , n2396 );
and ( n2398 , n2380 , n2397 );
and ( n2399 , n2378 , n2397 );
or ( n2400 , n2381 , n2398 , n2399 );
xor ( n2401 , n2345 , n2347 );
xor ( n2402 , n2401 , n2364 );
and ( n2403 , n2400 , n2402 );
buf ( n2404 , n1181 );
buf ( n2405 , n2404 );
buf ( n2406 , n2405 );
buf ( n2407 , n2406 );
and ( n2408 , n2407 , n1192 );
and ( n2409 , n2374 , n1190 );
nor ( n2410 , n2408 , n2409 );
not ( n2411 , n2410 );
xor ( n2412 , n2385 , n2389 );
xor ( n2413 , n2412 , n2394 );
and ( n2414 , n2411 , n2413 );
and ( n2415 , n2242 , n1304 );
and ( n2416 , n2209 , n1301 );
nor ( n2417 , n2415 , n2416 );
xnor ( n2418 , n2417 , n1199 );
and ( n2419 , n2308 , n1273 );
and ( n2420 , n2275 , n1271 );
nor ( n2421 , n2419 , n2420 );
xnor ( n2422 , n2421 , n1202 );
and ( n2423 , n2418 , n2422 );
and ( n2424 , n2374 , n1213 );
and ( n2425 , n2341 , n1211 );
nor ( n2426 , n2424 , n2425 );
xnor ( n2427 , n2426 , n1219 );
and ( n2428 , n2422 , n2427 );
and ( n2429 , n2418 , n2427 );
or ( n2430 , n2423 , n2428 , n2429 );
and ( n2431 , n2413 , n2430 );
and ( n2432 , n2411 , n2430 );
or ( n2433 , n2414 , n2431 , n2432 );
xor ( n2434 , n2378 , n2380 );
xor ( n2435 , n2434 , n2397 );
and ( n2436 , n2433 , n2435 );
buf ( n2437 , n1181 );
buf ( n2438 , n2437 );
buf ( n2439 , n2438 );
buf ( n2440 , n2439 );
and ( n2441 , n2440 , n1192 );
and ( n2442 , n2407 , n1190 );
nor ( n2443 , n2441 , n2442 );
not ( n2444 , n2443 );
xor ( n2445 , n2418 , n2422 );
xor ( n2446 , n2445 , n2427 );
and ( n2447 , n2444 , n2446 );
and ( n2448 , n2275 , n1304 );
and ( n2449 , n2242 , n1301 );
nor ( n2450 , n2448 , n2449 );
xnor ( n2451 , n2450 , n1199 );
and ( n2452 , n2341 , n1273 );
and ( n2453 , n2308 , n1271 );
nor ( n2454 , n2452 , n2453 );
xnor ( n2455 , n2454 , n1202 );
and ( n2456 , n2451 , n2455 );
and ( n2457 , n2407 , n1213 );
and ( n2458 , n2374 , n1211 );
nor ( n2459 , n2457 , n2458 );
xnor ( n2460 , n2459 , n1219 );
and ( n2461 , n2455 , n2460 );
and ( n2462 , n2451 , n2460 );
or ( n2463 , n2456 , n2461 , n2462 );
and ( n2464 , n2446 , n2463 );
and ( n2465 , n2444 , n2463 );
or ( n2466 , n2447 , n2464 , n2465 );
xor ( n2467 , n2411 , n2413 );
xor ( n2468 , n2467 , n2430 );
and ( n2469 , n2466 , n2468 );
buf ( n2470 , n1181 );
buf ( n2471 , n2470 );
buf ( n2472 , n2471 );
buf ( n2473 , n2472 );
and ( n2474 , n2473 , n1192 );
and ( n2475 , n2440 , n1190 );
nor ( n2476 , n2474 , n2475 );
not ( n2477 , n2476 );
xor ( n2478 , n2451 , n2455 );
xor ( n2479 , n2478 , n2460 );
and ( n2480 , n2477 , n2479 );
and ( n2481 , n2308 , n1304 );
and ( n2482 , n2275 , n1301 );
nor ( n2483 , n2481 , n2482 );
xnor ( n2484 , n2483 , n1199 );
and ( n2485 , n2374 , n1273 );
and ( n2486 , n2341 , n1271 );
nor ( n2487 , n2485 , n2486 );
xnor ( n2488 , n2487 , n1202 );
and ( n2489 , n2484 , n2488 );
and ( n2490 , n2440 , n1213 );
and ( n2491 , n2407 , n1211 );
nor ( n2492 , n2490 , n2491 );
xnor ( n2493 , n2492 , n1219 );
and ( n2494 , n2488 , n2493 );
and ( n2495 , n2484 , n2493 );
or ( n2496 , n2489 , n2494 , n2495 );
and ( n2497 , n2479 , n2496 );
and ( n2498 , n2477 , n2496 );
or ( n2499 , n2480 , n2497 , n2498 );
xor ( n2500 , n2444 , n2446 );
xor ( n2501 , n2500 , n2463 );
and ( n2502 , n2499 , n2501 );
buf ( n2503 , n1181 );
buf ( n2504 , n2503 );
buf ( n2505 , n2504 );
buf ( n2506 , n2505 );
and ( n2507 , n2506 , n1192 );
and ( n2508 , n2473 , n1190 );
nor ( n2509 , n2507 , n2508 );
not ( n2510 , n2509 );
xor ( n2511 , n2484 , n2488 );
xor ( n2512 , n2511 , n2493 );
and ( n2513 , n2510 , n2512 );
and ( n2514 , n2341 , n1304 );
and ( n2515 , n2308 , n1301 );
nor ( n2516 , n2514 , n2515 );
xnor ( n2517 , n2516 , n1199 );
and ( n2518 , n2407 , n1273 );
and ( n2519 , n2374 , n1271 );
nor ( n2520 , n2518 , n2519 );
xnor ( n2521 , n2520 , n1202 );
and ( n2522 , n2517 , n2521 );
and ( n2523 , n2473 , n1213 );
and ( n2524 , n2440 , n1211 );
nor ( n2525 , n2523 , n2524 );
xnor ( n2526 , n2525 , n1219 );
and ( n2527 , n2521 , n2526 );
and ( n2528 , n2517 , n2526 );
or ( n2529 , n2522 , n2527 , n2528 );
and ( n2530 , n2512 , n2529 );
and ( n2531 , n2510 , n2529 );
or ( n2532 , n2513 , n2530 , n2531 );
xor ( n2533 , n2477 , n2479 );
xor ( n2534 , n2533 , n2496 );
and ( n2535 , n2532 , n2534 );
buf ( n2536 , n1181 );
buf ( n2537 , n2536 );
buf ( n2538 , n2537 );
buf ( n2539 , n2538 );
and ( n2540 , n2539 , n1192 );
and ( n2541 , n2506 , n1190 );
nor ( n2542 , n2540 , n2541 );
not ( n2543 , n2542 );
xor ( n2544 , n2517 , n2521 );
xor ( n2545 , n2544 , n2526 );
and ( n2546 , n2543 , n2545 );
and ( n2547 , n2374 , n1304 );
and ( n2548 , n2341 , n1301 );
nor ( n2549 , n2547 , n2548 );
xnor ( n2550 , n2549 , n1199 );
and ( n2551 , n2440 , n1273 );
and ( n2552 , n2407 , n1271 );
nor ( n2553 , n2551 , n2552 );
xnor ( n2554 , n2553 , n1202 );
and ( n2555 , n2550 , n2554 );
and ( n2556 , n2506 , n1213 );
and ( n2557 , n2473 , n1211 );
nor ( n2558 , n2556 , n2557 );
xnor ( n2559 , n2558 , n1219 );
and ( n2560 , n2554 , n2559 );
and ( n2561 , n2550 , n2559 );
or ( n2562 , n2555 , n2560 , n2561 );
and ( n2563 , n2545 , n2562 );
and ( n2564 , n2543 , n2562 );
or ( n2565 , n2546 , n2563 , n2564 );
xor ( n2566 , n2510 , n2512 );
xor ( n2567 , n2566 , n2529 );
and ( n2568 , n2565 , n2567 );
buf ( n2569 , n1181 );
buf ( n2570 , n2569 );
buf ( n2571 , n2570 );
and ( n2572 , n2571 , n1192 );
and ( n2573 , n2539 , n1190 );
nor ( n2574 , n2572 , n2573 );
not ( n2575 , n2574 );
xor ( n2576 , n2550 , n2554 );
xor ( n2577 , n2576 , n2559 );
and ( n2578 , n2575 , n2577 );
and ( n2579 , n2407 , n1304 );
and ( n2580 , n2374 , n1301 );
nor ( n2581 , n2579 , n2580 );
xnor ( n2582 , n2581 , n1199 );
and ( n2583 , n2473 , n1273 );
and ( n2584 , n2440 , n1271 );
nor ( n2585 , n2583 , n2584 );
xnor ( n2586 , n2585 , n1202 );
and ( n2587 , n2582 , n2586 );
and ( n2588 , n2539 , n1213 );
and ( n2589 , n2506 , n1211 );
nor ( n2590 , n2588 , n2589 );
xnor ( n2591 , n2590 , n1219 );
and ( n2592 , n2586 , n2591 );
and ( n2593 , n2582 , n2591 );
or ( n2594 , n2587 , n2592 , n2593 );
and ( n2595 , n2577 , n2594 );
and ( n2596 , n2575 , n2594 );
or ( n2597 , n2578 , n2595 , n2596 );
xor ( n2598 , n2543 , n2545 );
xor ( n2599 , n2598 , n2562 );
and ( n2600 , n2597 , n2599 );
xor ( n2601 , n760 , n1178 );
buf ( n2602 , n2601 );
buf ( n2603 , n2602 );
buf ( n2604 , n2603 );
and ( n2605 , n2604 , n1192 );
and ( n2606 , n2571 , n1190 );
nor ( n2607 , n2605 , n2606 );
not ( n2608 , n2607 );
xor ( n2609 , n2582 , n2586 );
xor ( n2610 , n2609 , n2591 );
and ( n2611 , n2608 , n2610 );
and ( n2612 , n2440 , n1304 );
and ( n2613 , n2407 , n1301 );
nor ( n2614 , n2612 , n2613 );
xnor ( n2615 , n2614 , n1199 );
and ( n2616 , n2506 , n1273 );
and ( n2617 , n2473 , n1271 );
nor ( n2618 , n2616 , n2617 );
xnor ( n2619 , n2618 , n1202 );
and ( n2620 , n2615 , n2619 );
and ( n2621 , n2571 , n1213 );
and ( n2622 , n2539 , n1211 );
nor ( n2623 , n2621 , n2622 );
xnor ( n2624 , n2623 , n1219 );
and ( n2625 , n2619 , n2624 );
and ( n2626 , n2615 , n2624 );
or ( n2627 , n2620 , n2625 , n2626 );
and ( n2628 , n2610 , n2627 );
and ( n2629 , n2608 , n2627 );
or ( n2630 , n2611 , n2628 , n2629 );
xor ( n2631 , n2575 , n2577 );
xor ( n2632 , n2631 , n2594 );
and ( n2633 , n2630 , n2632 );
xor ( n2634 , n762 , n1176 );
buf ( n2635 , n2634 );
buf ( n2636 , n2635 );
buf ( n2637 , n2636 );
and ( n2638 , n2637 , n1192 );
and ( n2639 , n2604 , n1190 );
nor ( n2640 , n2638 , n2639 );
not ( n2641 , n2640 );
xor ( n2642 , n2615 , n2619 );
xor ( n2643 , n2642 , n2624 );
and ( n2644 , n2641 , n2643 );
and ( n2645 , n2473 , n1304 );
and ( n2646 , n2440 , n1301 );
nor ( n2647 , n2645 , n2646 );
xnor ( n2648 , n2647 , n1199 );
and ( n2649 , n2539 , n1273 );
and ( n2650 , n2506 , n1271 );
nor ( n2651 , n2649 , n2650 );
xnor ( n2652 , n2651 , n1202 );
and ( n2653 , n2648 , n2652 );
and ( n2654 , n2604 , n1213 );
and ( n2655 , n2571 , n1211 );
nor ( n2656 , n2654 , n2655 );
xnor ( n2657 , n2656 , n1219 );
and ( n2658 , n2652 , n2657 );
and ( n2659 , n2648 , n2657 );
or ( n2660 , n2653 , n2658 , n2659 );
and ( n2661 , n2643 , n2660 );
and ( n2662 , n2641 , n2660 );
or ( n2663 , n2644 , n2661 , n2662 );
xor ( n2664 , n2608 , n2610 );
xor ( n2665 , n2664 , n2627 );
and ( n2666 , n2663 , n2665 );
xor ( n2667 , n763 , n1175 );
buf ( n2668 , n2667 );
buf ( n2669 , n2668 );
buf ( n2670 , n2669 );
and ( n2671 , n2670 , n1192 );
and ( n2672 , n2637 , n1190 );
nor ( n2673 , n2671 , n2672 );
not ( n2674 , n2673 );
xor ( n2675 , n2648 , n2652 );
xor ( n2676 , n2675 , n2657 );
and ( n2677 , n2674 , n2676 );
and ( n2678 , n2506 , n1304 );
and ( n2679 , n2473 , n1301 );
nor ( n2680 , n2678 , n2679 );
xnor ( n2681 , n2680 , n1199 );
and ( n2682 , n2571 , n1273 );
and ( n2683 , n2539 , n1271 );
nor ( n2684 , n2682 , n2683 );
xnor ( n2685 , n2684 , n1202 );
and ( n2686 , n2681 , n2685 );
and ( n2687 , n2637 , n1213 );
and ( n2688 , n2604 , n1211 );
nor ( n2689 , n2687 , n2688 );
xnor ( n2690 , n2689 , n1219 );
and ( n2691 , n2685 , n2690 );
and ( n2692 , n2681 , n2690 );
or ( n2693 , n2686 , n2691 , n2692 );
and ( n2694 , n2676 , n2693 );
and ( n2695 , n2674 , n2693 );
or ( n2696 , n2677 , n2694 , n2695 );
xor ( n2697 , n2641 , n2643 );
xor ( n2698 , n2697 , n2660 );
and ( n2699 , n2696 , n2698 );
xor ( n2700 , n2674 , n2676 );
xor ( n2701 , n2700 , n2693 );
xor ( n2702 , n764 , n1174 );
buf ( n2703 , n2702 );
buf ( n2704 , n2703 );
buf ( n2705 , n2704 );
and ( n2706 , n2705 , n1192 );
and ( n2707 , n2670 , n1190 );
nor ( n2708 , n2706 , n2707 );
not ( n2709 , n2708 );
xor ( n2710 , n2681 , n2685 );
xor ( n2711 , n2710 , n2690 );
and ( n2712 , n2709 , n2711 );
buf ( n2713 , n372 );
buf ( n2714 , n2713 );
not ( n2715 , n2714 );
buf ( n2716 , n378 );
buf ( n2717 , n2716 );
not ( n2718 , n2717 );
and ( n2719 , n2718 , n2714 );
nor ( n2720 , n2715 , n2719 );
not ( n2721 , n2720 );
buf ( n2722 , n371 );
buf ( n2723 , n2722 );
buf ( n2724 , n379 );
buf ( n2725 , n2724 );
and ( n2726 , n2723 , n2725 );
not ( n2727 , n2726 );
and ( n2728 , n2721 , n2727 );
buf ( n2729 , n370 );
buf ( n2730 , n2729 );
not ( n2731 , n2730 );
buf ( n2732 , n380 );
buf ( n2733 , n2732 );
and ( n2734 , n2731 , n2733 );
not ( n2735 , n2733 );
nor ( n2736 , n2734 , n2735 );
not ( n2737 , n2736 );
and ( n2738 , n2727 , n2737 );
and ( n2739 , n2721 , n2737 );
or ( n2740 , n2728 , n2738 , n2739 );
not ( n2741 , n2723 );
and ( n2742 , n2718 , n2723 );
nor ( n2743 , n2741 , n2742 );
not ( n2744 , n2743 );
and ( n2745 , n2740 , n2744 );
and ( n2746 , n2731 , n2725 );
not ( n2747 , n2725 );
nor ( n2748 , n2746 , n2747 );
not ( n2749 , n2748 );
and ( n2750 , n2744 , n2749 );
and ( n2751 , n2740 , n2749 );
or ( n2752 , n2745 , n2750 , n2751 );
and ( n2753 , n2571 , n1304 );
and ( n2754 , n2539 , n1301 );
nor ( n2755 , n2753 , n2754 );
xnor ( n2756 , n2755 , n1199 );
and ( n2757 , n2752 , n2756 );
and ( n2758 , n2730 , n2717 );
not ( n2759 , n2758 );
and ( n2760 , n2756 , n2759 );
and ( n2761 , n2752 , n2759 );
or ( n2762 , n2757 , n2760 , n2761 );
and ( n2763 , n2539 , n1304 );
and ( n2764 , n2506 , n1301 );
nor ( n2765 , n2763 , n2764 );
xnor ( n2766 , n2765 , n1199 );
and ( n2767 , n2762 , n2766 );
and ( n2768 , n2604 , n1273 );
and ( n2769 , n2571 , n1271 );
nor ( n2770 , n2768 , n2769 );
xnor ( n2771 , n2770 , n1202 );
and ( n2772 , n2766 , n2771 );
and ( n2773 , n2762 , n2771 );
or ( n2774 , n2767 , n2772 , n2773 );
and ( n2775 , n2711 , n2774 );
and ( n2776 , n2709 , n2774 );
or ( n2777 , n2712 , n2775 , n2776 );
and ( n2778 , n2701 , n2777 );
and ( n2779 , n2670 , n1213 );
and ( n2780 , n2637 , n1211 );
nor ( n2781 , n2779 , n2780 );
xnor ( n2782 , n2781 , n1219 );
xor ( n2783 , n765 , n1173 );
buf ( n2784 , n2783 );
buf ( n2785 , n2784 );
buf ( n2786 , n2785 );
and ( n2787 , n2786 , n1192 );
and ( n2788 , n2705 , n1190 );
nor ( n2789 , n2787 , n2788 );
not ( n2790 , n2789 );
and ( n2791 , n2782 , n2790 );
xor ( n2792 , n2762 , n2766 );
xor ( n2793 , n2792 , n2771 );
and ( n2794 , n2790 , n2793 );
and ( n2795 , n2782 , n2793 );
or ( n2796 , n2791 , n2794 , n2795 );
xor ( n2797 , n2709 , n2711 );
xor ( n2798 , n2797 , n2774 );
and ( n2799 , n2796 , n2798 );
buf ( n2800 , n373 );
buf ( n2801 , n2800 );
not ( n2802 , n2801 );
and ( n2803 , n2718 , n2801 );
nor ( n2804 , n2802 , n2803 );
not ( n2805 , n2804 );
and ( n2806 , n2714 , n2725 );
not ( n2807 , n2806 );
and ( n2808 , n2805 , n2807 );
buf ( n2809 , n381 );
buf ( n2810 , n2809 );
and ( n2811 , n2731 , n2810 );
not ( n2812 , n2810 );
nor ( n2813 , n2811 , n2812 );
not ( n2814 , n2813 );
and ( n2815 , n2807 , n2814 );
and ( n2816 , n2805 , n2814 );
or ( n2817 , n2808 , n2815 , n2816 );
and ( n2818 , n2801 , n2725 );
not ( n2819 , n2818 );
and ( n2820 , n2723 , n2810 );
not ( n2821 , n2820 );
and ( n2822 , n2819 , n2821 );
buf ( n2823 , n382 );
buf ( n2824 , n2823 );
and ( n2825 , n2731 , n2824 );
not ( n2826 , n2824 );
nor ( n2827 , n2825 , n2826 );
not ( n2828 , n2827 );
and ( n2829 , n2821 , n2828 );
and ( n2830 , n2819 , n2828 );
or ( n2831 , n2822 , n2829 , n2830 );
and ( n2832 , n2723 , n2733 );
not ( n2833 , n2832 );
and ( n2834 , n2831 , n2833 );
xor ( n2835 , n2805 , n2807 );
xor ( n2836 , n2835 , n2814 );
and ( n2837 , n2833 , n2836 );
and ( n2838 , n2831 , n2836 );
or ( n2839 , n2834 , n2837 , n2838 );
and ( n2840 , n2817 , n2839 );
xor ( n2841 , n2721 , n2727 );
xor ( n2842 , n2841 , n2737 );
and ( n2843 , n2839 , n2842 );
and ( n2844 , n2817 , n2842 );
or ( n2845 , n2840 , n2843 , n2844 );
and ( n2846 , n2604 , n1304 );
and ( n2847 , n2571 , n1301 );
nor ( n2848 , n2846 , n2847 );
xnor ( n2849 , n2848 , n1199 );
and ( n2850 , n2845 , n2849 );
xor ( n2851 , n2740 , n2744 );
xor ( n2852 , n2851 , n2749 );
and ( n2853 , n2849 , n2852 );
and ( n2854 , n2845 , n2852 );
or ( n2855 , n2850 , n2853 , n2854 );
and ( n2856 , n2637 , n1273 );
and ( n2857 , n2604 , n1271 );
nor ( n2858 , n2856 , n2857 );
xnor ( n2859 , n2858 , n1202 );
and ( n2860 , n2855 , n2859 );
xor ( n2861 , n2752 , n2756 );
xor ( n2862 , n2861 , n2759 );
and ( n2863 , n2859 , n2862 );
and ( n2864 , n2855 , n2862 );
or ( n2865 , n2860 , n2863 , n2864 );
and ( n2866 , n2705 , n1213 );
and ( n2867 , n2670 , n1211 );
nor ( n2868 , n2866 , n2867 );
xnor ( n2869 , n2868 , n1219 );
xor ( n2870 , n942 , n1171 );
buf ( n2871 , n2870 );
buf ( n2872 , n2871 );
buf ( n2873 , n2872 );
and ( n2874 , n2873 , n1192 );
and ( n2875 , n2786 , n1190 );
nor ( n2876 , n2874 , n2875 );
not ( n2877 , n2876 );
and ( n2878 , n2869 , n2877 );
xor ( n2879 , n2855 , n2859 );
xor ( n2880 , n2879 , n2862 );
and ( n2881 , n2877 , n2880 );
and ( n2882 , n2869 , n2880 );
or ( n2883 , n2878 , n2881 , n2882 );
and ( n2884 , n2865 , n2883 );
xor ( n2885 , n2782 , n2790 );
xor ( n2886 , n2885 , n2793 );
and ( n2887 , n2883 , n2886 );
and ( n2888 , n2865 , n2886 );
or ( n2889 , n2884 , n2887 , n2888 );
and ( n2890 , n2798 , n2889 );
and ( n2891 , n2796 , n2889 );
or ( n2892 , n2799 , n2890 , n2891 );
and ( n2893 , n2777 , n2892 );
and ( n2894 , n2701 , n2892 );
or ( n2895 , n2778 , n2893 , n2894 );
and ( n2896 , n2698 , n2895 );
and ( n2897 , n2696 , n2895 );
or ( n2898 , n2699 , n2896 , n2897 );
and ( n2899 , n2665 , n2898 );
and ( n2900 , n2663 , n2898 );
or ( n2901 , n2666 , n2899 , n2900 );
and ( n2902 , n2632 , n2901 );
and ( n2903 , n2630 , n2901 );
or ( n2904 , n2633 , n2902 , n2903 );
and ( n2905 , n2599 , n2904 );
and ( n2906 , n2597 , n2904 );
or ( n2907 , n2600 , n2905 , n2906 );
and ( n2908 , n2567 , n2907 );
and ( n2909 , n2565 , n2907 );
or ( n2910 , n2568 , n2908 , n2909 );
and ( n2911 , n2534 , n2910 );
and ( n2912 , n2532 , n2910 );
or ( n2913 , n2535 , n2911 , n2912 );
and ( n2914 , n2501 , n2913 );
and ( n2915 , n2499 , n2913 );
or ( n2916 , n2502 , n2914 , n2915 );
and ( n2917 , n2468 , n2916 );
and ( n2918 , n2466 , n2916 );
or ( n2919 , n2469 , n2917 , n2918 );
and ( n2920 , n2435 , n2919 );
and ( n2921 , n2433 , n2919 );
or ( n2922 , n2436 , n2920 , n2921 );
and ( n2923 , n2402 , n2922 );
and ( n2924 , n2400 , n2922 );
or ( n2925 , n2403 , n2923 , n2924 );
and ( n2926 , n2369 , n2925 );
and ( n2927 , n2367 , n2925 );
or ( n2928 , n2370 , n2926 , n2927 );
and ( n2929 , n2336 , n2928 );
and ( n2930 , n2334 , n2928 );
or ( n2931 , n2337 , n2929 , n2930 );
and ( n2932 , n2303 , n2931 );
and ( n2933 , n2301 , n2931 );
or ( n2934 , n2304 , n2932 , n2933 );
and ( n2935 , n2270 , n2934 );
and ( n2936 , n2268 , n2934 );
or ( n2937 , n2271 , n2935 , n2936 );
and ( n2938 , n2237 , n2937 );
and ( n2939 , n2235 , n2937 );
or ( n2940 , n2238 , n2938 , n2939 );
and ( n2941 , n2204 , n2940 );
and ( n2942 , n2202 , n2940 );
or ( n2943 , n2205 , n2941 , n2942 );
and ( n2944 , n2171 , n2943 );
and ( n2945 , n2169 , n2943 );
or ( n2946 , n2172 , n2944 , n2945 );
and ( n2947 , n2138 , n2946 );
and ( n2948 , n2136 , n2946 );
or ( n2949 , n2139 , n2947 , n2948 );
and ( n2950 , n2105 , n2949 );
and ( n2951 , n2103 , n2949 );
or ( n2952 , n2106 , n2950 , n2951 );
and ( n2953 , n2072 , n2952 );
and ( n2954 , n2070 , n2952 );
or ( n2955 , n2073 , n2953 , n2954 );
and ( n2956 , n2039 , n2955 );
and ( n2957 , n2037 , n2955 );
or ( n2958 , n2040 , n2956 , n2957 );
and ( n2959 , n2006 , n2958 );
and ( n2960 , n2004 , n2958 );
or ( n2961 , n2007 , n2959 , n2960 );
and ( n2962 , n1973 , n2961 );
and ( n2963 , n1971 , n2961 );
or ( n2964 , n1974 , n2962 , n2963 );
and ( n2965 , n1940 , n2964 );
and ( n2966 , n1938 , n2964 );
or ( n2967 , n1941 , n2965 , n2966 );
and ( n2968 , n1907 , n2967 );
and ( n2969 , n1905 , n2967 );
or ( n2970 , n1908 , n2968 , n2969 );
and ( n2971 , n1874 , n2970 );
and ( n2972 , n1872 , n2970 );
or ( n2973 , n1875 , n2971 , n2972 );
and ( n2974 , n1841 , n2973 );
and ( n2975 , n1839 , n2973 );
or ( n2976 , n1842 , n2974 , n2975 );
and ( n2977 , n1808 , n2976 );
and ( n2978 , n1806 , n2976 );
or ( n2979 , n1809 , n2977 , n2978 );
and ( n2980 , n1775 , n2979 );
and ( n2981 , n1773 , n2979 );
or ( n2982 , n1776 , n2980 , n2981 );
and ( n2983 , n1742 , n2982 );
and ( n2984 , n1740 , n2982 );
or ( n2985 , n1743 , n2983 , n2984 );
and ( n2986 , n1709 , n2985 );
and ( n2987 , n1707 , n2985 );
or ( n2988 , n1710 , n2986 , n2987 );
and ( n2989 , n1676 , n2988 );
and ( n2990 , n1674 , n2988 );
or ( n2991 , n1677 , n2989 , n2990 );
and ( n2992 , n1643 , n2991 );
and ( n2993 , n1641 , n2991 );
or ( n2994 , n1644 , n2992 , n2993 );
and ( n2995 , n1610 , n2994 );
and ( n2996 , n1608 , n2994 );
or ( n2997 , n1611 , n2995 , n2996 );
and ( n2998 , n1577 , n2997 );
and ( n2999 , n1575 , n2997 );
or ( n3000 , n1578 , n2998 , n2999 );
and ( n3001 , n1544 , n3000 );
and ( n3002 , n1542 , n3000 );
or ( n3003 , n1545 , n3001 , n3002 );
and ( n3004 , n1511 , n3003 );
and ( n3005 , n1509 , n3003 );
or ( n3006 , n1512 , n3004 , n3005 );
and ( n3007 , n1478 , n3006 );
and ( n3008 , n1476 , n3006 );
or ( n3009 , n1479 , n3007 , n3008 );
and ( n3010 , n1445 , n3009 );
and ( n3011 , n1443 , n3009 );
or ( n3012 , n1446 , n3010 , n3011 );
and ( n3013 , n1412 , n3012 );
and ( n3014 , n1410 , n3012 );
or ( n3015 , n1413 , n3013 , n3014 );
and ( n3016 , n1409 , n3015 );
xor ( n3017 , n1410 , n1412 );
xor ( n3018 , n3017 , n3012 );
xor ( n3019 , n1443 , n1445 );
xor ( n3020 , n3019 , n3009 );
xor ( n3021 , n1476 , n1478 );
xor ( n3022 , n3021 , n3006 );
xor ( n3023 , n1509 , n1511 );
xor ( n3024 , n3023 , n3003 );
xor ( n3025 , n1542 , n1544 );
xor ( n3026 , n3025 , n3000 );
xor ( n3027 , n1575 , n1577 );
xor ( n3028 , n3027 , n2997 );
xor ( n3029 , n1608 , n1610 );
xor ( n3030 , n3029 , n2994 );
xor ( n3031 , n1641 , n1643 );
xor ( n3032 , n3031 , n2991 );
xor ( n3033 , n1674 , n1676 );
xor ( n3034 , n3033 , n2988 );
xor ( n3035 , n1707 , n1709 );
xor ( n3036 , n3035 , n2985 );
xor ( n3037 , n1740 , n1742 );
xor ( n3038 , n3037 , n2982 );
xor ( n3039 , n1773 , n1775 );
xor ( n3040 , n3039 , n2979 );
xor ( n3041 , n1806 , n1808 );
xor ( n3042 , n3041 , n2976 );
xor ( n3043 , n1839 , n1841 );
xor ( n3044 , n3043 , n2973 );
xor ( n3045 , n1872 , n1874 );
xor ( n3046 , n3045 , n2970 );
xor ( n3047 , n1905 , n1907 );
xor ( n3048 , n3047 , n2967 );
xor ( n3049 , n1938 , n1940 );
xor ( n3050 , n3049 , n2964 );
xor ( n3051 , n1971 , n1973 );
xor ( n3052 , n3051 , n2961 );
xor ( n3053 , n2004 , n2006 );
xor ( n3054 , n3053 , n2958 );
xor ( n3055 , n2037 , n2039 );
xor ( n3056 , n3055 , n2955 );
xor ( n3057 , n2070 , n2072 );
xor ( n3058 , n3057 , n2952 );
xor ( n3059 , n2103 , n2105 );
xor ( n3060 , n3059 , n2949 );
xor ( n3061 , n2136 , n2138 );
xor ( n3062 , n3061 , n2946 );
xor ( n3063 , n2169 , n2171 );
xor ( n3064 , n3063 , n2943 );
xor ( n3065 , n2202 , n2204 );
xor ( n3066 , n3065 , n2940 );
xor ( n3067 , n2235 , n2237 );
xor ( n3068 , n3067 , n2937 );
xor ( n3069 , n2268 , n2270 );
xor ( n3070 , n3069 , n2934 );
xor ( n3071 , n2301 , n2303 );
xor ( n3072 , n3071 , n2931 );
xor ( n3073 , n2334 , n2336 );
xor ( n3074 , n3073 , n2928 );
xor ( n3075 , n2367 , n2369 );
xor ( n3076 , n3075 , n2925 );
xor ( n3077 , n2400 , n2402 );
xor ( n3078 , n3077 , n2922 );
xor ( n3079 , n2433 , n2435 );
xor ( n3080 , n3079 , n2919 );
xor ( n3081 , n2466 , n2468 );
xor ( n3082 , n3081 , n2916 );
xor ( n3083 , n2499 , n2501 );
xor ( n3084 , n3083 , n2913 );
xor ( n3085 , n2532 , n2534 );
xor ( n3086 , n3085 , n2910 );
xor ( n3087 , n2565 , n2567 );
xor ( n3088 , n3087 , n2907 );
xor ( n3089 , n2597 , n2599 );
xor ( n3090 , n3089 , n2904 );
xor ( n3091 , n2630 , n2632 );
xor ( n3092 , n3091 , n2901 );
xor ( n3093 , n2663 , n2665 );
xor ( n3094 , n3093 , n2898 );
xor ( n3095 , n2696 , n2698 );
xor ( n3096 , n3095 , n2895 );
xor ( n3097 , n2701 , n2777 );
xor ( n3098 , n3097 , n2892 );
xor ( n3099 , n2796 , n2798 );
xor ( n3100 , n3099 , n2889 );
xor ( n3101 , n2865 , n2883 );
xor ( n3102 , n3101 , n2886 );
and ( n3103 , n2786 , n1213 );
and ( n3104 , n2705 , n1211 );
nor ( n3105 , n3103 , n3104 );
xnor ( n3106 , n3105 , n1219 );
and ( n3107 , n2637 , n1304 );
and ( n3108 , n2604 , n1301 );
nor ( n3109 , n3107 , n3108 );
xnor ( n3110 , n3109 , n1199 );
and ( n3111 , n2705 , n1273 );
and ( n3112 , n2670 , n1271 );
nor ( n3113 , n3111 , n3112 );
xnor ( n3114 , n3113 , n1202 );
and ( n3115 , n3110 , n3114 );
and ( n3116 , n2873 , n1213 );
and ( n3117 , n2786 , n1211 );
nor ( n3118 , n3116 , n3117 );
xnor ( n3119 , n3118 , n1219 );
and ( n3120 , n3114 , n3119 );
and ( n3121 , n3110 , n3119 );
or ( n3122 , n3115 , n3120 , n3121 );
and ( n3123 , n3106 , n3122 );
and ( n3124 , n2670 , n1304 );
and ( n3125 , n2637 , n1301 );
nor ( n3126 , n3124 , n3125 );
xnor ( n3127 , n3126 , n1199 );
and ( n3128 , n2786 , n1273 );
and ( n3129 , n2705 , n1271 );
nor ( n3130 , n3128 , n3129 );
xnor ( n3131 , n3130 , n1202 );
and ( n3132 , n3127 , n3131 );
xor ( n3133 , n945 , n1169 );
buf ( n3134 , n3133 );
buf ( n3135 , n3134 );
buf ( n3136 , n3135 );
and ( n3137 , n3136 , n1213 );
and ( n3138 , n2873 , n1211 );
nor ( n3139 , n3137 , n3138 );
xnor ( n3140 , n3139 , n1219 );
and ( n3141 , n3131 , n3140 );
and ( n3142 , n3127 , n3140 );
or ( n3143 , n3132 , n3141 , n3142 );
xor ( n3144 , n3110 , n3114 );
xor ( n3145 , n3144 , n3119 );
and ( n3146 , n3143 , n3145 );
xor ( n3147 , n1132 , n1165 );
buf ( n3148 , n3147 );
buf ( n3149 , n3148 );
buf ( n3150 , n3149 );
and ( n3151 , n3150 , n1192 );
xor ( n3152 , n1129 , n1167 );
buf ( n3153 , n3152 );
buf ( n3154 , n3153 );
buf ( n3155 , n3154 );
and ( n3156 , n3155 , n1190 );
nor ( n3157 , n3151 , n3156 );
not ( n3158 , n3157 );
and ( n3159 , n2705 , n1304 );
and ( n3160 , n2670 , n1301 );
nor ( n3161 , n3159 , n3160 );
xnor ( n3162 , n3161 , n1199 );
and ( n3163 , n2873 , n1273 );
and ( n3164 , n2786 , n1271 );
nor ( n3165 , n3163 , n3164 );
xnor ( n3166 , n3165 , n1202 );
and ( n3167 , n3162 , n3166 );
and ( n3168 , n3155 , n1213 );
and ( n3169 , n3136 , n1211 );
nor ( n3170 , n3168 , n3169 );
xnor ( n3171 , n3170 , n1219 );
and ( n3172 , n3166 , n3171 );
and ( n3173 , n3162 , n3171 );
or ( n3174 , n3167 , n3172 , n3173 );
and ( n3175 , n3158 , n3174 );
xor ( n3176 , n3127 , n3131 );
xor ( n3177 , n3176 , n3140 );
and ( n3178 , n3174 , n3177 );
and ( n3179 , n3158 , n3177 );
or ( n3180 , n3175 , n3178 , n3179 );
and ( n3181 , n3145 , n3180 );
and ( n3182 , n3143 , n3180 );
or ( n3183 , n3146 , n3181 , n3182 );
and ( n3184 , n3122 , n3183 );
and ( n3185 , n3106 , n3183 );
or ( n3186 , n3123 , n3184 , n3185 );
and ( n3187 , n2670 , n1273 );
and ( n3188 , n2637 , n1271 );
nor ( n3189 , n3187 , n3188 );
xnor ( n3190 , n3189 , n1202 );
and ( n3191 , n3136 , n1192 );
and ( n3192 , n2873 , n1190 );
nor ( n3193 , n3191 , n3192 );
not ( n3194 , n3193 );
and ( n3195 , n3190 , n3194 );
xor ( n3196 , n2845 , n2849 );
xor ( n3197 , n3196 , n2852 );
and ( n3198 , n3194 , n3197 );
and ( n3199 , n3190 , n3197 );
or ( n3200 , n3195 , n3198 , n3199 );
and ( n3201 , n3186 , n3200 );
xor ( n3202 , n2869 , n2877 );
xor ( n3203 , n3202 , n2880 );
and ( n3204 , n3200 , n3203 );
and ( n3205 , n3186 , n3203 );
or ( n3206 , n3201 , n3204 , n3205 );
and ( n3207 , n3102 , n3206 );
xor ( n3208 , n3106 , n3122 );
xor ( n3209 , n3208 , n3183 );
xor ( n3210 , n3190 , n3194 );
xor ( n3211 , n3210 , n3197 );
and ( n3212 , n3209 , n3211 );
and ( n3213 , n2801 , n2733 );
not ( n3214 , n3213 );
and ( n3215 , n2714 , n2810 );
not ( n3216 , n3215 );
and ( n3217 , n3214 , n3216 );
buf ( n3218 , n383 );
buf ( n3219 , n3218 );
and ( n3220 , n2731 , n3219 );
not ( n3221 , n3219 );
nor ( n3222 , n3220 , n3221 );
not ( n3223 , n3222 );
and ( n3224 , n3216 , n3223 );
and ( n3225 , n3214 , n3223 );
or ( n3226 , n3217 , n3224 , n3225 );
buf ( n3227 , n374 );
buf ( n3228 , n3227 );
not ( n3229 , n3228 );
and ( n3230 , n2718 , n3228 );
nor ( n3231 , n3229 , n3230 );
not ( n3232 , n3231 );
and ( n3233 , n3226 , n3232 );
and ( n3234 , n2714 , n2733 );
not ( n3235 , n3234 );
and ( n3236 , n3232 , n3235 );
and ( n3237 , n3226 , n3235 );
or ( n3238 , n3233 , n3236 , n3237 );
buf ( n3239 , n375 );
buf ( n3240 , n3239 );
not ( n3241 , n3240 );
and ( n3242 , n2718 , n3240 );
nor ( n3243 , n3241 , n3242 );
not ( n3244 , n3243 );
and ( n3245 , n3228 , n2725 );
not ( n3246 , n3245 );
and ( n3247 , n3244 , n3246 );
and ( n3248 , n2723 , n2824 );
not ( n3249 , n3248 );
and ( n3250 , n3246 , n3249 );
and ( n3251 , n3244 , n3249 );
or ( n3252 , n3247 , n3250 , n3251 );
xor ( n3253 , n2819 , n2821 );
xor ( n3254 , n3253 , n2828 );
and ( n3255 , n3252 , n3254 );
xor ( n3256 , n3226 , n3232 );
xor ( n3257 , n3256 , n3235 );
and ( n3258 , n3254 , n3257 );
and ( n3259 , n3252 , n3257 );
or ( n3260 , n3255 , n3258 , n3259 );
and ( n3261 , n3238 , n3260 );
xor ( n3262 , n2831 , n2833 );
xor ( n3263 , n3262 , n2836 );
and ( n3264 , n3260 , n3263 );
and ( n3265 , n3238 , n3263 );
or ( n3266 , n3261 , n3264 , n3265 );
xor ( n3267 , n2817 , n2839 );
xor ( n3268 , n3267 , n2842 );
or ( n3269 , n3266 , n3268 );
and ( n3270 , n3211 , n3269 );
and ( n3271 , n3209 , n3269 );
or ( n3272 , n3212 , n3270 , n3271 );
and ( n3273 , n3155 , n1192 );
and ( n3274 , n3136 , n1190 );
nor ( n3275 , n3273 , n3274 );
xnor ( n3276 , n3266 , n3268 );
and ( n3277 , n3275 , n3276 );
not ( n3278 , n3275 );
buf ( n3279 , n3278 );
and ( n3280 , n3277 , n3279 );
xor ( n3281 , n3143 , n3145 );
xor ( n3282 , n3281 , n3180 );
xor ( n3283 , n1134 , n1164 );
buf ( n3284 , n3283 );
buf ( n3285 , n3284 );
buf ( n3286 , n3285 );
and ( n3287 , n3286 , n1192 );
and ( n3288 , n3150 , n1190 );
nor ( n3289 , n3287 , n3288 );
not ( n3290 , n3289 );
and ( n3291 , n2786 , n1304 );
and ( n3292 , n2705 , n1301 );
nor ( n3293 , n3291 , n3292 );
xnor ( n3294 , n3293 , n1199 );
and ( n3295 , n3136 , n1273 );
and ( n3296 , n2873 , n1271 );
nor ( n3297 , n3295 , n3296 );
xnor ( n3298 , n3297 , n1202 );
and ( n3299 , n3294 , n3298 );
and ( n3300 , n3150 , n1213 );
and ( n3301 , n3155 , n1211 );
nor ( n3302 , n3300 , n3301 );
xnor ( n3303 , n3302 , n1219 );
and ( n3304 , n3298 , n3303 );
and ( n3305 , n3294 , n3303 );
or ( n3306 , n3299 , n3304 , n3305 );
and ( n3307 , n3290 , n3306 );
xor ( n3308 , n3162 , n3166 );
xor ( n3309 , n3308 , n3171 );
and ( n3310 , n3306 , n3309 );
and ( n3311 , n3290 , n3309 );
or ( n3312 , n3307 , n3310 , n3311 );
xor ( n3313 , n3158 , n3174 );
xor ( n3314 , n3313 , n3177 );
and ( n3315 , n3312 , n3314 );
xor ( n3316 , n1135 , n1163 );
buf ( n3317 , n3316 );
buf ( n3318 , n3317 );
buf ( n3319 , n3318 );
and ( n3320 , n3319 , n1192 );
and ( n3321 , n3286 , n1190 );
nor ( n3322 , n3320 , n3321 );
not ( n3323 , n3322 );
xor ( n3324 , n3214 , n3216 );
xor ( n3325 , n3324 , n3223 );
and ( n3326 , n3323 , n3325 );
buf ( n3327 , n376 );
buf ( n3328 , n3327 );
not ( n3329 , n3328 );
and ( n3330 , n2718 , n3328 );
nor ( n3331 , n3329 , n3330 );
not ( n3332 , n3331 );
and ( n3333 , n3228 , n2733 );
not ( n3334 , n3333 );
and ( n3335 , n3332 , n3334 );
and ( n3336 , n2723 , n3219 );
not ( n3337 , n3336 );
and ( n3338 , n3334 , n3337 );
and ( n3339 , n3332 , n3337 );
or ( n3340 , n3335 , n3338 , n3339 );
and ( n3341 , n3325 , n3340 );
and ( n3342 , n3323 , n3340 );
or ( n3343 , n3326 , n3341 , n3342 );
and ( n3344 , n2873 , n1304 );
and ( n3345 , n2786 , n1301 );
nor ( n3346 , n3344 , n3345 );
xnor ( n3347 , n3346 , n1199 );
and ( n3348 , n3155 , n1273 );
and ( n3349 , n3136 , n1271 );
nor ( n3350 , n3348 , n3349 );
xnor ( n3351 , n3350 , n1202 );
and ( n3352 , n3347 , n3351 );
and ( n3353 , n3286 , n1213 );
and ( n3354 , n3150 , n1211 );
nor ( n3355 , n3353 , n3354 );
xnor ( n3356 , n3355 , n1219 );
and ( n3357 , n3351 , n3356 );
and ( n3358 , n3347 , n3356 );
or ( n3359 , n3352 , n3357 , n3358 );
xor ( n3360 , n1137 , n1162 );
buf ( n3361 , n3360 );
buf ( n3362 , n3361 );
buf ( n3363 , n3362 );
and ( n3364 , n3363 , n1192 );
and ( n3365 , n3319 , n1190 );
nor ( n3366 , n3364 , n3365 );
not ( n3367 , n3366 );
and ( n3368 , n3240 , n2725 );
not ( n3369 , n3368 );
and ( n3370 , n3367 , n3369 );
and ( n3371 , n2801 , n2810 );
not ( n3372 , n3371 );
and ( n3373 , n3369 , n3372 );
and ( n3374 , n3367 , n3372 );
or ( n3375 , n3370 , n3373 , n3374 );
and ( n3376 , n3359 , n3375 );
xor ( n3377 , n3294 , n3298 );
xor ( n3378 , n3377 , n3303 );
and ( n3379 , n3375 , n3378 );
and ( n3380 , n3359 , n3378 );
or ( n3381 , n3376 , n3379 , n3380 );
and ( n3382 , n3343 , n3381 );
xor ( n3383 , n3290 , n3306 );
xor ( n3384 , n3383 , n3309 );
and ( n3385 , n3381 , n3384 );
and ( n3386 , n3343 , n3384 );
or ( n3387 , n3382 , n3385 , n3386 );
and ( n3388 , n3314 , n3387 );
and ( n3389 , n3312 , n3387 );
or ( n3390 , n3315 , n3388 , n3389 );
and ( n3391 , n3282 , n3390 );
xor ( n3392 , n3238 , n3260 );
xor ( n3393 , n3392 , n3263 );
xor ( n3394 , n3252 , n3254 );
xor ( n3395 , n3394 , n3257 );
buf ( n3396 , n377 );
buf ( n3397 , n3396 );
not ( n3398 , n3397 );
and ( n3399 , n2718 , n3397 );
nor ( n3400 , n3398 , n3399 );
not ( n3401 , n3400 );
and ( n3402 , n3328 , n2725 );
not ( n3403 , n3402 );
and ( n3404 , n3401 , n3403 );
and ( n3405 , n3240 , n2733 );
not ( n3406 , n3405 );
and ( n3407 , n3403 , n3406 );
and ( n3408 , n3401 , n3406 );
or ( n3409 , n3404 , n3407 , n3408 );
and ( n3410 , n2714 , n2824 );
not ( n3411 , n3410 );
and ( n3412 , n3409 , n3411 );
buf ( n3413 , n384 );
buf ( n3414 , n3413 );
and ( n3415 , n2731 , n3414 );
not ( n3416 , n3414 );
nor ( n3417 , n3415 , n3416 );
not ( n3418 , n3417 );
and ( n3419 , n3411 , n3418 );
and ( n3420 , n3409 , n3418 );
or ( n3421 , n3412 , n3419 , n3420 );
xor ( n3422 , n3244 , n3246 );
xor ( n3423 , n3422 , n3249 );
or ( n3424 , n3421 , n3423 );
and ( n3425 , n3395 , n3424 );
xor ( n3426 , n3332 , n3334 );
xor ( n3427 , n3426 , n3337 );
and ( n3428 , n3228 , n2810 );
not ( n3429 , n3428 );
and ( n3430 , n2801 , n2824 );
not ( n3431 , n3430 );
and ( n3432 , n3429 , n3431 );
buf ( n3433 , n385 );
buf ( n3434 , n3433 );
and ( n3435 , n2731 , n3434 );
not ( n3436 , n3434 );
nor ( n3437 , n3435 , n3436 );
not ( n3438 , n3437 );
and ( n3439 , n3431 , n3438 );
and ( n3440 , n3429 , n3438 );
or ( n3441 , n3432 , n3439 , n3440 );
and ( n3442 , n3427 , n3441 );
and ( n3443 , n3136 , n1304 );
and ( n3444 , n2873 , n1301 );
nor ( n3445 , n3443 , n3444 );
xnor ( n3446 , n3445 , n1199 );
and ( n3447 , n3150 , n1273 );
and ( n3448 , n3155 , n1271 );
nor ( n3449 , n3447 , n3448 );
xnor ( n3450 , n3449 , n1202 );
and ( n3451 , n3446 , n3450 );
and ( n3452 , n3319 , n1213 );
and ( n3453 , n3286 , n1211 );
nor ( n3454 , n3452 , n3453 );
xnor ( n3455 , n3454 , n1219 );
and ( n3456 , n3450 , n3455 );
and ( n3457 , n3446 , n3455 );
or ( n3458 , n3451 , n3456 , n3457 );
and ( n3459 , n3441 , n3458 );
and ( n3460 , n3427 , n3458 );
or ( n3461 , n3442 , n3459 , n3460 );
xor ( n3462 , n1140 , n1160 );
buf ( n3463 , n3462 );
buf ( n3464 , n3463 );
buf ( n3465 , n3464 );
and ( n3466 , n3465 , n1192 );
and ( n3467 , n3363 , n1190 );
nor ( n3468 , n3466 , n3467 );
not ( n3469 , n3468 );
and ( n3470 , n2714 , n3219 );
not ( n3471 , n3470 );
and ( n3472 , n3469 , n3471 );
and ( n3473 , n2723 , n3414 );
not ( n3474 , n3473 );
and ( n3475 , n3471 , n3474 );
and ( n3476 , n3469 , n3474 );
or ( n3477 , n3472 , n3475 , n3476 );
xor ( n3478 , n3347 , n3351 );
xor ( n3479 , n3478 , n3356 );
and ( n3480 , n3477 , n3479 );
xor ( n3481 , n3367 , n3369 );
xor ( n3482 , n3481 , n3372 );
and ( n3483 , n3479 , n3482 );
and ( n3484 , n3477 , n3482 );
or ( n3485 , n3480 , n3483 , n3484 );
and ( n3486 , n3461 , n3485 );
xor ( n3487 , n3323 , n3325 );
xor ( n3488 , n3487 , n3340 );
and ( n3489 , n3485 , n3488 );
and ( n3490 , n3461 , n3488 );
or ( n3491 , n3486 , n3489 , n3490 );
and ( n3492 , n3424 , n3491 );
and ( n3493 , n3395 , n3491 );
or ( n3494 , n3425 , n3492 , n3493 );
and ( n3495 , n3393 , n3494 );
xor ( n3496 , n3312 , n3314 );
xor ( n3497 , n3496 , n3387 );
and ( n3498 , n3494 , n3497 );
and ( n3499 , n3393 , n3497 );
or ( n3500 , n3495 , n3498 , n3499 );
and ( n3501 , n3390 , n3500 );
and ( n3502 , n3282 , n3500 );
or ( n3503 , n3391 , n3501 , n3502 );
and ( n3504 , n3279 , n3503 );
and ( n3505 , n3277 , n3503 );
or ( n3506 , n3280 , n3504 , n3505 );
and ( n3507 , n3272 , n3506 );
xor ( n3508 , n3186 , n3200 );
xor ( n3509 , n3508 , n3203 );
and ( n3510 , n3506 , n3509 );
and ( n3511 , n3272 , n3509 );
or ( n3512 , n3507 , n3510 , n3511 );
and ( n3513 , n3206 , n3512 );
and ( n3514 , n3102 , n3512 );
or ( n3515 , n3207 , n3513 , n3514 );
and ( n3516 , n3100 , n3515 );
xor ( n3517 , n3102 , n3206 );
xor ( n3518 , n3517 , n3512 );
xor ( n3519 , n3272 , n3506 );
xor ( n3520 , n3519 , n3509 );
xor ( n3521 , n3209 , n3211 );
xor ( n3522 , n3521 , n3269 );
xor ( n3523 , n3277 , n3279 );
xor ( n3524 , n3523 , n3503 );
and ( n3525 , n3522 , n3524 );
xor ( n3526 , n3275 , n3276 );
xor ( n3527 , n3282 , n3390 );
xor ( n3528 , n3527 , n3500 );
and ( n3529 , n3526 , n3528 );
xor ( n3530 , n3343 , n3381 );
xor ( n3531 , n3530 , n3384 );
xor ( n3532 , n3359 , n3375 );
xor ( n3533 , n3532 , n3378 );
xnor ( n3534 , n3421 , n3423 );
and ( n3535 , n3533 , n3534 );
xor ( n3536 , n3409 , n3411 );
xor ( n3537 , n3536 , n3418 );
xor ( n3538 , n3429 , n3431 );
xor ( n3539 , n3538 , n3438 );
xor ( n3540 , n3401 , n3403 );
xor ( n3541 , n3540 , n3406 );
and ( n3542 , n3539 , n3541 );
and ( n3543 , n3397 , n2725 );
not ( n3544 , n3543 );
and ( n3545 , n3240 , n2810 );
not ( n3546 , n3545 );
and ( n3547 , n3544 , n3546 );
and ( n3548 , n2714 , n3414 );
not ( n3549 , n3548 );
and ( n3550 , n3546 , n3549 );
and ( n3551 , n3544 , n3549 );
or ( n3552 , n3547 , n3550 , n3551 );
and ( n3553 , n3541 , n3552 );
and ( n3554 , n3539 , n3552 );
or ( n3555 , n3542 , n3553 , n3554 );
and ( n3556 , n3537 , n3555 );
and ( n3557 , n3155 , n1304 );
and ( n3558 , n3136 , n1301 );
nor ( n3559 , n3557 , n3558 );
xnor ( n3560 , n3559 , n1199 );
and ( n3561 , n3286 , n1273 );
and ( n3562 , n3150 , n1271 );
nor ( n3563 , n3561 , n3562 );
xnor ( n3564 , n3563 , n1202 );
and ( n3565 , n3560 , n3564 );
and ( n3566 , n3363 , n1213 );
and ( n3567 , n3319 , n1211 );
nor ( n3568 , n3566 , n3567 );
xnor ( n3569 , n3568 , n1219 );
and ( n3570 , n3564 , n3569 );
and ( n3571 , n3560 , n3569 );
or ( n3572 , n3565 , n3570 , n3571 );
and ( n3573 , n3465 , n1190 );
and ( n3574 , n3328 , n2733 );
not ( n3575 , n3574 );
and ( n3576 , n3573 , n3575 );
and ( n3577 , n3228 , n2824 );
not ( n3578 , n3577 );
and ( n3579 , n3575 , n3578 );
and ( n3580 , n3573 , n3578 );
or ( n3581 , n3576 , n3579 , n3580 );
and ( n3582 , n3572 , n3581 );
xor ( n3583 , n3446 , n3450 );
xor ( n3584 , n3583 , n3455 );
and ( n3585 , n3581 , n3584 );
and ( n3586 , n3572 , n3584 );
or ( n3587 , n3582 , n3585 , n3586 );
and ( n3588 , n3555 , n3587 );
and ( n3589 , n3537 , n3587 );
or ( n3590 , n3556 , n3588 , n3589 );
and ( n3591 , n3534 , n3590 );
and ( n3592 , n3533 , n3590 );
or ( n3593 , n3535 , n3591 , n3592 );
and ( n3594 , n3531 , n3593 );
xor ( n3595 , n3395 , n3424 );
xor ( n3596 , n3595 , n3491 );
and ( n3597 , n3593 , n3596 );
and ( n3598 , n3531 , n3596 );
or ( n3599 , n3594 , n3597 , n3598 );
xor ( n3600 , n3393 , n3494 );
xor ( n3601 , n3600 , n3497 );
and ( n3602 , n3599 , n3601 );
xor ( n3603 , n3461 , n3485 );
xor ( n3604 , n3603 , n3488 );
xor ( n3605 , n3427 , n3441 );
xor ( n3606 , n3605 , n3458 );
xor ( n3607 , n3477 , n3479 );
xor ( n3608 , n3607 , n3482 );
and ( n3609 , n3606 , n3608 );
xor ( n3610 , n3469 , n3471 );
xor ( n3611 , n3610 , n3474 );
and ( n3612 , n3397 , n2733 );
not ( n3613 , n3612 );
buf ( n3614 , n3613 );
and ( n3615 , n2801 , n3219 );
not ( n3616 , n3615 );
and ( n3617 , n3614 , n3616 );
and ( n3618 , n2723 , n3434 );
not ( n3619 , n3618 );
and ( n3620 , n3616 , n3619 );
and ( n3621 , n3614 , n3619 );
or ( n3622 , n3617 , n3620 , n3621 );
and ( n3623 , n3611 , n3622 );
and ( n3624 , n3328 , n2810 );
not ( n3625 , n3624 );
and ( n3626 , n3228 , n3219 );
not ( n3627 , n3626 );
and ( n3628 , n3625 , n3627 );
and ( n3629 , n2714 , n3434 );
not ( n3630 , n3629 );
and ( n3631 , n3627 , n3630 );
and ( n3632 , n3625 , n3630 );
or ( n3633 , n3628 , n3631 , n3632 );
xor ( n3634 , n3544 , n3546 );
xor ( n3635 , n3634 , n3549 );
or ( n3636 , n3633 , n3635 );
and ( n3637 , n3622 , n3636 );
and ( n3638 , n3611 , n3636 );
or ( n3639 , n3623 , n3637 , n3638 );
and ( n3640 , n3608 , n3639 );
and ( n3641 , n3606 , n3639 );
or ( n3642 , n3609 , n3640 , n3641 );
and ( n3643 , n3604 , n3642 );
xor ( n3644 , n3533 , n3534 );
xor ( n3645 , n3644 , n3590 );
and ( n3646 , n3642 , n3645 );
and ( n3647 , n3604 , n3645 );
or ( n3648 , n3643 , n3646 , n3647 );
xor ( n3649 , n3531 , n3593 );
xor ( n3650 , n3649 , n3596 );
and ( n3651 , n3648 , n3650 );
and ( n3652 , n3150 , n1304 );
and ( n3653 , n3155 , n1301 );
nor ( n3654 , n3652 , n3653 );
xnor ( n3655 , n3654 , n1199 );
and ( n3656 , n3319 , n1273 );
and ( n3657 , n3286 , n1271 );
nor ( n3658 , n3656 , n3657 );
xnor ( n3659 , n3658 , n1202 );
and ( n3660 , n3655 , n3659 );
and ( n3661 , n3465 , n1213 );
and ( n3662 , n3363 , n1211 );
nor ( n3663 , n3661 , n3662 );
xnor ( n3664 , n3663 , n1219 );
and ( n3665 , n3659 , n3664 );
and ( n3666 , n3655 , n3664 );
or ( n3667 , n3660 , n3665 , n3666 );
xor ( n3668 , n3560 , n3564 );
xor ( n3669 , n3668 , n3569 );
and ( n3670 , n3667 , n3669 );
xor ( n3671 , n3573 , n3575 );
xor ( n3672 , n3671 , n3578 );
and ( n3673 , n3669 , n3672 );
and ( n3674 , n3667 , n3672 );
or ( n3675 , n3670 , n3673 , n3674 );
xor ( n3676 , n3539 , n3541 );
xor ( n3677 , n3676 , n3552 );
and ( n3678 , n3675 , n3677 );
xor ( n3679 , n3572 , n3581 );
xor ( n3680 , n3679 , n3584 );
and ( n3681 , n3677 , n3680 );
and ( n3682 , n3675 , n3680 );
or ( n3683 , n3678 , n3681 , n3682 );
xor ( n3684 , n3537 , n3555 );
xor ( n3685 , n3684 , n3587 );
and ( n3686 , n3683 , n3685 );
and ( n3687 , n3240 , n2824 );
not ( n3688 , n3687 );
and ( n3689 , n3612 , n3688 );
and ( n3690 , n2801 , n3414 );
not ( n3691 , n3690 );
and ( n3692 , n3688 , n3691 );
and ( n3693 , n3612 , n3691 );
or ( n3694 , n3689 , n3692 , n3693 );
xor ( n3695 , n3614 , n3616 );
xor ( n3696 , n3695 , n3619 );
or ( n3697 , n3694 , n3696 );
xnor ( n3698 , n3633 , n3635 );
and ( n3699 , n3465 , n1211 );
not ( n3700 , n3699 );
and ( n3701 , n3700 , n1219 );
xor ( n3702 , n3625 , n3627 );
xor ( n3703 , n3702 , n3630 );
and ( n3704 , n3701 , n3703 );
xor ( n3705 , n3612 , n3688 );
xor ( n3706 , n3705 , n3691 );
and ( n3707 , n3703 , n3706 );
and ( n3708 , n3701 , n3706 );
or ( n3709 , n3704 , n3707 , n3708 );
and ( n3710 , n3698 , n3709 );
and ( n3711 , n3397 , n2810 );
not ( n3712 , n3711 );
and ( n3713 , n3240 , n3219 );
not ( n3714 , n3713 );
and ( n3715 , n3712 , n3714 );
and ( n3716 , n3228 , n3414 );
not ( n3717 , n3716 );
and ( n3718 , n3714 , n3717 );
and ( n3719 , n3712 , n3717 );
or ( n3720 , n3715 , n3718 , n3719 );
and ( n3721 , n3286 , n1304 );
and ( n3722 , n3150 , n1301 );
nor ( n3723 , n3721 , n3722 );
xnor ( n3724 , n3723 , n1199 );
and ( n3725 , n3363 , n1273 );
and ( n3726 , n3319 , n1271 );
nor ( n3727 , n3725 , n3726 );
xnor ( n3728 , n3727 , n1202 );
and ( n3729 , n3724 , n3728 );
and ( n3730 , n3728 , n3699 );
and ( n3731 , n3724 , n3699 );
or ( n3732 , n3729 , n3730 , n3731 );
and ( n3733 , n3720 , n3732 );
xor ( n3734 , n3655 , n3659 );
xor ( n3735 , n3734 , n3664 );
and ( n3736 , n3732 , n3735 );
and ( n3737 , n3720 , n3735 );
or ( n3738 , n3733 , n3736 , n3737 );
and ( n3739 , n3709 , n3738 );
and ( n3740 , n3698 , n3738 );
or ( n3741 , n3710 , n3739 , n3740 );
and ( n3742 , n3697 , n3741 );
xor ( n3743 , n3611 , n3622 );
xor ( n3744 , n3743 , n3636 );
and ( n3745 , n3741 , n3744 );
and ( n3746 , n3697 , n3744 );
or ( n3747 , n3742 , n3745 , n3746 );
and ( n3748 , n3685 , n3747 );
and ( n3749 , n3683 , n3747 );
or ( n3750 , n3686 , n3748 , n3749 );
xor ( n3751 , n3604 , n3642 );
xor ( n3752 , n3751 , n3645 );
and ( n3753 , n3750 , n3752 );
xor ( n3754 , n3606 , n3608 );
xor ( n3755 , n3754 , n3639 );
xor ( n3756 , n3675 , n3677 );
xor ( n3757 , n3756 , n3680 );
xor ( n3758 , n3667 , n3669 );
xor ( n3759 , n3758 , n3672 );
xnor ( n3760 , n3694 , n3696 );
and ( n3761 , n3759 , n3760 );
and ( n3762 , n3328 , n2824 );
not ( n3763 , n3762 );
and ( n3764 , n2801 , n3434 );
not ( n3765 , n3764 );
and ( n3766 , n3763 , n3765 );
xor ( n3767 , n3712 , n3714 );
xor ( n3768 , n3767 , n3717 );
and ( n3769 , n3765 , n3768 );
and ( n3770 , n3763 , n3768 );
or ( n3771 , n3766 , n3769 , n3770 );
and ( n3772 , n3397 , n2824 );
not ( n3773 , n3772 );
and ( n3774 , n3328 , n3219 );
not ( n3775 , n3774 );
and ( n3776 , n3773 , n3775 );
and ( n3777 , n3240 , n3414 );
not ( n3778 , n3777 );
and ( n3779 , n3775 , n3778 );
and ( n3780 , n3773 , n3778 );
or ( n3781 , n3776 , n3779 , n3780 );
and ( n3782 , n3319 , n1304 );
and ( n3783 , n3286 , n1301 );
nor ( n3784 , n3782 , n3783 );
xnor ( n3785 , n3784 , n1199 );
and ( n3786 , n3465 , n1273 );
and ( n3787 , n3363 , n1271 );
nor ( n3788 , n3786 , n3787 );
xnor ( n3789 , n3788 , n1202 );
and ( n3790 , n3785 , n3789 );
and ( n3791 , n3465 , n1271 );
not ( n3792 , n3791 );
and ( n3793 , n3792 , n1202 );
and ( n3794 , n3789 , n3793 );
and ( n3795 , n3785 , n3793 );
or ( n3796 , n3790 , n3794 , n3795 );
and ( n3797 , n3781 , n3796 );
xor ( n3798 , n3724 , n3728 );
xor ( n3799 , n3798 , n3699 );
and ( n3800 , n3796 , n3799 );
and ( n3801 , n3781 , n3799 );
or ( n3802 , n3797 , n3800 , n3801 );
and ( n3803 , n3771 , n3802 );
xor ( n3804 , n3701 , n3703 );
xor ( n3805 , n3804 , n3706 );
and ( n3806 , n3802 , n3805 );
and ( n3807 , n3771 , n3805 );
or ( n3808 , n3803 , n3806 , n3807 );
and ( n3809 , n3760 , n3808 );
and ( n3810 , n3759 , n3808 );
or ( n3811 , n3761 , n3809 , n3810 );
and ( n3812 , n3757 , n3811 );
xor ( n3813 , n3697 , n3741 );
xor ( n3814 , n3813 , n3744 );
and ( n3815 , n3811 , n3814 );
and ( n3816 , n3757 , n3814 );
or ( n3817 , n3812 , n3815 , n3816 );
or ( n3818 , n3755 , n3817 );
and ( n3819 , n3752 , n3818 );
and ( n3820 , n3750 , n3818 );
or ( n3821 , n3753 , n3819 , n3820 );
and ( n3822 , n3650 , n3821 );
and ( n3823 , n3648 , n3821 );
or ( n3824 , n3651 , n3822 , n3823 );
and ( n3825 , n3601 , n3824 );
and ( n3826 , n3599 , n3824 );
or ( n3827 , n3602 , n3825 , n3826 );
and ( n3828 , n3528 , n3827 );
and ( n3829 , n3526 , n3827 );
or ( n3830 , n3529 , n3828 , n3829 );
and ( n3831 , n3524 , n3830 );
and ( n3832 , n3522 , n3830 );
or ( n3833 , n3525 , n3831 , n3832 );
or ( n3834 , n3520 , n3833 );
or ( n3835 , n3518 , n3834 );
and ( n3836 , n3515 , n3835 );
and ( n3837 , n3100 , n3835 );
or ( n3838 , n3516 , n3836 , n3837 );
or ( n3839 , n3098 , n3838 );
or ( n3840 , n3096 , n3839 );
or ( n3841 , n3094 , n3840 );
or ( n3842 , n3092 , n3841 );
or ( n3843 , n3090 , n3842 );
or ( n3844 , n3088 , n3843 );
or ( n3845 , n3086 , n3844 );
or ( n3846 , n3084 , n3845 );
or ( n3847 , n3082 , n3846 );
or ( n3848 , n3080 , n3847 );
or ( n3849 , n3078 , n3848 );
or ( n3850 , n3076 , n3849 );
or ( n3851 , n3074 , n3850 );
or ( n3852 , n3072 , n3851 );
or ( n3853 , n3070 , n3852 );
or ( n3854 , n3068 , n3853 );
or ( n3855 , n3066 , n3854 );
or ( n3856 , n3064 , n3855 );
or ( n3857 , n3062 , n3856 );
or ( n3858 , n3060 , n3857 );
or ( n3859 , n3058 , n3858 );
or ( n3860 , n3056 , n3859 );
or ( n3861 , n3054 , n3860 );
or ( n3862 , n3052 , n3861 );
or ( n3863 , n3050 , n3862 );
or ( n3864 , n3048 , n3863 );
or ( n3865 , n3046 , n3864 );
or ( n3866 , n3044 , n3865 );
or ( n3867 , n3042 , n3866 );
or ( n3868 , n3040 , n3867 );
or ( n3869 , n3038 , n3868 );
or ( n3870 , n3036 , n3869 );
or ( n3871 , n3034 , n3870 );
or ( n3872 , n3032 , n3871 );
or ( n3873 , n3030 , n3872 );
or ( n3874 , n3028 , n3873 );
or ( n3875 , n3026 , n3874 );
or ( n3876 , n3024 , n3875 );
or ( n3877 , n3022 , n3876 );
or ( n3878 , n3020 , n3877 );
or ( n3879 , n3018 , n3878 );
and ( n3880 , n3015 , n3879 );
and ( n3881 , n1409 , n3879 );
or ( n3882 , n3016 , n3880 , n3881 );
or ( n3883 , n1407 , n3882 );
or ( n3884 , n1405 , n3883 );
and ( n3885 , n1403 , n3884 );
xor ( n3886 , n1403 , n3884 );
xnor ( n3887 , n1405 , n3883 );
xnor ( n3888 , n1407 , n3882 );
xor ( n3889 , n1409 , n3015 );
xor ( n3890 , n3889 , n3879 );
not ( n3891 , n3890 );
xnor ( n3892 , n3018 , n3878 );
xnor ( n3893 , n3020 , n3877 );
xnor ( n3894 , n3022 , n3876 );
xnor ( n3895 , n3024 , n3875 );
xnor ( n3896 , n3026 , n3874 );
xnor ( n3897 , n3028 , n3873 );
xnor ( n3898 , n3030 , n3872 );
xnor ( n3899 , n3032 , n3871 );
xnor ( n3900 , n3034 , n3870 );
xnor ( n3901 , n3036 , n3869 );
xnor ( n3902 , n3038 , n3868 );
xnor ( n3903 , n3040 , n3867 );
xnor ( n3904 , n3042 , n3866 );
xnor ( n3905 , n3044 , n3865 );
xnor ( n3906 , n3046 , n3864 );
xnor ( n3907 , n3048 , n3863 );
xnor ( n3908 , n3050 , n3862 );
xnor ( n3909 , n3052 , n3861 );
xnor ( n3910 , n3054 , n3860 );
xnor ( n3911 , n3056 , n3859 );
xnor ( n3912 , n3058 , n3858 );
xnor ( n3913 , n3060 , n3857 );
xnor ( n3914 , n3062 , n3856 );
xnor ( n3915 , n3064 , n3855 );
xnor ( n3916 , n3066 , n3854 );
xnor ( n3917 , n3068 , n3853 );
xnor ( n3918 , n3070 , n3852 );
xnor ( n3919 , n3072 , n3851 );
xnor ( n3920 , n3074 , n3850 );
xnor ( n3921 , n3076 , n3849 );
xnor ( n3922 , n3078 , n3848 );
xnor ( n3923 , n3080 , n3847 );
xnor ( n3924 , n3082 , n3846 );
xnor ( n3925 , n3084 , n3845 );
xnor ( n3926 , n3086 , n3844 );
xnor ( n3927 , n3088 , n3843 );
xnor ( n3928 , n3090 , n3842 );
xnor ( n3929 , n3092 , n3841 );
xnor ( n3930 , n3094 , n3840 );
xnor ( n3931 , n3096 , n3839 );
xnor ( n3932 , n3098 , n3838 );
xor ( n3933 , n3100 , n3515 );
xor ( n3934 , n3933 , n3835 );
xnor ( n3935 , n3518 , n3834 );
xnor ( n3936 , n3520 , n3833 );
xor ( n3937 , n3522 , n3524 );
xor ( n3938 , n3937 , n3830 );
xor ( n3939 , n3526 , n3528 );
xor ( n3940 , n3939 , n3827 );
not ( n3941 , n3940 );
xor ( n3942 , n3599 , n3601 );
xor ( n3943 , n3942 , n3824 );
not ( n3944 , n3943 );
xor ( n3945 , n3648 , n3650 );
xor ( n3946 , n3945 , n3821 );
not ( n3947 , n3946 );
xor ( n3948 , n3750 , n3752 );
xor ( n3949 , n3948 , n3818 );
not ( n3950 , n3949 );
xor ( n3951 , n3683 , n3685 );
xor ( n3952 , n3951 , n3747 );
xnor ( n3953 , n3755 , n3817 );
and ( n3954 , n3952 , n3953 );
xor ( n3955 , n3952 , n3953 );
xor ( n3956 , n3698 , n3709 );
xor ( n3957 , n3956 , n3738 );
xor ( n3958 , n3720 , n3732 );
xor ( n3959 , n3958 , n3735 );
and ( n3960 , n3228 , n3434 );
not ( n3961 , n3960 );
xor ( n3962 , n3773 , n3775 );
xor ( n3963 , n3962 , n3778 );
and ( n3964 , n3961 , n3963 );
and ( n3965 , n3363 , n1304 );
and ( n3966 , n3319 , n1301 );
nor ( n3967 , n3965 , n3966 );
xnor ( n3968 , n3967 , n1199 );
and ( n3969 , n3968 , n3791 );
and ( n3970 , n3328 , n3414 );
not ( n3971 , n3970 );
and ( n3972 , n3791 , n3971 );
and ( n3973 , n3968 , n3971 );
or ( n3974 , n3969 , n3972 , n3973 );
and ( n3975 , n3963 , n3974 );
and ( n3976 , n3961 , n3974 );
or ( n3977 , n3964 , n3975 , n3976 );
xor ( n3978 , n3763 , n3765 );
xor ( n3979 , n3978 , n3768 );
and ( n3980 , n3977 , n3979 );
xor ( n3981 , n3781 , n3796 );
xor ( n3982 , n3981 , n3799 );
and ( n3983 , n3979 , n3982 );
and ( n3984 , n3977 , n3982 );
or ( n3985 , n3980 , n3983 , n3984 );
and ( n3986 , n3959 , n3985 );
xor ( n3987 , n3771 , n3802 );
xor ( n3988 , n3987 , n3805 );
and ( n3989 , n3985 , n3988 );
and ( n3990 , n3959 , n3988 );
or ( n3991 , n3986 , n3989 , n3990 );
or ( n3992 , n3957 , n3991 );
xor ( n3993 , n3757 , n3811 );
xor ( n3994 , n3993 , n3814 );
and ( n3995 , n3992 , n3994 );
xor ( n3996 , n3992 , n3994 );
xor ( n3997 , n3759 , n3760 );
xor ( n3998 , n3997 , n3808 );
xnor ( n3999 , n3957 , n3991 );
and ( n4000 , n3998 , n3999 );
xor ( n4001 , n3998 , n3999 );
xor ( n4002 , n3959 , n3985 );
xor ( n4003 , n4002 , n3988 );
xor ( n4004 , n3785 , n3789 );
xor ( n4005 , n4004 , n3793 );
and ( n4006 , n3328 , n3434 );
not ( n4007 , n4006 );
buf ( n4008 , n4007 );
and ( n4009 , n3397 , n3219 );
not ( n4010 , n4009 );
or ( n4011 , n4008 , n4010 );
and ( n4012 , n4005 , n4011 );
and ( n4013 , n3240 , n3434 );
not ( n4014 , n4013 );
and ( n4015 , n3465 , n1301 );
not ( n4016 , n4015 );
and ( n4017 , n4016 , n1199 );
and ( n4018 , n3397 , n3414 );
not ( n4019 , n4018 );
and ( n4020 , n4017 , n4019 );
and ( n4021 , n4019 , n4006 );
and ( n4022 , n4017 , n4006 );
or ( n4023 , n4020 , n4021 , n4022 );
and ( n4024 , n4014 , n4023 );
xor ( n4025 , n3968 , n3791 );
xor ( n4026 , n4025 , n3971 );
and ( n4027 , n4023 , n4026 );
and ( n4028 , n4014 , n4026 );
or ( n4029 , n4024 , n4027 , n4028 );
and ( n4030 , n4011 , n4029 );
and ( n4031 , n4005 , n4029 );
or ( n4032 , n4012 , n4030 , n4031 );
xor ( n4033 , n3977 , n3979 );
xor ( n4034 , n4033 , n3982 );
and ( n4035 , n4032 , n4034 );
xor ( n4036 , n3961 , n3963 );
xor ( n4037 , n4036 , n3974 );
xnor ( n4038 , n4008 , n4010 );
and ( n4039 , n3465 , n1304 );
and ( n4040 , n3363 , n1301 );
nor ( n4041 , n4039 , n4040 );
xnor ( n4042 , n4041 , n1199 );
xor ( n4043 , n4017 , n4019 );
xor ( n4044 , n4043 , n4006 );
and ( n4045 , n4042 , n4044 );
and ( n4046 , n3397 , n3434 );
not ( n4047 , n4046 );
or ( n4048 , n4015 , n4047 );
and ( n4049 , n4044 , n4048 );
and ( n4050 , n4042 , n4048 );
or ( n4051 , n4045 , n4049 , n4050 );
and ( n4052 , n4038 , n4051 );
xor ( n4053 , n4014 , n4023 );
xor ( n4054 , n4053 , n4026 );
and ( n4055 , n4051 , n4054 );
and ( n4056 , n4038 , n4054 );
or ( n4057 , n4052 , n4055 , n4056 );
or ( n4058 , n4037 , n4057 );
and ( n4059 , n4034 , n4058 );
and ( n4060 , n4032 , n4058 );
or ( n4061 , n4035 , n4059 , n4060 );
and ( n4062 , n4003 , n4061 );
xor ( n4063 , n4003 , n4061 );
xor ( n4064 , n4032 , n4034 );
xor ( n4065 , n4064 , n4058 );
not ( n4066 , n4065 );
xor ( n4067 , n4005 , n4011 );
xor ( n4068 , n4067 , n4029 );
xnor ( n4069 , n4037 , n4057 );
and ( n4070 , n4068 , n4069 );
and ( n4071 , n4066 , n4070 );
or ( n4072 , n4065 , n4071 );
and ( n4073 , n4063 , n4072 );
or ( n4074 , n4062 , n4073 );
and ( n4075 , n4001 , n4074 );
or ( n4076 , n4000 , n4075 );
and ( n4077 , n3996 , n4076 );
or ( n4078 , n3995 , n4077 );
and ( n4079 , n3955 , n4078 );
or ( n4080 , n3954 , n4079 );
and ( n4081 , n3950 , n4080 );
or ( n4082 , n3949 , n4081 );
and ( n4083 , n3947 , n4082 );
or ( n4084 , n3946 , n4083 );
and ( n4085 , n3944 , n4084 );
or ( n4086 , n3943 , n4085 );
and ( n4087 , n3941 , n4086 );
or ( n4088 , n3940 , n4087 );
and ( n4089 , n3938 , n4088 );
and ( n4090 , n3936 , n4089 );
and ( n4091 , n3935 , n4090 );
and ( n4092 , n3934 , n4091 );
and ( n4093 , n3932 , n4092 );
and ( n4094 , n3931 , n4093 );
and ( n4095 , n3930 , n4094 );
and ( n4096 , n3929 , n4095 );
and ( n4097 , n3928 , n4096 );
and ( n4098 , n3927 , n4097 );
and ( n4099 , n3926 , n4098 );
and ( n4100 , n3925 , n4099 );
and ( n4101 , n3924 , n4100 );
and ( n4102 , n3923 , n4101 );
and ( n4103 , n3922 , n4102 );
and ( n4104 , n3921 , n4103 );
and ( n4105 , n3920 , n4104 );
and ( n4106 , n3919 , n4105 );
and ( n4107 , n3918 , n4106 );
and ( n4108 , n3917 , n4107 );
and ( n4109 , n3916 , n4108 );
and ( n4110 , n3915 , n4109 );
and ( n4111 , n3914 , n4110 );
and ( n4112 , n3913 , n4111 );
and ( n4113 , n3912 , n4112 );
and ( n4114 , n3911 , n4113 );
and ( n4115 , n3910 , n4114 );
and ( n4116 , n3909 , n4115 );
and ( n4117 , n3908 , n4116 );
and ( n4118 , n3907 , n4117 );
and ( n4119 , n3906 , n4118 );
and ( n4120 , n3905 , n4119 );
and ( n4121 , n3904 , n4120 );
and ( n4122 , n3903 , n4121 );
and ( n4123 , n3902 , n4122 );
and ( n4124 , n3901 , n4123 );
and ( n4125 , n3900 , n4124 );
and ( n4126 , n3899 , n4125 );
and ( n4127 , n3898 , n4126 );
and ( n4128 , n3897 , n4127 );
and ( n4129 , n3896 , n4128 );
and ( n4130 , n3895 , n4129 );
and ( n4131 , n3894 , n4130 );
and ( n4132 , n3893 , n4131 );
and ( n4133 , n3892 , n4132 );
and ( n4134 , n3891 , n4133 );
or ( n4135 , n3890 , n4134 );
and ( n4136 , n3888 , n4135 );
and ( n4137 , n3887 , n4136 );
and ( n4138 , n3886 , n4137 );
or ( n4139 , n3885 , n4138 );
and ( n4140 , n1401 , n4139 );
or ( n4141 , n1400 , n4140 );
xor ( n4142 , n1260 , n4141 );
buf ( n4143 , n4142 );
xor ( n4144 , n1401 , n4139 );
buf ( n4145 , n4144 );
xor ( n4146 , n3886 , n4137 );
buf ( n4147 , n4146 );
xor ( n4148 , n3887 , n4136 );
buf ( n4149 , n4148 );
xor ( n4150 , n3888 , n4135 );
buf ( n4151 , n4150 );
xor ( n4152 , n3891 , n4133 );
buf ( n4153 , n4152 );
xor ( n4154 , n3892 , n4132 );
buf ( n4155 , n4154 );
xor ( n4156 , n3893 , n4131 );
buf ( n4157 , n4156 );
xor ( n4158 , n3894 , n4130 );
buf ( n4159 , n4158 );
xor ( n4160 , n3895 , n4129 );
buf ( n4161 , n4160 );
xor ( n4162 , n3896 , n4128 );
buf ( n4163 , n4162 );
xor ( n4164 , n3897 , n4127 );
buf ( n4165 , n4164 );
xor ( n4166 , n3898 , n4126 );
buf ( n4167 , n4166 );
xor ( n4168 , n3899 , n4125 );
buf ( n4169 , n4168 );
xor ( n4170 , n3900 , n4124 );
buf ( n4171 , n4170 );
xor ( n4172 , n3901 , n4123 );
buf ( n4173 , n4172 );
xor ( n4174 , n3902 , n4122 );
buf ( n4175 , n4174 );
xor ( n4176 , n3903 , n4121 );
buf ( n4177 , n4176 );
xor ( n4178 , n3904 , n4120 );
buf ( n4179 , n4178 );
xor ( n4180 , n3905 , n4119 );
buf ( n4181 , n4180 );
xor ( n4182 , n3906 , n4118 );
buf ( n4183 , n4182 );
xor ( n4184 , n3907 , n4117 );
buf ( n4185 , n4184 );
xor ( n4186 , n3908 , n4116 );
buf ( n4187 , n4186 );
xor ( n4188 , n3909 , n4115 );
buf ( n4189 , n4188 );
xor ( n4190 , n3910 , n4114 );
buf ( n4191 , n4190 );
xor ( n4192 , n3911 , n4113 );
buf ( n4193 , n4192 );
xor ( n4194 , n3912 , n4112 );
buf ( n4195 , n4194 );
xor ( n4196 , n3913 , n4111 );
buf ( n4197 , n4196 );
xor ( n4198 , n3914 , n4110 );
buf ( n4199 , n4198 );
xor ( n4200 , n3915 , n4109 );
buf ( n4201 , n4200 );
xor ( n4202 , n3916 , n4108 );
buf ( n4203 , n4202 );
xor ( n4204 , n3917 , n4107 );
buf ( n4205 , n4204 );
xor ( n4206 , n3918 , n4106 );
buf ( n4207 , n4206 );
xor ( n4208 , n3919 , n4105 );
buf ( n4209 , n4208 );
xor ( n4210 , n3920 , n4104 );
buf ( n4211 , n4210 );
xor ( n4212 , n3921 , n4103 );
buf ( n4213 , n4212 );
xor ( n4214 , n3922 , n4102 );
buf ( n4215 , n4214 );
xor ( n4216 , n3923 , n4101 );
buf ( n4217 , n4216 );
xor ( n4218 , n3924 , n4100 );
buf ( n4219 , n4218 );
xor ( n4220 , n3925 , n4099 );
buf ( n4221 , n4220 );
xor ( n4222 , n3926 , n4098 );
buf ( n4223 , n4222 );
xor ( n4224 , n3927 , n4097 );
buf ( n4225 , n4224 );
xor ( n4226 , n3928 , n4096 );
buf ( n4227 , n4226 );
xor ( n4228 , n3929 , n4095 );
buf ( n4229 , n4228 );
xor ( n4230 , n3930 , n4094 );
buf ( n4231 , n4230 );
xor ( n4232 , n3931 , n4093 );
buf ( n4233 , n4232 );
xor ( n4234 , n3932 , n4092 );
buf ( n4235 , n4234 );
xor ( n4236 , n3934 , n4091 );
buf ( n4237 , n4236 );
xor ( n4238 , n3935 , n4090 );
buf ( n4239 , n4238 );
xor ( n4240 , n3936 , n4089 );
buf ( n4241 , n4240 );
xor ( n4242 , n3938 , n4088 );
buf ( n4243 , n4242 );
xor ( n4244 , n3941 , n4086 );
buf ( n4245 , n4244 );
xor ( n4246 , n3944 , n4084 );
buf ( n4247 , n4246 );
xor ( n4248 , n3947 , n4082 );
buf ( n4249 , n4248 );
xor ( n4250 , n3950 , n4080 );
buf ( n4251 , n4250 );
xor ( n4252 , n3955 , n4078 );
buf ( n4253 , n4252 );
xor ( n4254 , n3996 , n4076 );
buf ( n4255 , n4254 );
xor ( n4256 , n4001 , n4074 );
buf ( n4257 , n4256 );
xor ( n4258 , n4063 , n4072 );
buf ( n4259 , n4258 );
xor ( n4260 , n4066 , n4070 );
buf ( n4261 , n4260 );
xor ( n4262 , n4068 , n4069 );
buf ( n4263 , n4262 );
xor ( n4264 , n4038 , n4051 );
xor ( n4265 , n4264 , n4054 );
buf ( n4266 , n4265 );
xor ( n4267 , n4042 , n4044 );
xor ( n4268 , n4267 , n4048 );
buf ( n4269 , n4268 );
xnor ( n4270 , n4015 , n4047 );
buf ( n4271 , n4270 );
buf ( n4272 , n387 );
buf ( n4273 , n4272 );
buf ( n4274 , n386 );
buf ( n4275 , n4274 );
and ( n4276 , n4273 , n4275 );
buf ( n4277 , n386 );
buf ( n4278 , n4277 );
buf ( n4279 , n4278 );
and ( n4280 , n4276 , n4279 );
buf ( n4281 , n388 );
buf ( n4282 , n4281 );
and ( n4283 , n4282 , n4275 );
buf ( n4284 , n389 );
buf ( n4285 , n4284 );
and ( n4286 , n4285 , n4275 );
buf ( n4287 , n387 );
buf ( n4288 , n4287 );
and ( n4289 , n4282 , n4288 );
and ( n4290 , n4286 , n4289 );
buf ( n4291 , n4273 );
and ( n4292 , n4289 , n4291 );
and ( n4293 , n4286 , n4291 );
or ( n4294 , n4290 , n4292 , n4293 );
and ( n4295 , n4283 , n4294 );
xor ( n4296 , n4286 , n4289 );
xor ( n4297 , n4296 , n4291 );
buf ( n4298 , n391 );
buf ( n4299 , n4298 );
and ( n4300 , n4299 , n4275 );
buf ( n4301 , n388 );
buf ( n4302 , n4301 );
and ( n4303 , n4285 , n4302 );
and ( n4304 , n4300 , n4303 );
buf ( n4305 , n4282 );
and ( n4306 , n4303 , n4305 );
and ( n4307 , n4300 , n4305 );
or ( n4308 , n4304 , n4306 , n4307 );
buf ( n4309 , n390 );
buf ( n4310 , n4309 );
and ( n4311 , n4310 , n4275 );
and ( n4312 , n4308 , n4311 );
and ( n4313 , n4285 , n4288 );
and ( n4314 , n4311 , n4313 );
and ( n4315 , n4308 , n4313 );
or ( n4316 , n4312 , n4314 , n4315 );
and ( n4317 , n4297 , n4316 );
xor ( n4318 , n4308 , n4311 );
xor ( n4319 , n4318 , n4313 );
buf ( n4320 , n392 );
buf ( n4321 , n4320 );
and ( n4322 , n4321 , n4275 );
and ( n4323 , n4299 , n4288 );
and ( n4324 , n4322 , n4323 );
and ( n4325 , n4310 , n4302 );
and ( n4326 , n4323 , n4325 );
and ( n4327 , n4322 , n4325 );
or ( n4328 , n4324 , n4326 , n4327 );
and ( n4329 , n4310 , n4288 );
and ( n4330 , n4328 , n4329 );
xor ( n4331 , n4300 , n4303 );
xor ( n4332 , n4331 , n4305 );
and ( n4333 , n4329 , n4332 );
and ( n4334 , n4328 , n4332 );
or ( n4335 , n4330 , n4333 , n4334 );
and ( n4336 , n4319 , n4335 );
xor ( n4337 , n4328 , n4329 );
xor ( n4338 , n4337 , n4332 );
buf ( n4339 , n393 );
buf ( n4340 , n4339 );
and ( n4341 , n4340 , n4275 );
and ( n4342 , n4321 , n4288 );
and ( n4343 , n4341 , n4342 );
and ( n4344 , n4299 , n4302 );
and ( n4345 , n4342 , n4344 );
and ( n4346 , n4341 , n4344 );
or ( n4347 , n4343 , n4345 , n4346 );
buf ( n4348 , n389 );
buf ( n4349 , n4348 );
and ( n4350 , n4310 , n4349 );
buf ( n4351 , n4285 );
and ( n4352 , n4350 , n4351 );
and ( n4353 , n4347 , n4352 );
xor ( n4354 , n4322 , n4323 );
xor ( n4355 , n4354 , n4325 );
and ( n4356 , n4352 , n4355 );
and ( n4357 , n4347 , n4355 );
or ( n4358 , n4353 , n4356 , n4357 );
and ( n4359 , n4338 , n4358 );
xor ( n4360 , n4347 , n4352 );
xor ( n4361 , n4360 , n4355 );
xor ( n4362 , n4350 , n4351 );
and ( n4363 , n4321 , n4302 );
and ( n4364 , n4299 , n4349 );
and ( n4365 , n4363 , n4364 );
and ( n4366 , n4362 , n4365 );
xor ( n4367 , n4341 , n4342 );
xor ( n4368 , n4367 , n4344 );
and ( n4369 , n4365 , n4368 );
and ( n4370 , n4362 , n4368 );
or ( n4371 , n4366 , n4369 , n4370 );
and ( n4372 , n4361 , n4371 );
xor ( n4373 , n4362 , n4365 );
xor ( n4374 , n4373 , n4368 );
and ( n4375 , n4340 , n4288 );
xor ( n4376 , n4363 , n4364 );
and ( n4377 , n4375 , n4376 );
and ( n4378 , n4374 , n4377 );
and ( n4379 , n4340 , n4302 );
and ( n4380 , n4321 , n4349 );
and ( n4381 , n4379 , n4380 );
xor ( n4382 , n4375 , n4376 );
and ( n4383 , n4381 , n4382 );
buf ( n4384 , n390 );
buf ( n4385 , n4384 );
and ( n4386 , n4299 , n4385 );
buf ( n4387 , n4310 );
and ( n4388 , n4386 , n4387 );
xor ( n4389 , n4379 , n4380 );
and ( n4390 , n4387 , n4389 );
and ( n4391 , n4386 , n4389 );
or ( n4392 , n4388 , n4390 , n4391 );
and ( n4393 , n4382 , n4392 );
and ( n4394 , n4381 , n4392 );
or ( n4395 , n4383 , n4393 , n4394 );
and ( n4396 , n4377 , n4395 );
and ( n4397 , n4374 , n4395 );
or ( n4398 , n4378 , n4396 , n4397 );
and ( n4399 , n4371 , n4398 );
and ( n4400 , n4361 , n4398 );
or ( n4401 , n4372 , n4399 , n4400 );
and ( n4402 , n4358 , n4401 );
and ( n4403 , n4338 , n4401 );
or ( n4404 , n4359 , n4402 , n4403 );
and ( n4405 , n4335 , n4404 );
and ( n4406 , n4319 , n4404 );
or ( n4407 , n4336 , n4405 , n4406 );
and ( n4408 , n4316 , n4407 );
and ( n4409 , n4297 , n4407 );
or ( n4410 , n4317 , n4408 , n4409 );
and ( n4411 , n4294 , n4410 );
and ( n4412 , n4283 , n4410 );
or ( n4413 , n4295 , n4411 , n4412 );
and ( n4414 , n4279 , n4413 );
and ( n4415 , n4276 , n4413 );
or ( n4416 , n4280 , n4414 , n4415 );
xor ( n4417 , n4276 , n4279 );
xor ( n4418 , n4417 , n4413 );
xor ( n4419 , n4283 , n4294 );
xor ( n4420 , n4419 , n4410 );
xor ( n4421 , n4297 , n4316 );
xor ( n4422 , n4421 , n4407 );
xor ( n4423 , n4319 , n4335 );
xor ( n4424 , n4423 , n4404 );
xor ( n4425 , n4338 , n4358 );
xor ( n4426 , n4425 , n4401 );
xor ( n4427 , n4361 , n4371 );
xor ( n4428 , n4427 , n4398 );
xor ( n4429 , n4374 , n4377 );
xor ( n4430 , n4429 , n4395 );
xor ( n4431 , n4381 , n4382 );
xor ( n4432 , n4431 , n4392 );
and ( n4433 , n4340 , n4349 );
and ( n4434 , n4321 , n4385 );
and ( n4435 , n4433 , n4434 );
xor ( n4436 , n4386 , n4387 );
xor ( n4437 , n4436 , n4389 );
and ( n4438 , n4435 , n4437 );
xor ( n4439 , n4435 , n4437 );
xor ( n4440 , n4433 , n4434 );
and ( n4441 , n4340 , n4385 );
buf ( n4442 , n4299 );
and ( n4443 , n4441 , n4442 );
and ( n4444 , n4440 , n4443 );
xor ( n4445 , n4440 , n4443 );
buf ( n4446 , n391 );
buf ( n4447 , n4446 );
and ( n4448 , n4321 , n4447 );
xor ( n4449 , n4441 , n4442 );
and ( n4450 , n4448 , n4449 );
xor ( n4451 , n4448 , n4449 );
and ( n4452 , n4340 , n4447 );
buf ( n4453 , n392 );
buf ( n4454 , n4453 );
and ( n4455 , n4340 , n4454 );
buf ( n4456 , n4321 );
and ( n4457 , n4455 , n4456 );
and ( n4458 , n4452 , n4457 );
and ( n4459 , n4451 , n4458 );
or ( n4460 , n4450 , n4459 );
and ( n4461 , n4445 , n4460 );
or ( n4462 , n4444 , n4461 );
and ( n4463 , n4439 , n4462 );
or ( n4464 , n4438 , n4463 );
and ( n4465 , n4432 , n4464 );
and ( n4466 , n4430 , n4465 );
and ( n4467 , n4428 , n4466 );
and ( n4468 , n4426 , n4467 );
and ( n4469 , n4424 , n4468 );
and ( n4470 , n4422 , n4469 );
and ( n4471 , n4420 , n4470 );
and ( n4472 , n4418 , n4471 );
xor ( n4473 , n4416 , n4472 );
buf ( n4474 , n4473 );
and ( n4475 , n4474 , n392 );
buf ( n4476 , n4475 );
and ( n4477 , n4474 , n393 );
xor ( n4478 , n4418 , n4471 );
buf ( n4479 , n4478 );
and ( n4480 , n4479 , n392 );
and ( n4481 , n4477 , n4480 );
xor ( n4482 , n4477 , n4480 );
and ( n4483 , n4479 , n393 );
xor ( n4484 , n4420 , n4470 );
buf ( n4485 , n4484 );
and ( n4486 , n4485 , n392 );
and ( n4487 , n4483 , n4486 );
xor ( n4488 , n4483 , n4486 );
and ( n4489 , n4485 , n393 );
xor ( n4490 , n4422 , n4469 );
buf ( n4491 , n4490 );
and ( n4492 , n4491 , n392 );
and ( n4493 , n4489 , n4492 );
xor ( n4494 , n4489 , n4492 );
and ( n4495 , n4491 , n393 );
xor ( n4496 , n4424 , n4468 );
buf ( n4497 , n4496 );
and ( n4498 , n4497 , n392 );
and ( n4499 , n4495 , n4498 );
xor ( n4500 , n4495 , n4498 );
and ( n4501 , n4497 , n393 );
xor ( n4502 , n4426 , n4467 );
buf ( n4503 , n4502 );
and ( n4504 , n4503 , n392 );
and ( n4505 , n4501 , n4504 );
xor ( n4506 , n4501 , n4504 );
and ( n4507 , n4503 , n393 );
xor ( n4508 , n4428 , n4466 );
buf ( n4509 , n4508 );
and ( n4510 , n4509 , n392 );
and ( n4511 , n4507 , n4510 );
xor ( n4512 , n4507 , n4510 );
and ( n4513 , n4509 , n393 );
xor ( n4514 , n4430 , n4465 );
buf ( n4515 , n4514 );
and ( n4516 , n4515 , n392 );
and ( n4517 , n4513 , n4516 );
xor ( n4518 , n4513 , n4516 );
and ( n4519 , n4515 , n393 );
xor ( n4520 , n4432 , n4464 );
buf ( n4521 , n4520 );
and ( n4522 , n4521 , n392 );
and ( n4523 , n4519 , n4522 );
xor ( n4524 , n4519 , n4522 );
and ( n4525 , n4521 , n393 );
xor ( n4526 , n4439 , n4462 );
buf ( n4527 , n4526 );
and ( n4528 , n4527 , n392 );
and ( n4529 , n4525 , n4528 );
xor ( n4530 , n4525 , n4528 );
and ( n4531 , n4527 , n393 );
xor ( n4532 , n4445 , n4460 );
buf ( n4533 , n4532 );
and ( n4534 , n4533 , n392 );
and ( n4535 , n4531 , n4534 );
xor ( n4536 , n4531 , n4534 );
and ( n4537 , n4533 , n393 );
xor ( n4538 , n4451 , n4458 );
buf ( n4539 , n4538 );
and ( n4540 , n4539 , n392 );
and ( n4541 , n4537 , n4540 );
xor ( n4542 , n4537 , n4540 );
and ( n4543 , n4539 , n393 );
xor ( n4544 , n4452 , n4457 );
buf ( n4545 , n4544 );
and ( n4546 , n4545 , n392 );
and ( n4547 , n4543 , n4546 );
xor ( n4548 , n4543 , n4546 );
and ( n4549 , n4545 , n393 );
xor ( n4550 , n4455 , n4456 );
buf ( n4551 , n4550 );
and ( n4552 , n4551 , n392 );
and ( n4553 , n4549 , n4552 );
buf ( n4554 , n4553 );
and ( n4555 , n4548 , n4554 );
or ( n4556 , n4547 , n4555 );
and ( n4557 , n4542 , n4556 );
or ( n4558 , n4541 , n4557 );
and ( n4559 , n4536 , n4558 );
or ( n4560 , n4535 , n4559 );
and ( n4561 , n4530 , n4560 );
or ( n4562 , n4529 , n4561 );
and ( n4563 , n4524 , n4562 );
or ( n4564 , n4523 , n4563 );
and ( n4565 , n4518 , n4564 );
or ( n4566 , n4517 , n4565 );
and ( n4567 , n4512 , n4566 );
or ( n4568 , n4511 , n4567 );
and ( n4569 , n4506 , n4568 );
or ( n4570 , n4505 , n4569 );
and ( n4571 , n4500 , n4570 );
or ( n4572 , n4499 , n4571 );
and ( n4573 , n4494 , n4572 );
or ( n4574 , n4493 , n4573 );
and ( n4575 , n4488 , n4574 );
or ( n4576 , n4487 , n4575 );
and ( n4577 , n4482 , n4576 );
or ( n4578 , n4481 , n4577 );
and ( n4579 , n4476 , n4578 );
buf ( n4580 , n4579 );
buf ( n4581 , n4580 );
and ( n4582 , n4474 , n391 );
and ( n4583 , n4581 , n4582 );
xor ( n4584 , n4581 , n4582 );
xor ( n4585 , n4476 , n4578 );
and ( n4586 , n4479 , n391 );
and ( n4587 , n4585 , n4586 );
xor ( n4588 , n4585 , n4586 );
xor ( n4589 , n4482 , n4576 );
and ( n4590 , n4485 , n391 );
and ( n4591 , n4589 , n4590 );
xor ( n4592 , n4589 , n4590 );
xor ( n4593 , n4488 , n4574 );
and ( n4594 , n4491 , n391 );
and ( n4595 , n4593 , n4594 );
xor ( n4596 , n4593 , n4594 );
xor ( n4597 , n4494 , n4572 );
and ( n4598 , n4497 , n391 );
and ( n4599 , n4597 , n4598 );
xor ( n4600 , n4597 , n4598 );
xor ( n4601 , n4500 , n4570 );
and ( n4602 , n4503 , n391 );
and ( n4603 , n4601 , n4602 );
xor ( n4604 , n4601 , n4602 );
xor ( n4605 , n4506 , n4568 );
and ( n4606 , n4509 , n391 );
and ( n4607 , n4605 , n4606 );
xor ( n4608 , n4605 , n4606 );
xor ( n4609 , n4512 , n4566 );
and ( n4610 , n4515 , n391 );
and ( n4611 , n4609 , n4610 );
xor ( n4612 , n4609 , n4610 );
xor ( n4613 , n4518 , n4564 );
and ( n4614 , n4521 , n391 );
and ( n4615 , n4613 , n4614 );
xor ( n4616 , n4613 , n4614 );
xor ( n4617 , n4524 , n4562 );
and ( n4618 , n4527 , n391 );
and ( n4619 , n4617 , n4618 );
xor ( n4620 , n4617 , n4618 );
xor ( n4621 , n4530 , n4560 );
and ( n4622 , n4533 , n391 );
and ( n4623 , n4621 , n4622 );
xor ( n4624 , n4621 , n4622 );
xor ( n4625 , n4536 , n4558 );
and ( n4626 , n4539 , n391 );
and ( n4627 , n4625 , n4626 );
xor ( n4628 , n4625 , n4626 );
xor ( n4629 , n4542 , n4556 );
and ( n4630 , n4545 , n391 );
and ( n4631 , n4629 , n4630 );
xor ( n4632 , n4629 , n4630 );
xor ( n4633 , n4548 , n4554 );
and ( n4634 , n4551 , n391 );
and ( n4635 , n4633 , n4634 );
xor ( n4636 , n4633 , n4634 );
xor ( n4637 , n4549 , n4552 );
buf ( n4638 , n4637 );
buf ( n4639 , n4638 );
and ( n4640 , n4551 , n393 );
buf ( n4641 , n4640 );
buf ( n4642 , n4641 );
buf ( n4643 , n4340 );
buf ( n4644 , n4643 );
and ( n4645 , n4644 , n391 );
and ( n4646 , n4642 , n4645 );
and ( n4647 , n4639 , n4646 );
buf ( n4648 , n4647 );
and ( n4649 , n4636 , n4648 );
or ( n4650 , n4635 , n4649 );
and ( n4651 , n4632 , n4650 );
or ( n4652 , n4631 , n4651 );
and ( n4653 , n4628 , n4652 );
or ( n4654 , n4627 , n4653 );
and ( n4655 , n4624 , n4654 );
or ( n4656 , n4623 , n4655 );
and ( n4657 , n4620 , n4656 );
or ( n4658 , n4619 , n4657 );
and ( n4659 , n4616 , n4658 );
or ( n4660 , n4615 , n4659 );
and ( n4661 , n4612 , n4660 );
or ( n4662 , n4611 , n4661 );
and ( n4663 , n4608 , n4662 );
or ( n4664 , n4607 , n4663 );
and ( n4665 , n4604 , n4664 );
or ( n4666 , n4603 , n4665 );
and ( n4667 , n4600 , n4666 );
or ( n4668 , n4599 , n4667 );
and ( n4669 , n4596 , n4668 );
or ( n4670 , n4595 , n4669 );
and ( n4671 , n4592 , n4670 );
or ( n4672 , n4591 , n4671 );
and ( n4673 , n4588 , n4672 );
or ( n4674 , n4587 , n4673 );
and ( n4675 , n4584 , n4674 );
or ( n4676 , n4583 , n4675 );
buf ( n4677 , n4676 );
and ( n4678 , n4474 , n390 );
and ( n4679 , n4677 , n4678 );
xor ( n4680 , n4677 , n4678 );
xor ( n4681 , n4584 , n4674 );
and ( n4682 , n4479 , n390 );
and ( n4683 , n4681 , n4682 );
xor ( n4684 , n4681 , n4682 );
xor ( n4685 , n4588 , n4672 );
and ( n4686 , n4485 , n390 );
and ( n4687 , n4685 , n4686 );
xor ( n4688 , n4685 , n4686 );
xor ( n4689 , n4592 , n4670 );
and ( n4690 , n4491 , n390 );
and ( n4691 , n4689 , n4690 );
xor ( n4692 , n4689 , n4690 );
xor ( n4693 , n4596 , n4668 );
and ( n4694 , n4497 , n390 );
and ( n4695 , n4693 , n4694 );
xor ( n4696 , n4693 , n4694 );
xor ( n4697 , n4600 , n4666 );
and ( n4698 , n4503 , n390 );
and ( n4699 , n4697 , n4698 );
xor ( n4700 , n4697 , n4698 );
xor ( n4701 , n4604 , n4664 );
and ( n4702 , n4509 , n390 );
and ( n4703 , n4701 , n4702 );
xor ( n4704 , n4701 , n4702 );
xor ( n4705 , n4608 , n4662 );
and ( n4706 , n4515 , n390 );
and ( n4707 , n4705 , n4706 );
xor ( n4708 , n4705 , n4706 );
xor ( n4709 , n4612 , n4660 );
and ( n4710 , n4521 , n390 );
and ( n4711 , n4709 , n4710 );
xor ( n4712 , n4709 , n4710 );
xor ( n4713 , n4616 , n4658 );
and ( n4714 , n4527 , n390 );
and ( n4715 , n4713 , n4714 );
xor ( n4716 , n4713 , n4714 );
xor ( n4717 , n4620 , n4656 );
and ( n4718 , n4533 , n390 );
and ( n4719 , n4717 , n4718 );
xor ( n4720 , n4717 , n4718 );
xor ( n4721 , n4624 , n4654 );
and ( n4722 , n4539 , n390 );
and ( n4723 , n4721 , n4722 );
xor ( n4724 , n4721 , n4722 );
xor ( n4725 , n4628 , n4652 );
and ( n4726 , n4545 , n390 );
and ( n4727 , n4725 , n4726 );
xor ( n4728 , n4725 , n4726 );
xor ( n4729 , n4632 , n4650 );
and ( n4730 , n4551 , n390 );
and ( n4731 , n4729 , n4730 );
xor ( n4732 , n4729 , n4730 );
xor ( n4733 , n4636 , n4648 );
buf ( n4734 , n4733 );
xor ( n4735 , n4639 , n4646 );
and ( n4736 , n4644 , n390 );
and ( n4737 , n4735 , n4736 );
and ( n4738 , n4734 , n4737 );
buf ( n4739 , n4738 );
and ( n4740 , n4732 , n4739 );
or ( n4741 , n4731 , n4740 );
and ( n4742 , n4728 , n4741 );
or ( n4743 , n4727 , n4742 );
and ( n4744 , n4724 , n4743 );
or ( n4745 , n4723 , n4744 );
and ( n4746 , n4720 , n4745 );
or ( n4747 , n4719 , n4746 );
and ( n4748 , n4716 , n4747 );
or ( n4749 , n4715 , n4748 );
and ( n4750 , n4712 , n4749 );
or ( n4751 , n4711 , n4750 );
and ( n4752 , n4708 , n4751 );
or ( n4753 , n4707 , n4752 );
and ( n4754 , n4704 , n4753 );
or ( n4755 , n4703 , n4754 );
and ( n4756 , n4700 , n4755 );
or ( n4757 , n4699 , n4756 );
and ( n4758 , n4696 , n4757 );
or ( n4759 , n4695 , n4758 );
and ( n4760 , n4692 , n4759 );
or ( n4761 , n4691 , n4760 );
and ( n4762 , n4688 , n4761 );
or ( n4763 , n4687 , n4762 );
and ( n4764 , n4684 , n4763 );
or ( n4765 , n4683 , n4764 );
and ( n4766 , n4680 , n4765 );
or ( n4767 , n4679 , n4766 );
buf ( n4768 , n4767 );
and ( n4769 , n4474 , n389 );
and ( n4770 , n4768 , n4769 );
xor ( n4771 , n4768 , n4769 );
xor ( n4772 , n4680 , n4765 );
and ( n4773 , n4479 , n389 );
and ( n4774 , n4772 , n4773 );
xor ( n4775 , n4772 , n4773 );
xor ( n4776 , n4684 , n4763 );
and ( n4777 , n4485 , n389 );
and ( n4778 , n4776 , n4777 );
xor ( n4779 , n4776 , n4777 );
xor ( n4780 , n4688 , n4761 );
and ( n4781 , n4491 , n389 );
and ( n4782 , n4780 , n4781 );
xor ( n4783 , n4780 , n4781 );
xor ( n4784 , n4692 , n4759 );
and ( n4785 , n4497 , n389 );
and ( n4786 , n4784 , n4785 );
xor ( n4787 , n4784 , n4785 );
xor ( n4788 , n4696 , n4757 );
and ( n4789 , n4503 , n389 );
and ( n4790 , n4788 , n4789 );
xor ( n4791 , n4788 , n4789 );
xor ( n4792 , n4700 , n4755 );
and ( n4793 , n4509 , n389 );
and ( n4794 , n4792 , n4793 );
xor ( n4795 , n4792 , n4793 );
xor ( n4796 , n4704 , n4753 );
and ( n4797 , n4515 , n389 );
and ( n4798 , n4796 , n4797 );
xor ( n4799 , n4796 , n4797 );
xor ( n4800 , n4708 , n4751 );
and ( n4801 , n4521 , n389 );
and ( n4802 , n4800 , n4801 );
xor ( n4803 , n4800 , n4801 );
xor ( n4804 , n4712 , n4749 );
and ( n4805 , n4527 , n389 );
and ( n4806 , n4804 , n4805 );
xor ( n4807 , n4804 , n4805 );
xor ( n4808 , n4716 , n4747 );
and ( n4809 , n4533 , n389 );
and ( n4810 , n4808 , n4809 );
xor ( n4811 , n4808 , n4809 );
xor ( n4812 , n4720 , n4745 );
and ( n4813 , n4539 , n389 );
and ( n4814 , n4812 , n4813 );
xor ( n4815 , n4812 , n4813 );
xor ( n4816 , n4724 , n4743 );
and ( n4817 , n4545 , n389 );
and ( n4818 , n4816 , n4817 );
xor ( n4819 , n4816 , n4817 );
xor ( n4820 , n4728 , n4741 );
and ( n4821 , n4551 , n389 );
and ( n4822 , n4820 , n4821 );
xor ( n4823 , n4820 , n4821 );
xor ( n4824 , n4732 , n4739 );
buf ( n4825 , n4824 );
xor ( n4826 , n4734 , n4737 );
and ( n4827 , n4644 , n389 );
and ( n4828 , n4826 , n4827 );
and ( n4829 , n4825 , n4828 );
buf ( n4830 , n4829 );
and ( n4831 , n4823 , n4830 );
or ( n4832 , n4822 , n4831 );
and ( n4833 , n4819 , n4832 );
or ( n4834 , n4818 , n4833 );
and ( n4835 , n4815 , n4834 );
or ( n4836 , n4814 , n4835 );
and ( n4837 , n4811 , n4836 );
or ( n4838 , n4810 , n4837 );
and ( n4839 , n4807 , n4838 );
or ( n4840 , n4806 , n4839 );
and ( n4841 , n4803 , n4840 );
or ( n4842 , n4802 , n4841 );
and ( n4843 , n4799 , n4842 );
or ( n4844 , n4798 , n4843 );
and ( n4845 , n4795 , n4844 );
or ( n4846 , n4794 , n4845 );
and ( n4847 , n4791 , n4846 );
or ( n4848 , n4790 , n4847 );
and ( n4849 , n4787 , n4848 );
or ( n4850 , n4786 , n4849 );
and ( n4851 , n4783 , n4850 );
or ( n4852 , n4782 , n4851 );
and ( n4853 , n4779 , n4852 );
or ( n4854 , n4778 , n4853 );
and ( n4855 , n4775 , n4854 );
or ( n4856 , n4774 , n4855 );
and ( n4857 , n4771 , n4856 );
or ( n4858 , n4770 , n4857 );
buf ( n4859 , n4858 );
and ( n4860 , n4474 , n388 );
and ( n4861 , n4859 , n4860 );
xor ( n4862 , n4859 , n4860 );
xor ( n4863 , n4771 , n4856 );
and ( n4864 , n4479 , n388 );
and ( n4865 , n4863 , n4864 );
xor ( n4866 , n4863 , n4864 );
xor ( n4867 , n4775 , n4854 );
and ( n4868 , n4485 , n388 );
and ( n4869 , n4867 , n4868 );
xor ( n4870 , n4867 , n4868 );
xor ( n4871 , n4779 , n4852 );
and ( n4872 , n4491 , n388 );
and ( n4873 , n4871 , n4872 );
xor ( n4874 , n4871 , n4872 );
xor ( n4875 , n4783 , n4850 );
and ( n4876 , n4497 , n388 );
and ( n4877 , n4875 , n4876 );
xor ( n4878 , n4875 , n4876 );
xor ( n4879 , n4787 , n4848 );
and ( n4880 , n4503 , n388 );
and ( n4881 , n4879 , n4880 );
xor ( n4882 , n4879 , n4880 );
xor ( n4883 , n4791 , n4846 );
and ( n4884 , n4509 , n388 );
and ( n4885 , n4883 , n4884 );
xor ( n4886 , n4883 , n4884 );
xor ( n4887 , n4795 , n4844 );
and ( n4888 , n4515 , n388 );
and ( n4889 , n4887 , n4888 );
xor ( n4890 , n4887 , n4888 );
xor ( n4891 , n4799 , n4842 );
and ( n4892 , n4521 , n388 );
and ( n4893 , n4891 , n4892 );
xor ( n4894 , n4891 , n4892 );
xor ( n4895 , n4803 , n4840 );
and ( n4896 , n4527 , n388 );
and ( n4897 , n4895 , n4896 );
xor ( n4898 , n4895 , n4896 );
xor ( n4899 , n4807 , n4838 );
and ( n4900 , n4533 , n388 );
and ( n4901 , n4899 , n4900 );
xor ( n4902 , n4899 , n4900 );
xor ( n4903 , n4811 , n4836 );
and ( n4904 , n4539 , n388 );
and ( n4905 , n4903 , n4904 );
xor ( n4906 , n4903 , n4904 );
xor ( n4907 , n4815 , n4834 );
and ( n4908 , n4545 , n388 );
and ( n4909 , n4907 , n4908 );
xor ( n4910 , n4907 , n4908 );
xor ( n4911 , n4819 , n4832 );
and ( n4912 , n4551 , n388 );
and ( n4913 , n4911 , n4912 );
xor ( n4914 , n4911 , n4912 );
xor ( n4915 , n4823 , n4830 );
buf ( n4916 , n4915 );
xor ( n4917 , n4825 , n4828 );
and ( n4918 , n4644 , n388 );
and ( n4919 , n4917 , n4918 );
and ( n4920 , n4916 , n4919 );
buf ( n4921 , n4920 );
and ( n4922 , n4914 , n4921 );
or ( n4923 , n4913 , n4922 );
and ( n4924 , n4910 , n4923 );
or ( n4925 , n4909 , n4924 );
and ( n4926 , n4906 , n4925 );
or ( n4927 , n4905 , n4926 );
and ( n4928 , n4902 , n4927 );
or ( n4929 , n4901 , n4928 );
and ( n4930 , n4898 , n4929 );
or ( n4931 , n4897 , n4930 );
and ( n4932 , n4894 , n4931 );
or ( n4933 , n4893 , n4932 );
and ( n4934 , n4890 , n4933 );
or ( n4935 , n4889 , n4934 );
and ( n4936 , n4886 , n4935 );
or ( n4937 , n4885 , n4936 );
and ( n4938 , n4882 , n4937 );
or ( n4939 , n4881 , n4938 );
and ( n4940 , n4878 , n4939 );
or ( n4941 , n4877 , n4940 );
and ( n4942 , n4874 , n4941 );
or ( n4943 , n4873 , n4942 );
and ( n4944 , n4870 , n4943 );
or ( n4945 , n4869 , n4944 );
and ( n4946 , n4866 , n4945 );
or ( n4947 , n4865 , n4946 );
and ( n4948 , n4862 , n4947 );
or ( n4949 , n4861 , n4948 );
buf ( n4950 , n4949 );
and ( n4951 , n4474 , n387 );
and ( n4952 , n4950 , n4951 );
xor ( n4953 , n4950 , n4951 );
xor ( n4954 , n4862 , n4947 );
and ( n4955 , n4479 , n387 );
and ( n4956 , n4954 , n4955 );
xor ( n4957 , n4954 , n4955 );
xor ( n4958 , n4866 , n4945 );
and ( n4959 , n4485 , n387 );
and ( n4960 , n4958 , n4959 );
xor ( n4961 , n4958 , n4959 );
xor ( n4962 , n4870 , n4943 );
and ( n4963 , n4491 , n387 );
and ( n4964 , n4962 , n4963 );
xor ( n4965 , n4962 , n4963 );
xor ( n4966 , n4874 , n4941 );
and ( n4967 , n4497 , n387 );
and ( n4968 , n4966 , n4967 );
xor ( n4969 , n4966 , n4967 );
xor ( n4970 , n4878 , n4939 );
and ( n4971 , n4503 , n387 );
and ( n4972 , n4970 , n4971 );
xor ( n4973 , n4970 , n4971 );
xor ( n4974 , n4882 , n4937 );
and ( n4975 , n4509 , n387 );
and ( n4976 , n4974 , n4975 );
xor ( n4977 , n4974 , n4975 );
xor ( n4978 , n4886 , n4935 );
and ( n4979 , n4515 , n387 );
and ( n4980 , n4978 , n4979 );
xor ( n4981 , n4978 , n4979 );
xor ( n4982 , n4890 , n4933 );
and ( n4983 , n4521 , n387 );
and ( n4984 , n4982 , n4983 );
xor ( n4985 , n4982 , n4983 );
xor ( n4986 , n4894 , n4931 );
and ( n4987 , n4527 , n387 );
and ( n4988 , n4986 , n4987 );
xor ( n4989 , n4986 , n4987 );
xor ( n4990 , n4898 , n4929 );
and ( n4991 , n4533 , n387 );
and ( n4992 , n4990 , n4991 );
xor ( n4993 , n4990 , n4991 );
xor ( n4994 , n4902 , n4927 );
and ( n4995 , n4539 , n387 );
and ( n4996 , n4994 , n4995 );
xor ( n4997 , n4994 , n4995 );
xor ( n4998 , n4906 , n4925 );
and ( n4999 , n4545 , n387 );
and ( n5000 , n4998 , n4999 );
xor ( n5001 , n4998 , n4999 );
xor ( n5002 , n4910 , n4923 );
and ( n5003 , n4551 , n387 );
and ( n5004 , n5002 , n5003 );
xor ( n5005 , n5002 , n5003 );
xor ( n5006 , n4914 , n4921 );
buf ( n5007 , n5006 );
xor ( n5008 , n4916 , n4919 );
and ( n5009 , n4644 , n387 );
and ( n5010 , n5008 , n5009 );
and ( n5011 , n5007 , n5010 );
buf ( n5012 , n5011 );
and ( n5013 , n5005 , n5012 );
or ( n5014 , n5004 , n5013 );
and ( n5015 , n5001 , n5014 );
or ( n5016 , n5000 , n5015 );
and ( n5017 , n4997 , n5016 );
or ( n5018 , n4996 , n5017 );
and ( n5019 , n4993 , n5018 );
or ( n5020 , n4992 , n5019 );
and ( n5021 , n4989 , n5020 );
or ( n5022 , n4988 , n5021 );
and ( n5023 , n4985 , n5022 );
or ( n5024 , n4984 , n5023 );
and ( n5025 , n4981 , n5024 );
or ( n5026 , n4980 , n5025 );
and ( n5027 , n4977 , n5026 );
or ( n5028 , n4976 , n5027 );
and ( n5029 , n4973 , n5028 );
or ( n5030 , n4972 , n5029 );
and ( n5031 , n4969 , n5030 );
or ( n5032 , n4968 , n5031 );
and ( n5033 , n4965 , n5032 );
or ( n5034 , n4964 , n5033 );
and ( n5035 , n4961 , n5034 );
or ( n5036 , n4960 , n5035 );
and ( n5037 , n4957 , n5036 );
or ( n5038 , n4956 , n5037 );
and ( n5039 , n4953 , n5038 );
or ( n5040 , n4952 , n5039 );
buf ( n5041 , n5040 );
and ( n5042 , n4474 , n386 );
and ( n5043 , n5041 , n5042 );
xor ( n5044 , n5041 , n5042 );
xor ( n5045 , n4953 , n5038 );
and ( n5046 , n4479 , n386 );
and ( n5047 , n5045 , n5046 );
xor ( n5048 , n5045 , n5046 );
xor ( n5049 , n4957 , n5036 );
and ( n5050 , n4485 , n386 );
and ( n5051 , n5049 , n5050 );
xor ( n5052 , n5049 , n5050 );
xor ( n5053 , n4961 , n5034 );
and ( n5054 , n4491 , n386 );
and ( n5055 , n5053 , n5054 );
xor ( n5056 , n5053 , n5054 );
xor ( n5057 , n4965 , n5032 );
and ( n5058 , n4497 , n386 );
and ( n5059 , n5057 , n5058 );
xor ( n5060 , n5057 , n5058 );
xor ( n5061 , n4969 , n5030 );
and ( n5062 , n4503 , n386 );
and ( n5063 , n5061 , n5062 );
xor ( n5064 , n5061 , n5062 );
xor ( n5065 , n4973 , n5028 );
and ( n5066 , n4509 , n386 );
and ( n5067 , n5065 , n5066 );
xor ( n5068 , n5065 , n5066 );
xor ( n5069 , n4977 , n5026 );
and ( n5070 , n4515 , n386 );
and ( n5071 , n5069 , n5070 );
xor ( n5072 , n5069 , n5070 );
xor ( n5073 , n4981 , n5024 );
and ( n5074 , n4521 , n386 );
and ( n5075 , n5073 , n5074 );
xor ( n5076 , n5073 , n5074 );
xor ( n5077 , n4985 , n5022 );
and ( n5078 , n4527 , n386 );
and ( n5079 , n5077 , n5078 );
xor ( n5080 , n5077 , n5078 );
xor ( n5081 , n4989 , n5020 );
and ( n5082 , n4533 , n386 );
and ( n5083 , n5081 , n5082 );
xor ( n5084 , n5081 , n5082 );
xor ( n5085 , n4993 , n5018 );
and ( n5086 , n4539 , n386 );
and ( n5087 , n5085 , n5086 );
xor ( n5088 , n5085 , n5086 );
xor ( n5089 , n4997 , n5016 );
and ( n5090 , n4545 , n386 );
and ( n5091 , n5089 , n5090 );
xor ( n5092 , n5089 , n5090 );
xor ( n5093 , n5001 , n5014 );
and ( n5094 , n4551 , n386 );
and ( n5095 , n5093 , n5094 );
xor ( n5096 , n5093 , n5094 );
xor ( n5097 , n5005 , n5012 );
buf ( n5098 , n5097 );
xor ( n5099 , n5007 , n5010 );
and ( n5100 , n4644 , n386 );
and ( n5101 , n5099 , n5100 );
and ( n5102 , n5098 , n5101 );
buf ( n5103 , n5102 );
and ( n5104 , n5096 , n5103 );
or ( n5105 , n5095 , n5104 );
and ( n5106 , n5092 , n5105 );
or ( n5107 , n5091 , n5106 );
and ( n5108 , n5088 , n5107 );
or ( n5109 , n5087 , n5108 );
and ( n5110 , n5084 , n5109 );
or ( n5111 , n5083 , n5110 );
and ( n5112 , n5080 , n5111 );
or ( n5113 , n5079 , n5112 );
and ( n5114 , n5076 , n5113 );
or ( n5115 , n5075 , n5114 );
and ( n5116 , n5072 , n5115 );
or ( n5117 , n5071 , n5116 );
and ( n5118 , n5068 , n5117 );
or ( n5119 , n5067 , n5118 );
and ( n5120 , n5064 , n5119 );
or ( n5121 , n5063 , n5120 );
and ( n5122 , n5060 , n5121 );
or ( n5123 , n5059 , n5122 );
and ( n5124 , n5056 , n5123 );
or ( n5125 , n5055 , n5124 );
and ( n5126 , n5052 , n5125 );
or ( n5127 , n5051 , n5126 );
and ( n5128 , n5048 , n5127 );
or ( n5129 , n5047 , n5128 );
and ( n5130 , n5044 , n5129 );
or ( n5131 , n5043 , n5130 );
buf ( n5132 , n5131 );
buf ( n5133 , n5132 );
xor ( n5134 , n5044 , n5129 );
buf ( n5135 , n5134 );
xor ( n5136 , n5048 , n5127 );
buf ( n5137 , n5136 );
xor ( n5138 , n5052 , n5125 );
buf ( n5139 , n5138 );
xor ( n5140 , n5056 , n5123 );
buf ( n5141 , n5140 );
xor ( n5142 , n5060 , n5121 );
buf ( n5143 , n5142 );
xor ( n5144 , n5064 , n5119 );
buf ( n5145 , n5144 );
xor ( n5146 , n5068 , n5117 );
buf ( n5147 , n5146 );
xor ( n5148 , n5072 , n5115 );
buf ( n5149 , n5148 );
xor ( n5150 , n5076 , n5113 );
buf ( n5151 , n5150 );
xor ( n5152 , n5080 , n5111 );
buf ( n5153 , n5152 );
xor ( n5154 , n5084 , n5109 );
buf ( n5155 , n5154 );
xor ( n5156 , n5088 , n5107 );
buf ( n5157 , n5156 );
xor ( n5158 , n5092 , n5105 );
buf ( n5159 , n5158 );
xor ( n5160 , n5096 , n5103 );
buf ( n5161 , n5160 );
xor ( n5162 , n5098 , n5101 );
buf ( n5163 , n5162 );
xor ( n5164 , n5099 , n5100 );
buf ( n5165 , n5164 );
xor ( n5166 , n5008 , n5009 );
buf ( n5167 , n5166 );
xor ( n5168 , n4917 , n4918 );
buf ( n5169 , n5168 );
xor ( n5170 , n4826 , n4827 );
buf ( n5171 , n5170 );
xor ( n5172 , n4735 , n4736 );
buf ( n5173 , n5172 );
xor ( n5174 , n4642 , n4645 );
buf ( n5175 , n5174 );
and ( n5176 , n4644 , n392 );
buf ( n5177 , n5176 );
buf ( n5178 , n5177 );
buf ( n5179 , n4644 );
buf ( n5180 , n5179 );
buf ( n5181 , n402 );
buf ( n5182 , n416 );
buf ( n5183 , n417 );
buf ( n5184 , n403 );
buf ( n5185 , n404 );
buf ( n5186 , n405 );
buf ( n5187 , n406 );
buf ( n5188 , n407 );
buf ( n5189 , n408 );
buf ( n5190 , n409 );
buf ( n5191 , n415 );
buf ( n5192 , n414 );
buf ( n5193 , n413 );
buf ( n5194 , n412 );
buf ( n5195 , n411 );
buf ( n5196 , n410 );
buf ( n5197 , n5133 );
buf ( n5198 , n5135 );
buf ( n5199 , n5137 );
buf ( n5200 , n5139 );
buf ( n5201 , n5141 );
buf ( n5202 , n5143 );
buf ( n5203 , n5145 );
buf ( n5204 , n5147 );
buf ( n5205 , n5149 );
buf ( n5206 , n5181 );
buf ( n5207 , n5196 );
and ( n5208 , n5206 , n5207 );
buf ( n5209 , n5151 );
and ( n5210 , n5208 , n5209 );
buf ( n5211 , n5185 );
and ( n5212 , n5211 , n5207 );
buf ( n5213 , n5184 );
buf ( n5214 , n5195 );
and ( n5215 , n5213 , n5214 );
and ( n5216 , n5212 , n5215 );
buf ( n5217 , n5194 );
and ( n5218 , n5206 , n5217 );
and ( n5219 , n5215 , n5218 );
and ( n5220 , n5212 , n5218 );
or ( n5221 , n5216 , n5219 , n5220 );
and ( n5222 , n5213 , n5207 );
and ( n5223 , n5221 , n5222 );
and ( n5224 , n5206 , n5214 );
and ( n5225 , n5222 , n5224 );
and ( n5226 , n5221 , n5224 );
or ( n5227 , n5223 , n5225 , n5226 );
and ( n5228 , n5209 , n5227 );
and ( n5229 , n5208 , n5227 );
or ( n5230 , n5210 , n5228 , n5229 );
and ( n5231 , n5205 , n5230 );
xor ( n5232 , n5208 , n5209 );
xor ( n5233 , n5232 , n5227 );
buf ( n5234 , n5153 );
xor ( n5235 , n5221 , n5222 );
xor ( n5236 , n5235 , n5224 );
and ( n5237 , n5234 , n5236 );
and ( n5238 , n5211 , n5214 );
and ( n5239 , n5213 , n5217 );
and ( n5240 , n5238 , n5239 );
buf ( n5241 , n5193 );
and ( n5242 , n5206 , n5241 );
and ( n5243 , n5239 , n5242 );
and ( n5244 , n5238 , n5242 );
or ( n5245 , n5240 , n5243 , n5244 );
buf ( n5246 , n5187 );
and ( n5247 , n5246 , n5207 );
buf ( n5248 , n5186 );
and ( n5249 , n5248 , n5214 );
and ( n5250 , n5247 , n5249 );
and ( n5251 , n5211 , n5217 );
and ( n5252 , n5249 , n5251 );
and ( n5253 , n5247 , n5251 );
or ( n5254 , n5250 , n5252 , n5253 );
and ( n5255 , n5213 , n5241 );
buf ( n5256 , n5192 );
and ( n5257 , n5206 , n5256 );
and ( n5258 , n5255 , n5257 );
and ( n5259 , n5254 , n5258 );
and ( n5260 , n5248 , n5207 );
and ( n5261 , n5258 , n5260 );
and ( n5262 , n5254 , n5260 );
or ( n5263 , n5259 , n5261 , n5262 );
and ( n5264 , n5245 , n5263 );
xor ( n5265 , n5212 , n5215 );
xor ( n5266 , n5265 , n5218 );
and ( n5267 , n5263 , n5266 );
and ( n5268 , n5245 , n5266 );
or ( n5269 , n5264 , n5267 , n5268 );
and ( n5270 , n5236 , n5269 );
and ( n5271 , n5234 , n5269 );
or ( n5272 , n5237 , n5270 , n5271 );
and ( n5273 , n5233 , n5272 );
buf ( n5274 , n5155 );
xor ( n5275 , n5245 , n5263 );
xor ( n5276 , n5275 , n5266 );
and ( n5277 , n5274 , n5276 );
buf ( n5278 , n5157 );
xor ( n5279 , n5238 , n5239 );
xor ( n5280 , n5279 , n5242 );
and ( n5281 , n5278 , n5280 );
xor ( n5282 , n5254 , n5258 );
xor ( n5283 , n5282 , n5260 );
and ( n5284 , n5280 , n5283 );
and ( n5285 , n5278 , n5283 );
or ( n5286 , n5281 , n5284 , n5285 );
and ( n5287 , n5276 , n5286 );
and ( n5288 , n5274 , n5286 );
or ( n5289 , n5277 , n5287 , n5288 );
xor ( n5290 , n5234 , n5236 );
xor ( n5291 , n5290 , n5269 );
and ( n5292 , n5289 , n5291 );
and ( n5293 , n5246 , n5214 );
and ( n5294 , n5213 , n5256 );
and ( n5295 , n5293 , n5294 );
buf ( n5296 , n5191 );
and ( n5297 , n5206 , n5296 );
and ( n5298 , n5294 , n5297 );
and ( n5299 , n5293 , n5297 );
or ( n5300 , n5295 , n5298 , n5299 );
xor ( n5301 , n5247 , n5249 );
xor ( n5302 , n5301 , n5251 );
and ( n5303 , n5300 , n5302 );
buf ( n5304 , n5159 );
xor ( n5305 , n5255 , n5257 );
and ( n5306 , n5304 , n5305 );
buf ( n5307 , n5188 );
and ( n5308 , n5307 , n5207 );
and ( n5309 , n5248 , n5217 );
and ( n5310 , n5308 , n5309 );
and ( n5311 , n5211 , n5241 );
and ( n5312 , n5309 , n5311 );
and ( n5313 , n5308 , n5311 );
or ( n5314 , n5310 , n5312 , n5313 );
and ( n5315 , n5305 , n5314 );
and ( n5316 , n5304 , n5314 );
or ( n5317 , n5306 , n5315 , n5316 );
and ( n5318 , n5303 , n5317 );
xor ( n5319 , n5300 , n5302 );
buf ( n5320 , n5189 );
and ( n5321 , n5320 , n5207 );
and ( n5322 , n5211 , n5256 );
and ( n5323 , n5321 , n5322 );
and ( n5324 , n5213 , n5296 );
and ( n5325 , n5322 , n5324 );
and ( n5326 , n5321 , n5324 );
or ( n5327 , n5323 , n5325 , n5326 );
xor ( n5328 , n5293 , n5294 );
xor ( n5329 , n5328 , n5297 );
and ( n5330 , n5327 , n5329 );
xor ( n5331 , n5308 , n5309 );
xor ( n5332 , n5331 , n5311 );
and ( n5333 , n5329 , n5332 );
and ( n5334 , n5327 , n5332 );
or ( n5335 , n5330 , n5333 , n5334 );
and ( n5336 , n5319 , n5335 );
xor ( n5337 , n5304 , n5305 );
xor ( n5338 , n5337 , n5314 );
and ( n5339 , n5335 , n5338 );
and ( n5340 , n5319 , n5338 );
or ( n5341 , n5336 , n5339 , n5340 );
and ( n5342 , n5317 , n5341 );
and ( n5343 , n5303 , n5341 );
or ( n5344 , n5318 , n5342 , n5343 );
xor ( n5345 , n5274 , n5276 );
xor ( n5346 , n5345 , n5286 );
and ( n5347 , n5344 , n5346 );
xor ( n5348 , n5278 , n5280 );
xor ( n5349 , n5348 , n5283 );
xor ( n5350 , n5303 , n5317 );
xor ( n5351 , n5350 , n5341 );
and ( n5352 , n5349 , n5351 );
buf ( n5353 , n5161 );
and ( n5354 , n5307 , n5214 );
and ( n5355 , n5248 , n5241 );
and ( n5356 , n5354 , n5355 );
buf ( n5357 , n5182 );
and ( n5358 , n5206 , n5357 );
and ( n5359 , n5355 , n5358 );
and ( n5360 , n5354 , n5358 );
or ( n5361 , n5356 , n5359 , n5360 );
and ( n5362 , n5353 , n5361 );
xor ( n5363 , n5327 , n5329 );
xor ( n5364 , n5363 , n5332 );
and ( n5365 , n5361 , n5364 );
and ( n5366 , n5353 , n5364 );
or ( n5367 , n5362 , n5365 , n5366 );
xor ( n5368 , n5319 , n5335 );
xor ( n5369 , n5368 , n5338 );
and ( n5370 , n5367 , n5369 );
xor ( n5371 , n5321 , n5322 );
xor ( n5372 , n5371 , n5324 );
xor ( n5373 , n5354 , n5355 );
xor ( n5374 , n5373 , n5358 );
and ( n5375 , n5372 , n5374 );
and ( n5376 , n5246 , n5217 );
buf ( n5377 , n5163 );
and ( n5378 , n5376 , n5377 );
and ( n5379 , n5246 , n5241 );
and ( n5380 , n5211 , n5296 );
and ( n5381 , n5379 , n5380 );
and ( n5382 , n5213 , n5357 );
and ( n5383 , n5380 , n5382 );
and ( n5384 , n5379 , n5382 );
or ( n5385 , n5381 , n5383 , n5384 );
and ( n5386 , n5377 , n5385 );
and ( n5387 , n5376 , n5385 );
or ( n5388 , n5378 , n5386 , n5387 );
and ( n5389 , n5375 , n5388 );
buf ( n5390 , n5190 );
and ( n5391 , n5390 , n5207 );
and ( n5392 , n5307 , n5217 );
and ( n5393 , n5391 , n5392 );
and ( n5394 , n5248 , n5256 );
and ( n5395 , n5392 , n5394 );
and ( n5396 , n5391 , n5394 );
or ( n5397 , n5393 , n5395 , n5396 );
and ( n5398 , n5320 , n5214 );
buf ( n5399 , n5183 );
and ( n5400 , n5206 , n5399 );
and ( n5401 , n5398 , n5400 );
buf ( n5402 , n5165 );
and ( n5403 , n5400 , n5402 );
and ( n5404 , n5398 , n5402 );
or ( n5405 , n5401 , n5403 , n5404 );
and ( n5406 , n5397 , n5405 );
xor ( n5407 , n5372 , n5374 );
and ( n5408 , n5405 , n5407 );
and ( n5409 , n5397 , n5407 );
or ( n5410 , n5406 , n5408 , n5409 );
and ( n5411 , n5388 , n5410 );
and ( n5412 , n5375 , n5410 );
or ( n5413 , n5389 , n5411 , n5412 );
and ( n5414 , n5369 , n5413 );
and ( n5415 , n5367 , n5413 );
or ( n5416 , n5370 , n5414 , n5415 );
and ( n5417 , n5351 , n5416 );
and ( n5418 , n5349 , n5416 );
or ( n5419 , n5352 , n5417 , n5418 );
and ( n5420 , n5346 , n5419 );
and ( n5421 , n5344 , n5419 );
or ( n5422 , n5347 , n5420 , n5421 );
and ( n5423 , n5291 , n5422 );
and ( n5424 , n5289 , n5422 );
or ( n5425 , n5292 , n5423 , n5424 );
and ( n5426 , n5272 , n5425 );
and ( n5427 , n5233 , n5425 );
or ( n5428 , n5273 , n5426 , n5427 );
and ( n5429 , n5230 , n5428 );
and ( n5430 , n5205 , n5428 );
or ( n5431 , n5231 , n5429 , n5430 );
and ( n5432 , n5204 , n5431 );
xor ( n5433 , n5204 , n5431 );
xor ( n5434 , n5205 , n5230 );
xor ( n5435 , n5434 , n5428 );
xor ( n5436 , n5233 , n5272 );
xor ( n5437 , n5436 , n5425 );
xor ( n5438 , n5289 , n5291 );
xor ( n5439 , n5438 , n5422 );
xor ( n5440 , n5344 , n5346 );
xor ( n5441 , n5440 , n5419 );
xor ( n5442 , n5349 , n5351 );
xor ( n5443 , n5442 , n5416 );
and ( n5444 , n5320 , n5217 );
and ( n5445 , n5307 , n5241 );
and ( n5446 , n5444 , n5445 );
and ( n5447 , n5246 , n5256 );
and ( n5448 , n5445 , n5447 );
and ( n5449 , n5444 , n5447 );
or ( n5450 , n5446 , n5448 , n5449 );
xor ( n5451 , n5379 , n5380 );
xor ( n5452 , n5451 , n5382 );
and ( n5453 , n5450 , n5452 );
xor ( n5454 , n5391 , n5392 );
xor ( n5455 , n5454 , n5394 );
and ( n5456 , n5452 , n5455 );
and ( n5457 , n5450 , n5455 );
or ( n5458 , n5453 , n5456 , n5457 );
and ( n5459 , n5211 , n5357 );
and ( n5460 , n5213 , n5399 );
and ( n5461 , n5459 , n5460 );
and ( n5462 , n5390 , n5214 );
and ( n5463 , n5248 , n5296 );
and ( n5464 , n5462 , n5463 );
buf ( n5465 , n5167 );
and ( n5466 , n5463 , n5465 );
and ( n5467 , n5462 , n5465 );
or ( n5468 , n5464 , n5466 , n5467 );
and ( n5469 , n5461 , n5468 );
xor ( n5470 , n5398 , n5400 );
xor ( n5471 , n5470 , n5402 );
and ( n5472 , n5468 , n5471 );
and ( n5473 , n5461 , n5471 );
or ( n5474 , n5469 , n5472 , n5473 );
and ( n5475 , n5458 , n5474 );
xor ( n5476 , n5376 , n5377 );
xor ( n5477 , n5476 , n5385 );
and ( n5478 , n5474 , n5477 );
and ( n5479 , n5458 , n5477 );
or ( n5480 , n5475 , n5478 , n5479 );
xor ( n5481 , n5353 , n5361 );
xor ( n5482 , n5481 , n5364 );
and ( n5483 , n5480 , n5482 );
xor ( n5484 , n5450 , n5452 );
xor ( n5485 , n5484 , n5455 );
and ( n5486 , n5390 , n5217 );
and ( n5487 , n5320 , n5241 );
and ( n5488 , n5486 , n5487 );
and ( n5489 , n5307 , n5256 );
and ( n5490 , n5487 , n5489 );
and ( n5491 , n5486 , n5489 );
or ( n5492 , n5488 , n5490 , n5491 );
and ( n5493 , n5246 , n5296 );
and ( n5494 , n5248 , n5357 );
and ( n5495 , n5493 , n5494 );
and ( n5496 , n5492 , n5495 );
and ( n5497 , n5485 , n5496 );
xor ( n5498 , n5444 , n5445 );
xor ( n5499 , n5498 , n5447 );
xor ( n5500 , n5459 , n5460 );
and ( n5501 , n5499 , n5500 );
xor ( n5502 , n5462 , n5463 );
xor ( n5503 , n5502 , n5465 );
and ( n5504 , n5500 , n5503 );
and ( n5505 , n5499 , n5503 );
or ( n5506 , n5501 , n5504 , n5505 );
and ( n5507 , n5496 , n5506 );
and ( n5508 , n5485 , n5506 );
or ( n5509 , n5497 , n5507 , n5508 );
xor ( n5510 , n5397 , n5405 );
xor ( n5511 , n5510 , n5407 );
and ( n5512 , n5509 , n5511 );
xor ( n5513 , n5458 , n5474 );
xor ( n5514 , n5513 , n5477 );
and ( n5515 , n5511 , n5514 );
and ( n5516 , n5509 , n5514 );
or ( n5517 , n5512 , n5515 , n5516 );
and ( n5518 , n5482 , n5517 );
and ( n5519 , n5480 , n5517 );
or ( n5520 , n5483 , n5518 , n5519 );
xor ( n5521 , n5367 , n5369 );
xor ( n5522 , n5521 , n5413 );
and ( n5523 , n5520 , n5522 );
xor ( n5524 , n5520 , n5522 );
xor ( n5525 , n5375 , n5388 );
xor ( n5526 , n5525 , n5410 );
xor ( n5527 , n5480 , n5482 );
xor ( n5528 , n5527 , n5517 );
and ( n5529 , n5526 , n5528 );
xor ( n5530 , n5526 , n5528 );
xor ( n5531 , n5461 , n5468 );
xor ( n5532 , n5531 , n5471 );
xor ( n5533 , n5492 , n5495 );
and ( n5534 , n5390 , n5241 );
and ( n5535 , n5307 , n5296 );
and ( n5536 , n5534 , n5535 );
and ( n5537 , n5246 , n5357 );
and ( n5538 , n5535 , n5537 );
and ( n5539 , n5534 , n5537 );
or ( n5540 , n5536 , n5538 , n5539 );
xor ( n5541 , n5486 , n5487 );
xor ( n5542 , n5541 , n5489 );
and ( n5543 , n5540 , n5542 );
and ( n5544 , n5533 , n5543 );
and ( n5545 , n5211 , n5399 );
buf ( n5546 , n5169 );
and ( n5547 , n5545 , n5546 );
xor ( n5548 , n5493 , n5494 );
and ( n5549 , n5546 , n5548 );
and ( n5550 , n5545 , n5548 );
or ( n5551 , n5547 , n5549 , n5550 );
and ( n5552 , n5543 , n5551 );
and ( n5553 , n5533 , n5551 );
or ( n5554 , n5544 , n5552 , n5553 );
and ( n5555 , n5532 , n5554 );
xor ( n5556 , n5485 , n5496 );
xor ( n5557 , n5556 , n5506 );
and ( n5558 , n5554 , n5557 );
and ( n5559 , n5532 , n5557 );
or ( n5560 , n5555 , n5558 , n5559 );
xor ( n5561 , n5509 , n5511 );
xor ( n5562 , n5561 , n5514 );
and ( n5563 , n5560 , n5562 );
xor ( n5564 , n5560 , n5562 );
xor ( n5565 , n5499 , n5500 );
xor ( n5566 , n5565 , n5503 );
and ( n5567 , n5320 , n5256 );
and ( n5568 , n5248 , n5399 );
and ( n5569 , n5567 , n5568 );
buf ( n5570 , n5171 );
and ( n5571 , n5568 , n5570 );
and ( n5572 , n5567 , n5570 );
or ( n5573 , n5569 , n5571 , n5572 );
xor ( n5574 , n5540 , n5542 );
and ( n5575 , n5573 , n5574 );
xor ( n5576 , n5534 , n5535 );
xor ( n5577 , n5576 , n5537 );
and ( n5578 , n5320 , n5296 );
and ( n5579 , n5307 , n5357 );
and ( n5580 , n5578 , n5579 );
and ( n5581 , n5246 , n5399 );
and ( n5582 , n5579 , n5581 );
and ( n5583 , n5578 , n5581 );
or ( n5584 , n5580 , n5582 , n5583 );
and ( n5585 , n5577 , n5584 );
xor ( n5586 , n5567 , n5568 );
xor ( n5587 , n5586 , n5570 );
and ( n5588 , n5584 , n5587 );
and ( n5589 , n5577 , n5587 );
or ( n5590 , n5585 , n5588 , n5589 );
and ( n5591 , n5574 , n5590 );
and ( n5592 , n5573 , n5590 );
or ( n5593 , n5575 , n5591 , n5592 );
and ( n5594 , n5566 , n5593 );
xor ( n5595 , n5533 , n5543 );
xor ( n5596 , n5595 , n5551 );
and ( n5597 , n5593 , n5596 );
and ( n5598 , n5566 , n5596 );
or ( n5599 , n5594 , n5597 , n5598 );
xor ( n5600 , n5532 , n5554 );
xor ( n5601 , n5600 , n5557 );
and ( n5602 , n5599 , n5601 );
xor ( n5603 , n5599 , n5601 );
xor ( n5604 , n5566 , n5593 );
xor ( n5605 , n5604 , n5596 );
xor ( n5606 , n5545 , n5546 );
xor ( n5607 , n5606 , n5548 );
xor ( n5608 , n5573 , n5574 );
xor ( n5609 , n5608 , n5590 );
and ( n5610 , n5607 , n5609 );
and ( n5611 , n5390 , n5296 );
and ( n5612 , n5320 , n5357 );
and ( n5613 , n5611 , n5612 );
and ( n5614 , n5307 , n5399 );
and ( n5615 , n5612 , n5614 );
and ( n5616 , n5611 , n5614 );
or ( n5617 , n5613 , n5615 , n5616 );
xor ( n5618 , n5578 , n5579 );
xor ( n5619 , n5618 , n5581 );
and ( n5620 , n5617 , n5619 );
xor ( n5621 , n5577 , n5584 );
xor ( n5622 , n5621 , n5587 );
and ( n5623 , n5620 , n5622 );
and ( n5624 , n5390 , n5256 );
buf ( n5625 , n5173 );
and ( n5626 , n5624 , n5625 );
xor ( n5627 , n5617 , n5619 );
and ( n5628 , n5625 , n5627 );
and ( n5629 , n5624 , n5627 );
or ( n5630 , n5626 , n5628 , n5629 );
and ( n5631 , n5622 , n5630 );
and ( n5632 , n5620 , n5630 );
or ( n5633 , n5623 , n5631 , n5632 );
and ( n5634 , n5609 , n5633 );
and ( n5635 , n5607 , n5633 );
or ( n5636 , n5610 , n5634 , n5635 );
and ( n5637 , n5605 , n5636 );
xor ( n5638 , n5605 , n5636 );
xor ( n5639 , n5607 , n5609 );
xor ( n5640 , n5639 , n5633 );
xor ( n5641 , n5620 , n5622 );
xor ( n5642 , n5641 , n5630 );
buf ( n5643 , n5175 );
xor ( n5644 , n5611 , n5612 );
xor ( n5645 , n5644 , n5614 );
and ( n5646 , n5643 , n5645 );
and ( n5647 , n5390 , n5357 );
and ( n5648 , n5320 , n5399 );
and ( n5649 , n5647 , n5648 );
buf ( n5650 , n5178 );
and ( n5651 , n5648 , n5650 );
and ( n5652 , n5647 , n5650 );
or ( n5653 , n5649 , n5651 , n5652 );
and ( n5654 , n5645 , n5653 );
and ( n5655 , n5643 , n5653 );
or ( n5656 , n5646 , n5654 , n5655 );
xor ( n5657 , n5624 , n5625 );
xor ( n5658 , n5657 , n5627 );
and ( n5659 , n5656 , n5658 );
xor ( n5660 , n5656 , n5658 );
xor ( n5661 , n5643 , n5645 );
xor ( n5662 , n5661 , n5653 );
xor ( n5663 , n5647 , n5648 );
xor ( n5664 , n5663 , n5650 );
and ( n5665 , n5390 , n5399 );
buf ( n5666 , n5180 );
and ( n5667 , n5665 , n5666 );
and ( n5668 , n5664 , n5667 );
and ( n5669 , n5662 , n5668 );
and ( n5670 , n5660 , n5669 );
or ( n5671 , n5659 , n5670 );
and ( n5672 , n5642 , n5671 );
and ( n5673 , n5640 , n5672 );
and ( n5674 , n5638 , n5673 );
or ( n5675 , n5637 , n5674 );
and ( n5676 , n5603 , n5675 );
or ( n5677 , n5602 , n5676 );
and ( n5678 , n5564 , n5677 );
or ( n5679 , n5563 , n5678 );
and ( n5680 , n5530 , n5679 );
or ( n5681 , n5529 , n5680 );
and ( n5682 , n5524 , n5681 );
or ( n5683 , n5523 , n5682 );
and ( n5684 , n5443 , n5683 );
and ( n5685 , n5441 , n5684 );
and ( n5686 , n5439 , n5685 );
and ( n5687 , n5437 , n5686 );
and ( n5688 , n5435 , n5687 );
and ( n5689 , n5433 , n5688 );
or ( n5690 , n5432 , n5689 );
and ( n5691 , n5203 , n5690 );
and ( n5692 , n5202 , n5691 );
and ( n5693 , n5201 , n5692 );
and ( n5694 , n5200 , n5693 );
and ( n5695 , n5199 , n5694 );
and ( n5696 , n5198 , n5695 );
xor ( n5697 , n5197 , n5696 );
buf ( n5698 , n5697 );
xor ( n5699 , n5198 , n5695 );
buf ( n5700 , n5699 );
xor ( n5701 , n5199 , n5694 );
buf ( n5702 , n5701 );
xor ( n5703 , n5200 , n5693 );
buf ( n5704 , n5703 );
xor ( n5705 , n5201 , n5692 );
buf ( n5706 , n5705 );
xor ( n5707 , n5202 , n5691 );
buf ( n5708 , n5707 );
xor ( n5709 , n5203 , n5690 );
buf ( n5710 , n5709 );
xor ( n5711 , n5433 , n5688 );
buf ( n5712 , n5711 );
xor ( n5713 , n5435 , n5687 );
buf ( n5714 , n5713 );
xor ( n5715 , n5437 , n5686 );
buf ( n5716 , n5715 );
xor ( n5717 , n5439 , n5685 );
buf ( n5718 , n5717 );
xor ( n5719 , n5441 , n5684 );
buf ( n5720 , n5719 );
xor ( n5721 , n5443 , n5683 );
buf ( n5722 , n5721 );
xor ( n5723 , n5524 , n5681 );
buf ( n5724 , n5723 );
buf ( n5725 , n370 );
buf ( n5726 , n5725 );
buf ( n5727 , n5726 );
buf ( n5728 , n371 );
buf ( n5729 , n5728 );
buf ( n5730 , n370 );
buf ( n5731 , n5730 );
and ( n5732 , n5729 , n5731 );
buf ( n5733 , n371 );
buf ( n5734 , n5733 );
and ( n5735 , n5726 , n5734 );
and ( n5736 , n5732 , n5735 );
buf ( n5737 , n372 );
buf ( n5738 , n5737 );
and ( n5739 , n5726 , n5738 );
buf ( n5740 , n372 );
buf ( n5741 , n5740 );
and ( n5742 , n5741 , n5731 );
and ( n5743 , n5739 , n5742 );
and ( n5744 , n5735 , n5743 );
and ( n5745 , n5732 , n5743 );
or ( n5746 , n5736 , n5744 , n5745 );
and ( n5747 , n5727 , n5746 );
buf ( n5748 , n373 );
buf ( n5749 , n5748 );
and ( n5750 , n5749 , n5731 );
and ( n5751 , n5741 , n5734 );
or ( n5752 , n5750 , n5751 );
buf ( n5753 , n373 );
buf ( n5754 , n5753 );
and ( n5755 , n5726 , n5754 );
and ( n5756 , n5729 , n5738 );
or ( n5757 , n5755 , n5756 );
and ( n5758 , n5752 , n5757 );
xor ( n5759 , n5732 , n5735 );
xor ( n5760 , n5759 , n5743 );
and ( n5761 , n5758 , n5760 );
buf ( n5762 , n5729 );
xor ( n5763 , n5739 , n5742 );
and ( n5764 , n5762 , n5763 );
xor ( n5765 , n5752 , n5757 );
and ( n5766 , n5763 , n5765 );
and ( n5767 , n5762 , n5765 );
or ( n5768 , n5764 , n5766 , n5767 );
and ( n5769 , n5760 , n5768 );
and ( n5770 , n5758 , n5768 );
or ( n5771 , n5761 , n5769 , n5770 );
and ( n5772 , n5746 , n5771 );
and ( n5773 , n5727 , n5771 );
or ( n5774 , n5747 , n5772 , n5773 );
xor ( n5775 , n5727 , n5746 );
xor ( n5776 , n5775 , n5771 );
buf ( n5777 , n374 );
buf ( n5778 , n5777 );
and ( n5779 , n5778 , n5731 );
and ( n5780 , n5749 , n5734 );
or ( n5781 , n5779 , n5780 );
buf ( n5782 , n374 );
buf ( n5783 , n5782 );
and ( n5784 , n5726 , n5783 );
and ( n5785 , n5729 , n5754 );
or ( n5786 , n5784 , n5785 );
and ( n5787 , n5781 , n5786 );
xnor ( n5788 , n5750 , n5751 );
xnor ( n5789 , n5755 , n5756 );
and ( n5790 , n5788 , n5789 );
and ( n5791 , n5787 , n5790 );
xor ( n5792 , n5781 , n5786 );
xor ( n5793 , n5788 , n5789 );
and ( n5794 , n5792 , n5793 );
buf ( n5795 , n375 );
buf ( n5796 , n5795 );
and ( n5797 , n5726 , n5796 );
buf ( n5798 , n375 );
buf ( n5799 , n5798 );
and ( n5800 , n5799 , n5731 );
and ( n5801 , n5797 , n5800 );
and ( n5802 , n5741 , n5754 );
and ( n5803 , n5749 , n5738 );
and ( n5804 , n5802 , n5803 );
and ( n5805 , n5801 , n5804 );
buf ( n5806 , n5741 );
and ( n5807 , n5804 , n5806 );
and ( n5808 , n5801 , n5806 );
or ( n5809 , n5805 , n5807 , n5808 );
and ( n5810 , n5793 , n5809 );
and ( n5811 , n5792 , n5809 );
or ( n5812 , n5794 , n5810 , n5811 );
and ( n5813 , n5790 , n5812 );
and ( n5814 , n5787 , n5812 );
or ( n5815 , n5791 , n5813 , n5814 );
xor ( n5816 , n5758 , n5760 );
xor ( n5817 , n5816 , n5768 );
and ( n5818 , n5815 , n5817 );
xor ( n5819 , n5762 , n5763 );
xor ( n5820 , n5819 , n5765 );
xnor ( n5821 , n5779 , n5780 );
xnor ( n5822 , n5784 , n5785 );
and ( n5823 , n5821 , n5822 );
buf ( n5824 , n376 );
buf ( n5825 , n5824 );
and ( n5826 , n5825 , n5731 );
and ( n5827 , n5799 , n5734 );
and ( n5828 , n5826 , n5827 );
and ( n5829 , n5778 , n5738 );
and ( n5830 , n5827 , n5829 );
and ( n5831 , n5826 , n5829 );
or ( n5832 , n5828 , n5830 , n5831 );
buf ( n5833 , n376 );
buf ( n5834 , n5833 );
and ( n5835 , n5726 , n5834 );
and ( n5836 , n5729 , n5796 );
and ( n5837 , n5835 , n5836 );
and ( n5838 , n5741 , n5783 );
and ( n5839 , n5836 , n5838 );
and ( n5840 , n5835 , n5838 );
or ( n5841 , n5837 , n5839 , n5840 );
and ( n5842 , n5832 , n5841 );
and ( n5843 , n5729 , n5783 );
and ( n5844 , n5778 , n5734 );
and ( n5845 , n5843 , n5844 );
and ( n5846 , n5842 , n5845 );
xor ( n5847 , n5801 , n5804 );
xor ( n5848 , n5847 , n5806 );
and ( n5849 , n5845 , n5848 );
and ( n5850 , n5842 , n5848 );
or ( n5851 , n5846 , n5849 , n5850 );
and ( n5852 , n5823 , n5851 );
xor ( n5853 , n5792 , n5793 );
xor ( n5854 , n5853 , n5809 );
and ( n5855 , n5851 , n5854 );
and ( n5856 , n5823 , n5854 );
or ( n5857 , n5852 , n5855 , n5856 );
and ( n5858 , n5820 , n5857 );
xor ( n5859 , n5787 , n5790 );
xor ( n5860 , n5859 , n5812 );
and ( n5861 , n5857 , n5860 );
and ( n5862 , n5820 , n5860 );
or ( n5863 , n5858 , n5861 , n5862 );
and ( n5864 , n5817 , n5863 );
and ( n5865 , n5815 , n5863 );
or ( n5866 , n5818 , n5864 , n5865 );
or ( n5867 , n5776 , n5866 );
xnor ( n5868 , n5774 , n5867 );
xnor ( n5869 , n5776 , n5866 );
xor ( n5870 , n5815 , n5817 );
xor ( n5871 , n5870 , n5863 );
not ( n5872 , n5871 );
xor ( n5873 , n5820 , n5857 );
xor ( n5874 , n5873 , n5860 );
xor ( n5875 , n5821 , n5822 );
xor ( n5876 , n5797 , n5800 );
xor ( n5877 , n5843 , n5844 );
and ( n5878 , n5876 , n5877 );
xor ( n5879 , n5802 , n5803 );
and ( n5880 , n5877 , n5879 );
and ( n5881 , n5876 , n5879 );
or ( n5882 , n5878 , n5880 , n5881 );
and ( n5883 , n5875 , n5882 );
xor ( n5884 , n5842 , n5845 );
xor ( n5885 , n5884 , n5848 );
and ( n5886 , n5882 , n5885 );
and ( n5887 , n5875 , n5885 );
or ( n5888 , n5883 , n5886 , n5887 );
xor ( n5889 , n5823 , n5851 );
xor ( n5890 , n5889 , n5854 );
and ( n5891 , n5888 , n5890 );
xor ( n5892 , n5832 , n5841 );
and ( n5893 , n5825 , n5734 );
and ( n5894 , n5799 , n5738 );
or ( n5895 , n5893 , n5894 );
and ( n5896 , n5729 , n5834 );
and ( n5897 , n5741 , n5796 );
or ( n5898 , n5896 , n5897 );
and ( n5899 , n5895 , n5898 );
and ( n5900 , n5892 , n5899 );
xor ( n5901 , n5826 , n5827 );
xor ( n5902 , n5901 , n5829 );
xor ( n5903 , n5835 , n5836 );
xor ( n5904 , n5903 , n5838 );
and ( n5905 , n5902 , n5904 );
and ( n5906 , n5899 , n5905 );
and ( n5907 , n5892 , n5905 );
or ( n5908 , n5900 , n5906 , n5907 );
buf ( n5909 , n5749 );
buf ( n5910 , n377 );
buf ( n5911 , n5910 );
and ( n5912 , n5726 , n5911 );
buf ( n5913 , n377 );
buf ( n5914 , n5913 );
and ( n5915 , n5914 , n5731 );
and ( n5916 , n5912 , n5915 );
and ( n5917 , n5909 , n5916 );
and ( n5918 , n5749 , n5783 );
and ( n5919 , n5778 , n5754 );
and ( n5920 , n5918 , n5919 );
and ( n5921 , n5916 , n5920 );
and ( n5922 , n5909 , n5920 );
or ( n5923 , n5917 , n5921 , n5922 );
xor ( n5924 , n5876 , n5877 );
xor ( n5925 , n5924 , n5879 );
and ( n5926 , n5923 , n5925 );
xor ( n5927 , n5895 , n5898 );
xor ( n5928 , n5902 , n5904 );
and ( n5929 , n5927 , n5928 );
xnor ( n5930 , n5893 , n5894 );
xnor ( n5931 , n5896 , n5897 );
and ( n5932 , n5930 , n5931 );
and ( n5933 , n5928 , n5932 );
and ( n5934 , n5927 , n5932 );
or ( n5935 , n5929 , n5933 , n5934 );
and ( n5936 , n5925 , n5935 );
and ( n5937 , n5923 , n5935 );
or ( n5938 , n5926 , n5936 , n5937 );
and ( n5939 , n5908 , n5938 );
xor ( n5940 , n5875 , n5882 );
xor ( n5941 , n5940 , n5885 );
and ( n5942 , n5938 , n5941 );
and ( n5943 , n5908 , n5941 );
or ( n5944 , n5939 , n5942 , n5943 );
and ( n5945 , n5890 , n5944 );
and ( n5946 , n5888 , n5944 );
or ( n5947 , n5891 , n5945 , n5946 );
and ( n5948 , n5874 , n5947 );
xor ( n5949 , n5874 , n5947 );
xor ( n5950 , n5888 , n5890 );
xor ( n5951 , n5950 , n5944 );
xor ( n5952 , n5892 , n5899 );
xor ( n5953 , n5952 , n5905 );
xor ( n5954 , n5912 , n5915 );
xor ( n5955 , n5918 , n5919 );
and ( n5956 , n5954 , n5955 );
and ( n5957 , n5741 , n5834 );
and ( n5958 , n5825 , n5738 );
and ( n5959 , n5957 , n5958 );
and ( n5960 , n5955 , n5959 );
and ( n5961 , n5954 , n5959 );
or ( n5962 , n5956 , n5960 , n5961 );
xor ( n5963 , n5909 , n5916 );
xor ( n5964 , n5963 , n5920 );
and ( n5965 , n5962 , n5964 );
and ( n5966 , n5749 , n5796 );
and ( n5967 , n5799 , n5754 );
and ( n5968 , n5966 , n5967 );
xor ( n5969 , n5930 , n5931 );
and ( n5970 , n5968 , n5969 );
and ( n5971 , n5778 , n5796 );
and ( n5972 , n5799 , n5783 );
and ( n5973 , n5971 , n5972 );
and ( n5974 , n5729 , n5911 );
or ( n5975 , n5973 , n5974 );
and ( n5976 , n5969 , n5975 );
and ( n5977 , n5968 , n5975 );
or ( n5978 , n5970 , n5976 , n5977 );
and ( n5979 , n5964 , n5978 );
and ( n5980 , n5962 , n5978 );
or ( n5981 , n5965 , n5979 , n5980 );
and ( n5982 , n5953 , n5981 );
xor ( n5983 , n5923 , n5925 );
xor ( n5984 , n5983 , n5935 );
and ( n5985 , n5981 , n5984 );
and ( n5986 , n5953 , n5984 );
or ( n5987 , n5982 , n5985 , n5986 );
xor ( n5988 , n5908 , n5938 );
xor ( n5989 , n5988 , n5941 );
and ( n5990 , n5987 , n5989 );
and ( n5991 , n5914 , n5738 );
and ( n5992 , n5825 , n5754 );
or ( n5993 , n5991 , n5992 );
and ( n5994 , n5741 , n5911 );
and ( n5995 , n5749 , n5834 );
or ( n5996 , n5994 , n5995 );
and ( n5997 , n5993 , n5996 );
and ( n5998 , n5914 , n5734 );
buf ( n5999 , n5778 );
and ( n6000 , n5998 , n5999 );
xor ( n6001 , n5957 , n5958 );
and ( n6002 , n5999 , n6001 );
and ( n6003 , n5998 , n6001 );
or ( n6004 , n6000 , n6002 , n6003 );
and ( n6005 , n5997 , n6004 );
xor ( n6006 , n5954 , n5955 );
xor ( n6007 , n6006 , n5959 );
and ( n6008 , n6004 , n6007 );
and ( n6009 , n5997 , n6007 );
or ( n6010 , n6005 , n6008 , n6009 );
xor ( n6011 , n5927 , n5928 );
xor ( n6012 , n6011 , n5932 );
and ( n6013 , n6010 , n6012 );
xor ( n6014 , n5966 , n5967 );
xnor ( n6015 , n5973 , n5974 );
and ( n6016 , n6014 , n6015 );
xor ( n6017 , n5993 , n5996 );
and ( n6018 , n6015 , n6017 );
and ( n6019 , n6014 , n6017 );
or ( n6020 , n6016 , n6018 , n6019 );
and ( n6021 , n5914 , n5754 );
and ( n6022 , n5825 , n5783 );
or ( n6023 , n6021 , n6022 );
and ( n6024 , n5749 , n5911 );
and ( n6025 , n5778 , n5834 );
or ( n6026 , n6024 , n6025 );
and ( n6027 , n6023 , n6026 );
xnor ( n6028 , n5991 , n5992 );
xnor ( n6029 , n5994 , n5995 );
and ( n6030 , n6028 , n6029 );
and ( n6031 , n6027 , n6030 );
xor ( n6032 , n5998 , n5999 );
xor ( n6033 , n6032 , n6001 );
and ( n6034 , n6030 , n6033 );
and ( n6035 , n6027 , n6033 );
or ( n6036 , n6031 , n6034 , n6035 );
and ( n6037 , n6020 , n6036 );
xor ( n6038 , n5968 , n5969 );
xor ( n6039 , n6038 , n5975 );
and ( n6040 , n6036 , n6039 );
and ( n6041 , n6020 , n6039 );
or ( n6042 , n6037 , n6040 , n6041 );
and ( n6043 , n6012 , n6042 );
and ( n6044 , n6010 , n6042 );
or ( n6045 , n6013 , n6043 , n6044 );
xor ( n6046 , n5953 , n5981 );
xor ( n6047 , n6046 , n5984 );
and ( n6048 , n6045 , n6047 );
xor ( n6049 , n5962 , n5964 );
xor ( n6050 , n6049 , n5978 );
xor ( n6051 , n5997 , n6004 );
xor ( n6052 , n6051 , n6007 );
xor ( n6053 , n5971 , n5972 );
xor ( n6054 , n6023 , n6026 );
and ( n6055 , n6053 , n6054 );
xor ( n6056 , n6028 , n6029 );
and ( n6057 , n6054 , n6056 );
and ( n6058 , n6053 , n6056 );
or ( n6059 , n6055 , n6057 , n6058 );
xor ( n6060 , n6014 , n6015 );
xor ( n6061 , n6060 , n6017 );
and ( n6062 , n6059 , n6061 );
xor ( n6063 , n6027 , n6030 );
xor ( n6064 , n6063 , n6033 );
and ( n6065 , n6061 , n6064 );
and ( n6066 , n6059 , n6064 );
or ( n6067 , n6062 , n6065 , n6066 );
and ( n6068 , n6052 , n6067 );
xor ( n6069 , n6020 , n6036 );
xor ( n6070 , n6069 , n6039 );
and ( n6071 , n6067 , n6070 );
and ( n6072 , n6052 , n6070 );
or ( n6073 , n6068 , n6071 , n6072 );
and ( n6074 , n6050 , n6073 );
xor ( n6075 , n6010 , n6012 );
xor ( n6076 , n6075 , n6042 );
and ( n6077 , n6073 , n6076 );
and ( n6078 , n6050 , n6076 );
or ( n6079 , n6074 , n6077 , n6078 );
and ( n6080 , n6047 , n6079 );
and ( n6081 , n6045 , n6079 );
or ( n6082 , n6048 , n6080 , n6081 );
and ( n6083 , n5989 , n6082 );
and ( n6084 , n5987 , n6082 );
or ( n6085 , n5990 , n6083 , n6084 );
and ( n6086 , n5951 , n6085 );
xor ( n6087 , n5951 , n6085 );
xor ( n6088 , n5987 , n5989 );
xor ( n6089 , n6088 , n6082 );
not ( n6090 , n6089 );
xor ( n6091 , n6045 , n6047 );
xor ( n6092 , n6091 , n6079 );
not ( n6093 , n6092 );
xor ( n6094 , n6050 , n6073 );
xor ( n6095 , n6094 , n6076 );
xor ( n6096 , n6052 , n6067 );
xor ( n6097 , n6096 , n6070 );
xnor ( n6098 , n6021 , n6022 );
xnor ( n6099 , n6024 , n6025 );
and ( n6100 , n6098 , n6099 );
buf ( n6101 , n5799 );
and ( n6102 , n5778 , n5911 );
and ( n6103 , n5914 , n5783 );
and ( n6104 , n6102 , n6103 );
and ( n6105 , n6101 , n6104 );
and ( n6106 , n5799 , n5834 );
and ( n6107 , n5825 , n5796 );
and ( n6108 , n6106 , n6107 );
and ( n6109 , n6104 , n6108 );
and ( n6110 , n6101 , n6108 );
or ( n6111 , n6105 , n6109 , n6110 );
and ( n6112 , n6100 , n6111 );
xor ( n6113 , n6053 , n6054 );
xor ( n6114 , n6113 , n6056 );
and ( n6115 , n6111 , n6114 );
and ( n6116 , n6100 , n6114 );
or ( n6117 , n6112 , n6115 , n6116 );
xor ( n6118 , n6059 , n6061 );
xor ( n6119 , n6118 , n6064 );
and ( n6120 , n6117 , n6119 );
xor ( n6121 , n6098 , n6099 );
xor ( n6122 , n6101 , n6104 );
xor ( n6123 , n6122 , n6108 );
and ( n6124 , n6121 , n6123 );
xor ( n6125 , n6102 , n6103 );
xor ( n6126 , n6106 , n6107 );
and ( n6127 , n6125 , n6126 );
and ( n6128 , n5825 , n5911 );
and ( n6129 , n5914 , n5834 );
and ( n6130 , n6128 , n6129 );
and ( n6131 , n5799 , n5911 );
and ( n6132 , n6130 , n6131 );
and ( n6133 , n6126 , n6132 );
and ( n6134 , n6125 , n6132 );
or ( n6135 , n6127 , n6133 , n6134 );
and ( n6136 , n6123 , n6135 );
and ( n6137 , n6121 , n6135 );
or ( n6138 , n6124 , n6136 , n6137 );
xor ( n6139 , n6100 , n6111 );
xor ( n6140 , n6139 , n6114 );
or ( n6141 , n6138 , n6140 );
and ( n6142 , n6119 , n6141 );
and ( n6143 , n6117 , n6141 );
or ( n6144 , n6120 , n6142 , n6143 );
and ( n6145 , n6097 , n6144 );
xor ( n6146 , n6097 , n6144 );
xor ( n6147 , n6117 , n6119 );
xor ( n6148 , n6147 , n6141 );
not ( n6149 , n6148 );
xnor ( n6150 , n6138 , n6140 );
xor ( n6151 , n6121 , n6123 );
xor ( n6152 , n6151 , n6135 );
and ( n6153 , n5914 , n5796 );
buf ( n6154 , n5825 );
and ( n6155 , n6153 , n6154 );
xor ( n6156 , n6130 , n6131 );
and ( n6157 , n6154 , n6156 );
and ( n6158 , n6153 , n6156 );
or ( n6159 , n6155 , n6157 , n6158 );
xor ( n6160 , n6125 , n6126 );
xor ( n6161 , n6160 , n6132 );
and ( n6162 , n6159 , n6161 );
and ( n6163 , n6152 , n6162 );
and ( n6164 , n6150 , n6163 );
and ( n6165 , n6149 , n6164 );
or ( n6166 , n6148 , n6165 );
and ( n6167 , n6146 , n6166 );
or ( n6168 , n6145 , n6167 );
and ( n6169 , n6095 , n6168 );
and ( n6170 , n6093 , n6169 );
or ( n6171 , n6092 , n6170 );
and ( n6172 , n6090 , n6171 );
or ( n6173 , n6089 , n6172 );
and ( n6174 , n6087 , n6173 );
or ( n6175 , n6086 , n6174 );
and ( n6176 , n5949 , n6175 );
or ( n6177 , n5948 , n6176 );
and ( n6178 , n5872 , n6177 );
or ( n6179 , n5871 , n6178 );
and ( n6180 , n5869 , n6179 );
xor ( n6181 , n5868 , n6180 );
buf ( n6182 , n6181 );
and ( n6183 , n6182 , n376 );
buf ( n6184 , n6183 );
and ( n6185 , n6182 , n377 );
xor ( n6186 , n5869 , n6179 );
buf ( n6187 , n6186 );
and ( n6188 , n6187 , n376 );
and ( n6189 , n6185 , n6188 );
xor ( n6190 , n6185 , n6188 );
and ( n6191 , n6187 , n377 );
xor ( n6192 , n5872 , n6177 );
buf ( n6193 , n6192 );
and ( n6194 , n6193 , n376 );
and ( n6195 , n6191 , n6194 );
xor ( n6196 , n6191 , n6194 );
and ( n6197 , n6193 , n377 );
xor ( n6198 , n5949 , n6175 );
buf ( n6199 , n6198 );
and ( n6200 , n6199 , n376 );
and ( n6201 , n6197 , n6200 );
xor ( n6202 , n6197 , n6200 );
and ( n6203 , n6199 , n377 );
xor ( n6204 , n6087 , n6173 );
buf ( n6205 , n6204 );
and ( n6206 , n6205 , n376 );
and ( n6207 , n6203 , n6206 );
xor ( n6208 , n6203 , n6206 );
and ( n6209 , n6205 , n377 );
xor ( n6210 , n6090 , n6171 );
buf ( n6211 , n6210 );
and ( n6212 , n6211 , n376 );
and ( n6213 , n6209 , n6212 );
xor ( n6214 , n6209 , n6212 );
and ( n6215 , n6211 , n377 );
xor ( n6216 , n6093 , n6169 );
buf ( n6217 , n6216 );
and ( n6218 , n6217 , n376 );
and ( n6219 , n6215 , n6218 );
xor ( n6220 , n6215 , n6218 );
and ( n6221 , n6217 , n377 );
xor ( n6222 , n6095 , n6168 );
buf ( n6223 , n6222 );
and ( n6224 , n6223 , n376 );
and ( n6225 , n6221 , n6224 );
xor ( n6226 , n6221 , n6224 );
and ( n6227 , n6223 , n377 );
xor ( n6228 , n6146 , n6166 );
buf ( n6229 , n6228 );
and ( n6230 , n6229 , n376 );
and ( n6231 , n6227 , n6230 );
xor ( n6232 , n6227 , n6230 );
and ( n6233 , n6229 , n377 );
xor ( n6234 , n6149 , n6164 );
buf ( n6235 , n6234 );
and ( n6236 , n6235 , n376 );
and ( n6237 , n6233 , n6236 );
xor ( n6238 , n6233 , n6236 );
and ( n6239 , n6235 , n377 );
xor ( n6240 , n6150 , n6163 );
buf ( n6241 , n6240 );
and ( n6242 , n6241 , n376 );
and ( n6243 , n6239 , n6242 );
xor ( n6244 , n6239 , n6242 );
and ( n6245 , n6241 , n377 );
xor ( n6246 , n6152 , n6162 );
buf ( n6247 , n6246 );
and ( n6248 , n6247 , n376 );
and ( n6249 , n6245 , n6248 );
xor ( n6250 , n6245 , n6248 );
and ( n6251 , n6247 , n377 );
xor ( n6252 , n6159 , n6161 );
buf ( n6253 , n6252 );
and ( n6254 , n6253 , n376 );
and ( n6255 , n6251 , n6254 );
xor ( n6256 , n6251 , n6254 );
and ( n6257 , n6253 , n377 );
xor ( n6258 , n6153 , n6154 );
xor ( n6259 , n6258 , n6156 );
buf ( n6260 , n6259 );
and ( n6261 , n6260 , n376 );
and ( n6262 , n6257 , n6261 );
buf ( n6263 , n6262 );
and ( n6264 , n6256 , n6263 );
or ( n6265 , n6255 , n6264 );
and ( n6266 , n6250 , n6265 );
or ( n6267 , n6249 , n6266 );
and ( n6268 , n6244 , n6267 );
or ( n6269 , n6243 , n6268 );
and ( n6270 , n6238 , n6269 );
or ( n6271 , n6237 , n6270 );
and ( n6272 , n6232 , n6271 );
or ( n6273 , n6231 , n6272 );
and ( n6274 , n6226 , n6273 );
or ( n6275 , n6225 , n6274 );
and ( n6276 , n6220 , n6275 );
or ( n6277 , n6219 , n6276 );
and ( n6278 , n6214 , n6277 );
or ( n6279 , n6213 , n6278 );
and ( n6280 , n6208 , n6279 );
or ( n6281 , n6207 , n6280 );
and ( n6282 , n6202 , n6281 );
or ( n6283 , n6201 , n6282 );
and ( n6284 , n6196 , n6283 );
or ( n6285 , n6195 , n6284 );
and ( n6286 , n6190 , n6285 );
or ( n6287 , n6189 , n6286 );
and ( n6288 , n6184 , n6287 );
buf ( n6289 , n6288 );
buf ( n6290 , n6289 );
and ( n6291 , n6182 , n375 );
and ( n6292 , n6290 , n6291 );
xor ( n6293 , n6290 , n6291 );
xor ( n6294 , n6184 , n6287 );
and ( n6295 , n6187 , n375 );
and ( n6296 , n6294 , n6295 );
xor ( n6297 , n6294 , n6295 );
xor ( n6298 , n6190 , n6285 );
and ( n6299 , n6193 , n375 );
and ( n6300 , n6298 , n6299 );
xor ( n6301 , n6298 , n6299 );
xor ( n6302 , n6196 , n6283 );
and ( n6303 , n6199 , n375 );
and ( n6304 , n6302 , n6303 );
xor ( n6305 , n6302 , n6303 );
xor ( n6306 , n6202 , n6281 );
and ( n6307 , n6205 , n375 );
and ( n6308 , n6306 , n6307 );
xor ( n6309 , n6306 , n6307 );
xor ( n6310 , n6208 , n6279 );
and ( n6311 , n6211 , n375 );
and ( n6312 , n6310 , n6311 );
xor ( n6313 , n6310 , n6311 );
xor ( n6314 , n6214 , n6277 );
and ( n6315 , n6217 , n375 );
and ( n6316 , n6314 , n6315 );
xor ( n6317 , n6314 , n6315 );
xor ( n6318 , n6220 , n6275 );
and ( n6319 , n6223 , n375 );
and ( n6320 , n6318 , n6319 );
xor ( n6321 , n6318 , n6319 );
xor ( n6322 , n6226 , n6273 );
and ( n6323 , n6229 , n375 );
and ( n6324 , n6322 , n6323 );
xor ( n6325 , n6322 , n6323 );
xor ( n6326 , n6232 , n6271 );
and ( n6327 , n6235 , n375 );
and ( n6328 , n6326 , n6327 );
xor ( n6329 , n6326 , n6327 );
xor ( n6330 , n6238 , n6269 );
and ( n6331 , n6241 , n375 );
and ( n6332 , n6330 , n6331 );
xor ( n6333 , n6330 , n6331 );
xor ( n6334 , n6244 , n6267 );
and ( n6335 , n6247 , n375 );
and ( n6336 , n6334 , n6335 );
xor ( n6337 , n6334 , n6335 );
xor ( n6338 , n6250 , n6265 );
and ( n6339 , n6253 , n375 );
and ( n6340 , n6338 , n6339 );
xor ( n6341 , n6338 , n6339 );
xor ( n6342 , n6256 , n6263 );
and ( n6343 , n6260 , n375 );
and ( n6344 , n6342 , n6343 );
xor ( n6345 , n6342 , n6343 );
xor ( n6346 , n6257 , n6261 );
buf ( n6347 , n6346 );
buf ( n6348 , n6347 );
and ( n6349 , n6260 , n377 );
buf ( n6350 , n6349 );
buf ( n6351 , n6350 );
buf ( n6352 , n5914 );
buf ( n6353 , n6352 );
and ( n6354 , n6353 , n375 );
and ( n6355 , n6351 , n6354 );
and ( n6356 , n6348 , n6355 );
buf ( n6357 , n6356 );
and ( n6358 , n6345 , n6357 );
or ( n6359 , n6344 , n6358 );
and ( n6360 , n6341 , n6359 );
or ( n6361 , n6340 , n6360 );
and ( n6362 , n6337 , n6361 );
or ( n6363 , n6336 , n6362 );
and ( n6364 , n6333 , n6363 );
or ( n6365 , n6332 , n6364 );
and ( n6366 , n6329 , n6365 );
or ( n6367 , n6328 , n6366 );
and ( n6368 , n6325 , n6367 );
or ( n6369 , n6324 , n6368 );
and ( n6370 , n6321 , n6369 );
or ( n6371 , n6320 , n6370 );
and ( n6372 , n6317 , n6371 );
or ( n6373 , n6316 , n6372 );
and ( n6374 , n6313 , n6373 );
or ( n6375 , n6312 , n6374 );
and ( n6376 , n6309 , n6375 );
or ( n6377 , n6308 , n6376 );
and ( n6378 , n6305 , n6377 );
or ( n6379 , n6304 , n6378 );
and ( n6380 , n6301 , n6379 );
or ( n6381 , n6300 , n6380 );
and ( n6382 , n6297 , n6381 );
or ( n6383 , n6296 , n6382 );
and ( n6384 , n6293 , n6383 );
or ( n6385 , n6292 , n6384 );
buf ( n6386 , n6385 );
and ( n6387 , n6182 , n374 );
and ( n6388 , n6386 , n6387 );
xor ( n6389 , n6386 , n6387 );
xor ( n6390 , n6293 , n6383 );
and ( n6391 , n6187 , n374 );
and ( n6392 , n6390 , n6391 );
xor ( n6393 , n6390 , n6391 );
xor ( n6394 , n6297 , n6381 );
and ( n6395 , n6193 , n374 );
and ( n6396 , n6394 , n6395 );
xor ( n6397 , n6394 , n6395 );
xor ( n6398 , n6301 , n6379 );
and ( n6399 , n6199 , n374 );
and ( n6400 , n6398 , n6399 );
xor ( n6401 , n6398 , n6399 );
xor ( n6402 , n6305 , n6377 );
and ( n6403 , n6205 , n374 );
and ( n6404 , n6402 , n6403 );
xor ( n6405 , n6402 , n6403 );
xor ( n6406 , n6309 , n6375 );
and ( n6407 , n6211 , n374 );
and ( n6408 , n6406 , n6407 );
xor ( n6409 , n6406 , n6407 );
xor ( n6410 , n6313 , n6373 );
and ( n6411 , n6217 , n374 );
and ( n6412 , n6410 , n6411 );
xor ( n6413 , n6410 , n6411 );
xor ( n6414 , n6317 , n6371 );
and ( n6415 , n6223 , n374 );
and ( n6416 , n6414 , n6415 );
xor ( n6417 , n6414 , n6415 );
xor ( n6418 , n6321 , n6369 );
and ( n6419 , n6229 , n374 );
and ( n6420 , n6418 , n6419 );
xor ( n6421 , n6418 , n6419 );
xor ( n6422 , n6325 , n6367 );
and ( n6423 , n6235 , n374 );
and ( n6424 , n6422 , n6423 );
xor ( n6425 , n6422 , n6423 );
xor ( n6426 , n6329 , n6365 );
and ( n6427 , n6241 , n374 );
and ( n6428 , n6426 , n6427 );
xor ( n6429 , n6426 , n6427 );
xor ( n6430 , n6333 , n6363 );
and ( n6431 , n6247 , n374 );
and ( n6432 , n6430 , n6431 );
xor ( n6433 , n6430 , n6431 );
xor ( n6434 , n6337 , n6361 );
and ( n6435 , n6253 , n374 );
and ( n6436 , n6434 , n6435 );
xor ( n6437 , n6434 , n6435 );
xor ( n6438 , n6341 , n6359 );
and ( n6439 , n6260 , n374 );
and ( n6440 , n6438 , n6439 );
xor ( n6441 , n6438 , n6439 );
xor ( n6442 , n6345 , n6357 );
buf ( n6443 , n6442 );
xor ( n6444 , n6348 , n6355 );
and ( n6445 , n6353 , n374 );
and ( n6446 , n6444 , n6445 );
and ( n6447 , n6443 , n6446 );
buf ( n6448 , n6447 );
and ( n6449 , n6441 , n6448 );
or ( n6450 , n6440 , n6449 );
and ( n6451 , n6437 , n6450 );
or ( n6452 , n6436 , n6451 );
and ( n6453 , n6433 , n6452 );
or ( n6454 , n6432 , n6453 );
and ( n6455 , n6429 , n6454 );
or ( n6456 , n6428 , n6455 );
and ( n6457 , n6425 , n6456 );
or ( n6458 , n6424 , n6457 );
and ( n6459 , n6421 , n6458 );
or ( n6460 , n6420 , n6459 );
and ( n6461 , n6417 , n6460 );
or ( n6462 , n6416 , n6461 );
and ( n6463 , n6413 , n6462 );
or ( n6464 , n6412 , n6463 );
and ( n6465 , n6409 , n6464 );
or ( n6466 , n6408 , n6465 );
and ( n6467 , n6405 , n6466 );
or ( n6468 , n6404 , n6467 );
and ( n6469 , n6401 , n6468 );
or ( n6470 , n6400 , n6469 );
and ( n6471 , n6397 , n6470 );
or ( n6472 , n6396 , n6471 );
and ( n6473 , n6393 , n6472 );
or ( n6474 , n6392 , n6473 );
and ( n6475 , n6389 , n6474 );
or ( n6476 , n6388 , n6475 );
buf ( n6477 , n6476 );
and ( n6478 , n6182 , n373 );
and ( n6479 , n6477 , n6478 );
xor ( n6480 , n6477 , n6478 );
xor ( n6481 , n6389 , n6474 );
and ( n6482 , n6187 , n373 );
and ( n6483 , n6481 , n6482 );
xor ( n6484 , n6481 , n6482 );
xor ( n6485 , n6393 , n6472 );
and ( n6486 , n6193 , n373 );
and ( n6487 , n6485 , n6486 );
xor ( n6488 , n6485 , n6486 );
xor ( n6489 , n6397 , n6470 );
and ( n6490 , n6199 , n373 );
and ( n6491 , n6489 , n6490 );
xor ( n6492 , n6489 , n6490 );
xor ( n6493 , n6401 , n6468 );
and ( n6494 , n6205 , n373 );
and ( n6495 , n6493 , n6494 );
xor ( n6496 , n6493 , n6494 );
xor ( n6497 , n6405 , n6466 );
and ( n6498 , n6211 , n373 );
and ( n6499 , n6497 , n6498 );
xor ( n6500 , n6497 , n6498 );
xor ( n6501 , n6409 , n6464 );
and ( n6502 , n6217 , n373 );
and ( n6503 , n6501 , n6502 );
xor ( n6504 , n6501 , n6502 );
xor ( n6505 , n6413 , n6462 );
and ( n6506 , n6223 , n373 );
and ( n6507 , n6505 , n6506 );
xor ( n6508 , n6505 , n6506 );
xor ( n6509 , n6417 , n6460 );
and ( n6510 , n6229 , n373 );
and ( n6511 , n6509 , n6510 );
xor ( n6512 , n6509 , n6510 );
xor ( n6513 , n6421 , n6458 );
and ( n6514 , n6235 , n373 );
and ( n6515 , n6513 , n6514 );
xor ( n6516 , n6513 , n6514 );
xor ( n6517 , n6425 , n6456 );
and ( n6518 , n6241 , n373 );
and ( n6519 , n6517 , n6518 );
xor ( n6520 , n6517 , n6518 );
xor ( n6521 , n6429 , n6454 );
and ( n6522 , n6247 , n373 );
and ( n6523 , n6521 , n6522 );
xor ( n6524 , n6521 , n6522 );
xor ( n6525 , n6433 , n6452 );
and ( n6526 , n6253 , n373 );
and ( n6527 , n6525 , n6526 );
xor ( n6528 , n6525 , n6526 );
xor ( n6529 , n6437 , n6450 );
and ( n6530 , n6260 , n373 );
and ( n6531 , n6529 , n6530 );
xor ( n6532 , n6529 , n6530 );
xor ( n6533 , n6441 , n6448 );
buf ( n6534 , n6533 );
xor ( n6535 , n6443 , n6446 );
and ( n6536 , n6353 , n373 );
and ( n6537 , n6535 , n6536 );
and ( n6538 , n6534 , n6537 );
buf ( n6539 , n6538 );
and ( n6540 , n6532 , n6539 );
or ( n6541 , n6531 , n6540 );
and ( n6542 , n6528 , n6541 );
or ( n6543 , n6527 , n6542 );
and ( n6544 , n6524 , n6543 );
or ( n6545 , n6523 , n6544 );
and ( n6546 , n6520 , n6545 );
or ( n6547 , n6519 , n6546 );
and ( n6548 , n6516 , n6547 );
or ( n6549 , n6515 , n6548 );
and ( n6550 , n6512 , n6549 );
or ( n6551 , n6511 , n6550 );
and ( n6552 , n6508 , n6551 );
or ( n6553 , n6507 , n6552 );
and ( n6554 , n6504 , n6553 );
or ( n6555 , n6503 , n6554 );
and ( n6556 , n6500 , n6555 );
or ( n6557 , n6499 , n6556 );
and ( n6558 , n6496 , n6557 );
or ( n6559 , n6495 , n6558 );
and ( n6560 , n6492 , n6559 );
or ( n6561 , n6491 , n6560 );
and ( n6562 , n6488 , n6561 );
or ( n6563 , n6487 , n6562 );
and ( n6564 , n6484 , n6563 );
or ( n6565 , n6483 , n6564 );
and ( n6566 , n6480 , n6565 );
or ( n6567 , n6479 , n6566 );
buf ( n6568 , n6567 );
and ( n6569 , n6182 , n372 );
and ( n6570 , n6568 , n6569 );
xor ( n6571 , n6568 , n6569 );
xor ( n6572 , n6480 , n6565 );
and ( n6573 , n6187 , n372 );
and ( n6574 , n6572 , n6573 );
xor ( n6575 , n6572 , n6573 );
xor ( n6576 , n6484 , n6563 );
and ( n6577 , n6193 , n372 );
and ( n6578 , n6576 , n6577 );
xor ( n6579 , n6576 , n6577 );
xor ( n6580 , n6488 , n6561 );
and ( n6581 , n6199 , n372 );
and ( n6582 , n6580 , n6581 );
xor ( n6583 , n6580 , n6581 );
xor ( n6584 , n6492 , n6559 );
and ( n6585 , n6205 , n372 );
and ( n6586 , n6584 , n6585 );
xor ( n6587 , n6584 , n6585 );
xor ( n6588 , n6496 , n6557 );
and ( n6589 , n6211 , n372 );
and ( n6590 , n6588 , n6589 );
xor ( n6591 , n6588 , n6589 );
xor ( n6592 , n6500 , n6555 );
and ( n6593 , n6217 , n372 );
and ( n6594 , n6592 , n6593 );
xor ( n6595 , n6592 , n6593 );
xor ( n6596 , n6504 , n6553 );
and ( n6597 , n6223 , n372 );
and ( n6598 , n6596 , n6597 );
xor ( n6599 , n6596 , n6597 );
xor ( n6600 , n6508 , n6551 );
and ( n6601 , n6229 , n372 );
and ( n6602 , n6600 , n6601 );
xor ( n6603 , n6600 , n6601 );
xor ( n6604 , n6512 , n6549 );
and ( n6605 , n6235 , n372 );
and ( n6606 , n6604 , n6605 );
xor ( n6607 , n6604 , n6605 );
xor ( n6608 , n6516 , n6547 );
and ( n6609 , n6241 , n372 );
and ( n6610 , n6608 , n6609 );
xor ( n6611 , n6608 , n6609 );
xor ( n6612 , n6520 , n6545 );
and ( n6613 , n6247 , n372 );
and ( n6614 , n6612 , n6613 );
xor ( n6615 , n6612 , n6613 );
xor ( n6616 , n6524 , n6543 );
and ( n6617 , n6253 , n372 );
and ( n6618 , n6616 , n6617 );
xor ( n6619 , n6616 , n6617 );
xor ( n6620 , n6528 , n6541 );
and ( n6621 , n6260 , n372 );
and ( n6622 , n6620 , n6621 );
xor ( n6623 , n6620 , n6621 );
xor ( n6624 , n6532 , n6539 );
buf ( n6625 , n6624 );
xor ( n6626 , n6534 , n6537 );
and ( n6627 , n6353 , n372 );
and ( n6628 , n6626 , n6627 );
and ( n6629 , n6625 , n6628 );
buf ( n6630 , n6629 );
and ( n6631 , n6623 , n6630 );
or ( n6632 , n6622 , n6631 );
and ( n6633 , n6619 , n6632 );
or ( n6634 , n6618 , n6633 );
and ( n6635 , n6615 , n6634 );
or ( n6636 , n6614 , n6635 );
and ( n6637 , n6611 , n6636 );
or ( n6638 , n6610 , n6637 );
and ( n6639 , n6607 , n6638 );
or ( n6640 , n6606 , n6639 );
and ( n6641 , n6603 , n6640 );
or ( n6642 , n6602 , n6641 );
and ( n6643 , n6599 , n6642 );
or ( n6644 , n6598 , n6643 );
and ( n6645 , n6595 , n6644 );
or ( n6646 , n6594 , n6645 );
and ( n6647 , n6591 , n6646 );
or ( n6648 , n6590 , n6647 );
and ( n6649 , n6587 , n6648 );
or ( n6650 , n6586 , n6649 );
and ( n6651 , n6583 , n6650 );
or ( n6652 , n6582 , n6651 );
and ( n6653 , n6579 , n6652 );
or ( n6654 , n6578 , n6653 );
and ( n6655 , n6575 , n6654 );
or ( n6656 , n6574 , n6655 );
and ( n6657 , n6571 , n6656 );
or ( n6658 , n6570 , n6657 );
buf ( n6659 , n6658 );
and ( n6660 , n6182 , n371 );
and ( n6661 , n6659 , n6660 );
xor ( n6662 , n6659 , n6660 );
xor ( n6663 , n6571 , n6656 );
and ( n6664 , n6187 , n371 );
and ( n6665 , n6663 , n6664 );
xor ( n6666 , n6663 , n6664 );
xor ( n6667 , n6575 , n6654 );
and ( n6668 , n6193 , n371 );
and ( n6669 , n6667 , n6668 );
xor ( n6670 , n6667 , n6668 );
xor ( n6671 , n6579 , n6652 );
and ( n6672 , n6199 , n371 );
and ( n6673 , n6671 , n6672 );
xor ( n6674 , n6671 , n6672 );
xor ( n6675 , n6583 , n6650 );
and ( n6676 , n6205 , n371 );
and ( n6677 , n6675 , n6676 );
xor ( n6678 , n6675 , n6676 );
xor ( n6679 , n6587 , n6648 );
and ( n6680 , n6211 , n371 );
and ( n6681 , n6679 , n6680 );
xor ( n6682 , n6679 , n6680 );
xor ( n6683 , n6591 , n6646 );
and ( n6684 , n6217 , n371 );
and ( n6685 , n6683 , n6684 );
xor ( n6686 , n6683 , n6684 );
xor ( n6687 , n6595 , n6644 );
and ( n6688 , n6223 , n371 );
and ( n6689 , n6687 , n6688 );
xor ( n6690 , n6687 , n6688 );
xor ( n6691 , n6599 , n6642 );
and ( n6692 , n6229 , n371 );
and ( n6693 , n6691 , n6692 );
xor ( n6694 , n6691 , n6692 );
xor ( n6695 , n6603 , n6640 );
and ( n6696 , n6235 , n371 );
and ( n6697 , n6695 , n6696 );
xor ( n6698 , n6695 , n6696 );
xor ( n6699 , n6607 , n6638 );
and ( n6700 , n6241 , n371 );
and ( n6701 , n6699 , n6700 );
xor ( n6702 , n6699 , n6700 );
xor ( n6703 , n6611 , n6636 );
and ( n6704 , n6247 , n371 );
and ( n6705 , n6703 , n6704 );
xor ( n6706 , n6703 , n6704 );
xor ( n6707 , n6615 , n6634 );
and ( n6708 , n6253 , n371 );
and ( n6709 , n6707 , n6708 );
xor ( n6710 , n6707 , n6708 );
xor ( n6711 , n6619 , n6632 );
and ( n6712 , n6260 , n371 );
and ( n6713 , n6711 , n6712 );
xor ( n6714 , n6711 , n6712 );
xor ( n6715 , n6623 , n6630 );
buf ( n6716 , n6715 );
xor ( n6717 , n6625 , n6628 );
and ( n6718 , n6353 , n371 );
and ( n6719 , n6717 , n6718 );
and ( n6720 , n6716 , n6719 );
buf ( n6721 , n6720 );
and ( n6722 , n6714 , n6721 );
or ( n6723 , n6713 , n6722 );
and ( n6724 , n6710 , n6723 );
or ( n6725 , n6709 , n6724 );
and ( n6726 , n6706 , n6725 );
or ( n6727 , n6705 , n6726 );
and ( n6728 , n6702 , n6727 );
or ( n6729 , n6701 , n6728 );
and ( n6730 , n6698 , n6729 );
or ( n6731 , n6697 , n6730 );
and ( n6732 , n6694 , n6731 );
or ( n6733 , n6693 , n6732 );
and ( n6734 , n6690 , n6733 );
or ( n6735 , n6689 , n6734 );
and ( n6736 , n6686 , n6735 );
or ( n6737 , n6685 , n6736 );
and ( n6738 , n6682 , n6737 );
or ( n6739 , n6681 , n6738 );
and ( n6740 , n6678 , n6739 );
or ( n6741 , n6677 , n6740 );
and ( n6742 , n6674 , n6741 );
or ( n6743 , n6673 , n6742 );
and ( n6744 , n6670 , n6743 );
or ( n6745 , n6669 , n6744 );
and ( n6746 , n6666 , n6745 );
or ( n6747 , n6665 , n6746 );
and ( n6748 , n6662 , n6747 );
or ( n6749 , n6661 , n6748 );
buf ( n6750 , n6749 );
and ( n6751 , n6182 , n370 );
and ( n6752 , n6750 , n6751 );
xor ( n6753 , n6750 , n6751 );
xor ( n6754 , n6662 , n6747 );
and ( n6755 , n6187 , n370 );
and ( n6756 , n6754 , n6755 );
xor ( n6757 , n6754 , n6755 );
xor ( n6758 , n6666 , n6745 );
and ( n6759 , n6193 , n370 );
and ( n6760 , n6758 , n6759 );
xor ( n6761 , n6758 , n6759 );
xor ( n6762 , n6670 , n6743 );
and ( n6763 , n6199 , n370 );
and ( n6764 , n6762 , n6763 );
xor ( n6765 , n6762 , n6763 );
xor ( n6766 , n6674 , n6741 );
and ( n6767 , n6205 , n370 );
and ( n6768 , n6766 , n6767 );
xor ( n6769 , n6766 , n6767 );
xor ( n6770 , n6678 , n6739 );
and ( n6771 , n6211 , n370 );
and ( n6772 , n6770 , n6771 );
xor ( n6773 , n6770 , n6771 );
xor ( n6774 , n6682 , n6737 );
and ( n6775 , n6217 , n370 );
and ( n6776 , n6774 , n6775 );
xor ( n6777 , n6774 , n6775 );
xor ( n6778 , n6686 , n6735 );
and ( n6779 , n6223 , n370 );
and ( n6780 , n6778 , n6779 );
xor ( n6781 , n6778 , n6779 );
xor ( n6782 , n6690 , n6733 );
and ( n6783 , n6229 , n370 );
and ( n6784 , n6782 , n6783 );
xor ( n6785 , n6782 , n6783 );
xor ( n6786 , n6694 , n6731 );
and ( n6787 , n6235 , n370 );
and ( n6788 , n6786 , n6787 );
xor ( n6789 , n6786 , n6787 );
xor ( n6790 , n6698 , n6729 );
and ( n6791 , n6241 , n370 );
and ( n6792 , n6790 , n6791 );
xor ( n6793 , n6790 , n6791 );
xor ( n6794 , n6702 , n6727 );
and ( n6795 , n6247 , n370 );
and ( n6796 , n6794 , n6795 );
xor ( n6797 , n6794 , n6795 );
xor ( n6798 , n6706 , n6725 );
and ( n6799 , n6253 , n370 );
and ( n6800 , n6798 , n6799 );
xor ( n6801 , n6798 , n6799 );
xor ( n6802 , n6710 , n6723 );
and ( n6803 , n6260 , n370 );
and ( n6804 , n6802 , n6803 );
xor ( n6805 , n6802 , n6803 );
xor ( n6806 , n6714 , n6721 );
buf ( n6807 , n6806 );
xor ( n6808 , n6716 , n6719 );
and ( n6809 , n6353 , n370 );
and ( n6810 , n6808 , n6809 );
and ( n6811 , n6807 , n6810 );
buf ( n6812 , n6811 );
and ( n6813 , n6805 , n6812 );
or ( n6814 , n6804 , n6813 );
and ( n6815 , n6801 , n6814 );
or ( n6816 , n6800 , n6815 );
and ( n6817 , n6797 , n6816 );
or ( n6818 , n6796 , n6817 );
and ( n6819 , n6793 , n6818 );
or ( n6820 , n6792 , n6819 );
and ( n6821 , n6789 , n6820 );
or ( n6822 , n6788 , n6821 );
and ( n6823 , n6785 , n6822 );
or ( n6824 , n6784 , n6823 );
and ( n6825 , n6781 , n6824 );
or ( n6826 , n6780 , n6825 );
and ( n6827 , n6777 , n6826 );
or ( n6828 , n6776 , n6827 );
and ( n6829 , n6773 , n6828 );
or ( n6830 , n6772 , n6829 );
and ( n6831 , n6769 , n6830 );
or ( n6832 , n6768 , n6831 );
and ( n6833 , n6765 , n6832 );
or ( n6834 , n6764 , n6833 );
and ( n6835 , n6761 , n6834 );
or ( n6836 , n6760 , n6835 );
and ( n6837 , n6757 , n6836 );
or ( n6838 , n6756 , n6837 );
and ( n6839 , n6753 , n6838 );
or ( n6840 , n6752 , n6839 );
buf ( n6841 , n6840 );
and ( n6842 , n6841 , n376 );
buf ( n6843 , n6842 );
and ( n6844 , n6841 , n377 );
xor ( n6845 , n6753 , n6838 );
and ( n6846 , n6845 , n376 );
and ( n6847 , n6844 , n6846 );
xor ( n6848 , n6844 , n6846 );
and ( n6849 , n6845 , n377 );
xor ( n6850 , n6757 , n6836 );
and ( n6851 , n6850 , n376 );
and ( n6852 , n6849 , n6851 );
xor ( n6853 , n6849 , n6851 );
and ( n6854 , n6850 , n377 );
xor ( n6855 , n6761 , n6834 );
and ( n6856 , n6855 , n376 );
and ( n6857 , n6854 , n6856 );
xor ( n6858 , n6854 , n6856 );
and ( n6859 , n6855 , n377 );
xor ( n6860 , n6765 , n6832 );
and ( n6861 , n6860 , n376 );
and ( n6862 , n6859 , n6861 );
xor ( n6863 , n6859 , n6861 );
and ( n6864 , n6860 , n377 );
xor ( n6865 , n6769 , n6830 );
and ( n6866 , n6865 , n376 );
and ( n6867 , n6864 , n6866 );
xor ( n6868 , n6864 , n6866 );
and ( n6869 , n6865 , n377 );
xor ( n6870 , n6773 , n6828 );
and ( n6871 , n6870 , n376 );
and ( n6872 , n6869 , n6871 );
xor ( n6873 , n6869 , n6871 );
and ( n6874 , n6870 , n377 );
xor ( n6875 , n6777 , n6826 );
and ( n6876 , n6875 , n376 );
and ( n6877 , n6874 , n6876 );
xor ( n6878 , n6874 , n6876 );
and ( n6879 , n6875 , n377 );
xor ( n6880 , n6781 , n6824 );
and ( n6881 , n6880 , n376 );
and ( n6882 , n6879 , n6881 );
xor ( n6883 , n6879 , n6881 );
and ( n6884 , n6880 , n377 );
xor ( n6885 , n6785 , n6822 );
and ( n6886 , n6885 , n376 );
and ( n6887 , n6884 , n6886 );
xor ( n6888 , n6884 , n6886 );
and ( n6889 , n6885 , n377 );
xor ( n6890 , n6789 , n6820 );
and ( n6891 , n6890 , n376 );
and ( n6892 , n6889 , n6891 );
xor ( n6893 , n6889 , n6891 );
and ( n6894 , n6890 , n377 );
xor ( n6895 , n6793 , n6818 );
and ( n6896 , n6895 , n376 );
and ( n6897 , n6894 , n6896 );
xor ( n6898 , n6894 , n6896 );
and ( n6899 , n6895 , n377 );
xor ( n6900 , n6797 , n6816 );
and ( n6901 , n6900 , n376 );
and ( n6902 , n6899 , n6901 );
xor ( n6903 , n6899 , n6901 );
and ( n6904 , n6900 , n377 );
xor ( n6905 , n6801 , n6814 );
and ( n6906 , n6905 , n376 );
and ( n6907 , n6904 , n6906 );
xor ( n6908 , n6904 , n6906 );
and ( n6909 , n6905 , n377 );
xor ( n6910 , n6805 , n6812 );
and ( n6911 , n6910 , n376 );
and ( n6912 , n6909 , n6911 );
xor ( n6913 , n6909 , n6911 );
and ( n6914 , n6910 , n377 );
xor ( n6915 , n6807 , n6810 );
and ( n6916 , n6915 , n376 );
and ( n6917 , n6914 , n6916 );
xor ( n6918 , n6914 , n6916 );
and ( n6919 , n6915 , n377 );
xor ( n6920 , n6808 , n6809 );
and ( n6921 , n6920 , n376 );
and ( n6922 , n6919 , n6921 );
xor ( n6923 , n6919 , n6921 );
and ( n6924 , n6920 , n377 );
xor ( n6925 , n6717 , n6718 );
and ( n6926 , n6925 , n376 );
and ( n6927 , n6924 , n6926 );
xor ( n6928 , n6924 , n6926 );
and ( n6929 , n6925 , n377 );
xor ( n6930 , n6626 , n6627 );
and ( n6931 , n6930 , n376 );
and ( n6932 , n6929 , n6931 );
xor ( n6933 , n6929 , n6931 );
and ( n6934 , n6930 , n377 );
xor ( n6935 , n6535 , n6536 );
and ( n6936 , n6935 , n376 );
and ( n6937 , n6934 , n6936 );
xor ( n6938 , n6934 , n6936 );
and ( n6939 , n6935 , n377 );
xor ( n6940 , n6444 , n6445 );
and ( n6941 , n6940 , n376 );
and ( n6942 , n6939 , n6941 );
xor ( n6943 , n6939 , n6941 );
and ( n6944 , n6940 , n377 );
xor ( n6945 , n6351 , n6354 );
and ( n6946 , n6945 , n376 );
and ( n6947 , n6944 , n6946 );
xor ( n6948 , n6944 , n6946 );
and ( n6949 , n6945 , n377 );
and ( n6950 , n6353 , n376 );
buf ( n6951 , n6950 );
and ( n6952 , n6951 , n376 );
and ( n6953 , n6949 , n6952 );
xor ( n6954 , n6949 , n6952 );
and ( n6955 , n6951 , n377 );
buf ( n6956 , n6353 );
and ( n6957 , n6956 , n376 );
and ( n6958 , n6955 , n6957 );
and ( n6959 , n6954 , n6958 );
or ( n6960 , n6953 , n6959 );
and ( n6961 , n6948 , n6960 );
or ( n6962 , n6947 , n6961 );
and ( n6963 , n6943 , n6962 );
or ( n6964 , n6942 , n6963 );
and ( n6965 , n6938 , n6964 );
or ( n6966 , n6937 , n6965 );
and ( n6967 , n6933 , n6966 );
or ( n6968 , n6932 , n6967 );
and ( n6969 , n6928 , n6968 );
or ( n6970 , n6927 , n6969 );
and ( n6971 , n6923 , n6970 );
or ( n6972 , n6922 , n6971 );
and ( n6973 , n6918 , n6972 );
or ( n6974 , n6917 , n6973 );
and ( n6975 , n6913 , n6974 );
or ( n6976 , n6912 , n6975 );
and ( n6977 , n6908 , n6976 );
or ( n6978 , n6907 , n6977 );
and ( n6979 , n6903 , n6978 );
or ( n6980 , n6902 , n6979 );
and ( n6981 , n6898 , n6980 );
or ( n6982 , n6897 , n6981 );
and ( n6983 , n6893 , n6982 );
or ( n6984 , n6892 , n6983 );
and ( n6985 , n6888 , n6984 );
or ( n6986 , n6887 , n6985 );
and ( n6987 , n6883 , n6986 );
or ( n6988 , n6882 , n6987 );
and ( n6989 , n6878 , n6988 );
or ( n6990 , n6877 , n6989 );
and ( n6991 , n6873 , n6990 );
or ( n6992 , n6872 , n6991 );
and ( n6993 , n6868 , n6992 );
or ( n6994 , n6867 , n6993 );
and ( n6995 , n6863 , n6994 );
or ( n6996 , n6862 , n6995 );
and ( n6997 , n6858 , n6996 );
or ( n6998 , n6857 , n6997 );
and ( n6999 , n6853 , n6998 );
or ( n7000 , n6852 , n6999 );
and ( n7001 , n6848 , n7000 );
or ( n7002 , n6847 , n7001 );
and ( n7003 , n6843 , n7002 );
buf ( n7004 , n7003 );
buf ( n7005 , n7004 );
and ( n7006 , n6841 , n375 );
and ( n7007 , n7005 , n7006 );
xor ( n7008 , n7005 , n7006 );
xor ( n7009 , n6843 , n7002 );
and ( n7010 , n6845 , n375 );
and ( n7011 , n7009 , n7010 );
xor ( n7012 , n7009 , n7010 );
xor ( n7013 , n6848 , n7000 );
and ( n7014 , n6850 , n375 );
and ( n7015 , n7013 , n7014 );
xor ( n7016 , n7013 , n7014 );
xor ( n7017 , n6853 , n6998 );
and ( n7018 , n6855 , n375 );
and ( n7019 , n7017 , n7018 );
xor ( n7020 , n7017 , n7018 );
xor ( n7021 , n6858 , n6996 );
and ( n7022 , n6860 , n375 );
and ( n7023 , n7021 , n7022 );
xor ( n7024 , n7021 , n7022 );
xor ( n7025 , n6863 , n6994 );
and ( n7026 , n6865 , n375 );
and ( n7027 , n7025 , n7026 );
xor ( n7028 , n7025 , n7026 );
xor ( n7029 , n6868 , n6992 );
and ( n7030 , n6870 , n375 );
and ( n7031 , n7029 , n7030 );
xor ( n7032 , n7029 , n7030 );
xor ( n7033 , n6873 , n6990 );
and ( n7034 , n6875 , n375 );
and ( n7035 , n7033 , n7034 );
xor ( n7036 , n7033 , n7034 );
xor ( n7037 , n6878 , n6988 );
and ( n7038 , n6880 , n375 );
and ( n7039 , n7037 , n7038 );
xor ( n7040 , n7037 , n7038 );
xor ( n7041 , n6883 , n6986 );
and ( n7042 , n6885 , n375 );
and ( n7043 , n7041 , n7042 );
xor ( n7044 , n7041 , n7042 );
xor ( n7045 , n6888 , n6984 );
and ( n7046 , n6890 , n375 );
and ( n7047 , n7045 , n7046 );
xor ( n7048 , n7045 , n7046 );
xor ( n7049 , n6893 , n6982 );
and ( n7050 , n6895 , n375 );
and ( n7051 , n7049 , n7050 );
xor ( n7052 , n7049 , n7050 );
xor ( n7053 , n6898 , n6980 );
and ( n7054 , n6900 , n375 );
and ( n7055 , n7053 , n7054 );
xor ( n7056 , n7053 , n7054 );
xor ( n7057 , n6903 , n6978 );
and ( n7058 , n6905 , n375 );
and ( n7059 , n7057 , n7058 );
xor ( n7060 , n7057 , n7058 );
xor ( n7061 , n6908 , n6976 );
and ( n7062 , n6910 , n375 );
and ( n7063 , n7061 , n7062 );
xor ( n7064 , n7061 , n7062 );
xor ( n7065 , n6913 , n6974 );
and ( n7066 , n6915 , n375 );
and ( n7067 , n7065 , n7066 );
xor ( n7068 , n7065 , n7066 );
xor ( n7069 , n6918 , n6972 );
and ( n7070 , n6920 , n375 );
and ( n7071 , n7069 , n7070 );
xor ( n7072 , n7069 , n7070 );
xor ( n7073 , n6923 , n6970 );
and ( n7074 , n6925 , n375 );
and ( n7075 , n7073 , n7074 );
xor ( n7076 , n7073 , n7074 );
xor ( n7077 , n6928 , n6968 );
and ( n7078 , n6930 , n375 );
and ( n7079 , n7077 , n7078 );
xor ( n7080 , n7077 , n7078 );
xor ( n7081 , n6933 , n6966 );
and ( n7082 , n6935 , n375 );
and ( n7083 , n7081 , n7082 );
xor ( n7084 , n7081 , n7082 );
xor ( n7085 , n6938 , n6964 );
and ( n7086 , n6940 , n375 );
and ( n7087 , n7085 , n7086 );
xor ( n7088 , n7085 , n7086 );
xor ( n7089 , n6943 , n6962 );
and ( n7090 , n6945 , n375 );
and ( n7091 , n7089 , n7090 );
xor ( n7092 , n7089 , n7090 );
xor ( n7093 , n6948 , n6960 );
and ( n7094 , n6951 , n375 );
and ( n7095 , n7093 , n7094 );
xor ( n7096 , n7093 , n7094 );
xor ( n7097 , n6954 , n6958 );
and ( n7098 , n6956 , n375 );
and ( n7099 , n7097 , n7098 );
and ( n7100 , n7096 , n7099 );
or ( n7101 , n7095 , n7100 );
and ( n7102 , n7092 , n7101 );
or ( n7103 , n7091 , n7102 );
and ( n7104 , n7088 , n7103 );
or ( n7105 , n7087 , n7104 );
and ( n7106 , n7084 , n7105 );
or ( n7107 , n7083 , n7106 );
and ( n7108 , n7080 , n7107 );
or ( n7109 , n7079 , n7108 );
and ( n7110 , n7076 , n7109 );
or ( n7111 , n7075 , n7110 );
and ( n7112 , n7072 , n7111 );
or ( n7113 , n7071 , n7112 );
and ( n7114 , n7068 , n7113 );
or ( n7115 , n7067 , n7114 );
and ( n7116 , n7064 , n7115 );
or ( n7117 , n7063 , n7116 );
and ( n7118 , n7060 , n7117 );
or ( n7119 , n7059 , n7118 );
and ( n7120 , n7056 , n7119 );
or ( n7121 , n7055 , n7120 );
and ( n7122 , n7052 , n7121 );
or ( n7123 , n7051 , n7122 );
and ( n7124 , n7048 , n7123 );
or ( n7125 , n7047 , n7124 );
and ( n7126 , n7044 , n7125 );
or ( n7127 , n7043 , n7126 );
and ( n7128 , n7040 , n7127 );
or ( n7129 , n7039 , n7128 );
and ( n7130 , n7036 , n7129 );
or ( n7131 , n7035 , n7130 );
and ( n7132 , n7032 , n7131 );
or ( n7133 , n7031 , n7132 );
and ( n7134 , n7028 , n7133 );
or ( n7135 , n7027 , n7134 );
and ( n7136 , n7024 , n7135 );
or ( n7137 , n7023 , n7136 );
and ( n7138 , n7020 , n7137 );
or ( n7139 , n7019 , n7138 );
and ( n7140 , n7016 , n7139 );
or ( n7141 , n7015 , n7140 );
and ( n7142 , n7012 , n7141 );
or ( n7143 , n7011 , n7142 );
and ( n7144 , n7008 , n7143 );
or ( n7145 , n7007 , n7144 );
buf ( n7146 , n7145 );
and ( n7147 , n6841 , n374 );
and ( n7148 , n7146 , n7147 );
xor ( n7149 , n7146 , n7147 );
xor ( n7150 , n7008 , n7143 );
and ( n7151 , n6845 , n374 );
and ( n7152 , n7150 , n7151 );
xor ( n7153 , n7150 , n7151 );
xor ( n7154 , n7012 , n7141 );
and ( n7155 , n6850 , n374 );
and ( n7156 , n7154 , n7155 );
xor ( n7157 , n7154 , n7155 );
xor ( n7158 , n7016 , n7139 );
and ( n7159 , n6855 , n374 );
and ( n7160 , n7158 , n7159 );
xor ( n7161 , n7158 , n7159 );
xor ( n7162 , n7020 , n7137 );
and ( n7163 , n6860 , n374 );
and ( n7164 , n7162 , n7163 );
xor ( n7165 , n7162 , n7163 );
xor ( n7166 , n7024 , n7135 );
and ( n7167 , n6865 , n374 );
and ( n7168 , n7166 , n7167 );
xor ( n7169 , n7166 , n7167 );
xor ( n7170 , n7028 , n7133 );
and ( n7171 , n6870 , n374 );
and ( n7172 , n7170 , n7171 );
xor ( n7173 , n7170 , n7171 );
xor ( n7174 , n7032 , n7131 );
and ( n7175 , n6875 , n374 );
and ( n7176 , n7174 , n7175 );
xor ( n7177 , n7174 , n7175 );
xor ( n7178 , n7036 , n7129 );
and ( n7179 , n6880 , n374 );
and ( n7180 , n7178 , n7179 );
xor ( n7181 , n7178 , n7179 );
xor ( n7182 , n7040 , n7127 );
and ( n7183 , n6885 , n374 );
and ( n7184 , n7182 , n7183 );
xor ( n7185 , n7182 , n7183 );
xor ( n7186 , n7044 , n7125 );
and ( n7187 , n6890 , n374 );
and ( n7188 , n7186 , n7187 );
xor ( n7189 , n7186 , n7187 );
xor ( n7190 , n7048 , n7123 );
and ( n7191 , n6895 , n374 );
and ( n7192 , n7190 , n7191 );
xor ( n7193 , n7190 , n7191 );
xor ( n7194 , n7052 , n7121 );
and ( n7195 , n6900 , n374 );
and ( n7196 , n7194 , n7195 );
xor ( n7197 , n7194 , n7195 );
xor ( n7198 , n7056 , n7119 );
and ( n7199 , n6905 , n374 );
and ( n7200 , n7198 , n7199 );
xor ( n7201 , n7198 , n7199 );
xor ( n7202 , n7060 , n7117 );
and ( n7203 , n6910 , n374 );
and ( n7204 , n7202 , n7203 );
xor ( n7205 , n7202 , n7203 );
xor ( n7206 , n7064 , n7115 );
and ( n7207 , n6915 , n374 );
and ( n7208 , n7206 , n7207 );
xor ( n7209 , n7206 , n7207 );
xor ( n7210 , n7068 , n7113 );
and ( n7211 , n6920 , n374 );
and ( n7212 , n7210 , n7211 );
xor ( n7213 , n7210 , n7211 );
xor ( n7214 , n7072 , n7111 );
and ( n7215 , n6925 , n374 );
and ( n7216 , n7214 , n7215 );
xor ( n7217 , n7214 , n7215 );
xor ( n7218 , n7076 , n7109 );
and ( n7219 , n6930 , n374 );
and ( n7220 , n7218 , n7219 );
xor ( n7221 , n7218 , n7219 );
xor ( n7222 , n7080 , n7107 );
and ( n7223 , n6935 , n374 );
and ( n7224 , n7222 , n7223 );
xor ( n7225 , n7222 , n7223 );
xor ( n7226 , n7084 , n7105 );
and ( n7227 , n6940 , n374 );
and ( n7228 , n7226 , n7227 );
xor ( n7229 , n7226 , n7227 );
xor ( n7230 , n7088 , n7103 );
and ( n7231 , n6945 , n374 );
and ( n7232 , n7230 , n7231 );
xor ( n7233 , n7230 , n7231 );
xor ( n7234 , n7092 , n7101 );
and ( n7235 , n6951 , n374 );
and ( n7236 , n7234 , n7235 );
xor ( n7237 , n7234 , n7235 );
xor ( n7238 , n7096 , n7099 );
and ( n7239 , n6956 , n374 );
and ( n7240 , n7238 , n7239 );
and ( n7241 , n7237 , n7240 );
or ( n7242 , n7236 , n7241 );
and ( n7243 , n7233 , n7242 );
or ( n7244 , n7232 , n7243 );
and ( n7245 , n7229 , n7244 );
or ( n7246 , n7228 , n7245 );
and ( n7247 , n7225 , n7246 );
or ( n7248 , n7224 , n7247 );
and ( n7249 , n7221 , n7248 );
or ( n7250 , n7220 , n7249 );
and ( n7251 , n7217 , n7250 );
or ( n7252 , n7216 , n7251 );
and ( n7253 , n7213 , n7252 );
or ( n7254 , n7212 , n7253 );
and ( n7255 , n7209 , n7254 );
or ( n7256 , n7208 , n7255 );
and ( n7257 , n7205 , n7256 );
or ( n7258 , n7204 , n7257 );
and ( n7259 , n7201 , n7258 );
or ( n7260 , n7200 , n7259 );
and ( n7261 , n7197 , n7260 );
or ( n7262 , n7196 , n7261 );
and ( n7263 , n7193 , n7262 );
or ( n7264 , n7192 , n7263 );
and ( n7265 , n7189 , n7264 );
or ( n7266 , n7188 , n7265 );
and ( n7267 , n7185 , n7266 );
or ( n7268 , n7184 , n7267 );
and ( n7269 , n7181 , n7268 );
or ( n7270 , n7180 , n7269 );
and ( n7271 , n7177 , n7270 );
or ( n7272 , n7176 , n7271 );
and ( n7273 , n7173 , n7272 );
or ( n7274 , n7172 , n7273 );
and ( n7275 , n7169 , n7274 );
or ( n7276 , n7168 , n7275 );
and ( n7277 , n7165 , n7276 );
or ( n7278 , n7164 , n7277 );
and ( n7279 , n7161 , n7278 );
or ( n7280 , n7160 , n7279 );
and ( n7281 , n7157 , n7280 );
or ( n7282 , n7156 , n7281 );
and ( n7283 , n7153 , n7282 );
or ( n7284 , n7152 , n7283 );
and ( n7285 , n7149 , n7284 );
or ( n7286 , n7148 , n7285 );
buf ( n7287 , n7286 );
and ( n7288 , n6841 , n373 );
and ( n7289 , n7287 , n7288 );
xor ( n7290 , n7287 , n7288 );
xor ( n7291 , n7149 , n7284 );
and ( n7292 , n6845 , n373 );
and ( n7293 , n7291 , n7292 );
xor ( n7294 , n7291 , n7292 );
xor ( n7295 , n7153 , n7282 );
and ( n7296 , n6850 , n373 );
and ( n7297 , n7295 , n7296 );
xor ( n7298 , n7295 , n7296 );
xor ( n7299 , n7157 , n7280 );
and ( n7300 , n6855 , n373 );
and ( n7301 , n7299 , n7300 );
xor ( n7302 , n7299 , n7300 );
xor ( n7303 , n7161 , n7278 );
and ( n7304 , n6860 , n373 );
and ( n7305 , n7303 , n7304 );
xor ( n7306 , n7303 , n7304 );
xor ( n7307 , n7165 , n7276 );
and ( n7308 , n6865 , n373 );
and ( n7309 , n7307 , n7308 );
xor ( n7310 , n7307 , n7308 );
xor ( n7311 , n7169 , n7274 );
and ( n7312 , n6870 , n373 );
and ( n7313 , n7311 , n7312 );
xor ( n7314 , n7311 , n7312 );
xor ( n7315 , n7173 , n7272 );
and ( n7316 , n6875 , n373 );
and ( n7317 , n7315 , n7316 );
xor ( n7318 , n7315 , n7316 );
xor ( n7319 , n7177 , n7270 );
and ( n7320 , n6880 , n373 );
and ( n7321 , n7319 , n7320 );
xor ( n7322 , n7319 , n7320 );
xor ( n7323 , n7181 , n7268 );
and ( n7324 , n6885 , n373 );
and ( n7325 , n7323 , n7324 );
xor ( n7326 , n7323 , n7324 );
xor ( n7327 , n7185 , n7266 );
and ( n7328 , n6890 , n373 );
and ( n7329 , n7327 , n7328 );
xor ( n7330 , n7327 , n7328 );
xor ( n7331 , n7189 , n7264 );
and ( n7332 , n6895 , n373 );
and ( n7333 , n7331 , n7332 );
xor ( n7334 , n7331 , n7332 );
xor ( n7335 , n7193 , n7262 );
and ( n7336 , n6900 , n373 );
and ( n7337 , n7335 , n7336 );
xor ( n7338 , n7335 , n7336 );
xor ( n7339 , n7197 , n7260 );
and ( n7340 , n6905 , n373 );
and ( n7341 , n7339 , n7340 );
xor ( n7342 , n7339 , n7340 );
xor ( n7343 , n7201 , n7258 );
and ( n7344 , n6910 , n373 );
and ( n7345 , n7343 , n7344 );
xor ( n7346 , n7343 , n7344 );
xor ( n7347 , n7205 , n7256 );
and ( n7348 , n6915 , n373 );
and ( n7349 , n7347 , n7348 );
xor ( n7350 , n7347 , n7348 );
xor ( n7351 , n7209 , n7254 );
and ( n7352 , n6920 , n373 );
and ( n7353 , n7351 , n7352 );
xor ( n7354 , n7351 , n7352 );
xor ( n7355 , n7213 , n7252 );
and ( n7356 , n6925 , n373 );
and ( n7357 , n7355 , n7356 );
xor ( n7358 , n7355 , n7356 );
xor ( n7359 , n7217 , n7250 );
and ( n7360 , n6930 , n373 );
and ( n7361 , n7359 , n7360 );
xor ( n7362 , n7359 , n7360 );
xor ( n7363 , n7221 , n7248 );
and ( n7364 , n6935 , n373 );
and ( n7365 , n7363 , n7364 );
xor ( n7366 , n7363 , n7364 );
xor ( n7367 , n7225 , n7246 );
and ( n7368 , n6940 , n373 );
and ( n7369 , n7367 , n7368 );
xor ( n7370 , n7367 , n7368 );
xor ( n7371 , n7229 , n7244 );
and ( n7372 , n6945 , n373 );
and ( n7373 , n7371 , n7372 );
xor ( n7374 , n7371 , n7372 );
xor ( n7375 , n7233 , n7242 );
and ( n7376 , n6951 , n373 );
and ( n7377 , n7375 , n7376 );
xor ( n7378 , n7375 , n7376 );
xor ( n7379 , n7237 , n7240 );
and ( n7380 , n6956 , n373 );
and ( n7381 , n7379 , n7380 );
and ( n7382 , n7378 , n7381 );
or ( n7383 , n7377 , n7382 );
and ( n7384 , n7374 , n7383 );
or ( n7385 , n7373 , n7384 );
and ( n7386 , n7370 , n7385 );
or ( n7387 , n7369 , n7386 );
and ( n7388 , n7366 , n7387 );
or ( n7389 , n7365 , n7388 );
and ( n7390 , n7362 , n7389 );
or ( n7391 , n7361 , n7390 );
and ( n7392 , n7358 , n7391 );
or ( n7393 , n7357 , n7392 );
and ( n7394 , n7354 , n7393 );
or ( n7395 , n7353 , n7394 );
and ( n7396 , n7350 , n7395 );
or ( n7397 , n7349 , n7396 );
and ( n7398 , n7346 , n7397 );
or ( n7399 , n7345 , n7398 );
and ( n7400 , n7342 , n7399 );
or ( n7401 , n7341 , n7400 );
and ( n7402 , n7338 , n7401 );
or ( n7403 , n7337 , n7402 );
and ( n7404 , n7334 , n7403 );
or ( n7405 , n7333 , n7404 );
and ( n7406 , n7330 , n7405 );
or ( n7407 , n7329 , n7406 );
and ( n7408 , n7326 , n7407 );
or ( n7409 , n7325 , n7408 );
and ( n7410 , n7322 , n7409 );
or ( n7411 , n7321 , n7410 );
and ( n7412 , n7318 , n7411 );
or ( n7413 , n7317 , n7412 );
and ( n7414 , n7314 , n7413 );
or ( n7415 , n7313 , n7414 );
and ( n7416 , n7310 , n7415 );
or ( n7417 , n7309 , n7416 );
and ( n7418 , n7306 , n7417 );
or ( n7419 , n7305 , n7418 );
and ( n7420 , n7302 , n7419 );
or ( n7421 , n7301 , n7420 );
and ( n7422 , n7298 , n7421 );
or ( n7423 , n7297 , n7422 );
and ( n7424 , n7294 , n7423 );
or ( n7425 , n7293 , n7424 );
and ( n7426 , n7290 , n7425 );
or ( n7427 , n7289 , n7426 );
buf ( n7428 , n7427 );
and ( n7429 , n6841 , n372 );
and ( n7430 , n7428 , n7429 );
xor ( n7431 , n7428 , n7429 );
xor ( n7432 , n7290 , n7425 );
and ( n7433 , n6845 , n372 );
and ( n7434 , n7432 , n7433 );
xor ( n7435 , n7432 , n7433 );
xor ( n7436 , n7294 , n7423 );
and ( n7437 , n6850 , n372 );
and ( n7438 , n7436 , n7437 );
xor ( n7439 , n7436 , n7437 );
xor ( n7440 , n7298 , n7421 );
and ( n7441 , n6855 , n372 );
and ( n7442 , n7440 , n7441 );
xor ( n7443 , n7440 , n7441 );
xor ( n7444 , n7302 , n7419 );
and ( n7445 , n6860 , n372 );
and ( n7446 , n7444 , n7445 );
xor ( n7447 , n7444 , n7445 );
xor ( n7448 , n7306 , n7417 );
and ( n7449 , n6865 , n372 );
and ( n7450 , n7448 , n7449 );
xor ( n7451 , n7448 , n7449 );
xor ( n7452 , n7310 , n7415 );
and ( n7453 , n6870 , n372 );
and ( n7454 , n7452 , n7453 );
xor ( n7455 , n7452 , n7453 );
xor ( n7456 , n7314 , n7413 );
and ( n7457 , n6875 , n372 );
and ( n7458 , n7456 , n7457 );
xor ( n7459 , n7456 , n7457 );
xor ( n7460 , n7318 , n7411 );
and ( n7461 , n6880 , n372 );
and ( n7462 , n7460 , n7461 );
xor ( n7463 , n7460 , n7461 );
xor ( n7464 , n7322 , n7409 );
and ( n7465 , n6885 , n372 );
and ( n7466 , n7464 , n7465 );
xor ( n7467 , n7464 , n7465 );
xor ( n7468 , n7326 , n7407 );
and ( n7469 , n6890 , n372 );
and ( n7470 , n7468 , n7469 );
xor ( n7471 , n7468 , n7469 );
xor ( n7472 , n7330 , n7405 );
and ( n7473 , n6895 , n372 );
and ( n7474 , n7472 , n7473 );
xor ( n7475 , n7472 , n7473 );
xor ( n7476 , n7334 , n7403 );
and ( n7477 , n6900 , n372 );
and ( n7478 , n7476 , n7477 );
xor ( n7479 , n7476 , n7477 );
xor ( n7480 , n7338 , n7401 );
and ( n7481 , n6905 , n372 );
and ( n7482 , n7480 , n7481 );
xor ( n7483 , n7480 , n7481 );
xor ( n7484 , n7342 , n7399 );
and ( n7485 , n6910 , n372 );
and ( n7486 , n7484 , n7485 );
xor ( n7487 , n7484 , n7485 );
xor ( n7488 , n7346 , n7397 );
and ( n7489 , n6915 , n372 );
and ( n7490 , n7488 , n7489 );
xor ( n7491 , n7488 , n7489 );
xor ( n7492 , n7350 , n7395 );
and ( n7493 , n6920 , n372 );
and ( n7494 , n7492 , n7493 );
xor ( n7495 , n7492 , n7493 );
xor ( n7496 , n7354 , n7393 );
and ( n7497 , n6925 , n372 );
and ( n7498 , n7496 , n7497 );
xor ( n7499 , n7496 , n7497 );
xor ( n7500 , n7358 , n7391 );
and ( n7501 , n6930 , n372 );
and ( n7502 , n7500 , n7501 );
xor ( n7503 , n7500 , n7501 );
xor ( n7504 , n7362 , n7389 );
and ( n7505 , n6935 , n372 );
and ( n7506 , n7504 , n7505 );
xor ( n7507 , n7504 , n7505 );
xor ( n7508 , n7366 , n7387 );
and ( n7509 , n6940 , n372 );
and ( n7510 , n7508 , n7509 );
xor ( n7511 , n7508 , n7509 );
xor ( n7512 , n7370 , n7385 );
and ( n7513 , n6945 , n372 );
and ( n7514 , n7512 , n7513 );
xor ( n7515 , n7512 , n7513 );
xor ( n7516 , n7374 , n7383 );
and ( n7517 , n6951 , n372 );
and ( n7518 , n7516 , n7517 );
xor ( n7519 , n7516 , n7517 );
xor ( n7520 , n7378 , n7381 );
and ( n7521 , n6956 , n372 );
and ( n7522 , n7520 , n7521 );
and ( n7523 , n7519 , n7522 );
or ( n7524 , n7518 , n7523 );
and ( n7525 , n7515 , n7524 );
or ( n7526 , n7514 , n7525 );
and ( n7527 , n7511 , n7526 );
or ( n7528 , n7510 , n7527 );
and ( n7529 , n7507 , n7528 );
or ( n7530 , n7506 , n7529 );
and ( n7531 , n7503 , n7530 );
or ( n7532 , n7502 , n7531 );
and ( n7533 , n7499 , n7532 );
or ( n7534 , n7498 , n7533 );
and ( n7535 , n7495 , n7534 );
or ( n7536 , n7494 , n7535 );
and ( n7537 , n7491 , n7536 );
or ( n7538 , n7490 , n7537 );
and ( n7539 , n7487 , n7538 );
or ( n7540 , n7486 , n7539 );
and ( n7541 , n7483 , n7540 );
or ( n7542 , n7482 , n7541 );
and ( n7543 , n7479 , n7542 );
or ( n7544 , n7478 , n7543 );
and ( n7545 , n7475 , n7544 );
or ( n7546 , n7474 , n7545 );
and ( n7547 , n7471 , n7546 );
or ( n7548 , n7470 , n7547 );
and ( n7549 , n7467 , n7548 );
or ( n7550 , n7466 , n7549 );
and ( n7551 , n7463 , n7550 );
or ( n7552 , n7462 , n7551 );
and ( n7553 , n7459 , n7552 );
or ( n7554 , n7458 , n7553 );
and ( n7555 , n7455 , n7554 );
or ( n7556 , n7454 , n7555 );
and ( n7557 , n7451 , n7556 );
or ( n7558 , n7450 , n7557 );
and ( n7559 , n7447 , n7558 );
or ( n7560 , n7446 , n7559 );
and ( n7561 , n7443 , n7560 );
or ( n7562 , n7442 , n7561 );
and ( n7563 , n7439 , n7562 );
or ( n7564 , n7438 , n7563 );
and ( n7565 , n7435 , n7564 );
or ( n7566 , n7434 , n7565 );
and ( n7567 , n7431 , n7566 );
or ( n7568 , n7430 , n7567 );
buf ( n7569 , n7568 );
and ( n7570 , n6841 , n371 );
and ( n7571 , n7569 , n7570 );
xor ( n7572 , n7569 , n7570 );
xor ( n7573 , n7431 , n7566 );
and ( n7574 , n6845 , n371 );
and ( n7575 , n7573 , n7574 );
xor ( n7576 , n7573 , n7574 );
xor ( n7577 , n7435 , n7564 );
and ( n7578 , n6850 , n371 );
and ( n7579 , n7577 , n7578 );
xor ( n7580 , n7577 , n7578 );
xor ( n7581 , n7439 , n7562 );
and ( n7582 , n6855 , n371 );
and ( n7583 , n7581 , n7582 );
xor ( n7584 , n7581 , n7582 );
xor ( n7585 , n7443 , n7560 );
and ( n7586 , n6860 , n371 );
and ( n7587 , n7585 , n7586 );
xor ( n7588 , n7585 , n7586 );
xor ( n7589 , n7447 , n7558 );
and ( n7590 , n6865 , n371 );
and ( n7591 , n7589 , n7590 );
xor ( n7592 , n7589 , n7590 );
xor ( n7593 , n7451 , n7556 );
and ( n7594 , n6870 , n371 );
and ( n7595 , n7593 , n7594 );
xor ( n7596 , n7593 , n7594 );
xor ( n7597 , n7455 , n7554 );
and ( n7598 , n6875 , n371 );
and ( n7599 , n7597 , n7598 );
xor ( n7600 , n7597 , n7598 );
xor ( n7601 , n7459 , n7552 );
and ( n7602 , n6880 , n371 );
and ( n7603 , n7601 , n7602 );
xor ( n7604 , n7601 , n7602 );
xor ( n7605 , n7463 , n7550 );
and ( n7606 , n6885 , n371 );
and ( n7607 , n7605 , n7606 );
xor ( n7608 , n7605 , n7606 );
xor ( n7609 , n7467 , n7548 );
and ( n7610 , n6890 , n371 );
and ( n7611 , n7609 , n7610 );
xor ( n7612 , n7609 , n7610 );
xor ( n7613 , n7471 , n7546 );
and ( n7614 , n6895 , n371 );
and ( n7615 , n7613 , n7614 );
xor ( n7616 , n7613 , n7614 );
xor ( n7617 , n7475 , n7544 );
and ( n7618 , n6900 , n371 );
and ( n7619 , n7617 , n7618 );
xor ( n7620 , n7617 , n7618 );
xor ( n7621 , n7479 , n7542 );
and ( n7622 , n6905 , n371 );
and ( n7623 , n7621 , n7622 );
xor ( n7624 , n7621 , n7622 );
xor ( n7625 , n7483 , n7540 );
and ( n7626 , n6910 , n371 );
and ( n7627 , n7625 , n7626 );
xor ( n7628 , n7625 , n7626 );
xor ( n7629 , n7487 , n7538 );
and ( n7630 , n6915 , n371 );
and ( n7631 , n7629 , n7630 );
xor ( n7632 , n7629 , n7630 );
xor ( n7633 , n7491 , n7536 );
and ( n7634 , n6920 , n371 );
and ( n7635 , n7633 , n7634 );
xor ( n7636 , n7633 , n7634 );
xor ( n7637 , n7495 , n7534 );
and ( n7638 , n6925 , n371 );
and ( n7639 , n7637 , n7638 );
xor ( n7640 , n7637 , n7638 );
xor ( n7641 , n7499 , n7532 );
and ( n7642 , n6930 , n371 );
and ( n7643 , n7641 , n7642 );
xor ( n7644 , n7641 , n7642 );
xor ( n7645 , n7503 , n7530 );
and ( n7646 , n6935 , n371 );
and ( n7647 , n7645 , n7646 );
xor ( n7648 , n7645 , n7646 );
xor ( n7649 , n7507 , n7528 );
and ( n7650 , n6940 , n371 );
and ( n7651 , n7649 , n7650 );
xor ( n7652 , n7649 , n7650 );
xor ( n7653 , n7511 , n7526 );
and ( n7654 , n6945 , n371 );
and ( n7655 , n7653 , n7654 );
xor ( n7656 , n7653 , n7654 );
xor ( n7657 , n7515 , n7524 );
and ( n7658 , n6951 , n371 );
and ( n7659 , n7657 , n7658 );
xor ( n7660 , n7657 , n7658 );
xor ( n7661 , n7519 , n7522 );
and ( n7662 , n6956 , n371 );
and ( n7663 , n7661 , n7662 );
and ( n7664 , n7660 , n7663 );
or ( n7665 , n7659 , n7664 );
and ( n7666 , n7656 , n7665 );
or ( n7667 , n7655 , n7666 );
and ( n7668 , n7652 , n7667 );
or ( n7669 , n7651 , n7668 );
and ( n7670 , n7648 , n7669 );
or ( n7671 , n7647 , n7670 );
and ( n7672 , n7644 , n7671 );
or ( n7673 , n7643 , n7672 );
and ( n7674 , n7640 , n7673 );
or ( n7675 , n7639 , n7674 );
and ( n7676 , n7636 , n7675 );
or ( n7677 , n7635 , n7676 );
and ( n7678 , n7632 , n7677 );
or ( n7679 , n7631 , n7678 );
and ( n7680 , n7628 , n7679 );
or ( n7681 , n7627 , n7680 );
and ( n7682 , n7624 , n7681 );
or ( n7683 , n7623 , n7682 );
and ( n7684 , n7620 , n7683 );
or ( n7685 , n7619 , n7684 );
and ( n7686 , n7616 , n7685 );
or ( n7687 , n7615 , n7686 );
and ( n7688 , n7612 , n7687 );
or ( n7689 , n7611 , n7688 );
and ( n7690 , n7608 , n7689 );
or ( n7691 , n7607 , n7690 );
and ( n7692 , n7604 , n7691 );
or ( n7693 , n7603 , n7692 );
and ( n7694 , n7600 , n7693 );
or ( n7695 , n7599 , n7694 );
and ( n7696 , n7596 , n7695 );
or ( n7697 , n7595 , n7696 );
and ( n7698 , n7592 , n7697 );
or ( n7699 , n7591 , n7698 );
and ( n7700 , n7588 , n7699 );
or ( n7701 , n7587 , n7700 );
and ( n7702 , n7584 , n7701 );
or ( n7703 , n7583 , n7702 );
and ( n7704 , n7580 , n7703 );
or ( n7705 , n7579 , n7704 );
and ( n7706 , n7576 , n7705 );
or ( n7707 , n7575 , n7706 );
and ( n7708 , n7572 , n7707 );
or ( n7709 , n7571 , n7708 );
buf ( n7710 , n7709 );
and ( n7711 , n6841 , n370 );
and ( n7712 , n7710 , n7711 );
xor ( n7713 , n7710 , n7711 );
xor ( n7714 , n7572 , n7707 );
and ( n7715 , n6845 , n370 );
and ( n7716 , n7714 , n7715 );
xor ( n7717 , n7714 , n7715 );
xor ( n7718 , n7576 , n7705 );
and ( n7719 , n6850 , n370 );
and ( n7720 , n7718 , n7719 );
xor ( n7721 , n7718 , n7719 );
xor ( n7722 , n7580 , n7703 );
and ( n7723 , n6855 , n370 );
and ( n7724 , n7722 , n7723 );
xor ( n7725 , n7722 , n7723 );
xor ( n7726 , n7584 , n7701 );
and ( n7727 , n6860 , n370 );
and ( n7728 , n7726 , n7727 );
xor ( n7729 , n7726 , n7727 );
xor ( n7730 , n7588 , n7699 );
and ( n7731 , n6865 , n370 );
and ( n7732 , n7730 , n7731 );
xor ( n7733 , n7730 , n7731 );
xor ( n7734 , n7592 , n7697 );
and ( n7735 , n6870 , n370 );
and ( n7736 , n7734 , n7735 );
xor ( n7737 , n7734 , n7735 );
xor ( n7738 , n7596 , n7695 );
and ( n7739 , n6875 , n370 );
and ( n7740 , n7738 , n7739 );
xor ( n7741 , n7738 , n7739 );
xor ( n7742 , n7600 , n7693 );
and ( n7743 , n6880 , n370 );
and ( n7744 , n7742 , n7743 );
xor ( n7745 , n7742 , n7743 );
xor ( n7746 , n7604 , n7691 );
and ( n7747 , n6885 , n370 );
and ( n7748 , n7746 , n7747 );
xor ( n7749 , n7746 , n7747 );
xor ( n7750 , n7608 , n7689 );
and ( n7751 , n6890 , n370 );
and ( n7752 , n7750 , n7751 );
xor ( n7753 , n7750 , n7751 );
xor ( n7754 , n7612 , n7687 );
and ( n7755 , n6895 , n370 );
and ( n7756 , n7754 , n7755 );
xor ( n7757 , n7754 , n7755 );
xor ( n7758 , n7616 , n7685 );
and ( n7759 , n6900 , n370 );
and ( n7760 , n7758 , n7759 );
xor ( n7761 , n7758 , n7759 );
xor ( n7762 , n7620 , n7683 );
and ( n7763 , n6905 , n370 );
and ( n7764 , n7762 , n7763 );
xor ( n7765 , n7762 , n7763 );
xor ( n7766 , n7624 , n7681 );
and ( n7767 , n6910 , n370 );
and ( n7768 , n7766 , n7767 );
xor ( n7769 , n7766 , n7767 );
xor ( n7770 , n7628 , n7679 );
and ( n7771 , n6915 , n370 );
and ( n7772 , n7770 , n7771 );
xor ( n7773 , n7770 , n7771 );
xor ( n7774 , n7632 , n7677 );
and ( n7775 , n6920 , n370 );
and ( n7776 , n7774 , n7775 );
xor ( n7777 , n7774 , n7775 );
xor ( n7778 , n7636 , n7675 );
and ( n7779 , n6925 , n370 );
and ( n7780 , n7778 , n7779 );
xor ( n7781 , n7778 , n7779 );
xor ( n7782 , n7640 , n7673 );
and ( n7783 , n6930 , n370 );
and ( n7784 , n7782 , n7783 );
xor ( n7785 , n7782 , n7783 );
xor ( n7786 , n7644 , n7671 );
and ( n7787 , n6935 , n370 );
and ( n7788 , n7786 , n7787 );
xor ( n7789 , n7786 , n7787 );
xor ( n7790 , n7648 , n7669 );
and ( n7791 , n6940 , n370 );
and ( n7792 , n7790 , n7791 );
xor ( n7793 , n7790 , n7791 );
xor ( n7794 , n7652 , n7667 );
and ( n7795 , n6945 , n370 );
and ( n7796 , n7794 , n7795 );
xor ( n7797 , n7794 , n7795 );
xor ( n7798 , n7656 , n7665 );
and ( n7799 , n6951 , n370 );
and ( n7800 , n7798 , n7799 );
xor ( n7801 , n7798 , n7799 );
xor ( n7802 , n7660 , n7663 );
and ( n7803 , n6956 , n370 );
and ( n7804 , n7802 , n7803 );
and ( n7805 , n7801 , n7804 );
or ( n7806 , n7800 , n7805 );
and ( n7807 , n7797 , n7806 );
or ( n7808 , n7796 , n7807 );
and ( n7809 , n7793 , n7808 );
or ( n7810 , n7792 , n7809 );
and ( n7811 , n7789 , n7810 );
or ( n7812 , n7788 , n7811 );
and ( n7813 , n7785 , n7812 );
or ( n7814 , n7784 , n7813 );
and ( n7815 , n7781 , n7814 );
or ( n7816 , n7780 , n7815 );
and ( n7817 , n7777 , n7816 );
or ( n7818 , n7776 , n7817 );
and ( n7819 , n7773 , n7818 );
or ( n7820 , n7772 , n7819 );
and ( n7821 , n7769 , n7820 );
or ( n7822 , n7768 , n7821 );
and ( n7823 , n7765 , n7822 );
or ( n7824 , n7764 , n7823 );
and ( n7825 , n7761 , n7824 );
or ( n7826 , n7760 , n7825 );
and ( n7827 , n7757 , n7826 );
or ( n7828 , n7756 , n7827 );
and ( n7829 , n7753 , n7828 );
or ( n7830 , n7752 , n7829 );
and ( n7831 , n7749 , n7830 );
or ( n7832 , n7748 , n7831 );
and ( n7833 , n7745 , n7832 );
or ( n7834 , n7744 , n7833 );
and ( n7835 , n7741 , n7834 );
or ( n7836 , n7740 , n7835 );
and ( n7837 , n7737 , n7836 );
or ( n7838 , n7736 , n7837 );
and ( n7839 , n7733 , n7838 );
or ( n7840 , n7732 , n7839 );
and ( n7841 , n7729 , n7840 );
or ( n7842 , n7728 , n7841 );
and ( n7843 , n7725 , n7842 );
or ( n7844 , n7724 , n7843 );
and ( n7845 , n7721 , n7844 );
or ( n7846 , n7720 , n7845 );
and ( n7847 , n7717 , n7846 );
or ( n7848 , n7716 , n7847 );
and ( n7849 , n7713 , n7848 );
or ( n7850 , n7712 , n7849 );
buf ( n7851 , n7850 );
buf ( n7852 , n7851 );
xor ( n7853 , n7713 , n7848 );
buf ( n7854 , n7853 );
xor ( n7855 , n7717 , n7846 );
buf ( n7856 , n7855 );
xor ( n7857 , n7721 , n7844 );
buf ( n7858 , n7857 );
xor ( n7859 , n7725 , n7842 );
buf ( n7860 , n7859 );
xor ( n7861 , n7729 , n7840 );
buf ( n7862 , n7861 );
xor ( n7863 , n7733 , n7838 );
buf ( n7864 , n7863 );
xor ( n7865 , n7737 , n7836 );
buf ( n7866 , n7865 );
xor ( n7867 , n7741 , n7834 );
buf ( n7868 , n7867 );
xor ( n7869 , n7745 , n7832 );
buf ( n7870 , n7869 );
xor ( n7871 , n7749 , n7830 );
buf ( n7872 , n7871 );
xor ( n7873 , n7753 , n7828 );
buf ( n7874 , n7873 );
xor ( n7875 , n7757 , n7826 );
buf ( n7876 , n7875 );
xor ( n7877 , n7761 , n7824 );
buf ( n7878 , n7877 );
xor ( n7879 , n7765 , n7822 );
buf ( n7880 , n7879 );
xor ( n7881 , n7769 , n7820 );
buf ( n7882 , n7881 );
xor ( n7883 , n7773 , n7818 );
buf ( n7884 , n7883 );
xor ( n7885 , n7777 , n7816 );
buf ( n7886 , n7885 );
xor ( n7887 , n7781 , n7814 );
buf ( n7888 , n7887 );
xor ( n7889 , n7785 , n7812 );
buf ( n7890 , n7889 );
xor ( n7891 , n7789 , n7810 );
buf ( n7892 , n7891 );
xor ( n7893 , n7793 , n7808 );
buf ( n7894 , n7893 );
xor ( n7895 , n7797 , n7806 );
buf ( n7896 , n7895 );
xor ( n7897 , n7801 , n7804 );
buf ( n7898 , n7897 );
xor ( n7899 , n7802 , n7803 );
buf ( n7900 , n7899 );
xor ( n7901 , n7661 , n7662 );
buf ( n7902 , n7901 );
xor ( n7903 , n7520 , n7521 );
buf ( n7904 , n7903 );
xor ( n7905 , n7379 , n7380 );
buf ( n7906 , n7905 );
xor ( n7907 , n7238 , n7239 );
buf ( n7908 , n7907 );
xor ( n7909 , n7097 , n7098 );
buf ( n7910 , n7909 );
buf ( n7911 , n6956 );
buf ( n7912 , n7911 );
buf ( n7913 , n402 );
buf ( n7914 , n403 );
buf ( n7915 , n404 );
buf ( n7916 , n405 );
buf ( n7917 , n406 );
buf ( n7918 , n407 );
buf ( n7919 , n408 );
buf ( n7920 , n409 );
and ( n7921 , n7900 , n7913 );
and ( n7922 , n7902 , n7914 );
and ( n7923 , n7904 , n7915 );
and ( n7924 , n7906 , n7916 );
and ( n7925 , n7908 , n7917 );
and ( n7926 , n7910 , n7918 );
and ( n7927 , n7912 , n7920 );
and ( n7928 , n7919 , n7927 );
buf ( n7929 , n7928 );
and ( n7930 , n7918 , n7929 );
and ( n7931 , n7910 , n7929 );
or ( n7932 , n7926 , n7930 , n7931 );
and ( n7933 , n7917 , n7932 );
and ( n7934 , n7908 , n7932 );
or ( n7935 , n7925 , n7933 , n7934 );
and ( n7936 , n7916 , n7935 );
and ( n7937 , n7906 , n7935 );
or ( n7938 , n7924 , n7936 , n7937 );
and ( n7939 , n7915 , n7938 );
and ( n7940 , n7904 , n7938 );
or ( n7941 , n7923 , n7939 , n7940 );
and ( n7942 , n7914 , n7941 );
and ( n7943 , n7902 , n7941 );
or ( n7944 , n7922 , n7942 , n7943 );
and ( n7945 , n7913 , n7944 );
and ( n7946 , n7900 , n7944 );
or ( n7947 , n7921 , n7945 , n7946 );
and ( n7948 , n7898 , n7947 );
and ( n7949 , n7896 , n7948 );
and ( n7950 , n7894 , n7949 );
and ( n7951 , n7892 , n7950 );
and ( n7952 , n7890 , n7951 );
and ( n7953 , n7888 , n7952 );
and ( n7954 , n7886 , n7953 );
and ( n7955 , n7884 , n7954 );
and ( n7956 , n7882 , n7955 );
and ( n7957 , n7880 , n7956 );
and ( n7958 , n7878 , n7957 );
and ( n7959 , n7876 , n7958 );
and ( n7960 , n7874 , n7959 );
and ( n7961 , n7872 , n7960 );
and ( n7962 , n7870 , n7961 );
and ( n7963 , n7868 , n7962 );
and ( n7964 , n7866 , n7963 );
and ( n7965 , n7864 , n7964 );
and ( n7966 , n7862 , n7965 );
and ( n7967 , n7860 , n7966 );
and ( n7968 , n7858 , n7967 );
and ( n7969 , n7856 , n7968 );
and ( n7970 , n7854 , n7969 );
xor ( n7971 , n7852 , n7970 );
buf ( n7972 , n7971 );
xor ( n7973 , n7854 , n7969 );
buf ( n7974 , n7973 );
xor ( n7975 , n7856 , n7968 );
buf ( n7976 , n7975 );
xor ( n7977 , n7858 , n7967 );
buf ( n7978 , n7977 );
xor ( n7979 , n7860 , n7966 );
buf ( n7980 , n7979 );
xor ( n7981 , n7862 , n7965 );
buf ( n7982 , n7981 );
xor ( n7983 , n7864 , n7964 );
buf ( n7984 , n7983 );
xor ( n7985 , n7866 , n7963 );
buf ( n7986 , n7985 );
xor ( n7987 , n7868 , n7962 );
buf ( n7988 , n7987 );
xor ( n7989 , n7870 , n7961 );
buf ( n7990 , n7989 );
buf ( n7991 , n4143 );
buf ( n7992 , n4145 );
buf ( n7993 , n4147 );
buf ( n7994 , n4149 );
buf ( n7995 , n4151 );
buf ( n7996 , n4153 );
buf ( n7997 , n4155 );
buf ( n7998 , n4157 );
buf ( n7999 , n4159 );
buf ( n8000 , n4161 );
buf ( n8001 , n4163 );
buf ( n8002 , n4165 );
buf ( n8003 , n4167 );
buf ( n8004 , n4169 );
buf ( n8005 , n4171 );
buf ( n8006 , n4173 );
buf ( n8007 , n4175 );
buf ( n8008 , n4177 );
buf ( n8009 , n4179 );
buf ( n8010 , n4181 );
buf ( n8011 , n4183 );
buf ( n8012 , n4185 );
buf ( n8013 , n4187 );
buf ( n8014 , n4189 );
buf ( n8015 , n4191 );
buf ( n8016 , n4193 );
buf ( n8017 , n4195 );
buf ( n8018 , n4197 );
buf ( n8019 , n4199 );
buf ( n8020 , n4201 );
buf ( n8021 , n4203 );
buf ( n8022 , n4205 );
buf ( n8023 , n4207 );
buf ( n8024 , n4209 );
buf ( n8025 , n4211 );
buf ( n8026 , n4213 );
buf ( n8027 , n4215 );
buf ( n8028 , n4217 );
buf ( n8029 , n4219 );
buf ( n8030 , n4221 );
buf ( n8031 , n4223 );
buf ( n8032 , n4225 );
buf ( n8033 , n4227 );
buf ( n8034 , n4229 );
buf ( n8035 , n4231 );
buf ( n8036 , n4233 );
buf ( n8037 , n4235 );
buf ( n8038 , n4237 );
buf ( n8039 , n4239 );
buf ( n8040 , n4241 );
buf ( n8041 , n4243 );
buf ( n8042 , n4245 );
buf ( n8043 , n4247 );
buf ( n8044 , n4249 );
buf ( n8045 , n4251 );
buf ( n8046 , n4253 );
buf ( n8047 , n4255 );
buf ( n8048 , n4257 );
buf ( n8049 , n4259 );
buf ( n8050 , n4261 );
buf ( n8051 , n4263 );
buf ( n8052 , n4266 );
buf ( n8053 , n4269 );
buf ( n8054 , n4271 );
buf ( n8055 , n7991 );
buf ( n8056 , n7992 );
buf ( n8057 , n378 );
buf ( n8058 , n8057 );
buf ( n8059 , n379 );
buf ( n8060 , n8059 );
buf ( n8061 , n380 );
buf ( n8062 , n8061 );
and ( n8063 , n8060 , n8062 );
not ( n8064 , n8063 );
and ( n8065 , n8058 , n8064 );
not ( n8066 , n8065 );
buf ( n8067 , n7993 );
and ( n8068 , n8066 , n8067 );
buf ( n8069 , n7994 );
and ( n8070 , n8065 , n8069 );
buf ( n8071 , n381 );
buf ( n8072 , n8071 );
buf ( n8073 , n382 );
buf ( n8074 , n8073 );
and ( n8075 , n8072 , n8074 );
not ( n8076 , n8075 );
and ( n8077 , n8062 , n8076 );
not ( n8078 , n8077 );
and ( n8079 , n8078 , n8065 );
buf ( n8080 , n7995 );
and ( n8081 , n8065 , n8080 );
and ( n8082 , n8078 , n8080 );
or ( n8083 , n8079 , n8081 , n8082 );
and ( n8084 , n8069 , n8083 );
and ( n8085 , n8065 , n8083 );
or ( n8086 , n8070 , n8084 , n8085 );
and ( n8087 , n8067 , n8086 );
and ( n8088 , n8066 , n8086 );
or ( n8089 , n8068 , n8087 , n8088 );
or ( n8090 , n8056 , n8089 );
or ( n8091 , n8055 , n8090 );
not ( n8092 , n8091 );
xnor ( n8093 , n8055 , n8090 );
xnor ( n8094 , n8056 , n8089 );
xor ( n8095 , n8066 , n8067 );
xor ( n8096 , n8095 , n8086 );
xor ( n8097 , n8065 , n8069 );
xor ( n8098 , n8097 , n8083 );
and ( n8099 , n8077 , n8065 );
buf ( n8100 , n7996 );
and ( n8101 , n8065 , n8100 );
and ( n8102 , n8077 , n8100 );
or ( n8103 , n8099 , n8101 , n8102 );
xor ( n8104 , n8078 , n8065 );
xor ( n8105 , n8104 , n8080 );
and ( n8106 , n8103 , n8105 );
buf ( n8107 , n383 );
buf ( n8108 , n8107 );
buf ( n8109 , n384 );
buf ( n8110 , n8109 );
and ( n8111 , n8108 , n8110 );
not ( n8112 , n8111 );
and ( n8113 , n8074 , n8112 );
not ( n8114 , n8113 );
and ( n8115 , n8114 , n8077 );
xor ( n8116 , n8077 , n8065 );
xor ( n8117 , n8116 , n8100 );
and ( n8118 , n8115 , n8117 );
xor ( n8119 , n8114 , n8077 );
and ( n8120 , n8065 , n8119 );
and ( n8121 , n8117 , n8120 );
and ( n8122 , n8115 , n8120 );
or ( n8123 , n8118 , n8121 , n8122 );
and ( n8124 , n8105 , n8123 );
and ( n8125 , n8103 , n8123 );
or ( n8126 , n8106 , n8124 , n8125 );
or ( n8127 , n8098 , n8126 );
and ( n8128 , n8096 , n8127 );
xor ( n8129 , n8096 , n8127 );
xnor ( n8130 , n8098 , n8126 );
xor ( n8131 , n8103 , n8105 );
xor ( n8132 , n8131 , n8123 );
buf ( n8133 , n7997 );
and ( n8134 , n8113 , n8077 );
and ( n8135 , n8077 , n8065 );
and ( n8136 , n8113 , n8065 );
or ( n8137 , n8134 , n8135 , n8136 );
and ( n8138 , n8133 , n8137 );
xor ( n8139 , n8065 , n8119 );
and ( n8140 , n8137 , n8139 );
and ( n8141 , n8133 , n8139 );
or ( n8142 , n8138 , n8140 , n8141 );
xor ( n8143 , n8115 , n8117 );
xor ( n8144 , n8143 , n8120 );
and ( n8145 , n8142 , n8144 );
buf ( n8146 , n7998 );
xor ( n8147 , n8113 , n8077 );
xor ( n8148 , n8147 , n8065 );
and ( n8149 , n8146 , n8148 );
and ( n8150 , n8113 , n8077 );
and ( n8151 , n8077 , n8065 );
and ( n8152 , n8113 , n8065 );
or ( n8153 , n8150 , n8151 , n8152 );
and ( n8154 , n8148 , n8153 );
and ( n8155 , n8146 , n8153 );
or ( n8156 , n8149 , n8154 , n8155 );
and ( n8157 , n8110 , n8113 );
and ( n8158 , n8113 , n8065 );
and ( n8159 , n8110 , n8065 );
or ( n8160 , n8157 , n8158 , n8159 );
buf ( n8161 , n8000 );
and ( n8162 , n8077 , n8161 );
or ( n8163 , n8160 , n8162 );
not ( n8164 , n8110 );
buf ( n8165 , n7999 );
and ( n8166 , n8164 , n8165 );
xor ( n8167 , n8113 , n8077 );
xor ( n8168 , n8167 , n8065 );
and ( n8169 , n8165 , n8168 );
and ( n8170 , n8164 , n8168 );
or ( n8171 , n8166 , n8169 , n8170 );
and ( n8172 , n8163 , n8171 );
xor ( n8173 , n8146 , n8148 );
xor ( n8174 , n8173 , n8153 );
and ( n8175 , n8171 , n8174 );
and ( n8176 , n8163 , n8174 );
or ( n8177 , n8172 , n8175 , n8176 );
and ( n8178 , n8156 , n8177 );
xor ( n8179 , n8133 , n8137 );
xor ( n8180 , n8179 , n8139 );
and ( n8181 , n8177 , n8180 );
and ( n8182 , n8156 , n8180 );
or ( n8183 , n8178 , n8181 , n8182 );
and ( n8184 , n8144 , n8183 );
and ( n8185 , n8142 , n8183 );
or ( n8186 , n8145 , n8184 , n8185 );
and ( n8187 , n8132 , n8186 );
xor ( n8188 , n8132 , n8186 );
xor ( n8189 , n8142 , n8144 );
xor ( n8190 , n8189 , n8183 );
not ( n8191 , n8190 );
xor ( n8192 , n8156 , n8177 );
xor ( n8193 , n8192 , n8180 );
xnor ( n8194 , n8160 , n8162 );
xor ( n8195 , n8077 , n8161 );
and ( n8196 , n8110 , n8113 );
and ( n8197 , n8113 , n8065 );
and ( n8198 , n8110 , n8065 );
or ( n8199 , n8196 , n8197 , n8198 );
and ( n8200 , n8195 , n8199 );
buf ( n8201 , n8001 );
and ( n8202 , n8077 , n8201 );
and ( n8203 , n8199 , n8202 );
and ( n8204 , n8195 , n8202 );
or ( n8205 , n8200 , n8203 , n8204 );
and ( n8206 , n8194 , n8205 );
xor ( n8207 , n8164 , n8165 );
xor ( n8208 , n8207 , n8168 );
and ( n8209 , n8205 , n8208 );
and ( n8210 , n8194 , n8208 );
or ( n8211 , n8206 , n8209 , n8210 );
xor ( n8212 , n8163 , n8171 );
xor ( n8213 , n8212 , n8174 );
and ( n8214 , n8211 , n8213 );
xor ( n8215 , n8077 , n8201 );
and ( n8216 , n8110 , n8113 );
and ( n8217 , n8113 , n8065 );
and ( n8218 , n8110 , n8065 );
or ( n8219 , n8216 , n8217 , n8218 );
and ( n8220 , n8215 , n8219 );
buf ( n8221 , n8002 );
and ( n8222 , n8077 , n8221 );
and ( n8223 , n8219 , n8222 );
and ( n8224 , n8215 , n8222 );
or ( n8225 , n8220 , n8223 , n8224 );
xor ( n8226 , n8110 , n8113 );
xor ( n8227 , n8226 , n8065 );
and ( n8228 , n8225 , n8227 );
xor ( n8229 , n8195 , n8199 );
xor ( n8230 , n8229 , n8202 );
and ( n8231 , n8227 , n8230 );
and ( n8232 , n8225 , n8230 );
or ( n8233 , n8228 , n8231 , n8232 );
xor ( n8234 , n8194 , n8205 );
xor ( n8235 , n8234 , n8208 );
and ( n8236 , n8233 , n8235 );
xor ( n8237 , n8225 , n8227 );
xor ( n8238 , n8237 , n8230 );
xor ( n8239 , n8077 , n8221 );
and ( n8240 , n8110 , n8113 );
and ( n8241 , n8113 , n8065 );
and ( n8242 , n8110 , n8065 );
or ( n8243 , n8240 , n8241 , n8242 );
and ( n8244 , n8239 , n8243 );
buf ( n8245 , n8003 );
and ( n8246 , n8077 , n8245 );
and ( n8247 , n8243 , n8246 );
and ( n8248 , n8239 , n8246 );
or ( n8249 , n8244 , n8247 , n8248 );
xor ( n8250 , n8110 , n8113 );
xor ( n8251 , n8250 , n8065 );
and ( n8252 , n8249 , n8251 );
xor ( n8253 , n8215 , n8219 );
xor ( n8254 , n8253 , n8222 );
and ( n8255 , n8251 , n8254 );
and ( n8256 , n8249 , n8254 );
or ( n8257 , n8252 , n8255 , n8256 );
and ( n8258 , n8238 , n8257 );
xor ( n8259 , n8249 , n8251 );
xor ( n8260 , n8259 , n8254 );
xor ( n8261 , n8077 , n8245 );
and ( n8262 , n8110 , n8113 );
and ( n8263 , n8113 , n8065 );
and ( n8264 , n8110 , n8065 );
or ( n8265 , n8262 , n8263 , n8264 );
and ( n8266 , n8261 , n8265 );
buf ( n8267 , n8004 );
and ( n8268 , n8077 , n8267 );
and ( n8269 , n8265 , n8268 );
and ( n8270 , n8261 , n8268 );
or ( n8271 , n8266 , n8269 , n8270 );
xor ( n8272 , n8110 , n8113 );
xor ( n8273 , n8272 , n8065 );
and ( n8274 , n8271 , n8273 );
xor ( n8275 , n8239 , n8243 );
xor ( n8276 , n8275 , n8246 );
and ( n8277 , n8273 , n8276 );
and ( n8278 , n8271 , n8276 );
or ( n8279 , n8274 , n8277 , n8278 );
and ( n8280 , n8260 , n8279 );
xor ( n8281 , n8271 , n8273 );
xor ( n8282 , n8281 , n8276 );
xor ( n8283 , n8077 , n8267 );
and ( n8284 , n8110 , n8113 );
and ( n8285 , n8113 , n8065 );
and ( n8286 , n8110 , n8065 );
or ( n8287 , n8284 , n8285 , n8286 );
and ( n8288 , n8283 , n8287 );
buf ( n8289 , n8005 );
and ( n8290 , n8077 , n8289 );
and ( n8291 , n8287 , n8290 );
and ( n8292 , n8283 , n8290 );
or ( n8293 , n8288 , n8291 , n8292 );
xor ( n8294 , n8110 , n8113 );
xor ( n8295 , n8294 , n8065 );
and ( n8296 , n8293 , n8295 );
xor ( n8297 , n8261 , n8265 );
xor ( n8298 , n8297 , n8268 );
and ( n8299 , n8295 , n8298 );
and ( n8300 , n8293 , n8298 );
or ( n8301 , n8296 , n8299 , n8300 );
and ( n8302 , n8282 , n8301 );
xor ( n8303 , n8293 , n8295 );
xor ( n8304 , n8303 , n8298 );
xor ( n8305 , n8077 , n8289 );
and ( n8306 , n8110 , n8113 );
and ( n8307 , n8113 , n8065 );
and ( n8308 , n8110 , n8065 );
or ( n8309 , n8306 , n8307 , n8308 );
and ( n8310 , n8305 , n8309 );
buf ( n8311 , n8006 );
and ( n8312 , n8077 , n8311 );
and ( n8313 , n8309 , n8312 );
and ( n8314 , n8305 , n8312 );
or ( n8315 , n8310 , n8313 , n8314 );
xor ( n8316 , n8110 , n8113 );
xor ( n8317 , n8316 , n8065 );
and ( n8318 , n8315 , n8317 );
xor ( n8319 , n8283 , n8287 );
xor ( n8320 , n8319 , n8290 );
and ( n8321 , n8317 , n8320 );
and ( n8322 , n8315 , n8320 );
or ( n8323 , n8318 , n8321 , n8322 );
and ( n8324 , n8304 , n8323 );
xor ( n8325 , n8315 , n8317 );
xor ( n8326 , n8325 , n8320 );
xor ( n8327 , n8077 , n8311 );
and ( n8328 , n8110 , n8113 );
and ( n8329 , n8113 , n8065 );
and ( n8330 , n8110 , n8065 );
or ( n8331 , n8328 , n8329 , n8330 );
and ( n8332 , n8327 , n8331 );
buf ( n8333 , n8007 );
and ( n8334 , n8077 , n8333 );
and ( n8335 , n8331 , n8334 );
and ( n8336 , n8327 , n8334 );
or ( n8337 , n8332 , n8335 , n8336 );
xor ( n8338 , n8110 , n8113 );
xor ( n8339 , n8338 , n8065 );
and ( n8340 , n8337 , n8339 );
xor ( n8341 , n8305 , n8309 );
xor ( n8342 , n8341 , n8312 );
and ( n8343 , n8339 , n8342 );
and ( n8344 , n8337 , n8342 );
or ( n8345 , n8340 , n8343 , n8344 );
and ( n8346 , n8326 , n8345 );
xor ( n8347 , n8337 , n8339 );
xor ( n8348 , n8347 , n8342 );
xor ( n8349 , n8077 , n8333 );
and ( n8350 , n8110 , n8113 );
and ( n8351 , n8113 , n8065 );
and ( n8352 , n8110 , n8065 );
or ( n8353 , n8350 , n8351 , n8352 );
and ( n8354 , n8349 , n8353 );
buf ( n8355 , n8008 );
and ( n8356 , n8077 , n8355 );
and ( n8357 , n8353 , n8356 );
and ( n8358 , n8349 , n8356 );
or ( n8359 , n8354 , n8357 , n8358 );
xor ( n8360 , n8110 , n8113 );
xor ( n8361 , n8360 , n8065 );
and ( n8362 , n8359 , n8361 );
xor ( n8363 , n8327 , n8331 );
xor ( n8364 , n8363 , n8334 );
and ( n8365 , n8361 , n8364 );
and ( n8366 , n8359 , n8364 );
or ( n8367 , n8362 , n8365 , n8366 );
and ( n8368 , n8348 , n8367 );
xor ( n8369 , n8359 , n8361 );
xor ( n8370 , n8369 , n8364 );
xor ( n8371 , n8077 , n8355 );
and ( n8372 , n8110 , n8113 );
and ( n8373 , n8113 , n8065 );
and ( n8374 , n8110 , n8065 );
or ( n8375 , n8372 , n8373 , n8374 );
and ( n8376 , n8371 , n8375 );
buf ( n8377 , n8009 );
and ( n8378 , n8077 , n8377 );
and ( n8379 , n8375 , n8378 );
and ( n8380 , n8371 , n8378 );
or ( n8381 , n8376 , n8379 , n8380 );
xor ( n8382 , n8110 , n8113 );
xor ( n8383 , n8382 , n8065 );
and ( n8384 , n8381 , n8383 );
xor ( n8385 , n8349 , n8353 );
xor ( n8386 , n8385 , n8356 );
and ( n8387 , n8383 , n8386 );
and ( n8388 , n8381 , n8386 );
or ( n8389 , n8384 , n8387 , n8388 );
and ( n8390 , n8370 , n8389 );
xor ( n8391 , n8381 , n8383 );
xor ( n8392 , n8391 , n8386 );
xor ( n8393 , n8077 , n8377 );
and ( n8394 , n8110 , n8113 );
and ( n8395 , n8113 , n8065 );
and ( n8396 , n8110 , n8065 );
or ( n8397 , n8394 , n8395 , n8396 );
and ( n8398 , n8393 , n8397 );
buf ( n8399 , n8010 );
and ( n8400 , n8077 , n8399 );
and ( n8401 , n8397 , n8400 );
and ( n8402 , n8393 , n8400 );
or ( n8403 , n8398 , n8401 , n8402 );
xor ( n8404 , n8110 , n8113 );
xor ( n8405 , n8404 , n8065 );
and ( n8406 , n8403 , n8405 );
xor ( n8407 , n8371 , n8375 );
xor ( n8408 , n8407 , n8378 );
and ( n8409 , n8405 , n8408 );
and ( n8410 , n8403 , n8408 );
or ( n8411 , n8406 , n8409 , n8410 );
and ( n8412 , n8392 , n8411 );
xor ( n8413 , n8403 , n8405 );
xor ( n8414 , n8413 , n8408 );
xor ( n8415 , n8077 , n8399 );
and ( n8416 , n8110 , n8113 );
and ( n8417 , n8113 , n8065 );
and ( n8418 , n8110 , n8065 );
or ( n8419 , n8416 , n8417 , n8418 );
and ( n8420 , n8415 , n8419 );
buf ( n8421 , n8011 );
and ( n8422 , n8077 , n8421 );
and ( n8423 , n8419 , n8422 );
and ( n8424 , n8415 , n8422 );
or ( n8425 , n8420 , n8423 , n8424 );
xor ( n8426 , n8110 , n8113 );
xor ( n8427 , n8426 , n8065 );
and ( n8428 , n8425 , n8427 );
xor ( n8429 , n8393 , n8397 );
xor ( n8430 , n8429 , n8400 );
and ( n8431 , n8427 , n8430 );
and ( n8432 , n8425 , n8430 );
or ( n8433 , n8428 , n8431 , n8432 );
and ( n8434 , n8414 , n8433 );
xor ( n8435 , n8077 , n8421 );
and ( n8436 , n8110 , n8113 );
and ( n8437 , n8113 , n8065 );
and ( n8438 , n8110 , n8065 );
or ( n8439 , n8436 , n8437 , n8438 );
and ( n8440 , n8435 , n8439 );
buf ( n8441 , n8012 );
and ( n8442 , n8077 , n8441 );
and ( n8443 , n8439 , n8442 );
and ( n8444 , n8435 , n8442 );
or ( n8445 , n8440 , n8443 , n8444 );
xor ( n8446 , n8110 , n8113 );
xor ( n8447 , n8446 , n8065 );
and ( n8448 , n8445 , n8447 );
xor ( n8449 , n8415 , n8419 );
xor ( n8450 , n8449 , n8422 );
and ( n8451 , n8447 , n8450 );
and ( n8452 , n8445 , n8450 );
or ( n8453 , n8448 , n8451 , n8452 );
xor ( n8454 , n8425 , n8427 );
xor ( n8455 , n8454 , n8430 );
and ( n8456 , n8453 , n8455 );
xor ( n8457 , n8077 , n8441 );
and ( n8458 , n8110 , n8113 );
and ( n8459 , n8113 , n8065 );
and ( n8460 , n8110 , n8065 );
or ( n8461 , n8458 , n8459 , n8460 );
and ( n8462 , n8457 , n8461 );
buf ( n8463 , n8013 );
and ( n8464 , n8077 , n8463 );
and ( n8465 , n8461 , n8464 );
and ( n8466 , n8457 , n8464 );
or ( n8467 , n8462 , n8465 , n8466 );
xor ( n8468 , n8110 , n8113 );
xor ( n8469 , n8468 , n8065 );
and ( n8470 , n8467 , n8469 );
xor ( n8471 , n8435 , n8439 );
xor ( n8472 , n8471 , n8442 );
and ( n8473 , n8469 , n8472 );
and ( n8474 , n8467 , n8472 );
or ( n8475 , n8470 , n8473 , n8474 );
xor ( n8476 , n8445 , n8447 );
xor ( n8477 , n8476 , n8450 );
and ( n8478 , n8475 , n8477 );
xor ( n8479 , n8077 , n8463 );
and ( n8480 , n8110 , n8113 );
and ( n8481 , n8113 , n8065 );
and ( n8482 , n8110 , n8065 );
or ( n8483 , n8480 , n8481 , n8482 );
and ( n8484 , n8479 , n8483 );
buf ( n8485 , n8014 );
and ( n8486 , n8077 , n8485 );
and ( n8487 , n8483 , n8486 );
and ( n8488 , n8479 , n8486 );
or ( n8489 , n8484 , n8487 , n8488 );
xor ( n8490 , n8110 , n8113 );
xor ( n8491 , n8490 , n8065 );
and ( n8492 , n8489 , n8491 );
xor ( n8493 , n8457 , n8461 );
xor ( n8494 , n8493 , n8464 );
and ( n8495 , n8491 , n8494 );
and ( n8496 , n8489 , n8494 );
or ( n8497 , n8492 , n8495 , n8496 );
xor ( n8498 , n8467 , n8469 );
xor ( n8499 , n8498 , n8472 );
and ( n8500 , n8497 , n8499 );
xor ( n8501 , n8077 , n8485 );
and ( n8502 , n8110 , n8113 );
and ( n8503 , n8113 , n8065 );
and ( n8504 , n8110 , n8065 );
or ( n8505 , n8502 , n8503 , n8504 );
and ( n8506 , n8501 , n8505 );
buf ( n8507 , n8015 );
and ( n8508 , n8077 , n8507 );
and ( n8509 , n8505 , n8508 );
and ( n8510 , n8501 , n8508 );
or ( n8511 , n8506 , n8509 , n8510 );
xor ( n8512 , n8110 , n8113 );
xor ( n8513 , n8512 , n8065 );
and ( n8514 , n8511 , n8513 );
xor ( n8515 , n8479 , n8483 );
xor ( n8516 , n8515 , n8486 );
and ( n8517 , n8513 , n8516 );
and ( n8518 , n8511 , n8516 );
or ( n8519 , n8514 , n8517 , n8518 );
xor ( n8520 , n8489 , n8491 );
xor ( n8521 , n8520 , n8494 );
and ( n8522 , n8519 , n8521 );
xor ( n8523 , n8077 , n8507 );
and ( n8524 , n8110 , n8113 );
and ( n8525 , n8113 , n8065 );
and ( n8526 , n8110 , n8065 );
or ( n8527 , n8524 , n8525 , n8526 );
and ( n8528 , n8523 , n8527 );
buf ( n8529 , n8016 );
and ( n8530 , n8077 , n8529 );
and ( n8531 , n8527 , n8530 );
and ( n8532 , n8523 , n8530 );
or ( n8533 , n8528 , n8531 , n8532 );
xor ( n8534 , n8110 , n8113 );
xor ( n8535 , n8534 , n8065 );
and ( n8536 , n8533 , n8535 );
xor ( n8537 , n8501 , n8505 );
xor ( n8538 , n8537 , n8508 );
and ( n8539 , n8535 , n8538 );
and ( n8540 , n8533 , n8538 );
or ( n8541 , n8536 , n8539 , n8540 );
xor ( n8542 , n8511 , n8513 );
xor ( n8543 , n8542 , n8516 );
and ( n8544 , n8541 , n8543 );
xor ( n8545 , n8077 , n8529 );
and ( n8546 , n8110 , n8113 );
and ( n8547 , n8113 , n8065 );
and ( n8548 , n8110 , n8065 );
or ( n8549 , n8546 , n8547 , n8548 );
and ( n8550 , n8545 , n8549 );
buf ( n8551 , n8017 );
and ( n8552 , n8077 , n8551 );
and ( n8553 , n8549 , n8552 );
and ( n8554 , n8545 , n8552 );
or ( n8555 , n8550 , n8553 , n8554 );
xor ( n8556 , n8110 , n8113 );
xor ( n8557 , n8556 , n8065 );
and ( n8558 , n8555 , n8557 );
xor ( n8559 , n8523 , n8527 );
xor ( n8560 , n8559 , n8530 );
and ( n8561 , n8557 , n8560 );
and ( n8562 , n8555 , n8560 );
or ( n8563 , n8558 , n8561 , n8562 );
xor ( n8564 , n8533 , n8535 );
xor ( n8565 , n8564 , n8538 );
and ( n8566 , n8563 , n8565 );
xor ( n8567 , n8077 , n8551 );
and ( n8568 , n8110 , n8113 );
and ( n8569 , n8113 , n8065 );
and ( n8570 , n8110 , n8065 );
or ( n8571 , n8568 , n8569 , n8570 );
and ( n8572 , n8567 , n8571 );
buf ( n8573 , n8018 );
and ( n8574 , n8077 , n8573 );
and ( n8575 , n8571 , n8574 );
and ( n8576 , n8567 , n8574 );
or ( n8577 , n8572 , n8575 , n8576 );
xor ( n8578 , n8110 , n8113 );
xor ( n8579 , n8578 , n8065 );
and ( n8580 , n8577 , n8579 );
xor ( n8581 , n8545 , n8549 );
xor ( n8582 , n8581 , n8552 );
and ( n8583 , n8579 , n8582 );
and ( n8584 , n8577 , n8582 );
or ( n8585 , n8580 , n8583 , n8584 );
xor ( n8586 , n8555 , n8557 );
xor ( n8587 , n8586 , n8560 );
and ( n8588 , n8585 , n8587 );
xor ( n8589 , n8077 , n8573 );
and ( n8590 , n8110 , n8113 );
and ( n8591 , n8113 , n8065 );
and ( n8592 , n8110 , n8065 );
or ( n8593 , n8590 , n8591 , n8592 );
and ( n8594 , n8589 , n8593 );
buf ( n8595 , n8019 );
and ( n8596 , n8077 , n8595 );
and ( n8597 , n8593 , n8596 );
and ( n8598 , n8589 , n8596 );
or ( n8599 , n8594 , n8597 , n8598 );
xor ( n8600 , n8110 , n8113 );
xor ( n8601 , n8600 , n8065 );
and ( n8602 , n8599 , n8601 );
xor ( n8603 , n8567 , n8571 );
xor ( n8604 , n8603 , n8574 );
and ( n8605 , n8601 , n8604 );
and ( n8606 , n8599 , n8604 );
or ( n8607 , n8602 , n8605 , n8606 );
xor ( n8608 , n8577 , n8579 );
xor ( n8609 , n8608 , n8582 );
and ( n8610 , n8607 , n8609 );
xor ( n8611 , n8077 , n8595 );
and ( n8612 , n8110 , n8113 );
and ( n8613 , n8113 , n8065 );
and ( n8614 , n8110 , n8065 );
or ( n8615 , n8612 , n8613 , n8614 );
and ( n8616 , n8611 , n8615 );
buf ( n8617 , n8020 );
and ( n8618 , n8077 , n8617 );
and ( n8619 , n8615 , n8618 );
and ( n8620 , n8611 , n8618 );
or ( n8621 , n8616 , n8619 , n8620 );
xor ( n8622 , n8110 , n8113 );
xor ( n8623 , n8622 , n8065 );
and ( n8624 , n8621 , n8623 );
xor ( n8625 , n8589 , n8593 );
xor ( n8626 , n8625 , n8596 );
and ( n8627 , n8623 , n8626 );
and ( n8628 , n8621 , n8626 );
or ( n8629 , n8624 , n8627 , n8628 );
xor ( n8630 , n8599 , n8601 );
xor ( n8631 , n8630 , n8604 );
and ( n8632 , n8629 , n8631 );
xor ( n8633 , n8077 , n8617 );
and ( n8634 , n8110 , n8113 );
and ( n8635 , n8113 , n8065 );
and ( n8636 , n8110 , n8065 );
or ( n8637 , n8634 , n8635 , n8636 );
and ( n8638 , n8633 , n8637 );
buf ( n8639 , n8021 );
and ( n8640 , n8077 , n8639 );
and ( n8641 , n8637 , n8640 );
and ( n8642 , n8633 , n8640 );
or ( n8643 , n8638 , n8641 , n8642 );
xor ( n8644 , n8110 , n8113 );
xor ( n8645 , n8644 , n8065 );
and ( n8646 , n8643 , n8645 );
xor ( n8647 , n8611 , n8615 );
xor ( n8648 , n8647 , n8618 );
and ( n8649 , n8645 , n8648 );
and ( n8650 , n8643 , n8648 );
or ( n8651 , n8646 , n8649 , n8650 );
xor ( n8652 , n8621 , n8623 );
xor ( n8653 , n8652 , n8626 );
and ( n8654 , n8651 , n8653 );
xor ( n8655 , n8077 , n8639 );
and ( n8656 , n8110 , n8113 );
and ( n8657 , n8113 , n8065 );
and ( n8658 , n8110 , n8065 );
or ( n8659 , n8656 , n8657 , n8658 );
and ( n8660 , n8655 , n8659 );
buf ( n8661 , n8022 );
and ( n8662 , n8077 , n8661 );
and ( n8663 , n8659 , n8662 );
and ( n8664 , n8655 , n8662 );
or ( n8665 , n8660 , n8663 , n8664 );
xor ( n8666 , n8110 , n8113 );
xor ( n8667 , n8666 , n8065 );
and ( n8668 , n8665 , n8667 );
xor ( n8669 , n8633 , n8637 );
xor ( n8670 , n8669 , n8640 );
and ( n8671 , n8667 , n8670 );
and ( n8672 , n8665 , n8670 );
or ( n8673 , n8668 , n8671 , n8672 );
xor ( n8674 , n8643 , n8645 );
xor ( n8675 , n8674 , n8648 );
and ( n8676 , n8673 , n8675 );
xor ( n8677 , n8077 , n8661 );
and ( n8678 , n8110 , n8113 );
and ( n8679 , n8113 , n8065 );
and ( n8680 , n8110 , n8065 );
or ( n8681 , n8678 , n8679 , n8680 );
and ( n8682 , n8677 , n8681 );
buf ( n8683 , n8023 );
and ( n8684 , n8077 , n8683 );
and ( n8685 , n8681 , n8684 );
and ( n8686 , n8677 , n8684 );
or ( n8687 , n8682 , n8685 , n8686 );
xor ( n8688 , n8110 , n8113 );
xor ( n8689 , n8688 , n8065 );
and ( n8690 , n8687 , n8689 );
xor ( n8691 , n8655 , n8659 );
xor ( n8692 , n8691 , n8662 );
and ( n8693 , n8689 , n8692 );
and ( n8694 , n8687 , n8692 );
or ( n8695 , n8690 , n8693 , n8694 );
xor ( n8696 , n8665 , n8667 );
xor ( n8697 , n8696 , n8670 );
and ( n8698 , n8695 , n8697 );
xor ( n8699 , n8077 , n8683 );
and ( n8700 , n8110 , n8113 );
and ( n8701 , n8113 , n8065 );
and ( n8702 , n8110 , n8065 );
or ( n8703 , n8700 , n8701 , n8702 );
and ( n8704 , n8699 , n8703 );
buf ( n8705 , n8024 );
and ( n8706 , n8077 , n8705 );
and ( n8707 , n8703 , n8706 );
and ( n8708 , n8699 , n8706 );
or ( n8709 , n8704 , n8707 , n8708 );
xor ( n8710 , n8110 , n8113 );
xor ( n8711 , n8710 , n8065 );
and ( n8712 , n8709 , n8711 );
xor ( n8713 , n8677 , n8681 );
xor ( n8714 , n8713 , n8684 );
and ( n8715 , n8711 , n8714 );
and ( n8716 , n8709 , n8714 );
or ( n8717 , n8712 , n8715 , n8716 );
xor ( n8718 , n8687 , n8689 );
xor ( n8719 , n8718 , n8692 );
and ( n8720 , n8717 , n8719 );
xor ( n8721 , n8077 , n8705 );
and ( n8722 , n8110 , n8113 );
and ( n8723 , n8113 , n8065 );
and ( n8724 , n8110 , n8065 );
or ( n8725 , n8722 , n8723 , n8724 );
and ( n8726 , n8721 , n8725 );
buf ( n8727 , n8025 );
and ( n8728 , n8077 , n8727 );
and ( n8729 , n8725 , n8728 );
and ( n8730 , n8721 , n8728 );
or ( n8731 , n8726 , n8729 , n8730 );
xor ( n8732 , n8110 , n8113 );
xor ( n8733 , n8732 , n8065 );
and ( n8734 , n8731 , n8733 );
xor ( n8735 , n8699 , n8703 );
xor ( n8736 , n8735 , n8706 );
and ( n8737 , n8733 , n8736 );
and ( n8738 , n8731 , n8736 );
or ( n8739 , n8734 , n8737 , n8738 );
xor ( n8740 , n8709 , n8711 );
xor ( n8741 , n8740 , n8714 );
and ( n8742 , n8739 , n8741 );
xor ( n8743 , n8077 , n8727 );
and ( n8744 , n8110 , n8113 );
and ( n8745 , n8113 , n8065 );
and ( n8746 , n8110 , n8065 );
or ( n8747 , n8744 , n8745 , n8746 );
and ( n8748 , n8743 , n8747 );
buf ( n8749 , n8026 );
and ( n8750 , n8077 , n8749 );
and ( n8751 , n8747 , n8750 );
and ( n8752 , n8743 , n8750 );
or ( n8753 , n8748 , n8751 , n8752 );
xor ( n8754 , n8110 , n8113 );
xor ( n8755 , n8754 , n8065 );
and ( n8756 , n8753 , n8755 );
xor ( n8757 , n8721 , n8725 );
xor ( n8758 , n8757 , n8728 );
and ( n8759 , n8755 , n8758 );
and ( n8760 , n8753 , n8758 );
or ( n8761 , n8756 , n8759 , n8760 );
xor ( n8762 , n8731 , n8733 );
xor ( n8763 , n8762 , n8736 );
and ( n8764 , n8761 , n8763 );
xor ( n8765 , n8077 , n8749 );
and ( n8766 , n8110 , n8113 );
and ( n8767 , n8113 , n8065 );
and ( n8768 , n8110 , n8065 );
or ( n8769 , n8766 , n8767 , n8768 );
and ( n8770 , n8765 , n8769 );
buf ( n8771 , n8027 );
and ( n8772 , n8077 , n8771 );
and ( n8773 , n8769 , n8772 );
and ( n8774 , n8765 , n8772 );
or ( n8775 , n8770 , n8773 , n8774 );
xor ( n8776 , n8110 , n8113 );
xor ( n8777 , n8776 , n8065 );
and ( n8778 , n8775 , n8777 );
xor ( n8779 , n8743 , n8747 );
xor ( n8780 , n8779 , n8750 );
and ( n8781 , n8777 , n8780 );
and ( n8782 , n8775 , n8780 );
or ( n8783 , n8778 , n8781 , n8782 );
xor ( n8784 , n8753 , n8755 );
xor ( n8785 , n8784 , n8758 );
and ( n8786 , n8783 , n8785 );
xor ( n8787 , n8077 , n8771 );
and ( n8788 , n8110 , n8113 );
and ( n8789 , n8113 , n8065 );
and ( n8790 , n8110 , n8065 );
or ( n8791 , n8788 , n8789 , n8790 );
and ( n8792 , n8787 , n8791 );
buf ( n8793 , n8028 );
and ( n8794 , n8077 , n8793 );
and ( n8795 , n8791 , n8794 );
and ( n8796 , n8787 , n8794 );
or ( n8797 , n8792 , n8795 , n8796 );
xor ( n8798 , n8110 , n8113 );
xor ( n8799 , n8798 , n8065 );
and ( n8800 , n8797 , n8799 );
xor ( n8801 , n8765 , n8769 );
xor ( n8802 , n8801 , n8772 );
and ( n8803 , n8799 , n8802 );
and ( n8804 , n8797 , n8802 );
or ( n8805 , n8800 , n8803 , n8804 );
xor ( n8806 , n8775 , n8777 );
xor ( n8807 , n8806 , n8780 );
and ( n8808 , n8805 , n8807 );
xor ( n8809 , n8077 , n8793 );
and ( n8810 , n8110 , n8113 );
and ( n8811 , n8113 , n8065 );
and ( n8812 , n8110 , n8065 );
or ( n8813 , n8810 , n8811 , n8812 );
and ( n8814 , n8809 , n8813 );
buf ( n8815 , n8029 );
and ( n8816 , n8077 , n8815 );
and ( n8817 , n8813 , n8816 );
and ( n8818 , n8809 , n8816 );
or ( n8819 , n8814 , n8817 , n8818 );
xor ( n8820 , n8110 , n8113 );
xor ( n8821 , n8820 , n8065 );
and ( n8822 , n8819 , n8821 );
xor ( n8823 , n8787 , n8791 );
xor ( n8824 , n8823 , n8794 );
and ( n8825 , n8821 , n8824 );
and ( n8826 , n8819 , n8824 );
or ( n8827 , n8822 , n8825 , n8826 );
xor ( n8828 , n8797 , n8799 );
xor ( n8829 , n8828 , n8802 );
and ( n8830 , n8827 , n8829 );
xor ( n8831 , n8077 , n8815 );
and ( n8832 , n8110 , n8113 );
and ( n8833 , n8113 , n8065 );
and ( n8834 , n8110 , n8065 );
or ( n8835 , n8832 , n8833 , n8834 );
and ( n8836 , n8831 , n8835 );
buf ( n8837 , n8030 );
and ( n8838 , n8077 , n8837 );
and ( n8839 , n8835 , n8838 );
and ( n8840 , n8831 , n8838 );
or ( n8841 , n8836 , n8839 , n8840 );
xor ( n8842 , n8110 , n8113 );
xor ( n8843 , n8842 , n8065 );
and ( n8844 , n8841 , n8843 );
xor ( n8845 , n8809 , n8813 );
xor ( n8846 , n8845 , n8816 );
and ( n8847 , n8843 , n8846 );
and ( n8848 , n8841 , n8846 );
or ( n8849 , n8844 , n8847 , n8848 );
xor ( n8850 , n8819 , n8821 );
xor ( n8851 , n8850 , n8824 );
and ( n8852 , n8849 , n8851 );
xor ( n8853 , n8077 , n8837 );
and ( n8854 , n8110 , n8113 );
and ( n8855 , n8113 , n8065 );
and ( n8856 , n8110 , n8065 );
or ( n8857 , n8854 , n8855 , n8856 );
and ( n8858 , n8853 , n8857 );
buf ( n8859 , n8031 );
and ( n8860 , n8077 , n8859 );
and ( n8861 , n8857 , n8860 );
and ( n8862 , n8853 , n8860 );
or ( n8863 , n8858 , n8861 , n8862 );
xor ( n8864 , n8110 , n8113 );
xor ( n8865 , n8864 , n8065 );
and ( n8866 , n8863 , n8865 );
xor ( n8867 , n8831 , n8835 );
xor ( n8868 , n8867 , n8838 );
and ( n8869 , n8865 , n8868 );
and ( n8870 , n8863 , n8868 );
or ( n8871 , n8866 , n8869 , n8870 );
xor ( n8872 , n8841 , n8843 );
xor ( n8873 , n8872 , n8846 );
and ( n8874 , n8871 , n8873 );
xor ( n8875 , n8077 , n8859 );
and ( n8876 , n8110 , n8113 );
and ( n8877 , n8113 , n8065 );
and ( n8878 , n8110 , n8065 );
or ( n8879 , n8876 , n8877 , n8878 );
and ( n8880 , n8875 , n8879 );
buf ( n8881 , n8032 );
and ( n8882 , n8077 , n8881 );
and ( n8883 , n8879 , n8882 );
and ( n8884 , n8875 , n8882 );
or ( n8885 , n8880 , n8883 , n8884 );
xor ( n8886 , n8110 , n8113 );
xor ( n8887 , n8886 , n8065 );
and ( n8888 , n8885 , n8887 );
xor ( n8889 , n8853 , n8857 );
xor ( n8890 , n8889 , n8860 );
and ( n8891 , n8887 , n8890 );
and ( n8892 , n8885 , n8890 );
or ( n8893 , n8888 , n8891 , n8892 );
xor ( n8894 , n8863 , n8865 );
xor ( n8895 , n8894 , n8868 );
and ( n8896 , n8893 , n8895 );
xor ( n8897 , n8077 , n8881 );
and ( n8898 , n8110 , n8113 );
and ( n8899 , n8113 , n8065 );
and ( n8900 , n8110 , n8065 );
or ( n8901 , n8898 , n8899 , n8900 );
and ( n8902 , n8897 , n8901 );
buf ( n8903 , n8033 );
and ( n8904 , n8077 , n8903 );
and ( n8905 , n8901 , n8904 );
and ( n8906 , n8897 , n8904 );
or ( n8907 , n8902 , n8905 , n8906 );
xor ( n8908 , n8110 , n8113 );
xor ( n8909 , n8908 , n8065 );
and ( n8910 , n8907 , n8909 );
xor ( n8911 , n8875 , n8879 );
xor ( n8912 , n8911 , n8882 );
and ( n8913 , n8909 , n8912 );
and ( n8914 , n8907 , n8912 );
or ( n8915 , n8910 , n8913 , n8914 );
xor ( n8916 , n8885 , n8887 );
xor ( n8917 , n8916 , n8890 );
and ( n8918 , n8915 , n8917 );
xor ( n8919 , n8110 , n8113 );
xor ( n8920 , n8919 , n8065 );
xor ( n8921 , n8897 , n8901 );
xor ( n8922 , n8921 , n8904 );
and ( n8923 , n8920 , n8922 );
xor ( n8924 , n8920 , n8922 );
buf ( n8925 , n8034 );
and ( n8926 , n8077 , n8925 );
buf ( n8927 , n5698 );
buf ( n8928 , n8927 );
and ( n8929 , n8928 , n8058 );
and ( n8930 , n8926 , n8929 );
xor ( n8931 , n8110 , n8113 );
xor ( n8932 , n8931 , n8065 );
xor ( n8933 , n8077 , n8903 );
xor ( n8934 , n8932 , n8933 );
and ( n8935 , n8929 , n8934 );
and ( n8936 , n8926 , n8934 );
or ( n8937 , n8930 , n8935 , n8936 );
and ( n8938 , n8924 , n8937 );
and ( n8939 , n8932 , n8933 );
and ( n8940 , n8937 , n8939 );
and ( n8941 , n8924 , n8939 );
or ( n8942 , n8938 , n8940 , n8941 );
and ( n8943 , n8923 , n8942 );
xor ( n8944 , n8907 , n8909 );
xor ( n8945 , n8944 , n8912 );
and ( n8946 , n8942 , n8945 );
and ( n8947 , n8923 , n8945 );
or ( n8948 , n8943 , n8946 , n8947 );
and ( n8949 , n8917 , n8948 );
and ( n8950 , n8915 , n8948 );
or ( n8951 , n8918 , n8949 , n8950 );
and ( n8952 , n8895 , n8951 );
and ( n8953 , n8893 , n8951 );
or ( n8954 , n8896 , n8952 , n8953 );
and ( n8955 , n8873 , n8954 );
and ( n8956 , n8871 , n8954 );
or ( n8957 , n8874 , n8955 , n8956 );
and ( n8958 , n8851 , n8957 );
and ( n8959 , n8849 , n8957 );
or ( n8960 , n8852 , n8958 , n8959 );
and ( n8961 , n8829 , n8960 );
and ( n8962 , n8827 , n8960 );
or ( n8963 , n8830 , n8961 , n8962 );
and ( n8964 , n8807 , n8963 );
and ( n8965 , n8805 , n8963 );
or ( n8966 , n8808 , n8964 , n8965 );
and ( n8967 , n8785 , n8966 );
and ( n8968 , n8783 , n8966 );
or ( n8969 , n8786 , n8967 , n8968 );
and ( n8970 , n8763 , n8969 );
and ( n8971 , n8761 , n8969 );
or ( n8972 , n8764 , n8970 , n8971 );
and ( n8973 , n8741 , n8972 );
and ( n8974 , n8739 , n8972 );
or ( n8975 , n8742 , n8973 , n8974 );
and ( n8976 , n8719 , n8975 );
and ( n8977 , n8717 , n8975 );
or ( n8978 , n8720 , n8976 , n8977 );
and ( n8979 , n8697 , n8978 );
and ( n8980 , n8695 , n8978 );
or ( n8981 , n8698 , n8979 , n8980 );
and ( n8982 , n8675 , n8981 );
and ( n8983 , n8673 , n8981 );
or ( n8984 , n8676 , n8982 , n8983 );
and ( n8985 , n8653 , n8984 );
and ( n8986 , n8651 , n8984 );
or ( n8987 , n8654 , n8985 , n8986 );
and ( n8988 , n8631 , n8987 );
and ( n8989 , n8629 , n8987 );
or ( n8990 , n8632 , n8988 , n8989 );
and ( n8991 , n8609 , n8990 );
and ( n8992 , n8607 , n8990 );
or ( n8993 , n8610 , n8991 , n8992 );
and ( n8994 , n8587 , n8993 );
and ( n8995 , n8585 , n8993 );
or ( n8996 , n8588 , n8994 , n8995 );
and ( n8997 , n8565 , n8996 );
and ( n8998 , n8563 , n8996 );
or ( n8999 , n8566 , n8997 , n8998 );
and ( n9000 , n8543 , n8999 );
and ( n9001 , n8541 , n8999 );
or ( n9002 , n8544 , n9000 , n9001 );
and ( n9003 , n8521 , n9002 );
and ( n9004 , n8519 , n9002 );
or ( n9005 , n8522 , n9003 , n9004 );
and ( n9006 , n8499 , n9005 );
and ( n9007 , n8497 , n9005 );
or ( n9008 , n8500 , n9006 , n9007 );
and ( n9009 , n8477 , n9008 );
and ( n9010 , n8475 , n9008 );
or ( n9011 , n8478 , n9009 , n9010 );
and ( n9012 , n8455 , n9011 );
and ( n9013 , n8453 , n9011 );
or ( n9014 , n8456 , n9012 , n9013 );
and ( n9015 , n8433 , n9014 );
and ( n9016 , n8414 , n9014 );
or ( n9017 , n8434 , n9015 , n9016 );
and ( n9018 , n8411 , n9017 );
and ( n9019 , n8392 , n9017 );
or ( n9020 , n8412 , n9018 , n9019 );
and ( n9021 , n8389 , n9020 );
and ( n9022 , n8370 , n9020 );
or ( n9023 , n8390 , n9021 , n9022 );
and ( n9024 , n8367 , n9023 );
and ( n9025 , n8348 , n9023 );
or ( n9026 , n8368 , n9024 , n9025 );
and ( n9027 , n8345 , n9026 );
and ( n9028 , n8326 , n9026 );
or ( n9029 , n8346 , n9027 , n9028 );
and ( n9030 , n8323 , n9029 );
and ( n9031 , n8304 , n9029 );
or ( n9032 , n8324 , n9030 , n9031 );
and ( n9033 , n8301 , n9032 );
and ( n9034 , n8282 , n9032 );
or ( n9035 , n8302 , n9033 , n9034 );
and ( n9036 , n8279 , n9035 );
and ( n9037 , n8260 , n9035 );
or ( n9038 , n8280 , n9036 , n9037 );
and ( n9039 , n8257 , n9038 );
and ( n9040 , n8238 , n9038 );
or ( n9041 , n8258 , n9039 , n9040 );
and ( n9042 , n8235 , n9041 );
and ( n9043 , n8233 , n9041 );
or ( n9044 , n8236 , n9042 , n9043 );
and ( n9045 , n8213 , n9044 );
and ( n9046 , n8211 , n9044 );
or ( n9047 , n8214 , n9045 , n9046 );
and ( n9048 , n8193 , n9047 );
xor ( n9049 , n8193 , n9047 );
xor ( n9050 , n8211 , n8213 );
xor ( n9051 , n9050 , n9044 );
not ( n9052 , n9051 );
xor ( n9053 , n8233 , n8235 );
xor ( n9054 , n9053 , n9041 );
xor ( n9055 , n8238 , n8257 );
xor ( n9056 , n9055 , n9038 );
xor ( n9057 , n8260 , n8279 );
xor ( n9058 , n9057 , n9035 );
xor ( n9059 , n8282 , n8301 );
xor ( n9060 , n9059 , n9032 );
xor ( n9061 , n8304 , n8323 );
xor ( n9062 , n9061 , n9029 );
xor ( n9063 , n8326 , n8345 );
xor ( n9064 , n9063 , n9026 );
xor ( n9065 , n8348 , n8367 );
xor ( n9066 , n9065 , n9023 );
xor ( n9067 , n8370 , n8389 );
xor ( n9068 , n9067 , n9020 );
xor ( n9069 , n8392 , n8411 );
xor ( n9070 , n9069 , n9017 );
xor ( n9071 , n8414 , n8433 );
xor ( n9072 , n9071 , n9014 );
xor ( n9073 , n8453 , n8455 );
xor ( n9074 , n9073 , n9011 );
xor ( n9075 , n8475 , n8477 );
xor ( n9076 , n9075 , n9008 );
xor ( n9077 , n8497 , n8499 );
xor ( n9078 , n9077 , n9005 );
xor ( n9079 , n8519 , n8521 );
xor ( n9080 , n9079 , n9002 );
xor ( n9081 , n8541 , n8543 );
xor ( n9082 , n9081 , n8999 );
xor ( n9083 , n8563 , n8565 );
xor ( n9084 , n9083 , n8996 );
xor ( n9085 , n8585 , n8587 );
xor ( n9086 , n9085 , n8993 );
xor ( n9087 , n8607 , n8609 );
xor ( n9088 , n9087 , n8990 );
xor ( n9089 , n8629 , n8631 );
xor ( n9090 , n9089 , n8987 );
xor ( n9091 , n8651 , n8653 );
xor ( n9092 , n9091 , n8984 );
xor ( n9093 , n8673 , n8675 );
xor ( n9094 , n9093 , n8981 );
xor ( n9095 , n8695 , n8697 );
xor ( n9096 , n9095 , n8978 );
xor ( n9097 , n8717 , n8719 );
xor ( n9098 , n9097 , n8975 );
xor ( n9099 , n8739 , n8741 );
xor ( n9100 , n9099 , n8972 );
xor ( n9101 , n8761 , n8763 );
xor ( n9102 , n9101 , n8969 );
xor ( n9103 , n8783 , n8785 );
xor ( n9104 , n9103 , n8966 );
xor ( n9105 , n8805 , n8807 );
xor ( n9106 , n9105 , n8963 );
xor ( n9107 , n8827 , n8829 );
xor ( n9108 , n9107 , n8960 );
xor ( n9109 , n8849 , n8851 );
xor ( n9110 , n9109 , n8957 );
xor ( n9111 , n8871 , n8873 );
xor ( n9112 , n9111 , n8954 );
xor ( n9113 , n8893 , n8895 );
xor ( n9114 , n9113 , n8951 );
xor ( n9115 , n8915 , n8917 );
xor ( n9116 , n9115 , n8948 );
xor ( n9117 , n8923 , n8942 );
xor ( n9118 , n9117 , n8945 );
buf ( n9119 , n8035 );
and ( n9120 , n8077 , n9119 );
and ( n9121 , n9120 , n8110 );
and ( n9122 , n8110 , n8113 );
and ( n9123 , n9120 , n8113 );
or ( n9124 , n9121 , n9122 , n9123 );
buf ( n9125 , n5700 );
buf ( n9126 , n9125 );
and ( n9127 , n9126 , n8058 );
xor ( n9128 , n8077 , n8925 );
and ( n9129 , n9127 , n9128 );
and ( n9130 , n8110 , n8113 );
and ( n9131 , n9128 , n9130 );
and ( n9132 , n9127 , n9130 );
or ( n9133 , n9129 , n9131 , n9132 );
and ( n9134 , n9124 , n9133 );
xor ( n9135 , n8058 , n8060 );
xor ( n9136 , n8060 , n8062 );
not ( n9137 , n9136 );
and ( n9138 , n9135 , n9137 );
and ( n9139 , n8928 , n9138 );
not ( n9140 , n9139 );
xnor ( n9141 , n9140 , n8065 );
xor ( n9142 , n9120 , n8110 );
xor ( n9143 , n9142 , n8113 );
and ( n9144 , n9141 , n9143 );
buf ( n9145 , n5702 );
buf ( n9146 , n9145 );
and ( n9147 , n9146 , n8058 );
xor ( n9148 , n8110 , n8113 );
and ( n9149 , n9147 , n9148 );
xor ( n9150 , n8077 , n9119 );
and ( n9151 , n9148 , n9150 );
and ( n9152 , n9147 , n9150 );
or ( n9153 , n9149 , n9151 , n9152 );
and ( n9154 , n9143 , n9153 );
and ( n9155 , n9141 , n9153 );
or ( n9156 , n9144 , n9154 , n9155 );
and ( n9157 , n9133 , n9156 );
and ( n9158 , n9124 , n9156 );
or ( n9159 , n9134 , n9157 , n9158 );
xor ( n9160 , n8924 , n8937 );
xor ( n9161 , n9160 , n8939 );
and ( n9162 , n9159 , n9161 );
xor ( n9163 , n8926 , n8929 );
xor ( n9164 , n9163 , n8934 );
xor ( n9165 , n9127 , n9128 );
xor ( n9166 , n9165 , n9130 );
and ( n9167 , n8110 , n8113 );
and ( n9168 , n9126 , n9138 );
and ( n9169 , n8928 , n9136 );
nor ( n9170 , n9168 , n9169 );
xnor ( n9171 , n9170 , n8065 );
and ( n9172 , n9167 , n9171 );
buf ( n9173 , n5704 );
buf ( n9174 , n9173 );
and ( n9175 , n9174 , n8058 );
buf ( n9176 , n8036 );
and ( n9177 , n9175 , n9176 );
xor ( n9178 , n8110 , n8113 );
and ( n9179 , n9176 , n9178 );
and ( n9180 , n9175 , n9178 );
or ( n9181 , n9177 , n9179 , n9180 );
and ( n9182 , n9171 , n9181 );
and ( n9183 , n9167 , n9181 );
or ( n9184 , n9172 , n9182 , n9183 );
and ( n9185 , n9166 , n9184 );
xor ( n9186 , n9141 , n9143 );
xor ( n9187 , n9186 , n9153 );
and ( n9188 , n9184 , n9187 );
and ( n9189 , n9166 , n9187 );
or ( n9190 , n9185 , n9188 , n9189 );
and ( n9191 , n9164 , n9190 );
xor ( n9192 , n9124 , n9133 );
xor ( n9193 , n9192 , n9156 );
and ( n9194 , n9190 , n9193 );
and ( n9195 , n9164 , n9193 );
or ( n9196 , n9191 , n9194 , n9195 );
and ( n9197 , n9161 , n9196 );
and ( n9198 , n9159 , n9196 );
or ( n9199 , n9162 , n9197 , n9198 );
and ( n9200 , n9118 , n9199 );
xor ( n9201 , n9118 , n9199 );
xor ( n9202 , n9159 , n9161 );
xor ( n9203 , n9202 , n9196 );
xor ( n9204 , n9164 , n9190 );
xor ( n9205 , n9204 , n9193 );
xor ( n9206 , n9147 , n9148 );
xor ( n9207 , n9206 , n9150 );
xor ( n9208 , n8110 , n8113 );
buf ( n9209 , n5706 );
buf ( n9210 , n9209 );
and ( n9211 , n9210 , n8058 );
and ( n9212 , n9208 , n9211 );
buf ( n9213 , n8037 );
and ( n9214 , n9211 , n9213 );
and ( n9215 , n9208 , n9213 );
or ( n9216 , n9212 , n9214 , n9215 );
xor ( n9217 , n8062 , n8072 );
xor ( n9218 , n8072 , n8074 );
not ( n9219 , n9218 );
and ( n9220 , n9217 , n9219 );
and ( n9221 , n8928 , n9220 );
not ( n9222 , n9221 );
xnor ( n9223 , n9222 , n8077 );
and ( n9224 , n9216 , n9223 );
and ( n9225 , n9207 , n9224 );
and ( n9226 , n8110 , n8113 );
and ( n9227 , n9146 , n9138 );
and ( n9228 , n9126 , n9136 );
nor ( n9229 , n9227 , n9228 );
xnor ( n9230 , n9229 , n8065 );
and ( n9231 , n9226 , n9230 );
and ( n9232 , n9174 , n9138 );
and ( n9233 , n9146 , n9136 );
nor ( n9234 , n9232 , n9233 );
xnor ( n9235 , n9234 , n8065 );
buf ( n9236 , n8038 );
and ( n9237 , n8110 , n9236 );
and ( n9238 , n9235 , n9237 );
and ( n9239 , n9126 , n9220 );
and ( n9240 , n8928 , n9218 );
nor ( n9241 , n9239 , n9240 );
xnor ( n9242 , n9241 , n8077 );
and ( n9243 , n9237 , n9242 );
and ( n9244 , n9235 , n9242 );
or ( n9245 , n9238 , n9243 , n9244 );
and ( n9246 , n9230 , n9245 );
and ( n9247 , n9226 , n9245 );
or ( n9248 , n9231 , n9246 , n9247 );
and ( n9249 , n9224 , n9248 );
and ( n9250 , n9207 , n9248 );
or ( n9251 , n9225 , n9249 , n9250 );
xor ( n9252 , n9166 , n9184 );
xor ( n9253 , n9252 , n9187 );
and ( n9254 , n9251 , n9253 );
xor ( n9255 , n9167 , n9171 );
xor ( n9256 , n9255 , n9181 );
xor ( n9257 , n9175 , n9176 );
xor ( n9258 , n9257 , n9178 );
xor ( n9259 , n9216 , n9223 );
and ( n9260 , n9258 , n9259 );
xor ( n9261 , n9208 , n9211 );
xor ( n9262 , n9261 , n9213 );
xor ( n9263 , n8074 , n8108 );
xor ( n9264 , n8108 , n8110 );
not ( n9265 , n9264 );
and ( n9266 , n9263 , n9265 );
and ( n9267 , n8928 , n9266 );
not ( n9268 , n9267 );
xnor ( n9269 , n9268 , n8113 );
xor ( n9270 , n8110 , n9236 );
and ( n9271 , n9269 , n9270 );
and ( n9272 , n9262 , n9271 );
and ( n9273 , n9210 , n9138 );
and ( n9274 , n9174 , n9136 );
nor ( n9275 , n9273 , n9274 );
xnor ( n9276 , n9275 , n8065 );
buf ( n9277 , n5708 );
buf ( n9278 , n9277 );
and ( n9279 , n9278 , n8058 );
and ( n9280 , n9276 , n9279 );
and ( n9281 , n9126 , n9266 );
and ( n9282 , n8928 , n9264 );
nor ( n9283 , n9281 , n9282 );
xnor ( n9284 , n9283 , n8113 );
and ( n9285 , n9174 , n9220 );
and ( n9286 , n9146 , n9218 );
nor ( n9287 , n9285 , n9286 );
xnor ( n9288 , n9287 , n8077 );
and ( n9289 , n9284 , n9288 );
and ( n9290 , n9278 , n9138 );
and ( n9291 , n9210 , n9136 );
nor ( n9292 , n9290 , n9291 );
xnor ( n9293 , n9292 , n8065 );
and ( n9294 , n9288 , n9293 );
and ( n9295 , n9284 , n9293 );
or ( n9296 , n9289 , n9294 , n9295 );
and ( n9297 , n9279 , n9296 );
and ( n9298 , n9276 , n9296 );
or ( n9299 , n9280 , n9297 , n9298 );
and ( n9300 , n9271 , n9299 );
and ( n9301 , n9262 , n9299 );
or ( n9302 , n9272 , n9300 , n9301 );
and ( n9303 , n9259 , n9302 );
and ( n9304 , n9258 , n9302 );
or ( n9305 , n9260 , n9303 , n9304 );
and ( n9306 , n9256 , n9305 );
xor ( n9307 , n9207 , n9224 );
xor ( n9308 , n9307 , n9248 );
and ( n9309 , n9305 , n9308 );
and ( n9310 , n9256 , n9308 );
or ( n9311 , n9306 , n9309 , n9310 );
and ( n9312 , n9253 , n9311 );
and ( n9313 , n9251 , n9311 );
or ( n9314 , n9254 , n9312 , n9313 );
and ( n9315 , n9205 , n9314 );
xor ( n9316 , n9205 , n9314 );
xor ( n9317 , n9251 , n9253 );
xor ( n9318 , n9317 , n9311 );
xor ( n9319 , n9226 , n9230 );
xor ( n9320 , n9319 , n9245 );
xor ( n9321 , n9235 , n9237 );
xor ( n9322 , n9321 , n9242 );
and ( n9323 , n9146 , n9220 );
and ( n9324 , n9126 , n9218 );
nor ( n9325 , n9323 , n9324 );
xnor ( n9326 , n9325 , n8077 );
xor ( n9327 , n9269 , n9270 );
and ( n9328 , n9326 , n9327 );
buf ( n9329 , n5710 );
buf ( n9330 , n9329 );
and ( n9331 , n9330 , n8058 );
buf ( n9332 , n8039 );
and ( n9333 , n9331 , n9332 );
buf ( n9334 , n5712 );
buf ( n9335 , n9334 );
and ( n9336 , n9335 , n8058 );
buf ( n9337 , n8040 );
and ( n9338 , n9336 , n9337 );
and ( n9339 , n9332 , n9338 );
and ( n9340 , n9331 , n9338 );
or ( n9341 , n9333 , n9339 , n9340 );
and ( n9342 , n9327 , n9341 );
and ( n9343 , n9326 , n9341 );
or ( n9344 , n9328 , n9342 , n9343 );
and ( n9345 , n9322 , n9344 );
xor ( n9346 , n9262 , n9271 );
xor ( n9347 , n9346 , n9299 );
and ( n9348 , n9344 , n9347 );
and ( n9349 , n9322 , n9347 );
or ( n9350 , n9345 , n9348 , n9349 );
and ( n9351 , n9320 , n9350 );
xor ( n9352 , n9258 , n9259 );
xor ( n9353 , n9352 , n9302 );
and ( n9354 , n9350 , n9353 );
and ( n9355 , n9320 , n9353 );
or ( n9356 , n9351 , n9354 , n9355 );
xor ( n9357 , n9256 , n9305 );
xor ( n9358 , n9357 , n9308 );
and ( n9359 , n9356 , n9358 );
xor ( n9360 , n9356 , n9358 );
xor ( n9361 , n9320 , n9350 );
xor ( n9362 , n9361 , n9353 );
xor ( n9363 , n9276 , n9279 );
xor ( n9364 , n9363 , n9296 );
xor ( n9365 , n9284 , n9288 );
xor ( n9366 , n9365 , n9293 );
and ( n9367 , n8110 , n9366 );
and ( n9368 , n9210 , n9220 );
and ( n9369 , n9174 , n9218 );
nor ( n9370 , n9368 , n9369 );
xnor ( n9371 , n9370 , n8077 );
and ( n9372 , n9330 , n9138 );
and ( n9373 , n9278 , n9136 );
nor ( n9374 , n9372 , n9373 );
xnor ( n9375 , n9374 , n8065 );
and ( n9376 , n9371 , n9375 );
xor ( n9377 , n9336 , n9337 );
and ( n9378 , n9375 , n9377 );
and ( n9379 , n9371 , n9377 );
or ( n9380 , n9376 , n9378 , n9379 );
and ( n9381 , n9366 , n9380 );
and ( n9382 , n8110 , n9380 );
or ( n9383 , n9367 , n9381 , n9382 );
and ( n9384 , n9364 , n9383 );
xor ( n9385 , n9326 , n9327 );
xor ( n9386 , n9385 , n9341 );
and ( n9387 , n9383 , n9386 );
and ( n9388 , n9364 , n9386 );
or ( n9389 , n9384 , n9387 , n9388 );
xor ( n9390 , n9322 , n9344 );
xor ( n9391 , n9390 , n9347 );
and ( n9392 , n9389 , n9391 );
xor ( n9393 , n9331 , n9332 );
xor ( n9394 , n9393 , n9338 );
buf ( n9395 , n7972 );
buf ( n9396 , n9395 );
buf ( n9397 , n8042 );
and ( n9398 , n9396 , n9397 );
buf ( n9399 , n5714 );
buf ( n9400 , n9399 );
and ( n9401 , n9400 , n8058 );
and ( n9402 , n9398 , n9401 );
buf ( n9403 , n8041 );
and ( n9404 , n9401 , n9403 );
and ( n9405 , n9398 , n9403 );
or ( n9406 , n9402 , n9404 , n9405 );
buf ( n9407 , n385 );
buf ( n9408 , n9407 );
xor ( n9409 , n8110 , n9408 );
not ( n9410 , n9408 );
and ( n9411 , n9409 , n9410 );
and ( n9412 , n8928 , n9411 );
not ( n9413 , n9412 );
xnor ( n9414 , n9413 , n8110 );
and ( n9415 , n9406 , n9414 );
and ( n9416 , n9394 , n9415 );
and ( n9417 , n9146 , n9266 );
and ( n9418 , n9126 , n9264 );
nor ( n9419 , n9417 , n9418 );
xnor ( n9420 , n9419 , n8113 );
and ( n9421 , n9278 , n9220 );
and ( n9422 , n9210 , n9218 );
nor ( n9423 , n9421 , n9422 );
xnor ( n9424 , n9423 , n8077 );
and ( n9425 , n9330 , n9220 );
and ( n9426 , n9278 , n9218 );
nor ( n9427 , n9425 , n9426 );
xnor ( n9428 , n9427 , n8077 );
and ( n9429 , n9400 , n9138 );
and ( n9430 , n9335 , n9136 );
nor ( n9431 , n9429 , n9430 );
xnor ( n9432 , n9431 , n8065 );
and ( n9433 , n9428 , n9432 );
and ( n9434 , n9424 , n9433 );
and ( n9435 , n9146 , n9411 );
and ( n9436 , n9126 , n9408 );
nor ( n9437 , n9435 , n9436 );
xnor ( n9438 , n9437 , n8110 );
and ( n9439 , n9210 , n9266 );
and ( n9440 , n9174 , n9264 );
nor ( n9441 , n9439 , n9440 );
xnor ( n9442 , n9441 , n8113 );
and ( n9443 , n9438 , n9442 );
and ( n9444 , n9433 , n9443 );
and ( n9445 , n9424 , n9443 );
or ( n9446 , n9434 , n9444 , n9445 );
and ( n9447 , n9420 , n9446 );
xor ( n9448 , n9371 , n9375 );
xor ( n9449 , n9448 , n9377 );
and ( n9450 , n9446 , n9449 );
and ( n9451 , n9420 , n9449 );
or ( n9452 , n9447 , n9450 , n9451 );
and ( n9453 , n9415 , n9452 );
and ( n9454 , n9394 , n9452 );
or ( n9455 , n9416 , n9453 , n9454 );
xor ( n9456 , n9364 , n9383 );
xor ( n9457 , n9456 , n9386 );
and ( n9458 , n9455 , n9457 );
xor ( n9459 , n8110 , n9366 );
xor ( n9460 , n9459 , n9380 );
xor ( n9461 , n9406 , n9414 );
and ( n9462 , n9174 , n9266 );
and ( n9463 , n9146 , n9264 );
nor ( n9464 , n9462 , n9463 );
xnor ( n9465 , n9464 , n8113 );
xor ( n9466 , n9398 , n9401 );
xor ( n9467 , n9466 , n9403 );
and ( n9468 , n9465 , n9467 );
and ( n9469 , n9461 , n9468 );
xor ( n9470 , n9396 , n9397 );
buf ( n9471 , n5718 );
buf ( n9472 , n9471 );
and ( n9473 , n9472 , n8058 );
buf ( n9474 , n8043 );
and ( n9475 , n9473 , n9474 );
and ( n9476 , n9470 , n9475 );
buf ( n9477 , n5716 );
buf ( n9478 , n9477 );
and ( n9479 , n9478 , n8058 );
and ( n9480 , n9475 , n9479 );
and ( n9481 , n9470 , n9479 );
or ( n9482 , n9476 , n9480 , n9481 );
and ( n9483 , n9335 , n9138 );
and ( n9484 , n9330 , n9136 );
nor ( n9485 , n9483 , n9484 );
xnor ( n9486 , n9485 , n8065 );
and ( n9487 , n9482 , n9486 );
and ( n9488 , n9468 , n9487 );
and ( n9489 , n9461 , n9487 );
or ( n9490 , n9469 , n9488 , n9489 );
and ( n9491 , n9460 , n9490 );
xor ( n9492 , n9394 , n9415 );
xor ( n9493 , n9492 , n9452 );
and ( n9494 , n9490 , n9493 );
and ( n9495 , n9460 , n9493 );
or ( n9496 , n9491 , n9494 , n9495 );
and ( n9497 , n9457 , n9496 );
and ( n9498 , n9455 , n9496 );
or ( n9499 , n9458 , n9497 , n9498 );
and ( n9500 , n9391 , n9499 );
and ( n9501 , n9389 , n9499 );
or ( n9502 , n9392 , n9500 , n9501 );
and ( n9503 , n9362 , n9502 );
xor ( n9504 , n9362 , n9502 );
xor ( n9505 , n9389 , n9391 );
xor ( n9506 , n9505 , n9499 );
xor ( n9507 , n9455 , n9457 );
xor ( n9508 , n9507 , n9496 );
and ( n9509 , n9126 , n9411 );
and ( n9510 , n8928 , n9408 );
nor ( n9511 , n9509 , n9510 );
xnor ( n9512 , n9511 , n8110 );
xor ( n9513 , n9428 , n9432 );
and ( n9514 , n9174 , n9411 );
and ( n9515 , n9146 , n9408 );
nor ( n9516 , n9514 , n9515 );
xnor ( n9517 , n9516 , n8110 );
and ( n9518 , n9335 , n9220 );
and ( n9519 , n9330 , n9218 );
nor ( n9520 , n9518 , n9519 );
xnor ( n9521 , n9520 , n8077 );
and ( n9522 , n9517 , n9521 );
and ( n9523 , n9513 , n9522 );
xor ( n9524 , n9438 , n9442 );
and ( n9525 , n9522 , n9524 );
and ( n9526 , n9513 , n9524 );
or ( n9527 , n9523 , n9525 , n9526 );
and ( n9528 , n9512 , n9527 );
xor ( n9529 , n9424 , n9433 );
xor ( n9530 , n9529 , n9443 );
and ( n9531 , n9527 , n9530 );
and ( n9532 , n9512 , n9530 );
or ( n9533 , n9528 , n9531 , n9532 );
xor ( n9534 , n9420 , n9446 );
xor ( n9535 , n9534 , n9449 );
and ( n9536 , n9533 , n9535 );
xor ( n9537 , n9465 , n9467 );
xor ( n9538 , n9482 , n9486 );
and ( n9539 , n9537 , n9538 );
xor ( n9540 , n9473 , n9474 );
buf ( n9541 , n5720 );
buf ( n9542 , n9541 );
and ( n9543 , n9542 , n8058 );
buf ( n9544 , n8044 );
and ( n9545 , n9543 , n9544 );
and ( n9546 , n9540 , n9545 );
buf ( n9547 , n7974 );
buf ( n9548 , n9547 );
and ( n9549 , n9545 , n9548 );
and ( n9550 , n9540 , n9548 );
or ( n9551 , n9546 , n9549 , n9550 );
xor ( n9552 , n9470 , n9475 );
xor ( n9553 , n9552 , n9479 );
and ( n9554 , n9551 , n9553 );
and ( n9555 , n9538 , n9554 );
and ( n9556 , n9537 , n9554 );
or ( n9557 , n9539 , n9555 , n9556 );
and ( n9558 , n9535 , n9557 );
and ( n9559 , n9533 , n9557 );
or ( n9560 , n9536 , n9558 , n9559 );
xor ( n9561 , n9460 , n9490 );
xor ( n9562 , n9561 , n9493 );
and ( n9563 , n9560 , n9562 );
xor ( n9564 , n9461 , n9468 );
xor ( n9565 , n9564 , n9487 );
xor ( n9566 , n9512 , n9527 );
xor ( n9567 , n9566 , n9530 );
and ( n9568 , n9478 , n9138 );
and ( n9569 , n9400 , n9136 );
nor ( n9570 , n9568 , n9569 );
xnor ( n9571 , n9570 , n8065 );
buf ( n9572 , n7976 );
buf ( n9573 , n9572 );
and ( n9574 , n9210 , n9411 );
and ( n9575 , n9174 , n9408 );
nor ( n9576 , n9574 , n9575 );
xnor ( n9577 , n9576 , n8110 );
and ( n9578 , n9573 , n9577 );
and ( n9579 , n9571 , n9578 );
and ( n9580 , n9330 , n9266 );
and ( n9581 , n9278 , n9264 );
nor ( n9582 , n9580 , n9581 );
xnor ( n9583 , n9582 , n8113 );
and ( n9584 , n9400 , n9220 );
and ( n9585 , n9335 , n9218 );
nor ( n9586 , n9584 , n9585 );
xnor ( n9587 , n9586 , n8077 );
and ( n9588 , n9583 , n9587 );
and ( n9589 , n9472 , n9138 );
and ( n9590 , n9478 , n9136 );
nor ( n9591 , n9589 , n9590 );
xnor ( n9592 , n9591 , n8065 );
and ( n9593 , n9587 , n9592 );
and ( n9594 , n9583 , n9592 );
or ( n9595 , n9588 , n9593 , n9594 );
and ( n9596 , n9578 , n9595 );
and ( n9597 , n9571 , n9595 );
or ( n9598 , n9579 , n9596 , n9597 );
xor ( n9599 , n9513 , n9522 );
xor ( n9600 , n9599 , n9524 );
and ( n9601 , n9598 , n9600 );
xor ( n9602 , n9551 , n9553 );
and ( n9603 , n9600 , n9602 );
and ( n9604 , n9598 , n9602 );
or ( n9605 , n9601 , n9603 , n9604 );
and ( n9606 , n9567 , n9605 );
xor ( n9607 , n9537 , n9538 );
xor ( n9608 , n9607 , n9554 );
and ( n9609 , n9605 , n9608 );
and ( n9610 , n9567 , n9608 );
or ( n9611 , n9606 , n9609 , n9610 );
and ( n9612 , n9565 , n9611 );
xor ( n9613 , n9533 , n9535 );
xor ( n9614 , n9613 , n9557 );
and ( n9615 , n9611 , n9614 );
and ( n9616 , n9565 , n9614 );
or ( n9617 , n9612 , n9615 , n9616 );
and ( n9618 , n9562 , n9617 );
and ( n9619 , n9560 , n9617 );
or ( n9620 , n9563 , n9618 , n9619 );
and ( n9621 , n9508 , n9620 );
xor ( n9622 , n9508 , n9620 );
xor ( n9623 , n9560 , n9562 );
xor ( n9624 , n9623 , n9617 );
xor ( n9625 , n9565 , n9611 );
xor ( n9626 , n9625 , n9614 );
and ( n9627 , n9278 , n9266 );
and ( n9628 , n9210 , n9264 );
nor ( n9629 , n9627 , n9628 );
xnor ( n9630 , n9629 , n8113 );
xor ( n9631 , n9540 , n9545 );
xor ( n9632 , n9631 , n9548 );
and ( n9633 , n9630 , n9632 );
xor ( n9634 , n9517 , n9521 );
and ( n9635 , n9335 , n9266 );
and ( n9636 , n9330 , n9264 );
nor ( n9637 , n9635 , n9636 );
xnor ( n9638 , n9637 , n8113 );
and ( n9639 , n9542 , n9138 );
and ( n9640 , n9472 , n9136 );
nor ( n9641 , n9639 , n9640 );
xnor ( n9642 , n9641 , n8065 );
and ( n9643 , n9638 , n9642 );
xor ( n9644 , n9573 , n9577 );
and ( n9645 , n9643 , n9644 );
xor ( n9646 , n9583 , n9587 );
xor ( n9647 , n9646 , n9592 );
and ( n9648 , n9644 , n9647 );
and ( n9649 , n9643 , n9647 );
or ( n9650 , n9645 , n9648 , n9649 );
and ( n9651 , n9634 , n9650 );
xor ( n9652 , n9571 , n9578 );
xor ( n9653 , n9652 , n9595 );
and ( n9654 , n9650 , n9653 );
and ( n9655 , n9634 , n9653 );
or ( n9656 , n9651 , n9654 , n9655 );
and ( n9657 , n9633 , n9656 );
xor ( n9658 , n9630 , n9632 );
buf ( n9659 , n5724 );
buf ( n9660 , n9659 );
and ( n9661 , n9660 , n8058 );
buf ( n9662 , n8046 );
and ( n9663 , n9661 , n9662 );
buf ( n9664 , n8045 );
and ( n9665 , n9663 , n9664 );
xor ( n9666 , n9543 , n9544 );
and ( n9667 , n9665 , n9666 );
and ( n9668 , n9658 , n9667 );
xor ( n9669 , n9634 , n9650 );
xor ( n9670 , n9669 , n9653 );
and ( n9671 , n9667 , n9670 );
and ( n9672 , n9658 , n9670 );
or ( n9673 , n9668 , n9671 , n9672 );
and ( n9674 , n9656 , n9673 );
and ( n9675 , n9633 , n9673 );
or ( n9676 , n9657 , n9674 , n9675 );
xor ( n9677 , n9567 , n9605 );
xor ( n9678 , n9677 , n9608 );
and ( n9679 , n9676 , n9678 );
xor ( n9680 , n9598 , n9600 );
xor ( n9681 , n9680 , n9602 );
xor ( n9682 , n9633 , n9656 );
xor ( n9683 , n9682 , n9673 );
and ( n9684 , n9681 , n9683 );
xor ( n9685 , n9643 , n9644 );
xor ( n9686 , n9685 , n9647 );
xor ( n9687 , n9665 , n9666 );
and ( n9688 , n9686 , n9687 );
xor ( n9689 , n9661 , n9662 );
buf ( n9690 , n394 );
buf ( n9691 , n9690 );
buf ( n9692 , n8047 );
and ( n9693 , n9691 , n9692 );
and ( n9694 , n9689 , n9693 );
buf ( n9695 , n5722 );
buf ( n9696 , n9695 );
and ( n9697 , n9696 , n9138 );
and ( n9698 , n9542 , n9136 );
nor ( n9699 , n9697 , n9698 );
xnor ( n9700 , n9699 , n8065 );
and ( n9701 , n9693 , n9700 );
and ( n9702 , n9689 , n9700 );
or ( n9703 , n9694 , n9701 , n9702 );
buf ( n9704 , n7978 );
buf ( n9705 , n9704 );
and ( n9706 , n9703 , n9705 );
and ( n9707 , n9478 , n9220 );
and ( n9708 , n9400 , n9218 );
nor ( n9709 , n9707 , n9708 );
xnor ( n9710 , n9709 , n8077 );
and ( n9711 , n9705 , n9710 );
and ( n9712 , n9703 , n9710 );
or ( n9713 , n9706 , n9711 , n9712 );
and ( n9714 , n9687 , n9713 );
and ( n9715 , n9686 , n9713 );
or ( n9716 , n9688 , n9714 , n9715 );
xor ( n9717 , n9658 , n9667 );
xor ( n9718 , n9717 , n9670 );
and ( n9719 , n9716 , n9718 );
and ( n9720 , n9696 , n8058 );
xor ( n9721 , n9663 , n9664 );
and ( n9722 , n9720 , n9721 );
and ( n9723 , n9278 , n9411 );
and ( n9724 , n9210 , n9408 );
nor ( n9725 , n9723 , n9724 );
xnor ( n9726 , n9725 , n8110 );
xor ( n9727 , n9703 , n9705 );
xor ( n9728 , n9727 , n9710 );
and ( n9729 , n9726 , n9728 );
and ( n9730 , n9722 , n9729 );
xor ( n9731 , n9638 , n9642 );
xor ( n9732 , n9720 , n9721 );
and ( n9733 , n9731 , n9732 );
xor ( n9734 , n9691 , n9692 );
buf ( n9735 , n395 );
buf ( n9736 , n9735 );
and ( n9737 , n9660 , n9136 );
and ( n9738 , n9736 , n9737 );
buf ( n9739 , n8048 );
and ( n9740 , n9737 , n9739 );
and ( n9741 , n9736 , n9739 );
or ( n9742 , n9738 , n9740 , n9741 );
and ( n9743 , n9734 , n9742 );
not ( n9744 , n9737 );
and ( n9745 , n9744 , n8065 );
and ( n9746 , n9742 , n9745 );
and ( n9747 , n9734 , n9745 );
or ( n9748 , n9743 , n9746 , n9747 );
buf ( n9749 , n7980 );
buf ( n9750 , n9749 );
and ( n9751 , n9748 , n9750 );
and ( n9752 , n9472 , n9220 );
and ( n9753 , n9478 , n9218 );
nor ( n9754 , n9752 , n9753 );
xnor ( n9755 , n9754 , n8077 );
and ( n9756 , n9750 , n9755 );
and ( n9757 , n9748 , n9755 );
or ( n9758 , n9751 , n9756 , n9757 );
and ( n9759 , n9732 , n9758 );
and ( n9760 , n9731 , n9758 );
or ( n9761 , n9733 , n9759 , n9760 );
and ( n9762 , n9729 , n9761 );
and ( n9763 , n9722 , n9761 );
or ( n9764 , n9730 , n9762 , n9763 );
and ( n9765 , n9718 , n9764 );
and ( n9766 , n9716 , n9764 );
or ( n9767 , n9719 , n9765 , n9766 );
and ( n9768 , n9683 , n9767 );
and ( n9769 , n9681 , n9767 );
or ( n9770 , n9684 , n9768 , n9769 );
and ( n9771 , n9678 , n9770 );
and ( n9772 , n9676 , n9770 );
or ( n9773 , n9679 , n9771 , n9772 );
and ( n9774 , n9626 , n9773 );
xor ( n9775 , n9626 , n9773 );
xor ( n9776 , n9676 , n9678 );
xor ( n9777 , n9776 , n9770 );
xor ( n9778 , n9681 , n9683 );
xor ( n9779 , n9778 , n9767 );
xor ( n9780 , n9686 , n9687 );
xor ( n9781 , n9780 , n9713 );
and ( n9782 , n9400 , n9266 );
and ( n9783 , n9335 , n9264 );
nor ( n9784 , n9782 , n9783 );
xnor ( n9785 , n9784 , n8113 );
xor ( n9786 , n9689 , n9693 );
xor ( n9787 , n9786 , n9700 );
and ( n9788 , n9785 , n9787 );
xor ( n9789 , n9726 , n9728 );
and ( n9790 , n9788 , n9789 );
buf ( n9791 , n7982 );
buf ( n9792 , n9791 );
and ( n9793 , n9478 , n9266 );
and ( n9794 , n9400 , n9264 );
nor ( n9795 , n9793 , n9794 );
xnor ( n9796 , n9795 , n8113 );
and ( n9797 , n9792 , n9796 );
and ( n9798 , n9542 , n9220 );
and ( n9799 , n9472 , n9218 );
nor ( n9800 , n9798 , n9799 );
xnor ( n9801 , n9800 , n8077 );
and ( n9802 , n9796 , n9801 );
and ( n9803 , n9792 , n9801 );
or ( n9804 , n9797 , n9802 , n9803 );
and ( n9805 , n9330 , n9411 );
and ( n9806 , n9278 , n9408 );
nor ( n9807 , n9805 , n9806 );
xnor ( n9808 , n9807 , n8110 );
and ( n9809 , n9804 , n9808 );
xor ( n9810 , n9748 , n9750 );
xor ( n9811 , n9810 , n9755 );
and ( n9812 , n9808 , n9811 );
and ( n9813 , n9804 , n9811 );
or ( n9814 , n9809 , n9812 , n9813 );
and ( n9815 , n9789 , n9814 );
and ( n9816 , n9788 , n9814 );
or ( n9817 , n9790 , n9815 , n9816 );
and ( n9818 , n9781 , n9817 );
xor ( n9819 , n9722 , n9729 );
xor ( n9820 , n9819 , n9761 );
and ( n9821 , n9817 , n9820 );
and ( n9822 , n9781 , n9820 );
or ( n9823 , n9818 , n9821 , n9822 );
xor ( n9824 , n9716 , n9718 );
xor ( n9825 , n9824 , n9764 );
and ( n9826 , n9823 , n9825 );
xor ( n9827 , n9823 , n9825 );
and ( n9828 , n9335 , n9411 );
and ( n9829 , n9330 , n9408 );
nor ( n9830 , n9828 , n9829 );
xnor ( n9831 , n9830 , n8110 );
and ( n9832 , n9660 , n9138 );
and ( n9833 , n9696 , n9136 );
nor ( n9834 , n9832 , n9833 );
xnor ( n9835 , n9834 , n8065 );
and ( n9836 , n9831 , n9835 );
xor ( n9837 , n9792 , n9796 );
xor ( n9838 , n9837 , n9801 );
and ( n9839 , n9835 , n9838 );
and ( n9840 , n9831 , n9838 );
or ( n9841 , n9836 , n9839 , n9840 );
buf ( n9842 , n7984 );
buf ( n9843 , n9842 );
and ( n9844 , n9400 , n9411 );
and ( n9845 , n9335 , n9408 );
nor ( n9846 , n9844 , n9845 );
xnor ( n9847 , n9846 , n8110 );
and ( n9848 , n9843 , n9847 );
and ( n9849 , n9472 , n9266 );
and ( n9850 , n9478 , n9264 );
nor ( n9851 , n9849 , n9850 );
xnor ( n9852 , n9851 , n8113 );
and ( n9853 , n9847 , n9852 );
and ( n9854 , n9843 , n9852 );
or ( n9855 , n9848 , n9853 , n9854 );
xor ( n9856 , n9734 , n9742 );
xor ( n9857 , n9856 , n9745 );
and ( n9858 , n9855 , n9857 );
buf ( n9859 , n396 );
buf ( n9860 , n9859 );
buf ( n9861 , n8049 );
and ( n9862 , n9860 , n9861 );
xor ( n9863 , n9736 , n9737 );
xor ( n9864 , n9863 , n9739 );
and ( n9865 , n9862 , n9864 );
and ( n9866 , n9857 , n9865 );
and ( n9867 , n9855 , n9865 );
or ( n9868 , n9858 , n9866 , n9867 );
and ( n9869 , n9841 , n9868 );
xor ( n9870 , n9785 , n9787 );
and ( n9871 , n9868 , n9870 );
and ( n9872 , n9841 , n9870 );
or ( n9873 , n9869 , n9871 , n9872 );
xor ( n9874 , n9731 , n9732 );
xor ( n9875 , n9874 , n9758 );
and ( n9876 , n9873 , n9875 );
xor ( n9877 , n9804 , n9808 );
xor ( n9878 , n9877 , n9811 );
and ( n9879 , n9696 , n9220 );
and ( n9880 , n9542 , n9218 );
nor ( n9881 , n9879 , n9880 );
xnor ( n9882 , n9881 , n8077 );
buf ( n9883 , n7986 );
buf ( n9884 , n9883 );
and ( n9885 , n9542 , n9266 );
and ( n9886 , n9472 , n9264 );
nor ( n9887 , n9885 , n9886 );
xnor ( n9888 , n9887 , n8113 );
and ( n9889 , n9884 , n9888 );
and ( n9890 , n9882 , n9889 );
and ( n9891 , n9478 , n9411 );
and ( n9892 , n9400 , n9408 );
nor ( n9893 , n9891 , n9892 );
xnor ( n9894 , n9893 , n8110 );
and ( n9895 , n9660 , n9220 );
and ( n9896 , n9696 , n9218 );
nor ( n9897 , n9895 , n9896 );
xnor ( n9898 , n9897 , n8077 );
and ( n9899 , n9894 , n9898 );
and ( n9900 , n9660 , n9218 );
not ( n9901 , n9900 );
and ( n9902 , n9901 , n8077 );
and ( n9903 , n9898 , n9902 );
and ( n9904 , n9894 , n9902 );
or ( n9905 , n9899 , n9903 , n9904 );
and ( n9906 , n9889 , n9905 );
and ( n9907 , n9882 , n9905 );
or ( n9908 , n9890 , n9906 , n9907 );
xor ( n9909 , n9831 , n9835 );
xor ( n9910 , n9909 , n9838 );
and ( n9911 , n9908 , n9910 );
xor ( n9912 , n9843 , n9847 );
xor ( n9913 , n9912 , n9852 );
xor ( n9914 , n9862 , n9864 );
and ( n9915 , n9913 , n9914 );
xor ( n9916 , n9884 , n9888 );
xor ( n9917 , n9860 , n9861 );
and ( n9918 , n9916 , n9917 );
buf ( n9919 , n397 );
buf ( n9920 , n9919 );
buf ( n9921 , n7988 );
buf ( n9922 , n9921 );
and ( n9923 , n9920 , n9922 );
and ( n9924 , n9472 , n9411 );
and ( n9925 , n9478 , n9408 );
nor ( n9926 , n9924 , n9925 );
xnor ( n9927 , n9926 , n8110 );
and ( n9928 , n9922 , n9927 );
and ( n9929 , n9920 , n9927 );
or ( n9930 , n9923 , n9928 , n9929 );
and ( n9931 , n9917 , n9930 );
and ( n9932 , n9916 , n9930 );
or ( n9933 , n9918 , n9931 , n9932 );
and ( n9934 , n9914 , n9933 );
and ( n9935 , n9913 , n9933 );
or ( n9936 , n9915 , n9934 , n9935 );
and ( n9937 , n9910 , n9936 );
and ( n9938 , n9908 , n9936 );
or ( n9939 , n9911 , n9937 , n9938 );
and ( n9940 , n9878 , n9939 );
xor ( n9941 , n9841 , n9868 );
xor ( n9942 , n9941 , n9870 );
and ( n9943 , n9939 , n9942 );
and ( n9944 , n9878 , n9942 );
or ( n9945 , n9940 , n9943 , n9944 );
and ( n9946 , n9875 , n9945 );
and ( n9947 , n9873 , n9945 );
or ( n9948 , n9876 , n9946 , n9947 );
xor ( n9949 , n9781 , n9817 );
xor ( n9950 , n9949 , n9820 );
and ( n9951 , n9948 , n9950 );
xor ( n9952 , n9948 , n9950 );
xor ( n9953 , n9788 , n9789 );
xor ( n9954 , n9953 , n9814 );
xor ( n9955 , n9873 , n9875 );
xor ( n9956 , n9955 , n9945 );
and ( n9957 , n9954 , n9956 );
xor ( n9958 , n9954 , n9956 );
xor ( n9959 , n9855 , n9857 );
xor ( n9960 , n9959 , n9865 );
xor ( n9961 , n9882 , n9889 );
xor ( n9962 , n9961 , n9905 );
and ( n9963 , n9696 , n9266 );
and ( n9964 , n9542 , n9264 );
nor ( n9965 , n9963 , n9964 );
xnor ( n9966 , n9965 , n8113 );
and ( n9967 , n9966 , n9900 );
buf ( n9968 , n8050 );
and ( n9969 , n9900 , n9968 );
and ( n9970 , n9966 , n9968 );
or ( n9971 , n9967 , n9969 , n9970 );
xor ( n9972 , n9894 , n9898 );
xor ( n9973 , n9972 , n9902 );
and ( n9974 , n9971 , n9973 );
buf ( n9975 , n398 );
buf ( n9976 , n9975 );
buf ( n9977 , n7990 );
buf ( n9978 , n9977 );
and ( n9979 , n9976 , n9978 );
and ( n9980 , n9542 , n9411 );
and ( n9981 , n9472 , n9408 );
nor ( n9982 , n9980 , n9981 );
xnor ( n9983 , n9982 , n8110 );
and ( n9984 , n9978 , n9983 );
and ( n9985 , n9976 , n9983 );
or ( n9986 , n9979 , n9984 , n9985 );
and ( n9987 , n9660 , n9266 );
and ( n9988 , n9696 , n9264 );
nor ( n9989 , n9987 , n9988 );
xnor ( n9990 , n9989 , n8113 );
and ( n9991 , n9660 , n9264 );
not ( n9992 , n9991 );
and ( n9993 , n9992 , n8113 );
and ( n9994 , n9990 , n9993 );
buf ( n9995 , n8051 );
and ( n9996 , n9993 , n9995 );
and ( n9997 , n9990 , n9995 );
or ( n9998 , n9994 , n9996 , n9997 );
and ( n9999 , n9986 , n9998 );
xor ( n10000 , n9920 , n9922 );
xor ( n10001 , n10000 , n9927 );
and ( n10002 , n9998 , n10001 );
and ( n10003 , n9986 , n10001 );
or ( n10004 , n9999 , n10002 , n10003 );
and ( n10005 , n9973 , n10004 );
and ( n10006 , n9971 , n10004 );
or ( n10007 , n9974 , n10005 , n10006 );
and ( n10008 , n9962 , n10007 );
xor ( n10009 , n9913 , n9914 );
xor ( n10010 , n10009 , n9933 );
and ( n10011 , n10007 , n10010 );
and ( n10012 , n9962 , n10010 );
or ( n10013 , n10008 , n10011 , n10012 );
and ( n10014 , n9960 , n10013 );
xor ( n10015 , n9908 , n9910 );
xor ( n10016 , n10015 , n9936 );
and ( n10017 , n10013 , n10016 );
and ( n10018 , n9960 , n10016 );
or ( n10019 , n10014 , n10017 , n10018 );
xor ( n10020 , n9878 , n9939 );
xor ( n10021 , n10020 , n9942 );
and ( n10022 , n10019 , n10021 );
xor ( n10023 , n10019 , n10021 );
xor ( n10024 , n9960 , n10013 );
xor ( n10025 , n10024 , n10016 );
xor ( n10026 , n9916 , n9917 );
xor ( n10027 , n10026 , n9930 );
xor ( n10028 , n9966 , n9900 );
xor ( n10029 , n10028 , n9968 );
buf ( n10030 , n399 );
buf ( n10031 , n10030 );
and ( n10032 , n9696 , n9411 );
and ( n10033 , n9542 , n9408 );
nor ( n10034 , n10032 , n10033 );
xnor ( n10035 , n10034 , n8110 );
and ( n10036 , n10031 , n10035 );
xor ( n10037 , n9976 , n9978 );
xor ( n10038 , n10037 , n9983 );
and ( n10039 , n10036 , n10038 );
xor ( n10040 , n9990 , n9993 );
xor ( n10041 , n10040 , n9995 );
and ( n10042 , n10038 , n10041 );
and ( n10043 , n10036 , n10041 );
or ( n10044 , n10039 , n10042 , n10043 );
and ( n10045 , n10029 , n10044 );
xor ( n10046 , n9986 , n9998 );
xor ( n10047 , n10046 , n10001 );
and ( n10048 , n10044 , n10047 );
and ( n10049 , n10029 , n10047 );
or ( n10050 , n10045 , n10048 , n10049 );
and ( n10051 , n10027 , n10050 );
xor ( n10052 , n9971 , n9973 );
xor ( n10053 , n10052 , n10004 );
and ( n10054 , n10050 , n10053 );
and ( n10055 , n10027 , n10053 );
or ( n10056 , n10051 , n10054 , n10055 );
xor ( n10057 , n9962 , n10007 );
xor ( n10058 , n10057 , n10010 );
and ( n10059 , n10056 , n10058 );
xor ( n10060 , n10056 , n10058 );
xor ( n10061 , n10027 , n10050 );
xor ( n10062 , n10061 , n10053 );
xor ( n10063 , n10029 , n10044 );
xor ( n10064 , n10063 , n10047 );
buf ( n10065 , n8052 );
and ( n10066 , n9991 , n10065 );
buf ( n10067 , n400 );
buf ( n10068 , n10067 );
and ( n10069 , n9660 , n9408 );
not ( n10070 , n10069 );
and ( n10071 , n10070 , n8110 );
and ( n10072 , n10068 , n10071 );
buf ( n10073 , n8053 );
and ( n10074 , n10071 , n10073 );
and ( n10075 , n10068 , n10073 );
or ( n10076 , n10072 , n10074 , n10075 );
and ( n10077 , n10065 , n10076 );
and ( n10078 , n9991 , n10076 );
or ( n10079 , n10066 , n10077 , n10078 );
xor ( n10080 , n10036 , n10038 );
xor ( n10081 , n10080 , n10041 );
and ( n10082 , n10079 , n10081 );
xor ( n10083 , n10031 , n10035 );
buf ( n10084 , n401 );
buf ( n10085 , n10084 );
and ( n10086 , n10085 , n10069 );
buf ( n10087 , n8054 );
and ( n10088 , n10069 , n10087 );
and ( n10089 , n10085 , n10087 );
or ( n10090 , n10086 , n10088 , n10089 );
and ( n10091 , n9660 , n9411 );
and ( n10092 , n9696 , n9408 );
nor ( n10093 , n10091 , n10092 );
xnor ( n10094 , n10093 , n8110 );
and ( n10095 , n10090 , n10094 );
xor ( n10096 , n10068 , n10071 );
xor ( n10097 , n10096 , n10073 );
and ( n10098 , n10094 , n10097 );
and ( n10099 , n10090 , n10097 );
or ( n10100 , n10095 , n10098 , n10099 );
and ( n10101 , n10083 , n10100 );
xor ( n10102 , n9991 , n10065 );
xor ( n10103 , n10102 , n10076 );
and ( n10104 , n10100 , n10103 );
and ( n10105 , n10083 , n10103 );
or ( n10106 , n10101 , n10104 , n10105 );
and ( n10107 , n10081 , n10106 );
and ( n10108 , n10079 , n10106 );
or ( n10109 , n10082 , n10107 , n10108 );
and ( n10110 , n10064 , n10109 );
and ( n10111 , n10062 , n10110 );
and ( n10112 , n10060 , n10111 );
or ( n10113 , n10059 , n10112 );
and ( n10114 , n10025 , n10113 );
and ( n10115 , n10023 , n10114 );
or ( n10116 , n10022 , n10115 );
and ( n10117 , n9958 , n10116 );
or ( n10118 , n9957 , n10117 );
and ( n10119 , n9952 , n10118 );
or ( n10120 , n9951 , n10119 );
and ( n10121 , n9827 , n10120 );
or ( n10122 , n9826 , n10121 );
and ( n10123 , n9779 , n10122 );
and ( n10124 , n9777 , n10123 );
and ( n10125 , n9775 , n10124 );
or ( n10126 , n9774 , n10125 );
and ( n10127 , n9624 , n10126 );
and ( n10128 , n9622 , n10127 );
or ( n10129 , n9621 , n10128 );
and ( n10130 , n9506 , n10129 );
and ( n10131 , n9504 , n10130 );
or ( n10132 , n9503 , n10131 );
and ( n10133 , n9360 , n10132 );
or ( n10134 , n9359 , n10133 );
and ( n10135 , n9318 , n10134 );
and ( n10136 , n9316 , n10135 );
or ( n10137 , n9315 , n10136 );
and ( n10138 , n9203 , n10137 );
and ( n10139 , n9201 , n10138 );
or ( n10140 , n9200 , n10139 );
and ( n10141 , n9116 , n10140 );
and ( n10142 , n9114 , n10141 );
and ( n10143 , n9112 , n10142 );
and ( n10144 , n9110 , n10143 );
and ( n10145 , n9108 , n10144 );
and ( n10146 , n9106 , n10145 );
and ( n10147 , n9104 , n10146 );
and ( n10148 , n9102 , n10147 );
and ( n10149 , n9100 , n10148 );
and ( n10150 , n9098 , n10149 );
and ( n10151 , n9096 , n10150 );
and ( n10152 , n9094 , n10151 );
and ( n10153 , n9092 , n10152 );
and ( n10154 , n9090 , n10153 );
and ( n10155 , n9088 , n10154 );
and ( n10156 , n9086 , n10155 );
and ( n10157 , n9084 , n10156 );
and ( n10158 , n9082 , n10157 );
and ( n10159 , n9080 , n10158 );
and ( n10160 , n9078 , n10159 );
and ( n10161 , n9076 , n10160 );
and ( n10162 , n9074 , n10161 );
and ( n10163 , n9072 , n10162 );
and ( n10164 , n9070 , n10163 );
and ( n10165 , n9068 , n10164 );
and ( n10166 , n9066 , n10165 );
and ( n10167 , n9064 , n10166 );
and ( n10168 , n9062 , n10167 );
and ( n10169 , n9060 , n10168 );
and ( n10170 , n9058 , n10169 );
and ( n10171 , n9056 , n10170 );
and ( n10172 , n9054 , n10171 );
and ( n10173 , n9052 , n10172 );
or ( n10174 , n9051 , n10173 );
and ( n10175 , n9049 , n10174 );
or ( n10176 , n9048 , n10175 );
and ( n10177 , n8191 , n10176 );
or ( n10178 , n8190 , n10177 );
and ( n10179 , n8188 , n10178 );
or ( n10180 , n8187 , n10179 );
and ( n10181 , n8130 , n10180 );
and ( n10182 , n8129 , n10181 );
or ( n10183 , n8128 , n10182 );
and ( n10184 , n8094 , n10183 );
and ( n10185 , n8093 , n10184 );
xor ( n10186 , n8092 , n10185 );
buf ( n10187 , n10186 );
xor ( n10188 , n8093 , n10184 );
buf ( n10189 , n10188 );
xor ( n10190 , n8094 , n10183 );
buf ( n10191 , n10190 );
xor ( n10192 , n8129 , n10181 );
buf ( n10193 , n10192 );
xor ( n10194 , n8130 , n10180 );
buf ( n10195 , n10194 );
xor ( n10196 , n8188 , n10178 );
buf ( n10197 , n10196 );
xor ( n10198 , n8191 , n10176 );
buf ( n10199 , n10198 );
xor ( n10200 , n9049 , n10174 );
buf ( n10201 , n10200 );
xor ( n10202 , n9052 , n10172 );
buf ( n10203 , n10202 );
xor ( n10204 , n9054 , n10171 );
buf ( n10205 , n10204 );
xor ( n10206 , n9056 , n10170 );
buf ( n10207 , n10206 );
xor ( n10208 , n9058 , n10169 );
buf ( n10209 , n10208 );
xor ( n10210 , n9060 , n10168 );
buf ( n10211 , n10210 );
xor ( n10212 , n9062 , n10167 );
buf ( n10213 , n10212 );
xor ( n10214 , n9064 , n10166 );
buf ( n10215 , n10214 );
xor ( n10216 , n9066 , n10165 );
buf ( n10217 , n10216 );
xor ( n10218 , n9068 , n10164 );
buf ( n10219 , n10218 );
xor ( n10220 , n9070 , n10163 );
buf ( n10221 , n10220 );
xor ( n10222 , n9072 , n10162 );
buf ( n10223 , n10222 );
xor ( n10224 , n9074 , n10161 );
buf ( n10225 , n10224 );
xor ( n10226 , n9076 , n10160 );
buf ( n10227 , n10226 );
xor ( n10228 , n9078 , n10159 );
buf ( n10229 , n10228 );
xor ( n10230 , n9080 , n10158 );
buf ( n10231 , n10230 );
xor ( n10232 , n9082 , n10157 );
buf ( n10233 , n10232 );
xor ( n10234 , n9084 , n10156 );
buf ( n10235 , n10234 );
xor ( n10236 , n9086 , n10155 );
buf ( n10237 , n10236 );
xor ( n10238 , n9088 , n10154 );
buf ( n10239 , n10238 );
xor ( n10240 , n9090 , n10153 );
buf ( n10241 , n10240 );
xor ( n10242 , n9092 , n10152 );
buf ( n10243 , n10242 );
xor ( n10244 , n9094 , n10151 );
buf ( n10245 , n10244 );
xor ( n10246 , n9096 , n10150 );
buf ( n10247 , n10246 );
xor ( n10248 , n9098 , n10149 );
buf ( n10249 , n10248 );
xor ( n10250 , n9100 , n10148 );
buf ( n10251 , n10250 );
xor ( n10252 , n9102 , n10147 );
buf ( n10253 , n10252 );
xor ( n10254 , n9104 , n10146 );
buf ( n10255 , n10254 );
xor ( n10256 , n9106 , n10145 );
buf ( n10257 , n10256 );
xor ( n10258 , n9108 , n10144 );
buf ( n10259 , n10258 );
xor ( n10260 , n9110 , n10143 );
buf ( n10261 , n10260 );
xor ( n10262 , n9112 , n10142 );
buf ( n10263 , n10262 );
xor ( n10264 , n9114 , n10141 );
buf ( n10265 , n10264 );
xor ( n10266 , n9116 , n10140 );
buf ( n10267 , n10266 );
xor ( n10268 , n9201 , n10138 );
buf ( n10269 , n10268 );
xor ( n10270 , n9203 , n10137 );
buf ( n10271 , n10270 );
xor ( n10272 , n9316 , n10135 );
buf ( n10273 , n10272 );
xor ( n10274 , n9318 , n10134 );
buf ( n10275 , n10274 );
xor ( n10276 , n9360 , n10132 );
buf ( n10277 , n10276 );
xor ( n10278 , n9504 , n10130 );
buf ( n10279 , n10278 );
xor ( n10280 , n9506 , n10129 );
buf ( n10281 , n10280 );
xor ( n10282 , n9622 , n10127 );
buf ( n10283 , n10282 );
xor ( n10284 , n9624 , n10126 );
buf ( n10285 , n10284 );
xor ( n10286 , n9775 , n10124 );
buf ( n10287 , n10286 );
xor ( n10288 , n9777 , n10123 );
buf ( n10289 , n10288 );
xor ( n10290 , n9779 , n10122 );
buf ( n10291 , n10290 );
xor ( n10292 , n9827 , n10120 );
buf ( n10293 , n10292 );
xor ( n10294 , n9952 , n10118 );
buf ( n10295 , n10294 );
xor ( n10296 , n9958 , n10116 );
buf ( n10297 , n10296 );
xor ( n10298 , n10023 , n10114 );
buf ( n10299 , n10298 );
xor ( n10300 , n10025 , n10113 );
buf ( n10301 , n10300 );
xor ( n10302 , n10060 , n10111 );
buf ( n10303 , n10302 );
xor ( n10304 , n10062 , n10110 );
buf ( n10305 , n10304 );
xor ( n10306 , n10064 , n10109 );
buf ( n10307 , n10306 );
xor ( n10308 , n10079 , n10081 );
xor ( n10309 , n10308 , n10106 );
buf ( n10310 , n10309 );
xor ( n10311 , n10083 , n10100 );
xor ( n10312 , n10311 , n10103 );
buf ( n10313 , n10312 );
xor ( n10314 , n10090 , n10094 );
xor ( n10315 , n10314 , n10097 );
buf ( n10316 , n10315 );
buf ( n10317 , n10316 );
xor ( n10318 , n10085 , n10069 );
xor ( n10319 , n10318 , n10087 );
buf ( n10320 , n10319 );
buf ( n10321 , n10320 );
not ( C0n , n0 );
and ( C0 , C0n , n0 );
endmodule
