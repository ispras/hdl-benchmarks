// IWLS benchmark module "f51m" printed on Wed May 29 16:34:04 2002
module f51m(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \44 , \45 , \46 , \47 , \48 , \49 , \50 , \51 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ;
output
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ;
wire
  \[23] ,
  \[7] ,
  \[18] ,
  \[8] ,
  \[19] ,
  \[27] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[20] ,
  \[4] ,
  \[21] ,
  \[5] ,
  \[16] ,
  \[22] ,
  \[6] ,
  \[17] ;
assign
  \[23]  = ~\[6]  | ~\8 ,
  \[7]  = (~\8  & \7 ) | ~\[27] ,
  \[18]  = (~\5  & \3 ) | (\5  & ~\3 ),
  \[8]  = ~\8 ,
  \[19]  = \7  | \6 ,
  \[27]  = ~\8  | \7 ,
  \[1]  = (\[20]  & (~\[16]  & (\4  & \3 ))) | ((~\[21]  & (~\[16]  & \4 )) | ((~\[17]  & (\[16]  & ~\2 )) | ((\[17]  & (\[16]  & \[2] )) | (~\[16]  & (~\[2]  & \2 ))))),
  \[2]  = (\[21]  & (\[17]  & ~\3 )) | ((\[20]  & (~\[17]  & \3 )) | ((~\[21]  & ~\[17] ) | (~\[20]  & \[17] ))),
  \[3]  = (~\[18]  & (\[6]  & (\7  & \3 ))) | ((\[18]  & (~\[6]  & (~\8  & ~\5 ))) | ((~\[27]  & (~\[5]  & \3 )) | ((~\[23]  & (~\[18]  & ~\[7] )) | ((~\[18]  & (~\[4]  & \4 )) | ((\[18]  & (\[4]  & ~\4 )) | (~\[19]  & \[18] )))))),
  \[20]  = ~\[3]  | \5 ,
  \[4]  = (\[23]  & (\[19]  & (~\[7]  & ~\4 ))) | ((\[23]  & (\[5]  & (\6  & ~\4 ))) | ((\[7]  & (~\[5]  & (\6  & \4 ))) | ((\[7]  & (\[5]  & (~\6  & \4 ))) | ((~\[6]  & (~\[5]  & (\7  & ~\4 ))) | ((~\[23]  & \4 ) | (~\[19]  & \4 )))))),
  \[21]  = \[3]  | ~\5 ,
  \44  = \[1] ,
  \45  = \[2] ,
  \46  = \[3] ,
  \47  = \[4] ,
  \48  = \[5] ,
  \[5]  = (\[23]  & (\[7]  & ~\5 )) | ((~\[23]  & \5 ) | (~\[7]  & \5 )),
  \[16]  = (~\3  & \1 ) | (\3  & ~\1 ),
  \49  = \[6] ,
  \50  = \[7] ,
  \51  = \[8] ,
  \[22]  = 0,
  \[6]  = (\[27]  & \6 ) | (~\[19]  & \8 ),
  \[17]  = (~\4  & \2 ) | (\4  & ~\2 );
endmodule

