// IWLS benchmark module "sbc" printed on Wed May 29 21:45:20 2002
module sbc(ACKl, BUS_Inactive, GRANTi, LastRQSTi, SBCResetPCC, PCCReq, PCCReqCode0, PCCReqCode1, PCCReqCode2, PCCReqCode3, PCCConfirm, RQSTi, SingleStep, STARTi, TM0i, TM1i, VACKl, VTM0i, VSACKi, ACKi, RESETi, SlotSpace_Id_Match, PCCSawReset, CoherencyState1i, CoherencyState2i, NuBusActive, PCCAck, PCCsync, STARTo, Tag_Match, TM1l, VTM0l, VTM1l, PCCAckCode, VACKi, physrecXXXXstate0, physrecXXXXstate1, wdcntXXXXstate1, wdcntXXXXstate2, wdcntXXXXstate3, physrecXXXXNextState0, physrecXXXXNextState1, wdcntXXXXNextState1, wdcntXXXXNextState2, wdcntXXXXNextState3, masterXXXXArb_active, masterXXXXEn_ABufo, masterXXXXEn_PDBufi, masterXXXXL_PDBufi, masterXXXXEn_VDBufi, masterXXXXEn_PDBufo, masterXXXXL_DBufo_if_TM0, masterXXXXRQSTo, masterXXXXSBC_WriteCache, nubusXXXXNuBusActive, nubusXXXXL_PABufi, resetXXXXSBCResetPCC, resetXXXXReset, slaveXXXXL_VABufi, slaveXXXXSBCReq, slaveXXXXSBCReqCode0, slaveXXXXSBCReqCode1, slaveXXXXSBCReqCode2, slaveXXXXSnoopAddrFromProc, slaveXXXXSnoopVTag_W, slaveXXXXSnoopState_W, slaveXXXXGenerateNextState, slaveXXXXSnoopVTagState_R, virmachXXXXEn_VDBufo, virmachXXXXSBCsetDirty, virmachXXXXSBCCacheRelease, virmachXXXXSBCConfigure, wdcntXXXXwd_cnt0, wdcntXXXXwd_cnt1, wdcntXXXXwd_cnt2, encodemuxXXXXMX_AD_8, nextstateXXXXCoherencyState2o, orXXXXACKo, orXXXXEn_CNTL, orXXXXRESETo, orXXXXTM0o, orXXXXTM1o, orXXXXEn_START, orXXXXSBCAck, orXXXXSBCAckCodelatch, orXXXXSBCAckCode0, orXXXXSBCAckCode1, orXXXXSBCAckCode2, orXXXXSBCAckCode3, orXXXXSTARTo, orXXXXEn_VCNTL, orXXXXVSACKo, orXXXXVACKo, orXXXXVTM0o, orXXXXVTM1o, orXXXXL_DBufo);
input
  PCCsync,
  RQSTi,
  CoherencyState1i,
  CoherencyState2i,
  PCCReqCode0,
  PCCReqCode1,
  PCCReqCode2,
  PCCReqCode3,
  SlotSpace_Id_Match,
  wdcntXXXXstate1,
  wdcntXXXXstate2,
  wdcntXXXXstate3,
  STARTi,
  STARTo,
  BUS_Inactive,
  physrecXXXXstate0,
  physrecXXXXstate1,
  PCCReq,
  VACKi,
  VACKl,
  PCCSawReset,
  GRANTi,
  VTM0i,
  VTM0l,
  VTM1l,
  Tag_Match,
  SBCResetPCC,
  PCCAckCode,
  NuBusActive,
  SingleStep,
  PCCAck,
  PCCConfirm,
  ACKi,
  ACKl,
  LastRQSTi,
  VSACKi,
  RESETi,
  TM0i,
  TM1i,
  TM1l;
output
  physrecXXXXNextState0,
  physrecXXXXNextState1,
  orXXXXACKo,
  orXXXXSTARTo,
  masterXXXXEn_VDBufi,
  orXXXXVTM1o,
  orXXXXVTM0o,
  nubusXXXXNuBusActive,
  masterXXXXArb_active,
  slaveXXXXSnoopVTagState_R,
  orXXXXTM1o,
  orXXXXTM0o,
  slaveXXXXL_VABufi,
  orXXXXL_DBufo,
  masterXXXXL_DBufo_if_TM0,
  wdcntXXXXwd_cnt0,
  wdcntXXXXwd_cnt1,
  wdcntXXXXwd_cnt2,
  orXXXXEn_START,
  slaveXXXXGenerateNextState,
  masterXXXXL_PDBufi,
  slaveXXXXSBCReqCode0,
  slaveXXXXSBCReqCode1,
  slaveXXXXSBCReqCode2,
  virmachXXXXEn_VDBufo,
  resetXXXXReset,
  nextstateXXXXCoherencyState2o,
  nubusXXXXL_PABufi,
  orXXXXRESETo,
  masterXXXXEn_ABufo,
  orXXXXVSACKo,
  virmachXXXXSBCCacheRelease,
  virmachXXXXSBCConfigure,
  masterXXXXRQSTo,
  slaveXXXXSnoopAddrFromProc,
  orXXXXVACKo,
  orXXXXSBCAck,
  slaveXXXXSnoopVTag_W,
  masterXXXXEn_PDBufi,
  masterXXXXEn_PDBufo,
  wdcntXXXXNextState1,
  wdcntXXXXNextState2,
  wdcntXXXXNextState3,
  virmachXXXXSBCsetDirty,
  resetXXXXSBCResetPCC,
  orXXXXEn_VCNTL,
  orXXXXSBCAckCodelatch,
  orXXXXSBCAckCode0,
  orXXXXSBCAckCode1,
  orXXXXSBCAckCode2,
  orXXXXSBCAckCode3,
  orXXXXEn_CNTL,
  encodemuxXXXXMX_AD_8,
  slaveXXXXSBCReq,
  slaveXXXXSnoopState_W,
  masterXXXXSBC_WriteCache;
reg
  Set_ex_wd_cnt1,
  wd_cnt_test,
  wdcntXXXXstate0,
  V_transmit_begin,
  virmachXXXXstate0,
  virmachXXXXstate1,
  V_receive_begin,
  Reset_wd_cnt,
  Gen_Reset,
  resetXXXXstate0,
  resetXXXXstate1,
  resetXXXXstate2,
  UpdateReq,
  slaveXXXXstate0,
  slaveXXXXstate1,
  slaveXXXXstate2,
  P_receive_cancel,
  UpdateDone,
  masterXXXXstate0,
  masterXXXXstate1,
  masterXXXXstate2,
  masterXXXXstate3,
  Intr_done,
  P_receive_begin,
  Incr_wd_cnt,
  nubusXXXXstate0,
  nubusXXXXstate1,
  Intr_req;
wire
  \[14688]* ,
  \{masterXXXXSBC_WriteCache} ,
  \[14922] ,
  \[10624]_inv ,
  \[14541] ,
  \[14857]* ,
  \[15300]* ,
  \[15353]* ,
  \[14911]* ,
  \[15399]* ,
  \[14970]* ,
  \[10363] ,
  \[10889]_inv ,
  \[15526]* ,
  \[14928] ,
  \[10339]* ,
  \[14547] ,
  \[14737] ,
  \[10748]_inv ,
  \[14924] ,
  \[14543] ,
  \[14733] ,
  \[2836] ,
  \{resetXXXXSBCResetPCC} ,
  \[15017]* ,
  \[14603]* ,
  \[2838] ,
  \[10933]_inv ,
  \[15418]* ,
  \LastRQSTi* ,
  \[15510]* ,
  \[1] ,
  \[10375] ,
  \[14747] ,
  \[2] ,
  \[10190] ,
  \{orXXXXEn_CNTL} ,
  \[3] ,
  \[4] ,
  \[10894]_inv ,
  \[5] ,
  \[6] ,
  \[10657]_inv ,
  \[7] ,
  \[8] ,
  \[14571]* ,
  \[15037]* ,
  \[9] ,
  \[14940] ,
  \[14942] ,
  \[14751] ,
  \[10901]_inv* ,
  \[10932]_inv ,
  \[14897]* ,
  \[15302]* ,
  \[10911]_inv* ,
  \[15355]* ,
  \[15393]* ,
  \[10921]_inv* ,
  \[10126]* ,
  masterXXXXACKo,
  \PCCReqCode2* ,
  \[15545]* ,
  \[15566]* ,
  \PCCReqCode3* ,
  \[14567] ,
  \[14757] ,
  \[10580] ,
  \[10946]_inv ,
  \[15109] ,
  \[14944] ,
  \[10559]_inv* ,
  \{orXXXXRESETo} ,
  \{orXXXXIncr_wd_cnt} ,
  \PCCReqCode0* ,
  \[14946] ,
  \PCCReqCode1* ,
  \[15105] ,
  \[14760] ,
  \[14950] ,
  \[15300] ,
  \[14952] ,
  \[14781]* ,
  \[14571] ,
  \[15302] ,
  \[15247]* ,
  \[14879]* ,
  \NuBusActive* ,
  \[15396]* ,
  \[15512]* ,
  \[10586] ,
  \[15550]* ,
  \[14387] ,
  \[14767] ,
  \[15702]* ,
  \[14769] ,
  \[14959] ,
  \[14764] ,
  \[10591] ,
  \Reset_wd_cnt* ,
  \[15304] ,
  \[14575] ,
  \[14955] ,
  \[10889]_inv* ,
  \[15039]* ,
  \[10899]_inv* ,
  \[15120] ,
  \[15310] ,
  \[14771] ,
  \[15288]* ,
  \Intr_done* ,
  \[10651]_inv* ,
  \[10938]_inv ,
  \[10819]_inv* ,
  \[15508] ,
  \[15668]* ,
  \[15129] ,
  \[15319] ,
  \[14963] ,
  \[15123] ,
  \[14966] ,
  \[14517]* ,
  \[14585] ,
  \[15506] ,
  \[14970] ,
  \[15097]* ,
  \[14666]* ,
  \[15510] ,
  \[14972] ,
  \[14781] ,
  \[15512] ,
  \[15702] ,
  \[15362]* ,
  \[15439]* ,
  \[10923]_inv ,
  \[15137] ,
  \[15327] ,
  \[15707] ,
  \{orXXXXVSACKo} ,
  \[10749]_inv* ,
  \[15329] ,
  \[14593] ,
  \[10823]_inv ,
  \[15133] ,
  \[14496]* ,
  \[14976] ,
  \[14595] ,
  \[14537]* ,
  \[15135] ,
  \[14980] ,
  \[15079]* ,
  \[15710] ,
  \[15192]* ,
  \[14982] ,
  \[15206]* ,
  \[15223]* ,
  \[14802]* ,
  \[15712] ,
  \P_receive_begin* ,
  \[15141] ,
  \[15521] ,
  \[14917]* ,
  \[15382]* ,
  \[530]* ,
  \ACKi* ,
  \[10912]_inv* ,
  \[15572]* ,
  \[15148] ,
  \[14797] ,
  \[15338] ,
  \[15624]* ,
  \[14987] ,
  \[10932]_inv* ,
  \ACKl* ,
  \[14984] ,
  \[10586]* ,
  \[15529] ,
  \[10822]_inv ,
  \[15334] ,
  \[14421]* ,
  \[10936]_inv ,
  \[14480]* ,
  \[15143] ,
  \{virmachXXXXNextState1} ,
  \[15336] ,
  \[15526] ,
  \[14990] ,
  \[15074]* ,
  \[14709]* ,
  \[14747]* ,
  \[14860]* ,
  \{virmachXXXXNextState0} ,
  \[10821]_inv* ,
  \[15416]* ,
  \[14997] ,
  \[15538] ,
  \[15159] ,
  \[15349] ,
  \[14387]* ,
  \[15344] ,
  \[14993] ,
  \[10907]_inv* ,
  \[14539]* ,
  \VSACKi* ,
  \[15536] ,
  \[15035]* ,
  \[15056]* ,
  \[10937]_inv* ,
  \[14767]* ,
  \[10945]_inv ,
  \[14821]* ,
  \[15284]* ,
  \{orXXXXSBCAck} ,
  \[15541] ,
  \SlotSpace_Id_Match* ,
  \[10721]_inv* ,
  \{orXXXXReset_wd_cnt_x} ,
  \[15499]* ,
  \[10845]_inv ,
  \[15591]* ,
  \[15643]* ,
  \[15357] ,
  \[15169] ,
  \[10928]_inv ,
  \[10662]_inv* ,
  \resetXXXXstate2* ,
  \[15353] ,
  \[10682]_inv* ,
  \resetXXXXstate0* ,
  \[15355] ,
  \[15545] ,
  \resetXXXXstate1* ,
  \[15550] ,
  \[15230]* ,
  \[15362] ,
  \[15266]* ,
  \[14862]* ,
  \[15456]* ,
  \[10612]_inv* ,
  \[15558] ,
  \[15646]* ,
  \[15663]* ,
  \[15367] ,
  \[10497]* ,
  \[15369] ,
  \RESETi* ,
  \[15553] ,
  \[14533]* ,
  \[15176] ,
  \[10813]_inv ,
  \{orXXXXSBCAckCodelatch} ,
  \[15560] ,
  \[10937]_inv ,
  \[15137]* ,
  \[14723]* ,
  \[14769]* ,
  \[15182] ,
  \[10657]_inv* ,
  \PCCReq* ,
  \[15327]* ,
  \[14959]* ,
  \[13753]_inv* ,
  \[14997]* ,
  \[15538]* ,
  \[15377] ,
  \{slaveXXXXNextState1} ,
  \[15707]* ,
  \[10912]_inv ,
  \{slaveXXXXNextState2} ,
  \[15379] ,
  \[10483]_inv ,
  \[15569] ,
  \[15184] ,
  \{slaveXXXXNextState0} ,
  \[10612]_inv ,
  \[10882]_inv* ,
  \[15566] ,
  \[15021]* ,
  \[15190] ,
  \[14726]* ,
  \[14764]* ,
  \[15211]* ,
  \[15192] ,
  \[15232]* ,
  \[15382] ,
  \[15572] ,
  \[15558]* ,
  \[10822]_inv* ,
  \[15198] ,
  \[15665]* ,
  \[15686]* ,
  \[15577] ,
  \[14409] ,
  I105,
  \[10422] ,
  I108,
  I109,
  \[15389] ,
  \[10591]* ,
  \[15574] ,
  I126,
  I128,
  I130,
  I131,
  I139,
  \[10507]_inv* ,
  I140,
  \[15041]* ,
  \[10921]_inv ,
  I163,
  I164,
  I167,
  I172,
  \[10908]_inv* ,
  I173,
  I177,
  I179,
  \[14411] ,
  \[10918]_inv* ,
  \[15252]* ,
  \[14808]* ,
  \[15582] ,
  I187,
  I188,
  \[15290]* ,
  I192,
  \[10928]_inv* ,
  \[15391] ,
  I193,
  \[15304]* ,
  \[15329]* ,
  I199,
  \[14900]* ,
  \[15367]* ,
  \[14915]* ,
  \[10821]_inv ,
  \[10938]_inv* ,
  \[10682]_inv ,
  \[10877]_inv* ,
  \[10935]_inv ,
  \[10721]_inv ,
  \[15442]* ,
  \[15495]* ,
  \[10882]_inv ,
  \[10897]_inv* ,
  \[2838]* ,
  \[14417] ,
  \[15670]* ,
  \[15587] ,
  \[14419] ,
  I201,
  I207,
  I208,
  \[10696]_inv ,
  I211,
  \[15399] ,
  I214,
  I215,
  I219,
  \[14603] ,
  I220,
  I222,
  I223,
  \[14448]* ,
  I229,
  I231,
  I232,
  \[15393] ,
  I235,
  I236,
  \[15396] ,
  \[14593]* ,
  \[10918]_inv ,
  \[10817]_inv* ,
  \[10559]_inv ,
  \[14617]* ,
  \[15159]* ,
  \[14730]* ,
  \[14802] ,
  I273,
  I276,
  I279,
  \[14421] ,
  I280,
  I282,
  I284,
  I285,
  I287,
  I288,
  I292,
  I295,
  \[15591] ,
  I296,
  I299,
  \[15349]* ,
  \[14808] ,
  \[15577]* ,
  \[14617] ,
  \[14619] ,
  I300,
  I304,
  I305,
  \[10632] ,
  \[14804] ,
  \[10061] ,
  \[15599] ,
  \[14409]* ,
  I322,
  I323,
  I340,
  I341,
  \[14575]* ,
  I348,
  I354,
  \[15081]* ,
  I357,
  I361,
  I363,
  I364,
  I366,
  \[10750]_inv ,
  I368,
  \[15133]* ,
  I369,
  I373,
  I374,
  I377,
  \[15292]* ,
  \PCCAck* ,
  I398,
  I399,
  \[15344]* ,
  \[14902]* ,
  \[10703]_inv ,
  \[15369]* ,
  \[14940]* ,
  \[14955]* ,
  \[14993]* ,
  \TM0i* ,
  \{masterXXXXUpdateReq} ,
  \[10658]_inv* ,
  \[10483]_inv* ,
  \[14627] ,
  \[10640] ,
  \[10422]* ,
  \[10688]_inv ,
  \[10888]_inv ,
  I88,
  I91,
  \[14488]* ,
  \[14816] ,
  \[2536] ,
  \[14521]* ,
  \[14595]* ,
  \[2537] ,
  I450,
  I451,
  I453,
  \[14619]* ,
  \[10930]_inv* ,
  I465,
  \[14711]* ,
  \[10940]_inv* ,
  I475,
  I476,
  \[14441] ,
  \[14821] ,
  \[13378]_inv ,
  \physrecXXXXstate1* ,
  \[14922]* ,
  \[15389]* ,
  \physrecXXXXstate0* ,
  \TM1i* ,
  \[15481]* ,
  \{masterXXXXNextState1} ,
  \[14448] ,
  \{masterXXXXNextState2} ,
  \TM1l* ,
  \[10816]_inv ,
  \{masterXXXXNextState3} ,
  \[15692]* ,
  \PCCSawReset* ,
  \[10573]_inv ,
  \[14634] ,
  I515,
  I516,
  \[14443] ,
  \[14823] ,
  \{masterXXXXNextState0} ,
  I536,
  I537,
  \BUS_Inactive* ,
  I543,
  \[14450] ,
  \[14640] ,
  \[14830] ,
  \[14698]* ,
  \{orXXXXEn_START} ,
  \[15120]* ,
  \[15135]* ,
  \[10897]_inv ,
  \[14804]* ,
  \[10911]_inv ,
  \[10089] ,
  \[15310]* ,
  I599,
  \[14942]* ,
  \[14980]* ,
  \[10653] ,
  \[10511]_inv ,
  \[15536]* ,
  \[15553]* ,
  \[14838] ,
  \[15574]* ,
  \[15599]* ,
  \[10878]_inv* ,
  \{resetXXXXNextState1} ,
  \[10888]_inv* ,
  \{resetXXXXNextState2} ,
  \[10686]_inv ,
  \[14659]* ,
  \[10886]_inv ,
  \[15176]* ,
  \[14751]* ,
  \[10908]_inv ,
  \nubusXXXXstate0* ,
  \[10749]_inv ,
  \[15407]* ,
  \nubusXXXXstate1* ,
  \[14467] ,
  \{nubusXXXXL_PABufi} ,
  \[15710]* ,
  \[14469] ,
  \[14659] ,
  \{orXXXXACKo} ,
  \[14654] ,
  \{orXXXXVTM0o} ,
  \[14443]* ,
  \[15003] ,
  \[14846] ,
  \[10940]_inv ,
  \[15068]* ,
  \[10936]_inv* ,
  \[10946]_inv* ,
  \wd_cnt_test* ,
  \[14852] ,
  \[14771]* ,
  \{slaveXXXXL_VABufi} ,
  \[14661] ,
  \[14823]* ,
  \[2537]* ,
  \[15011] ,
  \[14982]* ,
  \[15427]* ,
  \[10748]_inv* ,
  \[10945]_inv* ,
  \[10296] ,
  \[14478] ,
  \[14668] ,
  \[14857] ,
  \[10854]_inv ,
  \[15017] ,
  \VACKi* ,
  \[10492] ,
  \[10533]* ,
  \[10817]_inv ,
  \[14484]* ,
  \[14666] ,
  \[14508]* ,
  \[15206] ,
  \[14480] ,
  \[10878]_inv ,
  \[14860] ,
  \Intr_req* ,
  \[14862] ,
  \[10497] ,
  \RQSTi* ,
  \[15219]* ,
  \[15021] ,
  \[15211] ,
  \[10935]_inv* ,
  \[10493] ,
  \[10890]_inv* ,
  \[14488] ,
  \[13378]_inv* ,
  \[15637]* ,
  \[15658]* ,
  \[15407] ,
  \[15712]* ,
  \[10506]_inv ,
  \[14484] ,
  \[14674] ,
  \[15219] ,
  \{wdcntXXXXwd_cnt_test} ,
  \[14676] ,
  \[15403] ,
  \[15026] ,
  \[10863]_inv ,
  \[15003]* ,
  \[14490] ,
  \[15215] ,
  \[15405] ,
  \[15030] ,
  \[15410] ,
  \[15141]* ,
  \[14492] ,
  \[10750]_inv* ,
  \[14681] ,
  \[14871] ,
  \[15412] ,
  \[1048]* ,
  \[15298]* ,
  \[14846]* ,
  \slaveXXXXstate2* ,
  \slaveXXXXstate1* ,
  \[10686]_inv* ,
  \slaveXXXXstate0* ,
  \[10696]_inv* ,
  \[10901]_inv ,
  \[15521]* ,
  \[14688] ,
  \[15228] ,
  \[15418] ,
  \[15037] ,
  \[14879] ,
  \[14494] ,
  \[15039] ,
  \wdcntXXXXstate3* ,
  \[10662]_inv ,
  \wdcntXXXXstate2* ,
  \[15604] ,
  \[14496] ,
  \[15223] ,
  \[1048] ,
  \[15416] ,
  \[10] ,
  \[15035] ,
  \PCCAckCode* ,
  \[14640]* ,
  \[11] ,
  \[14676]* ,
  \[15230] ,
  \[14693]* ,
  \[12] ,
  \[14717]* ,
  \wdcntXXXXstate1* ,
  \[15182]* ,
  \[13] ,
  \[10939]_inv ,
  \[15232] ,
  \[14830]* ,
  \[14] ,
  \[13753]_inv ,
  \[15041] ,
  \[15] ,
  \[16] ,
  \[15403]* ,
  \[17] ,
  \[15487]* ,
  \[18] ,
  \[15541]* ,
  \[14698] ,
  \[15614]* ,
  \[15427] ,
  \[10685]_inv* ,
  \[14693] ,
  \[14883] ,
  \[14411]* ,
  \[15614] ,
  \[15046] ,
  \[14547]* ,
  \[15026]* ,
  \[15235] ,
  \[15425] ,
  \[15064]* ,
  \[15089]* ,
  \[15050] ,
  \[15240] ,
  \[10930]_inv ,
  \[15052] ,
  \[10923]_inv* ,
  \[10866]_inv* ,
  \[10933]_inv* ,
  \[10943]_inv* ,
  \[10886]_inv* ,
  \[15444]* ,
  \[10685]_inv ,
  \[15582]* ,
  \[10944]_inv ,
  \[100] ,
  \[14897] ,
  \[101] ,
  \[15697]* ,
  \[15247] ,
  \[102] ,
  \{orXXXXSBCAckCode1} ,
  \[103] ,
  \{orXXXXSBCAckCode2} ,
  \[10907]_inv ,
  \[15439] ,
  \[10544]_inv ,
  \[104] ,
  \{orXXXXSBCAckCode3} ,
  \[15054] ,
  \[15624] ,
  \[105] ,
  \[14490]* ,
  \{orXXXXVACKo} ,
  \[10816]_inv* ,
  \[106] ,
  \[15056] ,
  \[107] ,
  \[10507]_inv ,
  \[15046]* ,
  \[108] ,
  \[109] ,
  \{orXXXXSBCAckCode0} ,
  \[14757]* ,
  \{slaveXXXXSBCReqCode0} ,
  \[15215]* ,
  \PCCsync* ,
  \[15252] ,
  \[15442] ,
  \[14909]* ,
  \[15391]* ,
  \[15405]* ,
  \[10845]_inv* ,
  \[15489]* ,
  \[110] ,
  \[15068] ,
  \[111] ,
  \{slaveXXXXSBCReqCode1} ,
  \[15637] ,
  \{orXXXXEn_VCNTL} ,
  \[10580]* ,
  \[15064] ,
  \[15444] ,
  \[14503]* ,
  \[15066] ,
  \masterXXXXstate3* ,
  \[15446] ,
  \[15030]* ,
  \masterXXXXstate2* ,
  \[15235]* ,
  \[15452] ,
  \[15294]* ,
  \[14852]* ,
  \{orXXXXL_DBufo} ,
  \masterXXXXstate1* ,
  \[15410]* ,
  \[15425]* ,
  \masterXXXXstate0* ,
  \[15446]* ,
  \{physrecXXXXNextState1} ,
  \[15508]* ,
  \[10877]_inv ,
  \[15653]* ,
  \[15674]* ,
  \[15079] ,
  \[15074] ,
  \[14492]* ,
  \[15643] ,
  \[15266] ,
  \[15456] ,
  \[15646] ,
  \[15050]* ,
  \[14661]* ,
  \[15148]* ,
  \[10307] ,
  \[14797]* ,
  \[15081] ,
  \[10089]* ,
  \[15338]* ,
  \[10643]_inv* ,
  \[14924]* ,
  \[14987]* ,
  \[10929]_inv ,
  \[10573]_inv* ,
  \[10866]_inv ,
  \PCCConfirm* ,
  \[15658] ,
  \[15089] ,
  \{nubusXXXXNuBusActive} ,
  \[15653] ,
  \[14505]* ,
  \[14543]* ,
  \[15276] ,
  \[15085] ,
  \[15465] ,
  \[15655] ,
  \[15085]* ,
  \{virmachXXXXSBCConfigure} ,
  \[15280] ,
  \[15109]* ,
  \[14733]* ,
  \[15296]* ,
  \[15091] ,
  \[14871]* ,
  \[15471] ,
  \[15661] ,
  \[14944]* ,
  \[15412]* ,
  \[10924]_inv* ,
  \[15465]* ,
  \[10863]_inv* ,
  \[10126] ,
  \[10934]_inv* ,
  \[10944]_inv* ,
  \Tag_Match* ,
  \[15288] ,
  \[15668] ,
  \[15097] ,
  \[10458]_inv ,
  \SingleStep* ,
  \[10934]_inv ,
  \VTM0l* ,
  \[15284] ,
  \[15663] ,
  \[14525]* ,
  \[15665] ,
  \[15290] ,
  \[15129]* ,
  \[15670] ,
  \[10327] ,
  \[10823]_inv* ,
  \[15292] ,
  \[10899]_inv ,
  \STARTi* ,
  \[15481] ,
  \[15319]* ,
  \[10658]_inv ,
  \[15357]* ,
  \[14508] ,
  \{nubusXXXXNextState0} ,
  \[530] ,
  \[15298] ,
  \STARTo* ,
  \[15487] ,
  \{nubusXXXXNextState1} ,
  \[15489] ,
  \VTM1l* ,
  \[14503] ,
  \[15294] ,
  \[15674] ,
  \[10653]* ,
  \[14505] ,
  \[15296] ,
  \[15676] ,
  \[10703]_inv* ,
  \[10943]_inv ,
  \[15680] ,
  \V_transmit_begin* ,
  \[10718] ,
  \[14512] ,
  \[10890]_inv ,
  \[15492] ,
  \[84] ,
  \[10643]_inv ,
  \[10339] ,
  \[85] ,
  \[15377]* ,
  \GRANTi* ,
  \[14946]* ,
  \[14963]* ,
  \[86] ,
  \[14984]* ,
  \[15452]* ,
  \[87] ,
  \{orXXXXTM1o} ,
  \[88] ,
  \[15529]* ,
  \{slaveXXXXSBCReq} ,
  \[10335] ,
  \[10525] ,
  \[89] ,
  masterXXXXVSACKo,
  \[14517] ,
  \[15680]* ,
  \[14709] ,
  \[15499] ,
  \[10718]* ,
  \[14512]* ,
  \[15686] ,
  \[90] ,
  \[14900] ,
  \[15495] ,
  \[14627]* ,
  \[91] ,
  \[15123]* ,
  \[92] ,
  \[14902] ,
  \[93] ,
  \[14521] ,
  \[14711] ,
  \[15692] ,
  \[14838]* ,
  \[94] ,
  \P_receive_cancel* ,
  \[95] ,
  \[14966]* ,
  \[96] ,
  \[10624]_inv* ,
  \[10533] ,
  \[97] ,
  \[98] ,
  \[10296]* ,
  \[15587]* ,
  \[99] ,
  \[14717] ,
  \SBCResetPCC* ,
  \[15697] ,
  \[14529] ,
  \[14909] ,
  \[14523] ,
  \[14419]* ,
  \[10640]* ,
  \[14478]* ,
  \masterXXXXVSACKo* ,
  \[14525] ,
  \[10819]_inv ,
  \[14585]* ,
  \{slaveXXXXSnoopState_W} ,
  \[15091]* ,
  \[14668]* ,
  \CoherencyState2i* ,
  \[15105]* ,
  \[15143]* ,
  \[14760]* ,
  \[14531] ,
  \[14911] ,
  \[15379]* ,
  \[14950]* ,
  \[15471]* ,
  \[15492]* ,
  \[15506]* ,
  \[15569]* ,
  \[10544]_inv* ,
  \[10651]_inv ,
  \[14537] ,
  \[14917] ,
  \[10854]_inv* ,
  \[15661]* ,
  \[10929]_inv* ,
  \[10939]_inv* ,
  \[14539] ,
  \[14533] ,
  \[14723] ,
  \[10894]_inv* ,
  \[14726] ,
  \virmachXXXXstate0* ,
  \[14535] ,
  \[14915] ,
  \[10924]_inv ,
  \virmachXXXXstate1* ,
  \[14730] ;
assign
  \[14688]*  = ~\[14688] ,
  \{masterXXXXSBC_WriteCache}  = \[10511]_inv  | \[14902] ,
  \[14922]  = \RQSTi*  & \[15074]* ,
  \[10624]_inv  = \[10750]_inv  | \TM1l* ,
  \[14541]  = \[10296]*  & SBCResetPCC,
  \[14857]*  = ~\[14857] ,
  \[15300]*  = ~\[15300] ,
  \[15353]*  = ~\[15353] ,
  \[14911]*  = ~\[14911] ,
  \[15399]*  = ~\[15399] ,
  \[14970]*  = ~\[14970] ,
  physrecXXXXNextState0 = \[14928] ,
  physrecXXXXNextState1 = \{physrecXXXXNextState1} ,
  \[10363]  = I398 | I399,
  \[10889]_inv  = SBCResetPCC | \masterXXXXstate0* ,
  \[15526]*  = ~\[15526] ,
  \[14928]  = \[10]  & \[10945]_inv* ,
  \[10339]*  = ~\[10339] ,
  \[14547]  = \[14897]*  & (\[14917]*  & (\[1048]*  & \[14982]* )),
  \[14737]  = \SBCResetPCC*  & (\[15026]*  & VTM0i),
  \[10748]_inv  = \[10813]_inv  | \PCCReqCode3* ,
  \[14924]  = \ACKl*  & \[15079]* ,
  \[14543]  = \slaveXXXXstate1*  & (\[10375]  & \[15553] ),
  \[14733]  = \[10640]*  & (\[10089]*  & (\[15382]*  & \[15362]* )),
  \[2836]  = \[14816]  | (\[15604]  | \[15052] ),
  \{resetXXXXSBCResetPCC}  = resetXXXXstate0 | (resetXXXXstate2 | (RESETi | \[15560] )),
  \[15017]*  = ~\[15017] ,
  \[14603]*  = ~\[14603] ,
  \[2838]  = \[1048]  | I201,
  orXXXXACKo = \{orXXXXACKo} ,
  \[10933]_inv  = STARTi | \NuBusActive* ,
  \[15418]*  = ~\[15418] ,
  \LastRQSTi*  = ~LastRQSTi,
  \[15510]*  = ~\[15510] ,
  \[1]  = \[10339]*  | \[14537]* ,
  \[10375]  = I231 | I232,
  \[14747]  = \[10497]*  & \[15182]* ,
  \[2]  = \[15465]*  | \[14911]* ,
  \[10190]  = I295 | I296,
  \{orXXXXEn_CNTL}  = I172 | I173,
  \[3]  = \[15396]*  | \[14823]* ,
  \[4]  = \[15074]*  | \[10924]_inv* ,
  \[10894]_inv  = PCCReqCode3 | \PCCReq* ,
  \[5]  = \[10819]_inv*  | \[15655] ,
  \[6]  = \[15109]*  | \[15247]* ,
  \[10657]_inv  = \[10813]_inv  | \masterXXXXstate3* ,
  \[7]  = \[15425]*  | NuBusActive,
  \[8]  = \[15382]*  | \[15017]* ,
  \[14571]*  = ~\[14571] ,
  \[15037]*  = ~\[15037] ,
  \[9]  = \masterXXXXstate2*  | \[15037]* ,
  \[14940]  = \[10816]_inv*  & (\[15344]  & PCCConfirm),
  \[14942]  = \[15097]*  & \[15577]* ,
  \[14751]  = \[10932]_inv*  & (\[15035]*  & \[15143] ),
  \[10901]_inv*  = ~\[10901]_inv ,
  \[10932]_inv  = \masterXXXXstate1*  | \masterXXXXstate2* ,
  \[14897]*  = ~\[14897] ,
  \[15302]*  = ~\[15302] ,
  \[10911]_inv*  = ~\[10911]_inv ,
  \[15355]*  = ~\[15355] ,
  \[15393]*  = ~\[15393] ,
  \[10921]_inv*  = ~\[10921]_inv ,
  \[10126]*  = ~\[10126] ,
  masterXXXXACKo = \[10506]_inv  | \[15041]* ,
  \PCCReqCode2*  = ~PCCReqCode2,
  \[15545]*  = ~\[15545] ,
  \[15566]*  = ~\[15566] ,
  \PCCReqCode3*  = ~PCCReqCode3,
  \[14567]  = \[10937]_inv*  & \[14619]* ,
  \[14757]  = \[10878]_inv*  & \[14909]* ,
  orXXXXSTARTo = \[14567] ,
  \[10580]  = \[10573]_inv*  | I282,
  \[10946]_inv  = SBCResetPCC | \virmachXXXXstate0* ,
  \[15109]  = \[10901]_inv*  & \[15399]* ,
  \[14944]  = \ACKl*  & \[15123]* ,
  \[10559]_inv*  = ~\[10559]_inv ,
  \{orXXXXRESETo}  = \[14972]  | (\[15276]  | \[14627]* ),
  \{orXXXXIncr_wd_cnt}  = \[15066]  | (\[15159]  | (\[14737]  | \[15054] )),
  \PCCReqCode0*  = ~PCCReqCode0,
  \[14946]  = \[15405]*  & (\[15577]*  & \[15471]* ),
  \PCCReqCode1*  = ~PCCReqCode1,
  \[15105]  = \[15338]*  & \[10817]_inv ,
  \[14760]  = \[10822]_inv*  & (\[15068]*  & masterXXXXstate2),
  \[14950]  = \[11]  & \[10908]_inv ,
  \[15300]  = \[15599]*  & \[15587]* ,
  \[14952]  = \[15192]*  & \PCCAck* ,
  \[14781]*  = ~\[14781] ,
  \[14571]  = \[10718]*  & \[15489]* ,
  masterXXXXEn_VDBufi = \[14902]* ,
  \[15302]  = \[15582]  & P_receive_begin,
  \[15247]*  = ~\[15247] ,
  \[14879]*  = ~\[14879] ,
  \NuBusActive*  = ~NuBusActive,
  \[15396]*  = ~\[15396] ,
  \[15512]*  = ~\[15512] ,
  \[10586]  = I304 | I305,
  \[15550]*  = ~\[15550] ,
  \[14387]  = \[14764]*  & (\[15159]*  & (\masterXXXXVSACKo*  & \[15192]* )),
  \[14767]  = \[5]  & \[15120]* ,
  \[15702]*  = ~\[15702] ,
  \[14769]  = \[6]  & \[10889]_inv ,
  \[14959]  = \[15223]  & STARTi,
  \[14764]  = \[10877]_inv*  & \[14915]* ,
  orXXXXVTM1o = \[14417] ,
  \[10591]  = I163 | I164,
  \Reset_wd_cnt*  = ~Reset_wd_cnt,
  \[15304]  = \slaveXXXXstate2*  & (\PCCAck*  & \[15553] ),
  orXXXXVTM0o = \{orXXXXVTM0o} ,
  \[14575]  = \[10882]_inv*  & (\masterXXXXstate1*  & \[14821]* ),
  \[14955]  = \[15393]*  & (\[15566]*  & \[15290]* ),
  \[10889]_inv*  = ~\[10889]_inv ,
  \[15039]*  = ~\[15039] ,
  \[10899]_inv*  = ~\[10899]_inv ,
  \[15120]  = \[15357]*  & \[15529]* ,
  \[15310]  = \PCCsync*  & \[15680]* ,
  \[14771]  = \[14955]*  & ACKl,
  \[15288]*  = ~\[15288] ,
  nubusXXXXNuBusActive = \{nubusXXXXNuBusActive} ,
  \Intr_done*  = ~Intr_done,
  \[10651]_inv*  = ~\[10651]_inv ,
  \[10938]_inv  = RESETi | \nubusXXXXstate0* ,
  \[10819]_inv*  = ~\[10819]_inv ,
  \[15508]  = \SBCResetPCC*  & (\wdcntXXXXstate1*  & (Reset_wd_cnt & Set_ex_wd_cnt1)),
  \[15668]*  = ~\[15668] ,
  masterXXXXArb_active = \[14529] ,
  \[15129]  = \resetXXXXstate2*  & \[15403]* ,
  \[15319]  = \STARTi*  & \[15566] ,
  slaveXXXXSnoopVTagState_R = \[14764] ,
  \[14963]  = \[15089]*  & Tag_Match,
  \[15123]  = \masterXXXXstate1*  & \[15338]* ,
  \[14966]  = \[12]  & \[10821]_inv* ,
  \[14517]*  = ~\[14517] ,
  \[14585]  = \[10882]_inv*  & (\masterXXXXstate2*  & \[14838]* ),
  \[15506]  = \ACKi*  & (\Intr_req*  & NuBusActive),
  \[14970]  = \[10899]_inv*  & (\[10894]_inv*  & \[15369]* ),
  \[15097]*  = ~\[15097] ,
  \[14666]*  = ~\[14666] ,
  \[15510]  = CoherencyState1i & (CoherencyState2i & TM1l),
  orXXXXTM1o = \{orXXXXTM1o} ,
  \[14972]  = \[10938]_inv*  & (\[15391]*  & STARTi),
  orXXXXTM0o = \[14862]* ,
  \[14781]  = \[14940]*  & GRANTi,
  \[15512]  = PCCReqCode1 & PCCReqCode2,
  \[15702]  = \SingleStep*  & \VSACKi* ,
  \[15362]*  = ~\[15362] ,
  \[15439]*  = ~\[15439] ,
  slaveXXXXL_VABufi = \{slaveXXXXL_VABufi} ,
  \[10923]_inv  = nubusXXXXstate0 | \SlotSpace_Id_Match* ,
  \[15137]  = \RQSTi*  & \[10821]_inv* ,
  \[15327]  = \[17]  & TM1l,
  \[15707]  = \ACKi*  & \slaveXXXXstate0* ,
  \{orXXXXVSACKo}  = \[14387]*  | \[14698]* ,
  \[10749]_inv*  = ~\[10749]_inv ,
  \[15329]  = \PCCReqCode2*  & \[15569] ,
  \[14593]  = \[14993]*  & (\[15223]*  & \[14693]* ),
  \[10823]_inv  = masterXXXXstate3 | \[10932]_inv ,
  \[15133]  = \[10854]_inv*  & \[15487]* ,
  \[14496]*  = ~\[14496] ,
  \[14976]  = \resetXXXXstate2*  & (\[15407]  & RESETi),
  \[14595]  = \[14959]*  & (\[15235]*  & \[14693]* ),
  \[14537]*  = ~\[14537] ,
  \[15135]  = \[15427]*  & \[15665]* ,
  \[14980]  = \[15135]*  & wd_cnt_test,
  \[15079]*  = ~\[15079] ,
  orXXXXL_DBufo = \{orXXXXL_DBufo} ,
  \[15710]  = wdcntXXXXstate3 & wdcntXXXXstate0,
  \[15192]*  = ~\[15192] ,
  \[14982]  = \[10943]_inv*  & (\VSACKi*  & \[15292]* ),
  \[15206]*  = ~\[15206] ,
  \[15223]*  = ~\[15223] ,
  masterXXXXL_DBufo_if_TM0 = \[15247] ,
  \[14802]*  = ~\[14802] ,
  \[15712]  = \TM1l*  & \VTM1l* ,
  \P_receive_begin*  = ~P_receive_begin,
  \[15141]  = \[15446]*  & \[15670]* ,
  \[15521]  = VACKl & masterXXXXstate1,
  \[14917]*  = ~\[14917] ,
  \[15382]*  = ~\[15382] ,
  \[530]*  = ~\[530] ,
  \ACKi*  = ~ACKi,
  \[10912]_inv*  = ~\[10912]_inv ,
  \[15572]*  = ~\[15572] ,
  \[15148]  = \[16]  & \[10901]_inv ,
  \[14797]  = \[15003]*  & \[15133]* ,
  \[15338]  = \[15599]*  & \masterXXXXstate2* ,
  \[15624]*  = ~\[15624] ,
  \[14987]  = \SBCResetPCC*  & \[15211]* ,
  \[10932]_inv*  = ~\[10932]_inv ,
  \ACKl*  = ~ACKl,
  \[14984]  = \[13]  & \[15085]* ,
  \[10586]*  = ~\[10586] ,
  \[15529]  = \CoherencyState2i*  & CoherencyState1i,
  \[10822]_inv  = \[15574]*  | \GRANTi* ,
  \[15334]  = \VTM1l*  & \[15655] ,
  \[14421]*  = ~\[14421] ,
  \[10936]_inv  = RESETi | slaveXXXXstate0,
  \[14480]*  = ~\[14480] ,
  \[15143]  = \[10816]_inv*  & GRANTi,
  \{virmachXXXXNextState1}  = \[14987]  | I273,
  \[15336]  = \[10935]_inv*  & \[15582]* ,
  \[15526]  = STARTo & VTM0l,
  \[14990]  = \[10907]_inv*  & (\STARTi*  & \[15389]* ),
  \[15074]*  = ~\[15074] ,
  \[14709]*  = ~\[14709] ,
  \[14747]*  = ~\[14747] ,
  \[14860]*  = ~\[14860] ,
  \{virmachXXXXNextState0}  = \[14808]*  | I199,
  \[10821]_inv*  = ~\[10821]_inv ,
  \[15416]*  = ~\[15416] ,
  wdcntXXXXwd_cnt0 = \[14984]* ,
  wdcntXXXXwd_cnt1 = \[14797]* ,
  wdcntXXXXwd_cnt2 = \[14857]* ,
  \[14997]  = \[15206]*  & \slaveXXXXstate2* ,
  \[15538]  = \TM0i*  & TM1i,
  \[15159]  = \wd_cnt_test*  & \[15452] ,
  \[15349]  = \physrecXXXXstate0*  & \[15665]* ,
  \[14387]*  = ~\[14387] ,
  \[15344]  = \[10894]_inv*  & \[15512]* ,
  \[14993]  = \[10823]_inv*  & \[15143]* ,
  \[10907]_inv*  = ~\[10907]_inv ,
  \[14539]*  = ~\[14539] ,
  \VSACKi*  = ~VSACKi,
  \[15536]  = VSACKi & slaveXXXXstate0,
  orXXXXEn_START = \{orXXXXEn_START} ,
  \[15035]*  = ~\[15035] ,
  \[15056]*  = ~\[15056] ,
  slaveXXXXGenerateNextState = \[14676]* ,
  \[10937]_inv*  = ~\[10937]_inv ,
  \[14767]*  = ~\[14767] ,
  \[10945]_inv  = SBCResetPCC | ACKi,
  masterXXXXL_PDBufi = \[10703]_inv* ,
  \[14821]*  = ~\[14821] ,
  \[15284]*  = ~\[15284] ,
  \{orXXXXSBCAck}  = \[2836]  | (masterXXXXACKo | (\[14494]  | \[14911] )),
  \[15541]  = \Intr_done*  & nubusXXXXstate1,
  \SlotSpace_Id_Match*  = ~SlotSpace_Id_Match,
  \[10721]_inv*  = ~\[10721]_inv ,
  \{orXXXXReset_wd_cnt_x}  = \[14496]  | (\[14512]  | (\[15011]  | \[15017] )),
  \[15499]*  = ~\[15499] ,
  \[10845]_inv  = SBCResetPCC | \P_receive_begin* ,
  \[15591]*  = ~\[15591] ,
  \[15643]*  = ~\[15643] ,
  \[15357]  = \[15529]*  & \[15712] ,
  \[15169]  = \[15452]  & wd_cnt_test,
  \[10928]_inv  = \masterXXXXstate2*  | \masterXXXXstate3* ,
  \[10662]_inv*  = ~\[10662]_inv ,
  \resetXXXXstate2*  = ~resetXXXXstate2,
  \[15353]  = \[15712]*  & CoherencyState1i,
  \[10682]_inv*  = ~\[10682]_inv ,
  \resetXXXXstate0*  = ~resetXXXXstate0,
  \[15355]  = \[10894]_inv*  & \[15661]* ,
  \[15545]  = masterXXXXstate1 & masterXXXXstate3,
  \resetXXXXstate1*  = ~resetXXXXstate1,
  \[15550]  = \PCCReqCode2*  & PCCReqCode1,
  slaveXXXXSBCReqCode0 = \{slaveXXXXSBCReqCode0} ,
  slaveXXXXSBCReqCode1 = \{slaveXXXXSBCReqCode1} ,
  slaveXXXXSBCReqCode2 = \[14654] ,
  \[15230]*  = ~\[15230] ,
  \[15362]  = \[10901]_inv*  & \[15558]* ,
  \[15266]*  = ~\[15266] ,
  \[14862]*  = ~\[14862] ,
  \[15456]*  = ~\[15456] ,
  \[10612]_inv*  = ~\[10612]_inv ,
  \[15558]  = \VSACKi*  & STARTi,
  \[15646]*  = ~\[15646] ,
  \[15663]*  = ~\[15663] ,
  \[15367]  = \[15680]*  & PCCsync,
  \[10497]*  = ~\[10497] ,
  \[15369]  = \[15550]*  & \[15697]* ,
  \RESETi*  = ~RESETi,
  \[15553]  = \RESETi*  & slaveXXXXstate0,
  \[14533]*  = ~\[14533] ,
  virmachXXXXEn_VDBufo = \[15452] ,
  \[15176]  = \[15412]*  & \[15574]* ,
  resetXXXXReset = \[15676] ,
  \[10813]_inv  = masterXXXXstate0 | (\[15646]*  | \PCCReq* ),
  \{orXXXXSBCAckCodelatch}  = \[2836]  | (\[15041]  | (\[14469]  | \[15336] )),
  \[15560]  = \PCCSawReset*  & resetXXXXstate1,
  \[10937]_inv  = SBCResetPCC | SingleStep,
  \[15137]*  = ~\[15137] ,
  \[14723]*  = ~\[14723] ,
  \[14769]*  = ~\[14769] ,
  \[15182]  = \[10918]_inv*  & \[15349]* ,
  nextstateXXXXCoherencyState2o = \[15334] ,
  \[10657]_inv*  = ~\[10657]_inv ,
  \PCCReq*  = ~PCCReq,
  \[15327]*  = ~\[15327] ,
  \[14959]*  = ~\[14959] ,
  \[13753]_inv*  = ~\[13753]_inv ,
  \[14997]*  = ~\[14997] ,
  \[15538]*  = ~\[15538] ,
  \[15377]  = \[15541]*  & \[10923]_inv ,
  \{slaveXXXXNextState1}  = I105 | \[14478]* ,
  \[15707]*  = ~\[15707] ,
  \[10912]_inv  = STARTi | ACKi,
  \{slaveXXXXNextState2}  = I126 | \[14484]* ,
  \[15379]  = \[15702]*  & \[15646] ,
  \[10483]_inv  = PCCReqCode1 | \[10507]_inv ,
  \[15569]  = \PCCReqCode1*  & PCCReqCode0,
  \[15184]  = \PCCAckCode*  & \[15452] ,
  \{slaveXXXXNextState0}  = I130 | I131,
  \[10612]_inv  = P_receive_cancel | (\[10945]_inv  | \[10911]_inv ),
  \[10882]_inv*  = ~\[10882]_inv ,
  \[15566]  = \VSACKi*  & masterXXXXstate2,
  \[15021]*  = ~\[15021] ,
  \[15190]  = \[15489]*  & \[10936]_inv ,
  \[14726]*  = ~\[14726] ,
  \[14764]*  = ~\[14764] ,
  \[15211]*  = ~\[15211] ,
  \[15192]  = \[15481]*  & \[13753]_inv* ,
  \[15232]*  = ~\[15232] ,
  \[15382]  = \[15574]*  & VACKl,
  \[15572]  = \physrecXXXXstate0*  & P_receive_cancel,
  \[15558]*  = ~\[15558] ,
  \[10822]_inv*  = ~\[10822]_inv ,
  \[15198]  = \PCCReqCode3*  & (\PCCReqCode2*  & \[15569]* ),
  \[15665]*  = ~\[15665] ,
  \[15686]*  = ~\[15686] ,
  \[15577]  = slaveXXXXstate1 & slaveXXXXstate2,
  \[14409]  = \[10580]*  & (\[14480]*  & (\[14751]*  & \[14959]* )),
  I105 = \RESETi*  & \[10696]_inv* ,
  \[10422]  = I515 | I516,
  I108 = \SBCResetPCC*  & \[14409]* ,
  I109 = \[10889]_inv*  & \[14490]* ,
  \[15389]  = \[15541]*  & \[15670]* ,
  \[10591]*  = ~\[10591] ,
  \[15574]  = \masterXXXXstate3*  & masterXXXXstate1,
  I126 = \RESETi*  & \[14571]* ,
  I128 = \SBCResetPCC*  & \[14525]* ,
  I130 = \[10682]_inv*  & \[10944]_inv* ,
  I131 = \[14539]*  & \[15553] ,
  I139 = \SBCResetPCC*  & \[14503]* ,
  \[10507]_inv*  = ~\[10507]_inv ,
  I140 = \resetXXXXstate1*  & \[15604] ,
  \[15041]*  = ~\[15041] ,
  \[10921]_inv  = slaveXXXXstate2 | \STARTi* ,
  I163 = \LastRQSTi*  & \[14659]* ,
  I164 = \ACKl*  & \[15545] ,
  I167 = \[10817]_inv*  & \[15148]* ,
  I172 = \SBCResetPCC*  & \[14661]* ,
  \[10908]_inv*  = ~\[10908]_inv ,
  I173 = \RESETi*  & \[10559]_inv* ,
  I177 = VSACKi & slaveXXXXstate1,
  I179 = \LastRQSTi*  & \[14830]* ,
  \[14411]  = \[14448]*  & \[14902] ,
  \[10918]_inv*  = ~\[10918]_inv ,
  \[15252]*  = ~\[15252] ,
  \[14808]*  = ~\[14808] ,
  \[15582]  = physrecXXXXstate0 & physrecXXXXstate1,
  I187 = \TM0i*  & \[14816] ,
  I188 = \[10935]_inv*  & \[10190] ,
  \[15290]*  = ~\[15290] ,
  I192 = \[14852]  & VTM1l,
  \[10928]_inv*  = ~\[10928]_inv ,
  \[15391]  = \[15541]*  & \[15692]* ,
  I193 = \[10624]_inv*  & \[15529] ,
  \[15304]*  = ~\[15304] ,
  \[15329]*  = ~\[15329] ,
  I199 = \[10866]_inv*  & PCCAck,
  \[14900]*  = ~\[14900] ,
  \[15367]*  = ~\[15367] ,
  \[14915]*  = ~\[14915] ,
  \[10821]_inv  = \[15646]*  | \masterXXXXstate3* ,
  \[10938]_inv*  = ~\[10938]_inv ,
  \[10682]_inv  = \[10907]_inv  | \[10921]_inv ,
  \[10877]_inv*  = ~\[10877]_inv ,
  \[10935]_inv  = SBCResetPCC | \ACKi* ,
  \[10721]_inv  = \STARTi*  | I543,
  \[15442]*  = ~\[15442] ,
  \[15495]*  = ~\[15495] ,
  \[10882]_inv  = masterXXXXstate0 | \masterXXXXstate3* ,
  \[10897]_inv*  = ~\[10897]_inv ,
  \[2838]*  = ~\[2838] ,
  \[14417]  = \[14443]  & PCCReqCode1,
  \[15670]*  = ~\[15670] ,
  \[15587]  = \STARTi*  & VSACKi,
  \[14419]  = \[14492]*  & (\[14757]*  & \[15105]* ),
  I201 = \[14897]  & masterXXXXstate3,
  I207 = \[10750]_inv*  & \[15357] ,
  I208 = \[10624]_inv*  & \[15529] ,
  \[10696]_inv  = \[10335]  | \[15707] ,
  I211 = \ACKi*  & \[10662]_inv* ,
  \[15399]  = \[15637]*  & \[15653]* ,
  I214 = \[10823]_inv*  & \[14781]* ,
  I215 = \STARTi*  & \[15223] ,
  I219 = \[10889]_inv*  & \[14733]* ,
  \[14603]  = \VSACKi*  & \[14711]* ,
  I220 = \[10937]_inv*  & \[14730] ,
  I222 = \[10935]_inv*  & \[14747]* ,
  I223 = \[14816]  & \[15538] ,
  \[14448]*  = ~\[14448] ,
  I229 = \[14944]*  & \[15109]* ,
  I231 = \slaveXXXXstate2*  & \PCCsync* ,
  I232 = slaveXXXXstate2 & \[14963]* ,
  \[15393]  = \masterXXXXstate3*  & \[15591] ,
  I235 = \slaveXXXXstate1*  & \[14963]* ,
  I236 = \[10944]_inv*  & \[15510]* ,
  \[15396]  = \RQSTi*  & \[15646] ,
  \[14593]*  = ~\[14593] ,
  \[10918]_inv  = TM1i | \TM0i* ,
  \[10817]_inv*  = ~\[10817]_inv ,
  \[10559]_inv  = \[10912]_inv  | I361,
  \[14617]*  = ~\[14617] ,
  \[15159]*  = ~\[15159] ,
  \[14730]*  = ~\[14730] ,
  \[14802]  = \[10685]_inv*  & \[10918]_inv* ,
  I273 = \PCCAck*  & \[10866]_inv* ,
  I276 = \TM1i*  & \[10863]_inv* ,
  I279 = \[10933]_inv*  & \[10907]_inv* ,
  \[14421]  = \[14862]*  & \[14450] ,
  I280 = \RESETi*  & \[14997]* ,
  I282 = \[10928]_inv*  & masterXXXXstate1,
  I284 = \[10921]_inv*  & \[15327]* ,
  I285 = \[15367]*  & slaveXXXXstate2,
  I287 = \[10945]_inv*  & \[15081]* ,
  I288 = \[10845]_inv*  & \[15582] ,
  I292 = \PCCSawReset*  & \[15129]* ,
  I295 = \TM0i*  & \[15349]* ,
  \[15591]  = \STARTi*  & masterXXXXstate2,
  I296 = \[15050]*  & physrecXXXXstate1,
  I299 = \[10657]_inv*  & \[10658]_inv* ,
  \[15349]*  = ~\[15349] ,
  \[14808]  = \[14987]*  & \[15159]* ,
  \[15577]*  = ~\[15577] ,
  \[14617]  = \[14666]*  & masterXXXXstate3,
  nubusXXXXL_PABufi = \{nubusXXXXL_PABufi} ,
  \[14619]  = \[14730]*  & \[15021]* ,
  I300 = \[10748]_inv*  & PCCReqCode1,
  orXXXXRESETo = \{orXXXXRESETo} ,
  I304 = \[10924]_inv*  & \[15176]* ,
  I305 = \masterXXXXstate0*  & \[10928]_inv* ,
  masterXXXXEn_ABufo = \[14535] ,
  \[10632]  = I219 | I220,
  \[14804]  = \[10750]_inv*  & \[15120]* ,
  \[10061]  = I235 | I236,
  \[15599]  = VTM0i & \VSACKi* ,
  \[14409]*  = ~\[14409] ,
  I322 = \[15206]*  & \[15577] ,
  I323 = \[10363]  & \[15707] ,
  I340 = \[10928]_inv*  & \[15300]* ,
  I341 = \[15379]  & masterXXXXstate3,
  \[14575]*  = ~\[14575] ,
  I348 = \[15393]*  & \[15545]* ,
  I354 = \[15407]*  & RESETi,
  \[15081]*  = ~\[15081] ,
  I357 = \RQSTi*  & \[15465]* ,
  I361 = \[15377]*  & \[15670]* ,
  I363 = \[10651]_inv*  & \[10943]_inv* ,
  I364 = \[10882]_inv*  & masterXXXXstate2,
  I366 = \[15418]*  & \[15456]* ,
  \[10750]_inv  = \[10819]_inv  | \slaveXXXXstate2* ,
  I368 = \[10939]_inv*  & \[15692] ,
  \[15133]*  = ~\[15133] ,
  I369 = \[2536]  & ACKi,
  I373 = \[15582]*  & \[15538] ,
  I374 = \[15266]*  & physrecXXXXstate1,
  I377 = \SlotSpace_Id_Match*  & \[10897]_inv* ,
  \[15292]*  = ~\[15292] ,
  \PCCAck*  = ~PCCAck,
  I398 = \[10721]_inv*  & \[10877]_inv* ,
  I399 = \[15310]*  & slaveXXXXstate2,
  \[15344]*  = ~\[15344] ,
  \[14902]*  = ~\[14902] ,
  \[10703]_inv  = \[10817]_inv  | I229,
  \[15369]*  = ~\[15369] ,
  \[14940]*  = ~\[14940] ,
  \[14955]*  = ~\[14955] ,
  \[14993]*  = ~\[14993] ,
  \TM0i*  = ~TM0i,
  \{masterXXXXUpdateReq}  = masterXXXXVSACKo | (\[14505]  | \[14757] ),
  \[10658]_inv*  = ~\[10658]_inv ,
  \[10483]_inv*  = ~\[10483]_inv ,
  \[14627]  = \[2]  & \[14879]* ,
  \[10640]  = I340 | I341,
  \[10422]*  = ~\[10422] ,
  \[10688]_inv  = \[10327]  | \Intr_done* ,
  \[10888]_inv  = RESETi | Intr_done,
  I88 = \[10483]_inv*  & PCCReqCode2,
  I91 = \[10889]_inv*  & \[10089] ,
  \[14488]*  = ~\[14488] ,
  orXXXXVSACKo = \{orXXXXVSACKo} ,
  \[14816]  = \SBCResetPCC*  & \[10685]_inv* ,
  virmachXXXXSBCCacheRelease = \[15169] ,
  \[2536]  = I450 | I451,
  virmachXXXXSBCConfigure = \{virmachXXXXSBCConfigure} ,
  \[14521]*  = ~\[14521] ,
  \[14595]*  = ~\[14595] ,
  \[2537]  = I599 | \wd_cnt_test* ,
  I450 = \nubusXXXXstate1*  & \[10940]_inv* ,
  I451 = \[10897]_inv*  & nubusXXXXstate0,
  I453 = \masterXXXXstate1*  & \[15591]* ,
  \[14619]*  = ~\[14619] ,
  \[10930]_inv*  = ~\[10930]_inv ,
  I465 = \V_transmit_begin*  & \virmachXXXXstate1* ,
  \[14711]*  = ~\[14711] ,
  \[10940]_inv*  = ~\[10940]_inv ,
  I475 = \[15574]  & VSACKi,
  I476 = \ACKl*  & masterXXXXstate1,
  \[14441]  = \[14496]*  & \PCCReqCode2* ,
  \[14821]  = \[15091]*  & (\[15643]*  & (\[15614]*  & PCCReq)),
  \[13378]_inv  = \[10061]  | I177,
  \physrecXXXXstate1*  = ~physrecXXXXstate1,
  \[14922]*  = ~\[14922] ,
  \[15389]*  = ~\[15389] ,
  \physrecXXXXstate0*  = ~physrecXXXXstate0,
  \TM1i*  = ~TM1i,
  \[15481]*  = ~\[15481] ,
  \{masterXXXXNextState1}  = \[14411]*  | I91,
  masterXXXXRQSTo = \[14531] ,
  \[14448]  = \SBCResetPCC*  & \[14488]* ,
  \{masterXXXXNextState2}  = \[14419]*  | \[14769]* ,
  \TM1l*  = ~TM1l,
  \[10816]_inv  = \[15702]*  | \BUS_Inactive* ,
  \{masterXXXXNextState3}  = I108 | I109,
  \[15692]*  = ~\[15692] ,
  \PCCSawReset*  = ~PCCSawReset,
  \[10573]_inv  = \[10929]_inv  | (\[15329]  | (masterXXXXstate1 | \[10882]_inv )),
  slaveXXXXSnoopAddrFromProc = \[14681] ,
  \[14634]  = \[10934]_inv*  & (\Intr_req*  & (\[14900]*  & slaveXXXXstate2)),
  I515 = STARTi & ACKi,
  I516 = \[10912]_inv*  & slaveXXXXstate0,
  \[14443]  = \[14512]*  & PCCReqCode0,
  \[14823]  = \[15021]  & PCCConfirm,
  \{masterXXXXNextState0}  = \[14541]  | (\[15247]  | \[10632] ),
  I536 = \PCCReqCode0*  & PCCReqCode2,
  I537 = PCCReqCode0 & \PCCReqCode2* ,
  \BUS_Inactive*  = ~BUS_Inactive,
  I543 = \STARTo*  & VTM0l,
  \[14450]  = \[14505]*  & \PCCReqCode0* ,
  \[14640]  = \[10643]_inv*  & (\[15344]*  & PCCConfirm),
  \[14830]  = \physrecXXXXstate0*  & \[14980]* ,
  \[14698]*  = ~\[14698] ,
  \{orXXXXEn_START}  = I128 | \[15046]* ,
  \[15120]*  = ~\[15120] ,
  \[15135]*  = ~\[15135] ,
  \[10897]_inv  = STARTi | \nubusXXXXstate1* ,
  \[14804]*  = ~\[14804] ,
  \[10911]_inv  = \TM0i*  | \physrecXXXXstate1* ,
  \[10089]  = I475 | I476,
  \[15310]*  = ~\[15310] ,
  I599 = \TM0i*  & \P_receive_cancel* ,
  \[14942]*  = ~\[14942] ,
  \[14980]*  = ~\[14980] ,
  \[10653]  = I363 | I364,
  \[10511]_inv  = \[15362]  | \[10817]_inv* ,
  \[15536]*  = ~\[15536] ,
  \[15553]*  = ~\[15553] ,
  \[14838]  = \masterXXXXstate1*  & \[14970]* ,
  \[15574]*  = ~\[15574] ,
  \[15599]*  = ~\[15599] ,
  \[10878]_inv*  = ~\[10878]_inv ,
  \{resetXXXXNextState1}  = \[15676]  | I292,
  \[10888]_inv*  = ~\[10888]_inv ,
  \{resetXXXXNextState2}  = \[15676]  | I354,
  \[10686]_inv  = I366 | \[15624]* ,
  \[14659]*  = ~\[14659] ,
  \[10886]_inv  = STARTo | (ACKi | \STARTi* ),
  \[15176]*  = ~\[15176] ,
  \[14751]*  = ~\[14751] ,
  \[10908]_inv  = slaveXXXXstate0 | slaveXXXXstate1,
  \nubusXXXXstate0*  = ~nubusXXXXstate0,
  \[10749]_inv  = SingleStep | \[15344]* ,
  \[15407]*  = ~\[15407] ,
  \nubusXXXXstate1*  = ~nubusXXXXstate1,
  \[14467]  = \[10126]*  & \[10483]_inv ,
  \{nubusXXXXL_PABufi}  = \[10688]_inv  | \RESETi* ,
  \[15710]*  = ~\[15710] ,
  \[14469]  = \SBCResetPCC*  & \[14508]* ,
  \[14659]  = \[14771]*  & \[15545]* ,
  \{orXXXXACKo}  = masterXXXXACKo | \[15219] ,
  orXXXXVACKo = \{orXXXXVACKo} ,
  \[14654]  = \[10907]_inv*  & (\[14950]*  & slaveXXXXstate2),
  \{orXXXXVTM0o}  = masterXXXXVSACKo | (\[15159]  | (\[14852]  | \[15184] )),
  \[14443]*  = ~\[14443] ,
  \[15003]  = \wdcntXXXXstate2*  & (\[15418]  & Incr_wd_cnt),
  orXXXXSBCAck = \{orXXXXSBCAck} ,
  \[14846]  = \[14922]*  & \[15545]* ,
  \[10940]_inv  = nubusXXXXstate0 | \STARTi* ,
  \[15068]*  = ~\[15068] ,
  \[10936]_inv*  = ~\[10936]_inv ,
  \[10946]_inv*  = ~\[10946]_inv ,
  \wd_cnt_test*  = ~wd_cnt_test,
  \[14852]  = \[10750]_inv*  & \[15655] ,
  \[14771]*  = ~\[14771] ,
  \{slaveXXXXL_VABufi}  = \[14634]  | (\[15280]  | (RESETi | \[14674] )),
  \[14661]  = \[14966]*  & (\[15039]*  & \[10653]* ),
  slaveXXXXSnoopVTag_W = \[14681] ,
  \[14823]*  = ~\[14823] ,
  \[2537]*  = ~\[2537] ,
  \[15011]  = \slaveXXXXstate2*  & (\[10944]_inv*  & (\[10886]_inv*  & \[10936]_inv* )),
  \[14982]*  = ~\[14982] ,
  \[15427]*  = ~\[15427] ,
  \[10748]_inv*  = ~\[10748]_inv ,
  \[10945]_inv*  = ~\[10945]_inv ,
  \[10296]  = I214 | I215,
  \[14478]  = \[1]  & \slaveXXXXstate1* ,
  \[14668]  = \[14823]*  & \[15137]* ,
  masterXXXXEn_PDBufi = \[10703]_inv* ,
  masterXXXXEn_PDBufo = \[15247] ,
  \[14857]  = \[15064]*  & \[15442]* ,
  \[10854]_inv  = \[10890]_inv  | \wdcntXXXXstate2* ,
  \[15017]  = \[10817]_inv*  & (\[15591]  & (VTM0i & VSACKi)),
  \VACKi*  = ~VACKi,
  \[10492]  = I139 | I140,
  \[10533]*  = ~\[10533] ,
  \[10817]_inv  = \[10889]_inv  | \masterXXXXstate3* ,
  \[14484]*  = ~\[14484] ,
  \[14666]  = \[14924]*  & (\[15396]*  & (\[15338]*  & \[15379]* )),
  \[14508]*  = ~\[14508] ,
  \[15206]  = \[15536]*  & (\[15707]*  & \[15506]* ),
  \[14480]  = \RQSTi*  & \[14517]* ,
  \[10878]_inv  = masterXXXXstate1 | (SBCResetPCC | masterXXXXstate0),
  \[14860]  = \[10907]_inv*  & (\[15215]*  & STARTi),
  \Intr_req*  = ~Intr_req,
  \[14862]  = \[15041]*  & \[15219]* ,
  \[10497]  = I373 | I374,
  \RQSTi*  = ~RQSTi,
  \[15219]*  = ~\[15219] ,
  \[15021]  = \[10822]_inv*  & (\[15566]  & BUS_Inactive),
  \[15211]  = \[15492]*  & \[15499]* ,
  \[10935]_inv*  = ~\[10935]_inv ,
  \[10493]  = I222 | I223,
  \[10890]_inv*  = ~\[10890]_inv ,
  \[14488]  = \[14726]*  & (\[14959]*  & \[14521]* ),
  \[13378]_inv*  = ~\[13378]_inv ,
  \[15637]*  = ~\[15637] ,
  \[15658]*  = ~\[15658] ,
  \[15407]  = Gen_Reset & \[15658] ,
  \[15712]*  = ~\[15712] ,
  \[10506]_inv  = \[14723]  | \SBCResetPCC* ,
  \[14484]  = \[14543]*  & \[14860]* ,
  \[14674]  = \slaveXXXXstate0*  & (\[14946]*  & ACKi),
  \[15219]  = \STARTi*  & (\[10938]_inv*  & (\[15692]  & Intr_done)),
  \{wdcntXXXXwd_cnt_test}  = \[10686]_inv*  | \[15030]* ,
  \[14676]  = \[14804]*  & \[14852]* ,
  \[15403]  = \RESETi*  & \[15658]* ,
  \[15026]  = \[14]  & V_transmit_begin,
  \[10863]_inv  = \[10940]_inv  | \[10907]_inv ,
  \[15003]*  = ~\[15003] ,
  \[14490]  = \[10591]*  & \[14617]* ,
  \[15215]  = \[15495]*  & \[15577]* ,
  \[15405]  = \[15680]*  & \slaveXXXXstate2* ,
  \[15030]  = \[15]  & \[15508]* ,
  \[15410]  = \[10890]_inv*  & wdcntXXXXstate0,
  \[15141]*  = ~\[15141] ,
  \[14492]  = \SBCResetPCC*  & \[14533]* ,
  \[10750]_inv*  = ~\[10750]_inv ,
  \[14681]  = \RESETi*  & (\[14942]*  & (\[15707]  & UpdateReq)),
  \[14871]  = \SingleStep*  & (\[15465]*  & (\[15232]  & BUS_Inactive)),
  \[15412]  = \masterXXXXstate3*  & \[10894]_inv* ,
  \[1048]*  = ~\[1048] ,
  \[15298]*  = ~\[15298] ,
  \[14846]*  = ~\[14846] ,
  \slaveXXXXstate2*  = ~slaveXXXXstate2,
  \slaveXXXXstate1*  = ~slaveXXXXstate1,
  \[10686]_inv*  = ~\[10686]_inv ,
  wdcntXXXXNextState1 = \[14857]* ,
  \slaveXXXXstate0*  = ~slaveXXXXstate0,
  wdcntXXXXNextState2 = \[14797]* ,
  wdcntXXXXNextState3 = \[14984]* ,
  \[10696]_inv*  = ~\[10696]_inv ,
  \[10901]_inv  = ACKl | \masterXXXXstate2* ,
  \[15521]*  = ~\[15521] ,
  \[14688]  = \[3]  & \[10882]_inv ,
  \[15228]  = \[10946]_inv*  & (VTM0i & (VACKi & virmachXXXXstate1)),
  \[15418]  = \[10890]_inv*  & wdcntXXXXstate3,
  \[15037]  = \PCCReqCode0*  & (\[10929]_inv*  & \[15686] ),
  \[14879]  = \SBCResetPCC*  & \[10748]_inv* ,
  \[14494]  = \SBCResetPCC*  & \[14547]* ,
  \[15039]  = \[15235]*  & \BUS_Inactive* ,
  \wdcntXXXXstate3*  = ~wdcntXXXXstate3,
  \[10662]_inv  = \[10307]  | \[10888]_inv* ,
  \wdcntXXXXstate2*  = ~wdcntXXXXstate2,
  \[15604]  = \RESETi*  & resetXXXXstate2,
  \[14496]  = \[15697]*  & \[10507]_inv ,
  \[15223]  = \masterXXXXstate3*  & (\[15646]  & masterXXXXstate0),
  \[1048]  = I299 | I300,
  \[15416]  = \P_receive_cancel*  & \[10918]_inv* ,
  \[10]  = \[15349]*  | \[15439] ,
  \[15035]  = \[530]*  & (\[15643]*  & (\[15614]*  & \[15686]* )),
  \PCCAckCode*  = ~PCCAckCode,
  \[14640]*  = ~\[14640] ,
  \[11]  = \[15310]*  | \[15252]* ,
  \[14676]*  = ~\[14676] ,
  \[15230]  = \[2537]*  & \[15663]* ,
  \[14693]*  = ~\[14693] ,
  \[12]  = \[15444]*  | \[15329]* ,
  \[14717]*  = ~\[14717] ,
  \wdcntXXXXstate1*  = ~wdcntXXXXstate1,
  \[15182]*  = ~\[15182] ,
  \[13]  = \[15710]*  | \[15456]* ,
  \[10939]_inv  = STARTi | nubusXXXXstate0,
  \[15232]  = \[530]*  & \[15512]* ,
  \[14830]*  = ~\[14830] ,
  \[14]  = \[15492]*  | \[15499]* ,
  \[13753]_inv  = SBCResetPCC | virmachXXXXstate0,
  \[15041]  = \[10821]_inv*  & (\[10889]_inv*  & \[15702] ),
  \[15]  = \[15668]*  | \[15410]* ,
  \[16]  = \[15637]*  | \[15646]* ,
  \[15403]*  = ~\[15403] ,
  \[17]  = \[15526]*  | VTM0l,
  \[15487]*  = ~\[15487] ,
  \[18]  = \V_transmit_begin*  | V_receive_begin,
  \[15541]*  = ~\[15541] ,
  \[14698]  = \[14767]*  & \[15304]* ,
  virmachXXXXSBCsetDirty = \[15228] ,
  \[15614]*  = ~\[15614] ,
  \[15427]  = \[10911]_inv*  & TM1i,
  \[10685]_inv*  = ~\[10685]_inv ,
  resetXXXXSBCResetPCC = \{resetXXXXSBCResetPCC} ,
  \[14693]  = \[10924]_inv*  & \[14846]* ,
  \[14883]  = \[10888]_inv*  & (\[10912]_inv*  & \[15141]* ),
  \[14411]*  = ~\[14411] ,
  \[15614]  = PCCReqCode0 & PCCReqCode2,
  \[15046]  = \[15296]*  & \[15247]* ,
  \[14547]*  = ~\[14547] ,
  \[15026]*  = ~\[15026] ,
  \[15235]  = \[10823]_inv*  & GRANTi,
  \[15425]  = \[10933]_inv*  & ACKi,
  \[15064]*  = ~\[15064] ,
  \[15089]*  = ~\[15089] ,
  \[15050]  = \physrecXXXXstate0*  & (\[15416]*  & (\[15538]*  & wd_cnt_test)),
  \[15240]  = \[10863]_inv*  & (\Intr_done*  & \nubusXXXXstate1* ),
  orXXXXEn_VCNTL = \{orXXXXEn_VCNTL} ,
  \[10930]_inv  = \PCCReq*  | \PCCReqCode3* ,
  \[15052]  = \[10878]_inv*  & (UpdateDone & masterXXXXstate2),
  \[10923]_inv*  = ~\[10923]_inv ,
  \[10866]_inv*  = ~\[10866]_inv ,
  \[10933]_inv*  = ~\[10933]_inv ,
  \[10943]_inv*  = ~\[10943]_inv ,
  \[10886]_inv*  = ~\[10886]_inv ,
  \[15444]*  = ~\[15444] ,
  \[10685]_inv  = \[10943]_inv  | I348,
  \[15582]*  = ~\[15582] ,
  \[10944]_inv  = slaveXXXXstate1 | \VTM0l* ,
  \[100]  = \[14883] ,
  \[14897]  = \[10748]_inv*  & PCCReqCode2,
  \[101]  = \[15190] ,
  \[15697]*  = ~\[15697] ,
  \[15247]  = \[10889]_inv*  & (\masterXXXXstate3*  & \[10901]_inv* ),
  \[102]  = \{masterXXXXUpdateReq} ,
  \{orXXXXSBCAckCode1}  = I187 | I188,
  \[103]  = \[14681] ,
  \{orXXXXSBCAckCode2}  = \[10492]  | \[10493] ,
  \[10907]_inv  = ACKi | RESETi,
  \[15439]  = \[10911]_inv*  & wd_cnt_test,
  \[10544]_inv  = \[10894]_inv  | I357,
  \[104]  = \{orXXXXReset_wd_cnt_x} ,
  \{orXXXXSBCAckCode3}  = \[15604]  | \[14627]* ,
  \[15054]  = \[10612]_inv*  & (\wd_cnt_test*  & \physrecXXXXstate0* ),
  \[15624]  = wdcntXXXXstate1 & wdcntXXXXstate2,
  \[105]  = \[14467] ,
  \[14490]*  = ~\[14490] ,
  \{orXXXXVACKo}  = \[15041]  | \[15169] ,
  \[10816]_inv*  = ~\[10816]_inv ,
  \[106]  = \{orXXXXIncr_wd_cnt} ,
  \[15056]  = \RESETi*  & (\[10886]_inv*  & VTM0l),
  \[107]  = \{wdcntXXXXwd_cnt_test} ,
  \[10507]_inv  = \[10894]_inv  | (\[14688]  | \[10937]_inv ),
  \[15046]*  = ~\[15046] ,
  \[108]  = \[14443] ,
  \[109]  = \[15017] ,
  \{orXXXXSBCAckCode0}  = \[14469]  | \[14911] ,
  \[14757]*  = ~\[14757] ,
  \{slaveXXXXSBCReqCode0}  = I192 | I193,
  \[15215]*  = ~\[15215] ,
  \PCCsync*  = ~PCCsync,
  \[15252]  = \[10933]_inv*  & (\[10934]_inv*  & (Intr_req & slaveXXXXstate0)),
  \[15442]  = \[10890]_inv*  & wdcntXXXXstate1,
  \[14909]*  = ~\[14909] ,
  \[15391]*  = ~\[15391] ,
  \[15405]*  = ~\[15405] ,
  \[10845]_inv*  = ~\[10845]_inv ,
  \[15489]*  = ~\[15489] ,
  \[110]  = \[15017] ,
  \[15068]  = \[530]*  & (\[10816]_inv*  & \[15569] ),
  \[111]  = \[14852] ,
  \{slaveXXXXSBCReqCode1}  = I207 | I208,
  orXXXXSBCAckCodelatch = \{orXXXXSBCAckCodelatch} ,
  \[15637]  = STARTi & VSACKi,
  \{orXXXXEn_VCNTL}  = \[14523]  | (\[15192]  | \[10525] ),
  \[10580]*  = ~\[10580] ,
  \[15064]  = \[10854]_inv*  & (Incr_wd_cnt & wdcntXXXXstate3),
  \[15444]  = \masterXXXXstate0*  & \[10930]_inv* ,
  \[14503]*  = ~\[14503] ,
  \[15066]  = \[15674]*  & \[15247] ,
  orXXXXSBCAckCode0 = \{orXXXXSBCAckCode0} ,
  orXXXXSBCAckCode1 = \{orXXXXSBCAckCode1} ,
  orXXXXSBCAckCode2 = \{orXXXXSBCAckCode2} ,
  \masterXXXXstate3*  = ~masterXXXXstate3,
  orXXXXSBCAckCode3 = \{orXXXXSBCAckCode3} ,
  \[15446]  = \[10923]_inv*  & nubusXXXXstate1,
  \[15030]*  = ~\[15030] ,
  \masterXXXXstate2*  = ~masterXXXXstate2,
  \[15235]*  = ~\[15235] ,
  \[15452]  = \virmachXXXXstate1*  & \[10946]_inv* ,
  \[15294]*  = ~\[15294] ,
  \[14852]*  = ~\[14852] ,
  \{orXXXXL_DBufo}  = \[14952]  | (\[15159]  | (\[14450]  | \[14441] )),
  \masterXXXXstate1*  = ~masterXXXXstate1,
  \[15410]*  = ~\[15410] ,
  \[15425]*  = ~\[15425] ,
  \masterXXXXstate0*  = ~masterXXXXstate0,
  \[15446]*  = ~\[15446] ,
  \{physrecXXXXNextState1}  = I287 | I288,
  orXXXXEn_CNTL = \{orXXXXEn_CNTL} ,
  \[15508]*  = ~\[15508] ,
  \[10877]_inv  = slaveXXXXstate1 | slaveXXXXstate2,
  \[15653]*  = ~\[15653] ,
  \[15674]*  = ~\[15674] ,
  \[15079]  = \[15319]*  & \[15637]* ,
  \[15074]  = \masterXXXXstate1*  & \[15355]* ,
  \[14492]*  = ~\[14492] ,
  \[15643]  = \PCCReqCode0*  & PCCReqCode1,
  \[15266]  = \physrecXXXXstate0*  & \[2537]* ,
  \[15456]  = \[10890]_inv*  & Incr_wd_cnt,
  \[15646]  = \masterXXXXstate1*  & \masterXXXXstate2* ,
  \[15050]*  = ~\[15050] ,
  \[14661]*  = ~\[14661] ,
  \[15148]*  = ~\[15148] ,
  \[10307]  = \[2536]  | I377,
  \[14797]*  = ~\[14797] ,
  \[15081]  = \[15298]*  & \[15439]* ,
  \[10089]*  = ~\[10089] ,
  \[15338]*  = ~\[15338] ,
  \[10643]_inv*  = ~\[10643]_inv ,
  \[14924]*  = ~\[14924] ,
  \[14987]*  = ~\[14987] ,
  \[10929]_inv  = masterXXXXstate2 | \[10930]_inv ,
  \[10573]_inv*  = ~\[10573]_inv ,
  \[10866]_inv  = \[13753]_inv  | I465,
  \PCCConfirm*  = ~PCCConfirm,
  \[15658]  = \resetXXXXstate0*  & \resetXXXXstate1* ,
  \[15089]  = \CoherencyState2i*  & \[15353]* ,
  \{nubusXXXXNuBusActive}  = \[14990]  | \[15240] ,
  \[15653]  = \STARTi*  & \VSACKi* ,
  \[14505]*  = ~\[14505] ,
  \[14543]*  = ~\[14543] ,
  \[15276]  = \nubusXXXXstate1*  & (\[10939]_inv*  & (\[10888]_inv*  & ACKi)),
  \[15085]  = \[15288]*  & \[15418] ,
  \[15465]  = \[15686]  & PCCReqCode0,
  \[15655]  = \TM1l*  & CoherencyState2i,
  \[15085]*  = ~\[15085] ,
  \{virmachXXXXSBCConfigure}  = \[14952]  | \[15452] ,
  \[15280]  = \[10912]_inv*  & (\slaveXXXXstate2*  & \[10908]_inv* ),
  \[15109]*  = ~\[15109] ,
  \[14733]*  = ~\[14733] ,
  \[15296]*  = ~\[15296] ,
  \[15091]  = \PCCReqCode3*  & \[15284]* ,
  \[14871]*  = ~\[14871] ,
  \[15471]  = \slaveXXXXstate1*  & \[10921]_inv* ,
  \[15661]  = \SingleStep*  & masterXXXXstate3,
  \[14944]*  = ~\[14944] ,
  \[15412]*  = ~\[15412] ,
  \[10924]_inv*  = ~\[10924]_inv ,
  \[15465]*  = ~\[15465] ,
  \[10863]_inv*  = ~\[10863]_inv ,
  \[10126]  = I536 | I537,
  \[10934]_inv*  = ~\[10934]_inv ,
  \[10944]_inv*  = ~\[10944]_inv ,
  \Tag_Match*  = ~Tag_Match,
  \[15288]  = \[15624]*  & Incr_wd_cnt,
  \[15668]  = \wdcntXXXXstate2*  & \wdcntXXXXstate3* ,
  \[15097]  = \[10877]_inv*  & \[15294]* ,
  \[10458]_inv  = \[15614]  | \[10483]_inv* ,
  \SingleStep*  = ~SingleStep,
  \[10934]_inv  = VSACKi | \slaveXXXXstate1* ,
  \VTM0l*  = ~VTM0l,
  \[15284]  = \SingleStep*  & \[15686]* ,
  \[15663]  = \TM1i*  & \P_receive_cancel* ,
  \[14525]*  = ~\[14525] ,
  \[15665]  = P_receive_cancel & physrecXXXXstate1,
  \[15290]  = \[15521]*  & VSACKi,
  \[15129]*  = ~\[15129] ,
  \[15670]  = \nubusXXXXstate1*  & nubusXXXXstate0,
  \[10327]  = I368 | I369,
  \[10823]_inv*  = ~\[10823]_inv ,
  \[15292]  = \[15591]*  & \[15521]* ,
  \[10899]_inv  = RQSTi | SingleStep,
  \STARTi*  = ~STARTi,
  \[15481]  = \[18]  & \virmachXXXXstate1* ,
  \[15319]*  = ~\[15319] ,
  \[10658]_inv  = \[15512]  | \[10899]_inv* ,
  \[15357]*  = ~\[15357] ,
  encodemuxXXXXMX_AD_8 = \[15198] ,
  \[14508]  = \[2838]*  & (\[14917]*  & \[14723]* ),
  \{nubusXXXXNextState0}  = \[14990]  | I276,
  \[530]  = \[10894]_inv  | \PCCConfirm* ,
  \[15298]  = \[15572]*  & physrecXXXXstate1,
  \STARTo*  = ~STARTo,
  \[15487]  = \wdcntXXXXstate1*  & (Incr_wd_cnt & wdcntXXXXstate3),
  \{nubusXXXXNextState1}  = \[15219]  | I211,
  \[15489]  = \slaveXXXXstate2*  & (PCCAck & slaveXXXXstate1),
  \VTM1l*  = ~VTM1l,
  \[14503]  = \[14640]*  & (\[14717]*  & (\[2838]*  & \[14802]* )),
  \[15294]  = \[15526]*  & STARTi,
  \[15674]  = \STARTi*  & \TM0i* ,
  \[10653]*  = ~\[10653] ,
  \[14505]  = \[15550]*  & \[10507]_inv ,
  \[15296]  = \[10945]_inv*  & \[15582]* ,
  \[15676]  = RESETi & resetXXXXstate2,
  \[10703]_inv*  = ~\[10703]_inv ,
  \[10943]_inv  = \ACKl*  | \masterXXXXstate0* ,
  \[15680]  = \SlotSpace_Id_Match*  & \Intr_req* ,
  \V_transmit_begin*  = ~V_transmit_begin,
  \[10718]  = I322 | I323,
  \[14512]  = \PCCReqCode2*  & \[10507]_inv* ,
  \[10890]_inv  = \SBCResetPCC*  | \Reset_wd_cnt* ,
  \[15492]  = \virmachXXXXstate1*  & (\virmachXXXXstate0*  & V_receive_begin),
  \[84]  = \{masterXXXXNextState0} ,
  \[10643]_inv  = SingleStep | \[15021]* ,
  \[10339]  = I279 | I280,
  \[85]  = \{masterXXXXNextState1} ,
  \[15377]*  = ~\[15377] ,
  \GRANTi*  = ~GRANTi,
  \[14946]*  = ~\[14946] ,
  \[14963]*  = ~\[14963] ,
  \[86]  = \{masterXXXXNextState2} ,
  \[14984]*  = ~\[14984] ,
  \[15452]*  = ~\[15452] ,
  \[87]  = \{masterXXXXNextState3} ,
  \{orXXXXTM1o}  = \[14421]*  | I88,
  \[88]  = \{nubusXXXXNextState0} ,
  \[15529]*  = ~\[15529] ,
  \{slaveXXXXSBCReq}  = \[14654]  | \[14676]* ,
  \[10335]  = I284 | I285,
  \[10525]  = I167 | \[14709]* ,
  \[89]  = \{nubusXXXXNextState1} ,
  masterXXXXVSACKo = \[10458]_inv  | \[14443]* ,
  \[14517]  = \[10586]*  & \[14575]* ,
  \[15680]*  = ~\[15680] ,
  \[14709]  = \[14852]*  & \[15452]* ,
  \[15499]  = \VACKi*  & (virmachXXXXstate0 & virmachXXXXstate1),
  \[10718]*  = ~\[10718] ,
  \[14512]*  = ~\[14512] ,
  \[15686]  = \PCCReqCode1*  & \PCCReqCode2* ,
  \[90]  = \{slaveXXXXNextState0} ,
  \[14900]  = \[7]  & \[10422]* ,
  \[15495]  = \PCCsync*  & \[10877]_inv* ,
  \[14627]*  = ~\[14627] ,
  \[91]  = \{slaveXXXXNextState1} ,
  \[15123]*  = ~\[15123] ,
  \[92]  = \{slaveXXXXNextState2} ,
  \[14902]  = \[8]  & \[10889]_inv ,
  \[93]  = \[14976] ,
  \[14521]  = \[10822]_inv*  & \[14603]* ,
  \[14711]  = \[14871]*  & masterXXXXstate2,
  \[15692]  = \ACKi*  & \nubusXXXXstate1* ,
  \[14838]*  = ~\[14838] ,
  \[94]  = \{resetXXXXNextState1} ,
  \P_receive_cancel*  = ~P_receive_cancel,
  \[95]  = \{resetXXXXNextState2} ,
  \[14966]*  = ~\[14966] ,
  \[96]  = \{virmachXXXXNextState0} ,
  slaveXXXXSBCReq = \{slaveXXXXSBCReq} ,
  \[10624]_inv*  = ~\[10624]_inv ,
  \[10533]  = I179 | \[14661]* ,
  \[97]  = \{virmachXXXXNextState1} ,
  \[98]  = \[15030]* ,
  \[10296]*  = ~\[10296] ,
  \[15587]*  = ~\[15587] ,
  \[99]  = \[14627]* ,
  \[14717]  = \[14897]  & PCCReqCode0,
  \SBCResetPCC*  = ~SBCResetPCC,
  \[15697]  = \PCCReqCode0*  & \PCCReqCode1* ,
  \[14529]  = \SBCResetPCC*  & \[14595]* ,
  slaveXXXXSnoopState_W = \{slaveXXXXSnoopState_W} ,
  \[14909]  = \[9]  & UpdateDone,
  \[14523]  = \[10749]_inv*  & (\SBCResetPCC*  & \[14668]* ),
  \[14419]*  = ~\[14419] ,
  \[10640]*  = ~\[10640] ,
  \[14478]*  = ~\[14478] ,
  \masterXXXXVSACKo*  = ~masterXXXXVSACKo,
  \[14525]  = \[10533]*  & \[15302]* ,
  \[10819]_inv  = \[10944]_inv  | (\[15553]*  | \Tag_Match* ),
  \[14585]*  = ~\[14585] ,
  \{slaveXXXXSnoopState_W}  = \[14681]  | \[14676]* ,
  \[15091]*  = ~\[15091] ,
  \[14668]*  = ~\[14668] ,
  \CoherencyState2i*  = ~CoherencyState2i,
  \[15105]*  = ~\[15105] ,
  \[15143]*  = ~\[15143] ,
  \[14760]*  = ~\[14760] ,
  \[14531]  = \SBCResetPCC*  & \[14593]* ,
  \[14911]  = \physrecXXXXstate0*  & (\[15230]*  & (\[10935]_inv*  & physrecXXXXstate1)),
  \[15379]*  = ~\[15379] ,
  masterXXXXSBC_WriteCache = \{masterXXXXSBC_WriteCache} ,
  \[14950]*  = ~\[14950] ,
  \[15471]*  = ~\[15471] ,
  \[15492]*  = ~\[15492] ,
  \[15506]*  = ~\[15506] ,
  \[15569]*  = ~\[15569] ,
  \[10544]_inv*  = ~\[10544]_inv ,
  \[10651]_inv  = LastRQSTi | I453,
  \[14537]  = \[10061]  & (\[15553]  & slaveXXXXstate2),
  \[14917]  = \[10748]_inv*  & PCCReqCode0,
  \[10854]_inv*  = ~\[10854]_inv ,
  \[15661]*  = ~\[15661] ,
  \[10929]_inv*  = ~\[10929]_inv ,
  \[10939]_inv*  = ~\[10939]_inv ,
  \[14539]  = \[13378]_inv*  & slaveXXXXstate2,
  \[14533]  = \[14585]*  & \[14760]* ,
  \[14723]  = \[10643]_inv*  & \[15232]* ,
  \[10894]_inv*  = ~\[10894]_inv ,
  \[14726]  = \[4]  & \[10544]_inv* ,
  \virmachXXXXstate0*  = ~virmachXXXXstate0,
  \[14535]  = \[10749]_inv*  & (\SBCResetPCC*  & \[14688]* ),
  \[14915]  = \[15056]*  & \[15553]* ,
  \[10924]_inv  = masterXXXXstate0 | masterXXXXstate2,
  \virmachXXXXstate1*  = ~virmachXXXXstate1,
  \[14730]  = \PCCReqCode3*  & (\RQSTi*  & (\[10657]_inv*  & \[15512]* ));
always begin
  Set_ex_wd_cnt1 = \[105] ;
  wd_cnt_test = \[107] ;
  wdcntXXXXstate0 = \[98] ;
  V_transmit_begin = \[111] ;
  virmachXXXXstate0 = \[96] ;
  virmachXXXXstate1 = \[97] ;
  V_receive_begin = \[110] ;
  Reset_wd_cnt = \[104] ;
  Gen_Reset = \[99] ;
  resetXXXXstate0 = \[93] ;
  resetXXXXstate1 = \[94] ;
  resetXXXXstate2 = \[95] ;
  UpdateReq = \[102] ;
  slaveXXXXstate0 = \[90] ;
  slaveXXXXstate1 = \[91] ;
  slaveXXXXstate2 = \[92] ;
  P_receive_cancel = \[109] ;
  UpdateDone = \[103] ;
  masterXXXXstate0 = \[84] ;
  masterXXXXstate1 = \[85] ;
  masterXXXXstate2 = \[86] ;
  masterXXXXstate3 = \[87] ;
  Intr_done = \[101] ;
  P_receive_begin = \[108] ;
  Incr_wd_cnt = \[106] ;
  nubusXXXXstate0 = \[88] ;
  nubusXXXXstate1 = \[89] ;
  Intr_req = \[100] ;
end
initial begin
  Set_ex_wd_cnt1 = 0;
  wd_cnt_test = 0;
  wdcntXXXXstate0 = 0;
  V_transmit_begin = 0;
  virmachXXXXstate0 = 0;
  virmachXXXXstate1 = 0;
  V_receive_begin = 0;
  Reset_wd_cnt = 0;
  Gen_Reset = 0;
  resetXXXXstate0 = 0;
  resetXXXXstate1 = 0;
  resetXXXXstate2 = 0;
  UpdateReq = 0;
  slaveXXXXstate0 = 0;
  slaveXXXXstate1 = 0;
  slaveXXXXstate2 = 0;
  P_receive_cancel = 0;
  UpdateDone = 0;
  masterXXXXstate0 = 0;
  masterXXXXstate1 = 0;
  masterXXXXstate2 = 0;
  masterXXXXstate3 = 0;
  Intr_done = 0;
  P_receive_begin = 0;
  Incr_wd_cnt = 0;
  nubusXXXXstate0 = 0;
  nubusXXXXstate1 = 0;
  Intr_req = 0;
end
endmodule

