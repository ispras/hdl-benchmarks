module lut_output(result, out);
  output result;
  output out;
endmodule