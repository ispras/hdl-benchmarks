//NOTE: no-implementation module stub

module GTECH_OR_NOT (
    input wire A,
    input wire B,
    output wire Z
);

endmodule
