module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 ;
output g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( g245 , n246 );
buf ( g246 , n247 );
buf ( g247 , n248 );
buf ( g248 , n249 );
buf ( g249 , n250 );
buf ( g250 , n251 );
buf ( g251 , n252 );
buf ( g252 , n253 );
buf ( g253 , n254 );
buf ( g254 , n255 );
buf ( g255 , n256 );
buf ( g256 , n257 );
buf ( g257 , n258 );
buf ( g258 , n259 );
buf ( g259 , n260 );
buf ( g260 , n261 );
buf ( g261 , n262 );
buf ( g262 , n263 );
buf ( g263 , n264 );
buf ( g264 , n265 );
buf ( g265 , n266 );
buf ( g266 , n267 );
buf ( g267 , n268 );
buf ( g268 , n269 );
buf ( g269 , n270 );
buf ( g270 , n271 );
buf ( g271 , n272 );
buf ( g272 , n273 );
buf ( g273 , n274 );
buf ( g274 , n275 );
buf ( g275 , n276 );
buf ( g276 , n277 );
buf ( g277 , n278 );
buf ( g278 , n279 );
buf ( g279 , n280 );
buf ( g280 , n281 );
buf ( g281 , n282 );
buf ( g282 , n283 );
buf ( g283 , n284 );
buf ( g284 , n285 );
buf ( g285 , n286 );
buf ( g286 , n287 );
buf ( g287 , n288 );
buf ( g288 , n289 );
buf ( g289 , n290 );
buf ( g290 , n291 );
buf ( g291 , n292 );
buf ( g292 , n293 );
buf ( g293 , n294 );
buf ( g294 , n295 );
buf ( g295 , n296 );
buf ( g296 , n297 );
buf ( g297 , n298 );
buf ( g298 , n299 );
buf ( g299 , n300 );
buf ( g300 , n301 );
buf ( g301 , n302 );
buf ( g302 , n303 );
buf ( g303 , n304 );
buf ( g304 , n305 );
buf ( g305 , n306 );
buf ( g306 , n307 );
buf ( g307 , n308 );
buf ( g308 , n309 );
buf ( g309 , n310 );
buf ( g310 , n311 );
buf ( g311 , n312 );
buf ( g312 , n313 );
buf ( g313 , n314 );
buf ( g314 , n315 );
buf ( g315 , n316 );
buf ( g316 , n317 );
buf ( g317 , n318 );
buf ( g318 , n319 );
buf ( g319 , n320 );
buf ( g320 , n321 );
buf ( g321 , n322 );
buf ( g322 , n323 );
buf ( g323 , n324 );
buf ( g324 , n325 );
buf ( g325 , n326 );
buf ( g326 , n327 );
buf ( g327 , n328 );
buf ( g328 , n329 );
buf ( g329 , n330 );
buf ( g330 , n331 );
buf ( g331 , n332 );
buf ( g332 , n333 );
buf ( g333 , n334 );
buf ( g334 , n335 );
buf ( g335 , n336 );
buf ( g336 , n337 );
buf ( g337 , n338 );
buf ( g338 , n339 );
buf ( g339 , n340 );
buf ( g340 , n341 );
buf ( g341 , n342 );
buf ( g342 , n343 );
buf ( g343 , n344 );
buf ( g344 , n345 );
buf ( n246 , n2365 );
buf ( n247 , n2838 );
buf ( n248 , n2872 );
buf ( n249 , n2414 );
buf ( n250 , n2905 );
buf ( n251 , n2962 );
buf ( n252 , n3173 );
buf ( n253 , n3285 );
buf ( n254 , n3150 );
buf ( n255 , n3213 );
buf ( n256 , n3295 );
buf ( n257 , n3157 );
buf ( n258 , n3336 );
buf ( n259 , n2970 );
buf ( n260 , n3067 );
buf ( n261 , n3001 );
buf ( n262 , n3187 );
buf ( n263 , n3223 );
buf ( n264 , n3258 );
buf ( n265 , n3232 );
buf ( n266 , n3238 );
buf ( n267 , n3246 );
buf ( n268 , n3101 );
buf ( n269 , n3035 );
buf ( n270 , n3132 );
buf ( n271 , n3594 );
buf ( n272 , n3616 );
buf ( n273 , n3778 );
buf ( n274 , n3783 );
buf ( n275 , n3613 );
buf ( n276 , n3587 );
buf ( n277 , n3590 );
buf ( n278 , n3610 );
buf ( n279 , n3675 );
buf ( n280 , n3631 );
buf ( n281 , n2074 );
buf ( n282 , n3607 );
buf ( n283 , n3619 );
buf ( n284 , n3774 );
buf ( n285 , n3622 );
buf ( n286 , n3770 );
buf ( n287 , n3598 );
buf ( n288 , n3604 );
buf ( n289 , n3634 );
buf ( n290 , n3601 );
buf ( n291 , n3637 );
buf ( n292 , n3640 );
buf ( n293 , n3643 );
buf ( n294 , n3646 );
buf ( n295 , n3649 );
buf ( n296 , n3652 );
buf ( n297 , n3655 );
buf ( n298 , n3658 );
buf ( n299 , n3661 );
buf ( n300 , n3664 );
buf ( n301 , n2797 );
buf ( n302 , n2982 );
buf ( n303 , n3200 );
buf ( n304 , n3275 );
buf ( n305 , n3358 );
buf ( n306 , n3395 );
buf ( n307 , n3416 );
buf ( n308 , n3433 );
buf ( n309 , n3467 );
buf ( n310 , n3563 );
buf ( n311 , n3477 );
buf ( n312 , n3374 );
buf ( n313 , n3485 );
buf ( n314 , n3505 );
buf ( n315 , n3571 );
buf ( n316 , n3539 );
buf ( n317 , n3554 );
buf ( n318 , n3582 );
buf ( n319 , n3316 );
buf ( n320 , n3332 );
buf ( n321 , n3665 );
buf ( n322 , n3666 );
buf ( n323 , n3625 );
buf ( n324 , n3669 );
buf ( n325 , n3672 );
buf ( n326 , n3628 );
buf ( n327 , n3678 );
buf ( n328 , n3716 );
buf ( n329 , n3735 );
buf ( n330 , n3721 );
buf ( n331 , n3701 );
buf ( n332 , n3706 );
buf ( n333 , n3711 );
buf ( n334 , n3745 );
buf ( n335 , n3761 );
buf ( n336 , n3726 );
buf ( n337 , n3750 );
buf ( n338 , n3755 );
buf ( n339 , n3682 );
buf ( n340 , n3691 );
buf ( n341 , n3687 );
buf ( n342 , n3696 );
buf ( n343 , n3730 );
buf ( n344 , n3740 );
buf ( n345 , n3766 );
not ( n348 , n27 );
nor ( n349 , n28 , n30 );
nor ( n350 , n29 , n32 );
nand ( n351 , n349 , n350 );
not ( n352 , n351 );
nor ( n353 , n18 , n20 );
nor ( n354 , n19 , n31 );
and ( n355 , n352 , n353 , n354 );
not ( n356 , n6 );
nor ( n357 , n8 , n7 , n9 );
nor ( n358 , n24 , n25 , n26 );
nand ( n359 , n356 , n357 , n358 );
nor ( n360 , n2 , n5 );
nor ( n361 , n12 , n14 );
nor ( n362 , n16 , n17 );
nor ( n363 , n10 , n22 );
nand ( n364 , n360 , n361 , n362 , n363 );
nor ( n365 , n359 , n364 );
nor ( n366 , n13 , n21 );
not ( n367 , n15 );
nand ( n368 , n366 , n367 );
nor ( n369 , n3 , n4 );
nor ( n370 , n11 , n23 );
nand ( n371 , n369 , n370 );
nor ( n372 , n368 , n371 );
nand ( n373 , n355 , n365 , n372 );
nand ( n374 , n373 , n1 );
not ( n375 , n374 );
or ( n376 , n348 , n375 );
nand ( n377 , n355 , n365 , n372 );
not ( n378 , n27 );
nand ( n379 , n377 , n378 , n1 );
nand ( n380 , n376 , n379 );
not ( n381 , n380 );
not ( n382 , n25 );
not ( n383 , n382 );
not ( n384 , n374 );
or ( n385 , n383 , n384 );
nand ( n386 , n1 , n26 );
not ( n387 , n386 );
nor ( n388 , n13 , n21 );
nor ( n389 , n8 , n9 );
not ( n390 , n3 );
nand ( n391 , n388 , n389 , n390 );
nor ( n392 , n19 , n31 );
nand ( n393 , n392 , n367 );
nor ( n394 , n391 , n393 , n351 );
not ( n395 , n364 );
nor ( n396 , n18 , n20 );
nor ( n397 , n6 , n7 );
nor ( n398 , n4 , n24 );
and ( n399 , n396 , n397 , n370 , n398 );
nand ( n400 , n394 , n395 , n399 );
nand ( n401 , n400 , n1 );
not ( n402 , n401 );
or ( n403 , n387 , n402 );
nand ( n404 , n403 , n25 );
nand ( n405 , n385 , n404 );
nand ( n406 , n381 , n405 );
not ( n407 , n406 );
buf ( n408 , n407 );
and ( n409 , n408 , n96 );
not ( n410 , n380 );
not ( n411 , n410 );
not ( n412 , n405 );
not ( n413 , n412 );
nand ( n414 , n411 , n413 );
buf ( n415 , n414 );
not ( n416 , n415 );
and ( n417 , n416 , n93 );
nor ( n418 , n409 , n417 );
not ( n419 , n405 );
nand ( n420 , n419 , n410 );
not ( n421 , n420 );
and ( n422 , n421 , n94 );
not ( n423 , n95 );
not ( n424 , n405 );
not ( n425 , n410 );
nand ( n426 , n424 , n425 );
not ( n427 , n426 );
not ( n428 , n427 );
nor ( n429 , n423 , n428 );
nor ( n430 , n422 , n429 );
nand ( n431 , n418 , n430 );
not ( n432 , n431 );
not ( n433 , n432 );
nand ( n434 , n419 , n410 );
buf ( n435 , n434 );
not ( n436 , n435 );
not ( n437 , n436 );
not ( n438 , n437 );
not ( n439 , n125 );
not ( n440 , n439 );
and ( n441 , n438 , n440 );
not ( n442 , n415 );
not ( n443 , n442 );
not ( n444 , n443 );
and ( n445 , n444 , n124 );
nor ( n446 , n441 , n445 );
not ( n447 , n406 );
not ( n448 , n447 );
not ( n449 , n448 );
and ( n450 , n449 , n126 );
not ( n451 , n127 );
buf ( n452 , n426 );
not ( n453 , n452 );
not ( n454 , n453 );
nor ( n455 , n451 , n454 );
nor ( n456 , n450 , n455 );
nand ( n457 , n446 , n456 );
not ( n458 , n443 );
not ( n459 , n140 );
not ( n460 , n459 );
and ( n461 , n458 , n460 );
and ( n462 , n449 , n141 );
nor ( n463 , n461 , n462 );
not ( n464 , n427 );
not ( n465 , n464 );
and ( n466 , n465 , n142 );
not ( n467 , n139 );
nor ( n468 , n467 , n437 );
nor ( n469 , n466 , n468 );
nand ( n470 , n463 , n469 );
not ( n471 , n407 );
not ( n472 , n471 );
and ( n473 , n472 , n102 );
not ( n474 , n452 );
and ( n475 , n474 , n103 );
nor ( n476 , n473 , n475 );
not ( n477 , n415 );
and ( n478 , n477 , n100 );
and ( n479 , n421 , n101 );
nor ( n480 , n478 , n479 );
nand ( n481 , n476 , n480 );
and ( n482 , n457 , n470 , n481 );
nand ( n483 , n407 , n44 );
not ( n484 , n483 );
and ( n485 , n465 , n43 );
nor ( n486 , n484 , n485 );
not ( n487 , n415 );
nand ( n488 , n487 , n42 );
not ( n489 , n488 );
not ( n490 , n434 );
buf ( n491 , n490 );
and ( n492 , n491 , n41 );
nor ( n493 , n489 , n492 );
nand ( n494 , n486 , n493 );
not ( n495 , n49 );
not ( n496 , n410 );
buf ( n497 , n405 );
nand ( n498 , n496 , n497 );
not ( n499 , n498 );
not ( n500 , n499 );
or ( n501 , n495 , n500 );
nand ( n502 , n419 , n410 );
not ( n503 , n502 );
nand ( n504 , n503 , n50 );
nand ( n505 , n501 , n504 );
not ( n506 , n52 );
not ( n507 , n407 );
or ( n508 , n506 , n507 );
nand ( n509 , n412 , n425 );
not ( n510 , n509 );
nand ( n511 , n510 , n51 );
nand ( n512 , n508 , n511 );
nor ( n513 , n505 , n512 );
not ( n514 , n513 );
nand ( n515 , n494 , n514 );
not ( n516 , n515 );
not ( n517 , n415 );
not ( n518 , n69 );
not ( n519 , n518 );
and ( n520 , n517 , n519 );
not ( n521 , n448 );
and ( n522 , n521 , n72 );
nor ( n523 , n520 , n522 );
and ( n524 , n491 , n70 );
not ( n525 , n71 );
not ( n526 , n427 );
nor ( n527 , n525 , n526 );
nor ( n528 , n524 , n527 );
nand ( n529 , n523 , n528 );
not ( n530 , n464 );
not ( n531 , n75 );
not ( n532 , n531 );
and ( n533 , n530 , n532 );
and ( n534 , n472 , n76 );
nor ( n535 , n533 , n534 );
not ( n536 , n435 );
not ( n537 , n74 );
not ( n538 , n537 );
and ( n539 , n536 , n538 );
and ( n540 , n487 , n73 );
nor ( n541 , n539 , n540 );
nand ( n542 , n535 , n541 );
and ( n543 , n529 , n542 );
not ( n544 , n121 );
not ( n545 , n442 );
or ( n546 , n544 , n545 );
nand ( n547 , n449 , n120 );
nand ( n548 , n546 , n547 );
not ( n549 , n122 );
not ( n550 , n436 );
or ( n551 , n549 , n550 );
nand ( n552 , n474 , n123 );
nand ( n553 , n551 , n552 );
nor ( n554 , n548 , n553 );
not ( n555 , n66 );
not ( n556 , n436 );
or ( n557 , n555 , n556 );
nand ( n558 , n499 , n65 );
nand ( n559 , n557 , n558 );
not ( n560 , n67 );
not ( n561 , n427 );
or ( n562 , n560 , n561 );
nand ( n563 , n447 , n68 );
nand ( n564 , n562 , n563 );
nor ( n565 , n559 , n564 );
nor ( n566 , n554 , n565 );
nand ( n567 , n482 , n516 , n543 , n566 );
not ( n568 , n129 );
not ( n569 , n421 );
or ( n570 , n568 , n569 );
not ( n571 , n415 );
nand ( n572 , n571 , n130 );
nand ( n573 , n570 , n572 );
not ( n574 , n449 );
not ( n575 , n131 );
or ( n576 , n574 , n575 );
not ( n577 , n428 );
nand ( n578 , n577 , n128 );
nand ( n579 , n576 , n578 );
nor ( n580 , n573 , n579 );
not ( n581 , n109 );
not ( n582 , n442 );
or ( n583 , n581 , n582 );
nand ( n584 , n421 , n110 );
nand ( n585 , n583 , n584 );
not ( n586 , n108 );
not ( n587 , n407 );
or ( n588 , n586 , n587 );
nand ( n589 , n474 , n111 );
nand ( n590 , n588 , n589 );
nor ( n591 , n585 , n590 );
nor ( n592 , n580 , n591 );
not ( n593 , n133 );
not ( n594 , n490 );
not ( n595 , n594 );
not ( n596 , n595 );
or ( n597 , n593 , n596 );
nand ( n598 , n416 , n132 );
nand ( n599 , n597 , n598 );
not ( n600 , n134 );
not ( n601 , n453 );
or ( n602 , n600 , n601 );
nand ( n603 , n521 , n135 );
nand ( n604 , n602 , n603 );
nor ( n605 , n599 , n604 );
not ( n606 , n105 );
not ( n607 , n421 );
or ( n608 , n606 , n607 );
nand ( n609 , n477 , n106 );
nand ( n610 , n608 , n609 );
not ( n611 , n104 );
not ( n612 , n465 );
or ( n613 , n611 , n612 );
nand ( n614 , n472 , n107 );
nand ( n615 , n613 , n614 );
nor ( n616 , n610 , n615 );
nor ( n617 , n605 , n616 );
not ( n618 , n57 );
not ( n619 , n477 );
or ( n620 , n618 , n619 );
nand ( n621 , n436 , n58 );
nand ( n622 , n620 , n621 );
not ( n623 , n60 );
not ( n624 , n447 );
or ( n625 , n623 , n624 );
nand ( n626 , n427 , n59 );
nand ( n627 , n625 , n626 );
nor ( n628 , n622 , n627 );
nand ( n629 , n427 , n47 );
nand ( n630 , n490 , n46 );
nand ( n631 , n499 , n48 );
nand ( n632 , n447 , n45 );
nand ( n633 , n629 , n630 , n631 , n632 );
not ( n634 , n633 );
nor ( n635 , n628 , n634 );
and ( n636 , n592 , n617 , n635 );
not ( n637 , n113 );
not ( n638 , n421 );
or ( n639 , n637 , n638 );
nand ( n640 , n571 , n112 );
nand ( n641 , n639 , n640 );
not ( n642 , n115 );
not ( n643 , n428 );
not ( n644 , n643 );
or ( n645 , n642 , n644 );
nand ( n646 , n449 , n114 );
nand ( n647 , n645 , n646 );
nor ( n648 , n641 , n647 );
not ( n649 , n117 );
not ( n650 , n436 );
or ( n651 , n649 , n650 );
nand ( n652 , n416 , n118 );
nand ( n653 , n651 , n652 );
not ( n654 , n116 );
not ( n655 , n521 );
or ( n656 , n654 , n655 );
nand ( n657 , n474 , n119 );
nand ( n658 , n656 , n657 );
nor ( n659 , n653 , n658 );
nor ( n660 , n648 , n659 );
not ( n661 , n660 );
and ( n662 , n421 , n79 );
and ( n663 , n474 , n77 );
nor ( n664 , n662 , n663 );
and ( n665 , n416 , n78 );
not ( n666 , n80 );
nor ( n667 , n666 , n448 );
nor ( n668 , n665 , n667 );
nand ( n669 , n664 , n668 );
not ( n670 , n420 );
not ( n671 , n82 );
not ( n672 , n671 );
and ( n673 , n670 , n672 );
and ( n674 , n487 , n81 );
nor ( n675 , n673 , n674 );
not ( n676 , n428 );
not ( n677 , n83 );
not ( n678 , n677 );
and ( n679 , n676 , n678 );
and ( n680 , n449 , n84 );
nor ( n681 , n679 , n680 );
nand ( n682 , n675 , n681 );
nand ( n683 , n669 , n682 );
nor ( n684 , n661 , n683 );
nand ( n685 , n595 , n54 );
not ( n686 , n526 );
nand ( n687 , n686 , n55 );
nand ( n688 , n407 , n56 );
nand ( n689 , n416 , n53 );
nand ( n690 , n685 , n687 , n688 , n689 );
not ( n691 , n34 );
not ( n692 , n490 );
or ( n693 , n691 , n692 );
nand ( n694 , n499 , n33 );
nand ( n695 , n693 , n694 );
not ( n696 , n35 );
not ( n697 , n427 );
or ( n698 , n696 , n697 );
nand ( n699 , n447 , n36 );
nand ( n700 , n698 , n699 );
nor ( n701 , n695 , n700 );
not ( n702 , n701 );
nand ( n703 , n690 , n702 );
not ( n704 , n415 );
not ( n705 , n62 );
not ( n706 , n705 );
and ( n707 , n704 , n706 );
not ( n708 , n64 );
nor ( n709 , n708 , n448 );
nor ( n710 , n707 , n709 );
not ( n711 , n61 );
nor ( n712 , n711 , n452 );
not ( n713 , n63 );
nor ( n714 , n713 , n435 );
nor ( n715 , n712 , n714 );
nand ( n716 , n710 , n715 );
nand ( n717 , n686 , n39 );
not ( n718 , n717 );
nand ( n719 , n716 , n718 );
nor ( n720 , n703 , n719 );
nand ( n721 , n636 , n684 , n720 );
nor ( n722 , n567 , n721 );
not ( n723 , n86 );
not ( n724 , n571 );
nor ( n725 , n723 , n724 );
and ( n726 , n421 , n85 );
nor ( n727 , n725 , n726 );
not ( n728 , n454 );
not ( n729 , n87 );
not ( n730 , n729 );
and ( n731 , n728 , n730 );
and ( n732 , n449 , n88 );
nor ( n733 , n731 , n732 );
nand ( n734 , n727 , n733 );
and ( n735 , n722 , n734 );
not ( n736 , n90 );
nor ( n737 , n736 , n437 );
not ( n738 , n737 );
not ( n739 , n724 );
nand ( n740 , n739 , n89 );
not ( n741 , n454 );
not ( n742 , n92 );
not ( n743 , n742 );
and ( n744 , n741 , n743 );
and ( n745 , n472 , n91 );
nor ( n746 , n744 , n745 );
nand ( n747 , n738 , n740 , n746 );
buf ( n748 , n747 );
nand ( n749 , n735 , n748 );
not ( n750 , n749 );
not ( n751 , n750 );
or ( n752 , n433 , n751 );
nand ( n753 , n749 , n431 );
nand ( n754 , n752 , n753 );
not ( n755 , n24 );
not ( n756 , n23 );
not ( n757 , n1 );
or ( n758 , n756 , n757 );
nor ( n759 , n6 , n8 );
nor ( n760 , n7 , n9 );
nand ( n761 , n759 , n760 );
not ( n762 , n761 );
not ( n763 , n11 );
and ( n764 , n369 , n763 );
and ( n765 , n353 , n354 );
nand ( n766 , n762 , n764 , n765 );
not ( n767 , n368 );
buf ( n768 , n352 );
and ( n769 , n361 , n362 );
and ( n770 , n360 , n363 );
nand ( n771 , n767 , n768 , n769 , n770 );
or ( n772 , n766 , n771 );
nand ( n773 , n772 , n1 );
nand ( n774 , n758 , n773 );
not ( n775 , n774 );
or ( n776 , n755 , n775 );
not ( n777 , n24 );
nand ( n778 , n777 , n401 );
nand ( n779 , n776 , n778 );
not ( n780 , n401 );
not ( n781 , n26 );
xor ( n782 , n780 , n781 );
nand ( n783 , n779 , n782 );
buf ( n784 , n783 );
nand ( n785 , n784 , n188 );
or ( n786 , n754 , n785 );
nand ( n787 , n784 , n187 );
not ( n788 , n431 );
not ( n789 , n750 );
or ( n790 , n788 , n789 );
not ( n791 , n99 );
not ( n792 , n444 );
or ( n793 , n791 , n792 );
and ( n794 , n595 , n98 );
not ( n795 , n97 );
nor ( n796 , n795 , n448 );
nor ( n797 , n794 , n796 );
nand ( n798 , n793 , n797 );
not ( n799 , n798 );
nand ( n800 , n790 , n799 );
or ( n801 , n787 , n800 );
nand ( n802 , n786 , n801 );
not ( n803 , n802 );
nand ( n804 , n800 , n787 );
not ( n805 , n785 );
nor ( n806 , n798 , n787 );
nor ( n807 , n805 , n806 );
nand ( n808 , n754 , n807 );
nand ( n809 , n804 , n808 );
nor ( n810 , n803 , n809 );
nand ( n811 , n487 , n145 );
nand ( n812 , n421 , n143 );
nand ( n813 , n407 , n144 );
nand ( n814 , n811 , n812 , n813 );
nand ( n815 , n444 , n137 );
nand ( n816 , n595 , n136 );
nand ( n817 , n408 , n138 );
nand ( n818 , n815 , n816 , n817 );
and ( n819 , n784 , n190 );
and ( n820 , n814 , n818 , n819 );
not ( n821 , n819 );
nand ( n822 , n821 , n814 );
nand ( n823 , n784 , n189 );
and ( n824 , n822 , n823 );
nor ( n825 , n820 , n824 );
not ( n826 , n825 );
not ( n827 , n28 );
not ( n828 , n6 );
nor ( n829 , n2 , n8 );
nor ( n830 , n4 , n11 );
nand ( n831 , n828 , n829 , n830 );
nor ( n832 , n3 , n7 );
nor ( n833 , n5 , n9 );
nand ( n834 , n832 , n833 );
nor ( n835 , n831 , n834 );
not ( n836 , n10 );
and ( n837 , n835 , n836 );
not ( n838 , n13 );
nand ( n839 , n837 , n838 );
nor ( n840 , n839 , n12 );
not ( n841 , n14 );
and ( n842 , n840 , n841 );
not ( n843 , n16 );
nand ( n844 , n842 , n843 );
nor ( n845 , n844 , n17 );
not ( n846 , n19 );
and ( n847 , n353 , n367 , n846 );
and ( n848 , n845 , n847 );
not ( n849 , n29 );
nand ( n850 , n848 , n849 );
nor ( n851 , n850 , n32 );
nand ( n852 , n827 , n851 );
not ( n853 , n852 );
not ( n854 , n30 );
nand ( n855 , n853 , n854 );
nor ( n856 , n855 , n31 );
buf ( n857 , n856 );
not ( n858 , n31 );
not ( n859 , n855 );
or ( n860 , n858 , n859 );
nand ( n861 , n860 , n1 );
or ( n862 , n857 , n861 );
not ( n863 , n1 );
nand ( n864 , n863 , n31 );
nand ( n865 , n862 , n864 );
not ( n866 , n865 );
buf ( n867 , n866 );
not ( n868 , n851 );
and ( n869 , n868 , n28 );
not ( n870 , n1 );
nor ( n871 , n869 , n870 );
not ( n872 , n871 );
not ( n873 , n853 );
not ( n874 , n873 );
or ( n875 , n872 , n874 );
not ( n876 , n1 );
nand ( n877 , n876 , n28 );
nand ( n878 , n875 , n877 );
not ( n879 , n878 );
nor ( n880 , n867 , n879 );
not ( n881 , n849 );
not ( n882 , n876 );
or ( n883 , n881 , n882 );
buf ( n884 , n848 );
or ( n885 , n884 , n849 );
buf ( n886 , n850 );
nand ( n887 , n885 , n886 );
nand ( n888 , n887 , n1 );
nand ( n889 , n883 , n888 );
buf ( n890 , n889 );
not ( n891 , n868 );
and ( n892 , n886 , n32 );
not ( n893 , n1 );
nor ( n894 , n892 , n893 );
not ( n895 , n894 );
or ( n896 , n891 , n895 );
nand ( n897 , n876 , n32 );
nand ( n898 , n896 , n897 );
nand ( n899 , n161 , n898 );
nor ( n900 , n890 , n899 );
nand ( n901 , n880 , n900 );
not ( n902 , n855 );
and ( n903 , n852 , n30 );
nor ( n904 , n903 , n870 );
not ( n905 , n904 );
or ( n906 , n902 , n905 );
nand ( n907 , n876 , n30 );
nand ( n908 , n906 , n907 );
buf ( n909 , n908 );
nand ( n910 , n909 , n158 );
nand ( n911 , n826 , n901 , n910 );
nor ( n912 , n810 , n911 );
not ( n913 , n912 );
nand ( n914 , n784 , n194 );
not ( n915 , n914 );
not ( n916 , n915 );
not ( n917 , n457 );
not ( n918 , n917 );
nand ( n919 , n566 , n543 );
not ( n920 , n683 );
not ( n921 , n719 );
nand ( n922 , n920 , n921 );
nor ( n923 , n919 , n922 );
nand ( n924 , n488 , n483 );
not ( n925 , n924 );
not ( n926 , n41 );
not ( n927 , n491 );
or ( n928 , n926 , n927 );
not ( n929 , n464 );
nand ( n930 , n929 , n43 );
nand ( n931 , n928 , n930 );
not ( n932 , n931 );
and ( n933 , n925 , n932 );
nand ( n934 , n687 , n685 );
nand ( n935 , n689 , n688 );
nor ( n936 , n934 , n935 );
nor ( n937 , n933 , n936 );
nand ( n938 , n937 , n592 , n660 );
not ( n939 , n505 );
not ( n940 , n512 );
and ( n941 , n939 , n940 );
nor ( n942 , n941 , n701 );
nand ( n943 , n942 , n635 );
nor ( n944 , n938 , n943 );
nand ( n945 , n923 , n944 );
not ( n946 , n945 );
buf ( n947 , n617 );
nand ( n948 , n946 , n947 );
not ( n949 , n481 );
nor ( n950 , n948 , n949 );
buf ( n951 , n470 );
nand ( n952 , n950 , n951 );
not ( n953 , n952 );
or ( n954 , n918 , n953 );
not ( n955 , n722 );
nand ( n956 , n954 , n955 );
not ( n957 , n956 );
or ( n958 , n916 , n957 );
nor ( n959 , n950 , n951 );
not ( n960 , n959 );
nand ( n961 , n960 , n952 );
buf ( n962 , n784 );
nand ( n963 , n962 , n193 );
not ( n964 , n963 );
nand ( n965 , n961 , n964 );
nand ( n966 , n958 , n965 );
nand ( n967 , n784 , n191 );
not ( n968 , n967 );
not ( n969 , n968 );
xnor ( n970 , n735 , n748 );
not ( n971 , n970 );
or ( n972 , n969 , n971 );
nand ( n973 , n784 , n192 );
not ( n974 , n973 );
and ( n975 , n722 , n734 );
not ( n976 , n975 );
not ( n977 , n734 );
nand ( n978 , n977 , n955 );
nand ( n979 , n976 , n978 );
nand ( n980 , n974 , n979 );
nand ( n981 , n972 , n980 );
buf ( n982 , n981 );
nor ( n983 , n966 , n982 );
nor ( n984 , n983 , n809 );
not ( n985 , n984 );
not ( n986 , n634 );
not ( n987 , n718 );
not ( n988 , n987 );
or ( n989 , n986 , n988 );
not ( n990 , n717 );
not ( n991 , n990 );
nor ( n992 , n991 , n634 );
not ( n993 , n992 );
nand ( n994 , n989 , n993 );
not ( n995 , n994 );
not ( n996 , n995 );
and ( n997 , n783 , n168 );
not ( n998 , n783 );
not ( n999 , n762 );
nand ( n1000 , n999 , n1 );
not ( n1001 , n2 );
and ( n1002 , n1000 , n1001 );
not ( n1003 , n1000 );
and ( n1004 , n1003 , n2 );
nor ( n1005 , n1002 , n1004 );
and ( n1006 , n998 , n1005 );
or ( n1007 , n997 , n1006 );
not ( n1008 , n1007 );
not ( n1009 , n1008 );
and ( n1010 , n996 , n1009 );
nor ( n1011 , n514 , n992 );
not ( n1012 , n1011 );
nand ( n1013 , n992 , n514 );
nand ( n1014 , n1012 , n1013 );
not ( n1015 , n784 );
not ( n1016 , n1001 );
not ( n1017 , n762 );
or ( n1018 , n1016 , n1017 );
nand ( n1019 , n1018 , n1 );
buf ( n1020 , n1019 );
and ( n1021 , n1020 , n390 );
not ( n1022 , n1020 );
and ( n1023 , n1022 , n3 );
nor ( n1024 , n1021 , n1023 );
not ( n1025 , n1024 );
and ( n1026 , n1015 , n1025 );
not ( n1027 , n167 );
and ( n1028 , n784 , n1027 );
nor ( n1029 , n1026 , n1028 );
and ( n1030 , n1014 , n1029 );
nor ( n1031 , n1010 , n1030 );
not ( n1032 , n1031 );
not ( n1033 , n415 );
not ( n1034 , n155 );
not ( n1035 , n1034 );
and ( n1036 , n1033 , n1035 );
not ( n1037 , n156 );
nor ( n1038 , n448 , n1037 );
nor ( n1039 , n1036 , n1038 );
not ( n1040 , n452 );
not ( n1041 , n154 );
not ( n1042 , n1041 );
and ( n1043 , n1040 , n1042 );
not ( n1044 , n157 );
nor ( n1045 , n594 , n1044 );
nor ( n1046 , n1043 , n1045 );
nand ( n1047 , n1039 , n1046 );
not ( n1048 , n1 );
nor ( n1049 , n397 , n1048 );
and ( n1050 , n1049 , n8 );
not ( n1051 , n1049 );
not ( n1052 , n8 );
and ( n1053 , n1051 , n1052 );
nor ( n1054 , n1050 , n1053 );
or ( n1055 , n784 , n1054 );
not ( n1056 , n170 );
nand ( n1057 , n1056 , n783 );
nand ( n1058 , n1055 , n1057 );
and ( n1059 , n1047 , n1058 );
not ( n1060 , n1059 );
not ( n1061 , n1047 );
not ( n1062 , n1058 );
nand ( n1063 , n1061 , n1062 );
nand ( n1064 , n1060 , n1063 );
not ( n1065 , n1064 );
not ( n1066 , n502 );
not ( n1067 , n148 );
not ( n1068 , n1067 );
and ( n1069 , n1066 , n1068 );
and ( n1070 , n499 , n147 );
nor ( n1071 , n1069 , n1070 );
not ( n1072 , n149 );
nor ( n1073 , n1072 , n448 );
not ( n1074 , n146 );
nor ( n1075 , n1074 , n509 );
nor ( n1076 , n1073 , n1075 );
nand ( n1077 , n1071 , n1076 );
not ( n1078 , n1077 );
and ( n1079 , n779 , n782 );
and ( n1080 , n1079 , n6 );
not ( n1081 , n1079 );
and ( n1082 , n1081 , n172 );
nor ( n1083 , n1080 , n1082 );
not ( n1084 , n1083 );
nand ( n1085 , n1078 , n1084 );
not ( n1086 , n1085 );
not ( n1087 , n151 );
not ( n1088 , n447 );
or ( n1089 , n1087 , n1088 );
nand ( n1090 , n510 , n150 );
nand ( n1091 , n1089 , n1090 );
not ( n1092 , n153 );
not ( n1093 , n499 );
or ( n1094 , n1092 , n1093 );
not ( n1095 , n502 );
nand ( n1096 , n1095 , n152 );
nand ( n1097 , n1094 , n1096 );
nor ( n1098 , n1091 , n1097 );
not ( n1099 , n1098 );
not ( n1100 , n1079 );
not ( n1101 , n7 );
not ( n1102 , n1101 );
not ( n1103 , n1049 );
not ( n1104 , n1103 );
or ( n1105 , n1102 , n1104 );
nand ( n1106 , n1 , n6 , n7 );
nand ( n1107 , n1105 , n1106 );
not ( n1108 , n1107 );
or ( n1109 , n1100 , n1108 );
not ( n1110 , n171 );
nand ( n1111 , n1110 , n783 );
nand ( n1112 , n1109 , n1111 );
not ( n1113 , n1112 );
or ( n1114 , n1099 , n1113 );
or ( n1115 , n1098 , n1112 );
nand ( n1116 , n1114 , n1115 );
not ( n1117 , n1116 );
or ( n1118 , n1086 , n1117 );
not ( n1119 , n1113 );
not ( n1120 , n1099 );
not ( n1121 , n1120 );
or ( n1122 , n1119 , n1121 );
not ( n1123 , n1112 );
not ( n1124 , n1099 );
or ( n1125 , n1123 , n1124 );
nand ( n1126 , n1077 , n1083 );
nand ( n1127 , n1125 , n1126 );
nand ( n1128 , n1122 , n1127 );
nand ( n1129 , n1118 , n1128 );
nand ( n1130 , n1065 , n1129 );
not ( n1131 , n1059 );
nand ( n1132 , n1130 , n1131 );
not ( n1133 , n987 );
not ( n1134 , n37 );
not ( n1135 , n1134 );
not ( n1136 , n442 );
or ( n1137 , n1135 , n1136 );
not ( n1138 , n40 );
not ( n1139 , n1138 );
buf ( n1140 , n497 );
not ( n1141 , n1140 );
or ( n1142 , n1139 , n1141 );
or ( n1143 , n38 , n1140 );
nand ( n1144 , n1142 , n1143 );
nand ( n1145 , n1144 , n410 );
nand ( n1146 , n1137 , n1145 );
nor ( n1147 , n1133 , n1146 );
buf ( n1148 , n1079 );
or ( n1149 , n1148 , n169 );
nand ( n1150 , n1 , n8 );
not ( n1151 , n1150 );
not ( n1152 , n1103 );
or ( n1153 , n1151 , n1152 );
nand ( n1154 , n1153 , n9 );
not ( n1155 , n1 );
not ( n1156 , n9 );
and ( n1157 , n1155 , n1156 );
nor ( n1158 , n1157 , n762 );
nand ( n1159 , n1154 , n1158 );
not ( n1160 , n1159 );
not ( n1161 , n1160 );
nand ( n1162 , n1161 , n1079 );
nand ( n1163 , n1149 , n1162 );
nor ( n1164 , n1147 , n1163 );
not ( n1165 , n1164 );
nand ( n1166 , n1147 , n1163 );
nand ( n1167 , n1165 , n1166 );
not ( n1168 , n1167 );
and ( n1169 , n1132 , n1168 );
not ( n1170 , n1169 );
or ( n1171 , n1032 , n1170 );
not ( n1172 , n702 );
not ( n1173 , n1172 );
not ( n1174 , n1013 );
or ( n1175 , n1173 , n1174 );
nand ( n1176 , n992 , n942 );
nand ( n1177 , n1175 , n1176 );
not ( n1178 , n1177 );
not ( n1179 , n390 );
not ( n1180 , n1019 );
or ( n1181 , n1179 , n1180 );
nand ( n1182 , n1181 , n1 );
not ( n1183 , n5 );
and ( n1184 , n1182 , n1183 );
not ( n1185 , n1182 );
and ( n1186 , n1185 , n5 );
nor ( n1187 , n1184 , n1186 );
and ( n1188 , n1148 , n1187 );
not ( n1189 , n1148 );
and ( n1190 , n1189 , n166 );
nor ( n1191 , n1188 , n1190 );
not ( n1192 , n1191 );
not ( n1193 , n1192 );
and ( n1194 , n1178 , n1193 );
not ( n1195 , n1014 );
not ( n1196 , n1029 );
and ( n1197 , n1195 , n1196 );
nor ( n1198 , n1194 , n1197 );
and ( n1199 , n1128 , n1131 );
not ( n1200 , n1063 );
nor ( n1201 , n1199 , n1164 , n1200 );
nor ( n1202 , n994 , n1007 );
not ( n1203 , n1166 );
or ( n1204 , n1201 , n1202 , n1203 );
nand ( n1205 , n1204 , n1031 );
nand ( n1206 , n1198 , n1205 );
not ( n1207 , n1176 );
not ( n1208 , n494 );
not ( n1209 , n1208 );
or ( n1210 , n1207 , n1209 );
not ( n1211 , n1176 );
not ( n1212 , n1208 );
nand ( n1213 , n1211 , n1212 );
nand ( n1214 , n1210 , n1213 );
not ( n1215 , n1214 );
not ( n1216 , n1215 );
not ( n1217 , n1183 );
not ( n1218 , n1182 );
or ( n1219 , n1217 , n1218 );
nand ( n1220 , n1219 , n1 );
not ( n1221 , n1220 );
not ( n1222 , n4 );
and ( n1223 , n1221 , n1222 );
and ( n1224 , n1220 , n4 );
nor ( n1225 , n1223 , n1224 );
and ( n1226 , n1148 , n1225 );
not ( n1227 , n1148 );
not ( n1228 , n165 );
and ( n1229 , n1227 , n1228 );
or ( n1230 , n1226 , n1229 );
not ( n1231 , n1230 );
or ( n1232 , n1216 , n1231 );
buf ( n1233 , n628 );
not ( n1234 , n1233 );
not ( n1235 , n1213 );
or ( n1236 , n1234 , n1235 );
nor ( n1237 , n1208 , n1233 );
nand ( n1238 , n1211 , n1237 );
nand ( n1239 , n1236 , n1238 );
not ( n1240 , n1148 );
not ( n1241 , n762 );
nand ( n1242 , n369 , n360 );
or ( n1243 , n1241 , n1242 );
and ( n1244 , n1 , n11 );
nand ( n1245 , n1243 , n1244 );
not ( n1246 , n835 );
nand ( n1247 , n876 , n763 );
nand ( n1248 , n1245 , n1246 , n1247 );
not ( n1249 , n1248 );
or ( n1250 , n1240 , n1249 );
not ( n1251 , n164 );
nand ( n1252 , n1251 , n784 );
nand ( n1253 , n1250 , n1252 );
not ( n1254 , n1253 );
or ( n1255 , n1239 , n1254 );
nand ( n1256 , n1232 , n1255 );
nor ( n1257 , n1206 , n1256 );
nand ( n1258 , n1171 , n1257 );
not ( n1259 , n1256 );
not ( n1260 , n1192 );
not ( n1261 , n1177 );
or ( n1262 , n1260 , n1261 );
not ( n1263 , n1230 );
nand ( n1264 , n1214 , n1263 );
nand ( n1265 , n1262 , n1264 );
and ( n1266 , n1259 , n1265 );
not ( n1267 , n690 );
not ( n1268 , n1267 );
not ( n1269 , n1268 );
not ( n1270 , n1238 );
or ( n1271 , n1269 , n1270 );
not ( n1272 , n1238 );
nand ( n1273 , n1272 , n1267 );
nand ( n1274 , n1271 , n1273 );
not ( n1275 , n10 );
not ( n1276 , n876 );
or ( n1277 , n1275 , n1276 );
and ( n1278 , n1246 , n10 );
not ( n1279 , n1 );
nor ( n1280 , n1278 , n1279 );
not ( n1281 , n837 );
nand ( n1282 , n1280 , n1281 );
nand ( n1283 , n1277 , n1282 );
and ( n1284 , n1148 , n1283 );
not ( n1285 , n1148 );
and ( n1286 , n1285 , n163 );
or ( n1287 , n1284 , n1286 );
not ( n1288 , n1287 );
or ( n1289 , n1274 , n1288 );
not ( n1290 , n1239 );
or ( n1291 , n1290 , n1253 );
nand ( n1292 , n1289 , n1291 );
nor ( n1293 , n1266 , n1292 );
and ( n1294 , n1258 , n1293 );
and ( n1295 , n784 , n162 );
not ( n1296 , n784 );
not ( n1297 , n13 );
not ( n1298 , n1 );
not ( n1299 , n1298 );
or ( n1300 , n1297 , n1299 );
buf ( n1301 , n839 );
and ( n1302 , n1281 , n13 );
nor ( n1303 , n1302 , n1048 );
nand ( n1304 , n1301 , n1303 );
nand ( n1305 , n1300 , n1304 );
not ( n1306 , n1305 );
not ( n1307 , n1306 );
and ( n1308 , n1296 , n1307 );
nor ( n1309 , n1295 , n1308 );
not ( n1310 , n1309 );
not ( n1311 , n1268 );
not ( n1312 , n1272 );
or ( n1313 , n1311 , n1312 );
buf ( n1314 , n716 );
not ( n1315 , n1314 );
nand ( n1316 , n1313 , n1315 );
nand ( n1317 , n937 , n921 );
nor ( n1318 , n1317 , n943 );
not ( n1319 , n1318 );
nand ( n1320 , n1316 , n1319 );
not ( n1321 , n1320 );
not ( n1322 , n1321 );
or ( n1323 , n1310 , n1322 );
not ( n1324 , n565 );
and ( n1325 , n1318 , n1324 );
not ( n1326 , n1325 );
not ( n1327 , n1324 );
nand ( n1328 , n1319 , n1327 );
nand ( n1329 , n1326 , n1328 );
not ( n1330 , n1329 );
and ( n1331 , n1301 , n12 );
nor ( n1332 , n1331 , n893 );
not ( n1333 , n1332 );
not ( n1334 , n840 );
not ( n1335 , n1334 );
or ( n1336 , n1333 , n1335 );
not ( n1337 , n1 );
nand ( n1338 , n1337 , n12 );
nand ( n1339 , n1336 , n1338 );
not ( n1340 , n1339 );
not ( n1341 , n1340 );
not ( n1342 , n1148 );
or ( n1343 , n1341 , n1342 );
not ( n1344 , n186 );
nand ( n1345 , n1344 , n784 );
nand ( n1346 , n1343 , n1345 );
not ( n1347 , n1346 );
not ( n1348 , n1347 );
and ( n1349 , n1330 , n1348 );
and ( n1350 , n1274 , n1288 );
nor ( n1351 , n1349 , n1350 );
nand ( n1352 , n1323 , n1351 );
nor ( n1353 , n1294 , n1352 );
not ( n1354 , n842 );
and ( n1355 , n1334 , n14 );
nor ( n1356 , n1355 , n876 );
nand ( n1357 , n1354 , n1356 );
nand ( n1358 , n876 , n14 );
and ( n1359 , n1357 , n1358 );
not ( n1360 , n1359 );
not ( n1361 , n1148 );
or ( n1362 , n1360 , n1361 );
not ( n1363 , n185 );
nand ( n1364 , n1363 , n784 );
nand ( n1365 , n1362 , n1364 );
not ( n1366 , n1365 );
not ( n1367 , n1366 );
buf ( n1368 , n1325 );
not ( n1369 , n1368 );
buf ( n1370 , n542 );
not ( n1371 , n1370 );
not ( n1372 , n1371 );
and ( n1373 , n1369 , n1372 );
and ( n1374 , n1368 , n1371 );
nor ( n1375 , n1373 , n1374 );
not ( n1376 , n1375 );
or ( n1377 , n1367 , n1376 );
nand ( n1378 , n1325 , n543 );
not ( n1379 , n1370 );
not ( n1380 , n1325 );
or ( n1381 , n1379 , n1380 );
not ( n1382 , n529 );
nand ( n1383 , n1381 , n1382 );
and ( n1384 , n1378 , n1383 );
not ( n1385 , n1384 );
and ( n1386 , n784 , n184 );
not ( n1387 , n784 );
not ( n1388 , n16 );
not ( n1389 , n876 );
or ( n1390 , n1388 , n1389 );
buf ( n1391 , n844 );
and ( n1392 , n1354 , n16 );
nor ( n1393 , n1392 , n876 );
nand ( n1394 , n1391 , n1393 );
nand ( n1395 , n1390 , n1394 );
and ( n1396 , n1387 , n1395 );
nor ( n1397 , n1386 , n1396 );
not ( n1398 , n1397 );
nand ( n1399 , n1385 , n1398 );
nand ( n1400 , n1377 , n1399 );
or ( n1401 , n1353 , n1400 );
nand ( n1402 , n1384 , n1397 );
not ( n1403 , n1402 );
not ( n1404 , n1375 );
nand ( n1405 , n1404 , n1365 );
not ( n1406 , n1405 );
or ( n1407 , n1403 , n1406 );
nand ( n1408 , n1407 , n1399 );
nand ( n1409 , n1401 , n1408 );
buf ( n1410 , n648 );
not ( n1411 , n1410 );
not ( n1412 , n937 );
not ( n1413 , n543 );
nor ( n1414 , n1412 , n1413 );
nand ( n1415 , n1324 , n942 );
not ( n1416 , n635 );
nor ( n1417 , n1415 , n1416 );
not ( n1418 , n922 );
nand ( n1419 , n1414 , n1417 , n1418 );
not ( n1420 , n1419 );
buf ( n1421 , n554 );
not ( n1422 , n1421 );
nand ( n1423 , n1420 , n1422 );
not ( n1424 , n1423 );
not ( n1425 , n659 );
nand ( n1426 , n1424 , n1425 );
not ( n1427 , n1426 );
or ( n1428 , n1411 , n1427 );
not ( n1429 , n566 );
nor ( n1430 , n1429 , n1416 );
nor ( n1431 , n1413 , n719 );
nor ( n1432 , n515 , n703 );
and ( n1433 , n1430 , n1431 , n1432 , n684 );
not ( n1434 , n1433 );
nand ( n1435 , n1428 , n1434 );
not ( n1436 , n201 );
and ( n1437 , n962 , n1436 );
not ( n1438 , n962 );
buf ( n1439 , n845 );
nand ( n1440 , n1439 , n367 );
not ( n1441 , n1440 );
nand ( n1442 , n1441 , n846 );
not ( n1443 , n1442 );
not ( n1444 , n18 );
nand ( n1445 , n1443 , n1444 );
and ( n1446 , n1445 , n20 );
not ( n1447 , n884 );
nand ( n1448 , n1447 , n1 );
nor ( n1449 , n1446 , n1448 );
not ( n1450 , n20 );
nor ( n1451 , n1450 , n1 );
nor ( n1452 , n1449 , n1451 );
and ( n1453 , n1438 , n1452 );
nor ( n1454 , n1437 , n1453 );
nand ( n1455 , n1435 , n1454 );
nand ( n1456 , n784 , n196 );
not ( n1457 , n1456 );
buf ( n1458 , n616 );
not ( n1459 , n1458 );
not ( n1460 , n945 );
not ( n1461 , n605 );
nand ( n1462 , n1460 , n1461 );
not ( n1463 , n1462 );
or ( n1464 , n1459 , n1463 );
nand ( n1465 , n1464 , n948 );
nand ( n1466 , n1457 , n1465 );
not ( n1467 , n1433 );
buf ( n1468 , n591 );
nand ( n1469 , n1467 , n1468 );
not ( n1470 , n1468 );
nand ( n1471 , n1470 , n1433 );
nand ( n1472 , n1469 , n1471 );
and ( n1473 , n889 , n1148 );
not ( n1474 , n202 );
and ( n1475 , n962 , n1474 );
nor ( n1476 , n1473 , n1475 );
nand ( n1477 , n1472 , n1476 );
not ( n1478 , n1419 );
not ( n1479 , n1478 );
nand ( n1480 , n1479 , n1421 );
nand ( n1481 , n1480 , n1423 );
or ( n1482 , n1441 , n846 );
nand ( n1483 , n1482 , n1442 );
and ( n1484 , n1 , n1483 );
not ( n1485 , n1 );
and ( n1486 , n1485 , n846 );
or ( n1487 , n1484 , n1486 );
and ( n1488 , n1487 , n1148 );
nor ( n1489 , n1148 , n199 );
nor ( n1490 , n1488 , n1489 );
nand ( n1491 , n1481 , n1490 );
and ( n1492 , n1477 , n1491 );
nand ( n1493 , n1455 , n1466 , n1492 );
or ( n1494 , n1424 , n1425 );
nand ( n1495 , n1494 , n1426 );
and ( n1496 , n962 , n200 );
not ( n1497 , n962 );
nand ( n1498 , n1442 , n1 );
and ( n1499 , n1498 , n1444 );
not ( n1500 , n1498 );
and ( n1501 , n1500 , n18 );
nor ( n1502 , n1499 , n1501 );
and ( n1503 , n1497 , n1502 );
nor ( n1504 , n1496 , n1503 );
not ( n1505 , n1504 );
nand ( n1506 , n1495 , n1505 );
nand ( n1507 , n784 , n198 );
not ( n1508 , n1507 );
not ( n1509 , n580 );
not ( n1510 , n1509 );
not ( n1511 , n1510 );
not ( n1512 , n1471 );
or ( n1513 , n1511 , n1512 );
not ( n1514 , n945 );
not ( n1515 , n1514 );
nand ( n1516 , n1513 , n1515 );
nand ( n1517 , n1508 , n1516 );
nand ( n1518 , n784 , n197 );
not ( n1519 , n1518 );
or ( n1520 , n1514 , n1461 );
nand ( n1521 , n1520 , n1462 );
nand ( n1522 , n1519 , n1521 );
nand ( n1523 , n784 , n195 );
not ( n1524 , n1523 );
nand ( n1525 , n949 , n1524 );
and ( n1526 , n948 , n1525 );
not ( n1527 , n948 );
not ( n1528 , n949 );
nand ( n1529 , n1528 , n1524 );
and ( n1530 , n1527 , n1529 );
or ( n1531 , n1526 , n1530 );
nand ( n1532 , n1506 , n1517 , n1522 , n1531 );
nor ( n1533 , n1493 , n1532 );
not ( n1534 , n1148 );
not ( n1535 , n367 );
not ( n1536 , n1 );
and ( n1537 , n1535 , n1536 );
not ( n1538 , n1439 );
and ( n1539 , n1538 , n15 );
nor ( n1540 , n1539 , n1279 );
and ( n1541 , n1440 , n1540 );
nor ( n1542 , n1537 , n1541 );
not ( n1543 , n1542 );
or ( n1544 , n1534 , n1543 );
not ( n1545 , n182 );
nand ( n1546 , n1545 , n784 );
nand ( n1547 , n1544 , n1546 );
not ( n1548 , n1547 );
not ( n1549 , n1478 );
buf ( n1550 , n682 );
buf ( n1551 , n1550 );
not ( n1552 , n1551 );
not ( n1553 , n1378 );
not ( n1554 , n1553 );
or ( n1555 , n1552 , n1554 );
buf ( n1556 , n669 );
not ( n1557 , n1556 );
nand ( n1558 , n1555 , n1557 );
nand ( n1559 , n1549 , n1558 );
nand ( n1560 , n1548 , n1559 );
and ( n1561 , n784 , n183 );
not ( n1562 , n784 );
not ( n1563 , n1538 );
and ( n1564 , n1391 , n17 );
nor ( n1565 , n1564 , n863 );
not ( n1566 , n1565 );
or ( n1567 , n1563 , n1566 );
not ( n1568 , n1 );
nand ( n1569 , n1568 , n17 );
nand ( n1570 , n1567 , n1569 );
and ( n1571 , n1562 , n1570 );
nor ( n1572 , n1561 , n1571 );
not ( n1573 , n1572 );
xnor ( n1574 , n1553 , n1551 );
nand ( n1575 , n1573 , n1574 );
and ( n1576 , n1560 , n1575 );
not ( n1577 , n1309 );
not ( n1578 , n1577 );
not ( n1579 , n1320 );
or ( n1580 , n1578 , n1579 );
nand ( n1581 , n1580 , n1346 );
nor ( n1582 , n1346 , n1309 );
not ( n1583 , n1582 );
not ( n1584 , n1320 );
or ( n1585 , n1583 , n1584 );
not ( n1586 , n1329 );
nand ( n1587 , n1585 , n1586 );
nand ( n1588 , n1581 , n1587 );
not ( n1589 , n1588 );
nand ( n1590 , n1589 , n1408 );
nand ( n1591 , n1409 , n1533 , n1576 , n1590 );
not ( n1592 , n1559 );
nand ( n1593 , n1592 , n1547 );
not ( n1594 , n1574 );
nand ( n1595 , n1594 , n1572 );
nand ( n1596 , n1593 , n1595 );
and ( n1597 , n1533 , n1596 , n1560 );
not ( n1598 , n948 );
not ( n1599 , n1528 );
and ( n1600 , n1598 , n1599 );
and ( n1601 , n948 , n1528 );
nor ( n1602 , n1600 , n1601 );
not ( n1603 , n1602 );
nand ( n1604 , n1603 , n1523 );
nand ( n1605 , n808 , n804 , n1604 );
nor ( n1606 , n1597 , n1605 );
not ( n1607 , n1507 );
nor ( n1608 , n1607 , n1516 );
not ( n1609 , n1608 );
or ( n1610 , n1472 , n1476 );
nand ( n1611 , n1609 , n1610 );
not ( n1612 , n1456 );
not ( n1613 , n1465 );
not ( n1614 , n1613 );
or ( n1615 , n1612 , n1614 );
not ( n1616 , n1521 );
nand ( n1617 , n1616 , n1518 );
nand ( n1618 , n1615 , n1617 );
nor ( n1619 , n1611 , n1618 );
or ( n1620 , n1505 , n1495 );
or ( n1621 , n1481 , n1490 );
nand ( n1622 , n1620 , n1621 );
nand ( n1623 , n1455 , n1622 , n1506 );
nor ( n1624 , n1435 , n1454 );
not ( n1625 , n1624 );
nand ( n1626 , n1619 , n1623 , n1625 );
not ( n1627 , n1477 );
not ( n1628 , n1516 );
nand ( n1629 , n1628 , n1507 );
nand ( n1630 , n1627 , n1629 );
nand ( n1631 , n1630 , n1517 , n1522 );
not ( n1632 , n1618 );
and ( n1633 , n1631 , n1632 );
not ( n1634 , n1524 );
not ( n1635 , n1602 );
or ( n1636 , n1634 , n1635 );
nand ( n1637 , n1636 , n1466 );
nor ( n1638 , n1633 , n1637 );
nand ( n1639 , n1626 , n1638 );
nand ( n1640 , n1591 , n1606 , n1639 );
nand ( n1641 , n985 , n1640 );
not ( n1642 , n970 );
nand ( n1643 , n1642 , n967 );
and ( n1644 , n981 , n1643 );
not ( n1645 , n1644 );
not ( n1646 , n966 );
not ( n1647 , n1646 );
nor ( n1648 , n961 , n964 );
not ( n1649 , n1648 );
or ( n1650 , n1647 , n1649 );
not ( n1651 , n956 );
nand ( n1652 , n1651 , n914 );
not ( n1653 , n979 );
nand ( n1654 , n1653 , n973 );
and ( n1655 , n1652 , n1643 , n1654 );
nand ( n1656 , n1650 , n1655 );
nand ( n1657 , n1645 , n1656 );
nand ( n1658 , n1641 , n1657 );
not ( n1659 , n1658 );
or ( n1660 , n913 , n1659 );
not ( n1661 , n890 );
nor ( n1662 , n1661 , n899 );
nand ( n1663 , n880 , n1662 );
not ( n1664 , n823 );
not ( n1665 , n818 );
or ( n1666 , n1664 , n1665 );
not ( n1667 , n814 );
nand ( n1668 , n1667 , n819 );
nand ( n1669 , n1666 , n1668 );
nand ( n1670 , n1669 , n819 );
and ( n1671 , n1663 , n910 , n1670 );
and ( n1672 , n1641 , n1657 , n1671 );
not ( n1673 , n1671 );
not ( n1674 , n810 );
or ( n1675 , n1673 , n1674 );
and ( n1676 , n1671 , n825 );
not ( n1677 , n1670 );
not ( n1678 , n1677 );
not ( n1679 , n910 );
or ( n1680 , n1678 , n1679 );
not ( n1681 , n1663 );
nand ( n1682 , n1680 , n1681 );
and ( n1683 , n1682 , n901 );
nor ( n1684 , n1676 , n1683 );
nand ( n1685 , n1675 , n1684 );
nor ( n1686 , n1672 , n1685 );
nand ( n1687 , n1660 , n1686 );
not ( n1688 , n810 );
not ( n1689 , n818 );
or ( n1690 , n1689 , n814 );
nand ( n1691 , n1690 , n825 );
nand ( n1692 , n1688 , n1691 );
buf ( n1693 , n867 );
not ( n1694 , n1693 );
nand ( n1695 , n1694 , n879 );
not ( n1696 , n1695 );
not ( n1697 , n161 );
nor ( n1698 , n898 , n890 , n1697 );
nand ( n1699 , n1696 , n1698 );
nor ( n1700 , n1692 , n1699 );
and ( n1701 , n1658 , n1700 );
nand ( n1702 , n702 , n1191 );
nor ( n1703 , n494 , n1230 );
not ( n1704 , n1703 );
nand ( n1705 , n494 , n1230 );
nand ( n1706 , n1704 , n1705 );
xor ( n1707 , n1702 , n1706 );
not ( n1708 , n1254 );
not ( n1709 , n1233 );
or ( n1710 , n1708 , n1709 );
not ( n1711 , n1233 );
nand ( n1712 , n1711 , n1253 );
nand ( n1713 , n1710 , n1712 );
not ( n1714 , n1713 );
and ( n1715 , n1705 , n1714 );
not ( n1716 , n1705 );
and ( n1717 , n1716 , n1713 );
or ( n1718 , n1715 , n1717 );
or ( n1719 , n1550 , n1572 );
nand ( n1720 , n1550 , n1572 );
nand ( n1721 , n1719 , n1720 );
not ( n1722 , n1721 );
nand ( n1723 , n529 , n1397 );
not ( n1724 , n1723 );
and ( n1725 , n1722 , n1724 );
and ( n1726 , n1721 , n1723 );
nor ( n1727 , n1725 , n1726 );
and ( n1728 , n1707 , n1718 , n1727 );
not ( n1729 , n915 );
not ( n1730 , n917 );
or ( n1731 , n1729 , n1730 );
nand ( n1732 , n457 , n914 );
nand ( n1733 , n1731 , n1732 );
and ( n1734 , n951 , n1733 );
not ( n1735 , n951 );
and ( n1736 , n1735 , n964 );
nor ( n1737 , n1734 , n1736 );
nand ( n1738 , n481 , n1523 );
not ( n1739 , n1738 );
and ( n1740 , n1737 , n1739 );
not ( n1741 , n1458 );
nand ( n1742 , n1741 , n1456 );
not ( n1743 , n1742 );
nand ( n1744 , n1525 , n1738 );
not ( n1745 , n1744 );
or ( n1746 , n1743 , n1745 );
or ( n1747 , n431 , n785 );
nand ( n1748 , n431 , n785 );
nand ( n1749 , n1747 , n1748 );
nand ( n1750 , n747 , n967 );
and ( n1751 , n1749 , n1750 );
not ( n1752 , n1749 );
not ( n1753 , n1750 );
and ( n1754 , n1752 , n1753 );
nor ( n1755 , n1751 , n1754 );
nand ( n1756 , n1746 , n1755 );
not ( n1757 , n454 );
nand ( n1758 , n1757 , n1163 );
not ( n1759 , n1758 );
nor ( n1760 , n634 , n1007 );
not ( n1761 , n1760 );
nand ( n1762 , n634 , n1007 );
nand ( n1763 , n1761 , n1762 );
not ( n1764 , n1763 );
or ( n1765 , n1759 , n1764 );
or ( n1766 , n1763 , n1758 );
nand ( n1767 , n1765 , n1766 );
nor ( n1768 , n1740 , n1756 , n1767 );
nor ( n1769 , n1287 , n1267 );
not ( n1770 , n1769 );
nand ( n1771 , n1267 , n1287 );
nand ( n1772 , n1770 , n1771 );
and ( n1773 , n1772 , n1712 );
not ( n1774 , n1772 );
not ( n1775 , n1712 );
and ( n1776 , n1774 , n1775 );
nor ( n1777 , n1773 , n1776 );
nor ( n1778 , n1461 , n1518 );
nand ( n1779 , n1509 , n1507 );
and ( n1780 , n1778 , n1779 );
nor ( n1781 , n1744 , n1742 );
nor ( n1782 , n1739 , n951 , n963 );
nor ( n1783 , n1780 , n1781 , n1782 );
nand ( n1784 , n1728 , n1768 , n1777 , n1783 );
not ( n1785 , n1410 );
not ( n1786 , n1454 );
or ( n1787 , n1785 , n1786 );
or ( n1788 , n1454 , n1410 );
nand ( n1789 , n1787 , n1788 );
nand ( n1790 , n1504 , n1425 );
nor ( n1791 , n1789 , n1790 );
or ( n1792 , n818 , n823 );
not ( n1793 , n787 );
or ( n1794 , n1793 , n799 );
nand ( n1795 , n1792 , n1794 , n822 );
not ( n1796 , n1795 );
not ( n1797 , n1769 );
nor ( n1798 , n1314 , n1309 );
not ( n1799 , n1798 );
nand ( n1800 , n1314 , n1309 );
nand ( n1801 , n1799 , n1800 );
not ( n1802 , n1801 );
or ( n1803 , n1797 , n1802 );
or ( n1804 , n1801 , n1769 );
nand ( n1805 , n1803 , n1804 );
nand ( n1806 , n1461 , n1518 );
or ( n1807 , n1779 , n1806 );
nor ( n1808 , n1741 , n1456 );
not ( n1809 , n1808 );
nand ( n1810 , n1809 , n1742 );
nand ( n1811 , n1807 , n1810 );
nand ( n1812 , n1796 , n1805 , n1811 );
nor ( n1813 , n702 , n1191 );
not ( n1814 , n1813 );
nand ( n1815 , n1814 , n1702 );
nor ( n1816 , n513 , n1029 );
not ( n1817 , n1816 );
xnor ( n1818 , n1815 , n1817 );
nor ( n1819 , n1812 , n1818 );
not ( n1820 , n1816 );
nand ( n1821 , n513 , n1029 );
nand ( n1822 , n1820 , n1821 );
xor ( n1823 , n1822 , n1760 );
nand ( n1824 , n1370 , n1365 );
not ( n1825 , n1824 );
not ( n1826 , n1398 );
not ( n1827 , n1382 );
or ( n1828 , n1826 , n1827 );
nand ( n1829 , n1828 , n1723 );
not ( n1830 , n1829 );
or ( n1831 , n1825 , n1830 );
or ( n1832 , n1829 , n1824 );
nand ( n1833 , n1831 , n1832 );
nor ( n1834 , n1823 , n1833 );
not ( n1835 , n1810 );
or ( n1836 , n1779 , n1778 );
nand ( n1837 , n1836 , n1806 );
and ( n1838 , n1835 , n1837 );
nand ( n1839 , n951 , n963 );
and ( n1840 , n1733 , n1839 );
not ( n1841 , n968 );
not ( n1842 , n747 );
not ( n1843 , n1842 );
or ( n1844 , n1841 , n1843 );
nand ( n1845 , n1844 , n1750 );
nand ( n1846 , n734 , n973 );
nor ( n1847 , n1845 , n1846 );
nor ( n1848 , n1838 , n1840 , n1847 );
and ( n1849 , n1845 , n1846 );
nor ( n1850 , n1849 , n1167 , n1669 );
nand ( n1851 , n1819 , n1834 , n1848 , n1850 );
nor ( n1852 , n1784 , n1791 , n1851 );
not ( n1853 , n1790 );
not ( n1854 , n1789 );
or ( n1855 , n1853 , n1854 );
or ( n1856 , n1370 , n1365 );
nand ( n1857 , n1856 , n1824 );
not ( n1858 , n1857 );
and ( n1859 , n1858 , n1324 );
and ( n1860 , n1327 , n1346 );
nor ( n1861 , n1859 , n1860 );
or ( n1862 , n1861 , n1800 );
not ( n1863 , n1739 );
not ( n1864 , n1839 );
and ( n1865 , n1863 , n1864 );
not ( n1866 , n1748 );
not ( n1867 , n806 );
or ( n1868 , n1866 , n1867 );
or ( n1869 , n806 , n1748 );
nand ( n1870 , n1868 , n1869 );
nor ( n1871 , n1865 , n1870 );
or ( n1872 , n734 , n973 );
nand ( n1873 , n1872 , n1846 );
not ( n1874 , n1873 );
not ( n1875 , n1732 );
and ( n1876 , n1874 , n1875 );
and ( n1877 , n1873 , n1732 );
nor ( n1878 , n1876 , n1877 );
nand ( n1879 , n1862 , n1871 , n1878 );
not ( n1880 , n1720 );
or ( n1881 , n1547 , n1556 );
nand ( n1882 , n1547 , n1556 );
nand ( n1883 , n1881 , n1882 );
not ( n1884 , n1883 );
or ( n1885 , n1880 , n1884 );
or ( n1886 , n1883 , n1720 );
nand ( n1887 , n1885 , n1886 );
nand ( n1888 , n1324 , n1346 );
and ( n1889 , n1857 , n1888 );
not ( n1890 , n1347 );
not ( n1891 , n1327 );
or ( n1892 , n1890 , n1891 );
nand ( n1893 , n1892 , n1888 );
and ( n1894 , n1893 , n1800 );
nor ( n1895 , n1889 , n1894 );
nand ( n1896 , n1895 , n1128 );
nor ( n1897 , n1879 , n1130 , n1887 , n1896 );
nand ( n1898 , n1855 , n1897 );
or ( n1899 , n1504 , n1425 );
nand ( n1900 , n1899 , n1790 );
or ( n1901 , n1490 , n1421 );
or ( n1902 , n1900 , n1901 );
not ( n1903 , n1421 );
not ( n1904 , n1490 );
or ( n1905 , n1903 , n1904 );
nand ( n1906 , n1905 , n1901 );
or ( n1907 , n1882 , n1906 );
nand ( n1908 , n1906 , n1882 );
nand ( n1909 , n1902 , n1907 , n1908 );
nor ( n1910 , n1898 , n1909 );
not ( n1911 , n1468 );
not ( n1912 , n1476 );
or ( n1913 , n1911 , n1912 );
or ( n1914 , n1476 , n1468 );
nand ( n1915 , n1913 , n1914 );
not ( n1916 , n1915 );
not ( n1917 , n1788 );
and ( n1918 , n1916 , n1917 );
and ( n1919 , n1915 , n1788 );
nor ( n1920 , n1918 , n1919 );
and ( n1921 , n1900 , n1901 );
not ( n1922 , n1507 );
not ( n1923 , n1922 );
not ( n1924 , n1510 );
or ( n1925 , n1923 , n1924 );
nand ( n1926 , n1925 , n1779 );
not ( n1927 , n1926 );
not ( n1928 , n1914 );
or ( n1929 , n1927 , n1928 );
or ( n1930 , n1914 , n1926 );
nand ( n1931 , n1929 , n1930 );
nor ( n1932 , n1921 , n1931 );
nand ( n1933 , n1852 , n1910 , n1920 , n1932 );
not ( n1934 , n1933 );
and ( n1935 , n1934 , n1662 );
and ( n1936 , n1669 , n822 );
and ( n1937 , n1936 , n1698 );
nor ( n1938 , n1935 , n1937 );
or ( n1939 , n1938 , n1695 );
and ( n1940 , n1933 , n900 );
not ( n1941 , n910 );
and ( n1942 , n1941 , n161 );
nor ( n1943 , n1940 , n1942 );
or ( n1944 , n1695 , n1943 );
nand ( n1945 , n908 , n878 );
buf ( n1946 , n1945 );
buf ( n1947 , n1946 );
not ( n1948 , n1947 );
not ( n1949 , n889 );
nor ( n1950 , n1949 , n898 );
buf ( n1951 , n1950 );
not ( n1952 , n1951 );
not ( n1953 , n1952 );
nand ( n1954 , n1948 , n1953 );
or ( n1955 , n1954 , n1693 );
not ( n1956 , n782 );
not ( n1957 , n1954 );
nand ( n1958 , n1956 , n1957 );
buf ( n1959 , n779 );
or ( n1960 , n1958 , n1959 );
nand ( n1961 , n1960 , n1693 );
not ( n1962 , n866 );
not ( n1963 , n22 );
not ( n1964 , n1298 );
or ( n1965 , n1963 , n1964 );
not ( n1966 , n22 );
or ( n1967 , n856 , n1966 );
not ( n1968 , n765 );
not ( n1969 , n768 );
nor ( n1970 , n1968 , n1969 , n22 );
nand ( n1971 , n1441 , n1970 );
not ( n1972 , n1971 );
nor ( n1973 , n1972 , n876 );
nand ( n1974 , n1967 , n1973 );
nand ( n1975 , n1965 , n1974 );
not ( n1976 , n21 );
not ( n1977 , n1971 );
or ( n1978 , n1976 , n1977 );
not ( n1979 , n773 );
nand ( n1980 , n1978 , n1979 );
nand ( n1981 , n876 , n21 );
nand ( n1982 , n1980 , n1981 );
not ( n1983 , n1982 );
xnor ( n1984 , n23 , n1979 );
nor ( n1985 , n1983 , n1984 );
and ( n1986 , n1975 , n1985 );
not ( n1987 , n1986 );
or ( n1988 , n1962 , n1987 );
nand ( n1989 , n1988 , n161 );
not ( n1990 , n1989 );
nand ( n1991 , n1955 , n1961 , n1990 );
nand ( n1992 , n1991 , n158 );
nand ( n1993 , n1939 , n1944 , n1992 );
nor ( n1994 , n1701 , n1993 );
not ( n1995 , n1692 );
not ( n1996 , n1995 );
not ( n1997 , n1658 );
or ( n1998 , n1996 , n1997 );
buf ( n1999 , n1953 );
not ( n2000 , n1999 );
nor ( n2001 , n2000 , n1697 );
not ( n2002 , n2001 );
nor ( n2003 , n1695 , n1936 , n2002 );
nand ( n2004 , n1998 , n2003 );
not ( n2005 , n1533 );
not ( n2006 , n2005 );
not ( n2007 , n1639 );
or ( n2008 , n2006 , n2007 );
not ( n2009 , n1257 );
not ( n2010 , n2009 );
not ( n2011 , n1293 );
or ( n2012 , n2010 , n2011 );
not ( n2013 , n1352 );
nand ( n2014 , n2012 , n2013 );
not ( n2015 , n2014 );
not ( n2016 , n1588 );
or ( n2017 , n2015 , n2016 );
nand ( n2018 , n2017 , n1405 );
not ( n2019 , n1400 );
nand ( n2020 , n2018 , n1576 , n2019 );
not ( n2021 , n1402 );
not ( n2022 , n1595 );
or ( n2023 , n2021 , n2022 );
nand ( n2024 , n2023 , n1576 );
nor ( n2025 , n1624 , n1622 );
and ( n2026 , n1619 , n1593 , n2025 );
nand ( n2027 , n2020 , n2024 , n2026 );
nand ( n2028 , n2008 , n2027 );
not ( n2029 , n1655 );
nor ( n2030 , n809 , n1669 );
nand ( n2031 , n880 , n2001 );
and ( n2032 , n2031 , n910 );
nand ( n2033 , n2030 , n2032 );
not ( n2034 , n1648 );
nand ( n2035 , n2034 , n1604 );
nor ( n2036 , n2029 , n2033 , n2035 );
and ( n2037 , n2028 , n2036 );
not ( n2038 , n2028 );
nor ( n2039 , n1644 , n802 );
and ( n2040 , n880 , n1698 );
not ( n2041 , n1668 );
nor ( n2042 , n2041 , n1691 );
nor ( n2043 , n2040 , n2042 );
nand ( n2044 , n2039 , n2043 );
nor ( n2045 , n2044 , n966 );
and ( n2046 , n2038 , n2045 );
nor ( n2047 , n2037 , n2046 );
not ( n2048 , n2035 );
not ( n2049 , n2045 );
or ( n2050 , n2048 , n2049 );
not ( n2051 , n2044 );
not ( n2052 , n1655 );
and ( n2053 , n2051 , n2052 );
not ( n2054 , n2042 );
or ( n2055 , n1941 , n2054 );
nand ( n2056 , n2055 , n2040 );
not ( n2057 , n2056 );
not ( n2058 , n2031 );
or ( n2059 , n2057 , n2058 );
not ( n2060 , n2043 );
or ( n2061 , n2060 , n2030 );
nand ( n2062 , n2059 , n2061 );
nor ( n2063 , n2053 , n2062 );
nand ( n2064 , n2050 , n2063 );
not ( n2065 , n2039 );
not ( n2066 , n2065 );
not ( n2067 , n2033 );
not ( n2068 , n2067 );
or ( n2069 , n2066 , n2068 );
nand ( n2070 , n2067 , n1655 , n966 );
nand ( n2071 , n2069 , n2070 );
nor ( n2072 , n2064 , n2071 );
nand ( n2073 , n2047 , n2072 );
nand ( n2074 , n1687 , n1994 , n2004 , n2073 );
not ( n2075 , n1586 );
nand ( n2076 , n814 , n1077 );
nor ( n2077 , n2076 , n1120 );
and ( n2078 , n2077 , n1047 );
and ( n2079 , n2078 , n1147 );
not ( n2080 , n634 );
nand ( n2081 , n2079 , n2080 );
nor ( n2082 , n2081 , n1014 );
not ( n2083 , n1172 );
nand ( n2084 , n2082 , n2083 );
not ( n2085 , n2084 );
buf ( n2086 , n1214 );
not ( n2087 , n2086 );
nand ( n2088 , n2085 , n2087 );
nor ( n2089 , n2088 , n1233 );
nand ( n2090 , n2089 , n1274 );
not ( n2091 , n2090 );
nand ( n2092 , n2091 , n1314 );
not ( n2093 , n2092 );
or ( n2094 , n2075 , n2093 );
or ( n2095 , n2092 , n1586 );
nand ( n2096 , n2094 , n2095 );
not ( n2097 , n1984 );
nand ( n2098 , n2097 , n158 );
and ( n2099 , n1975 , n2098 );
not ( n2100 , n2099 );
not ( n2101 , n1975 );
not ( n2102 , n158 );
nor ( n2103 , n1982 , n2102 );
nand ( n2104 , n2101 , n2103 );
buf ( n2105 , n2104 );
not ( n2106 , n2102 );
not ( n2107 , n1975 );
or ( n2108 , n2106 , n2107 );
nor ( n2109 , n1984 , n160 );
nand ( n2110 , n2108 , n2109 );
not ( n2111 , n2110 );
nand ( n2112 , n2100 , n2105 , n2111 );
not ( n2113 , n2099 );
not ( n2114 , n159 );
nand ( n2115 , n2113 , n2105 , n2114 );
not ( n2116 , n2099 );
nand ( n2117 , n2116 , n1984 );
not ( n2118 , n1986 );
nor ( n2119 , n865 , n1697 );
nand ( n2120 , n1983 , n1984 );
and ( n2121 , n2118 , n2119 , n2120 );
and ( n2122 , n2112 , n2115 , n2117 , n2121 );
buf ( n2123 , n2122 );
not ( n2124 , n782 );
not ( n2125 , n2124 );
and ( n2126 , n2123 , n1957 , n2125 );
and ( n2127 , n2096 , n2126 );
buf ( n2128 , n2122 );
not ( n2129 , n2128 );
nor ( n2130 , n1958 , n2129 );
buf ( n2131 , n2130 );
not ( n2132 , n2131 );
not ( n2133 , n1274 );
nor ( n2134 , n2132 , n2133 );
nor ( n2135 , n2127 , n2134 );
not ( n2136 , n1805 );
not ( n2137 , n2136 );
or ( n2138 , n1713 , n1705 );
not ( n2139 , n1822 );
nand ( n2140 , n2139 , n1760 );
and ( n2141 , n2138 , n2140 );
buf ( n2142 , n987 );
nand ( n2143 , n1166 , n2142 );
not ( n2144 , n1763 );
nand ( n2145 , n2143 , n2144 );
nor ( n2146 , n1706 , n1702 );
not ( n2147 , n2146 );
nor ( n2148 , n1815 , n1817 );
not ( n2149 , n2148 );
and ( n2150 , n2141 , n2145 , n2147 , n2149 );
not ( n2151 , n2150 );
nor ( n2152 , n2143 , n2144 );
not ( n2153 , n2152 );
nand ( n2154 , n2153 , n2145 );
not ( n2155 , n2154 );
nand ( n2156 , n1169 , n2155 );
not ( n2157 , n2156 );
or ( n2158 , n2151 , n2157 );
not ( n2159 , n2146 );
not ( n2160 , n2138 );
not ( n2161 , n2160 );
nand ( n2162 , n2159 , n2161 , n1818 , n2149 );
nor ( n2163 , n2146 , n2148 );
nand ( n2164 , n2141 , n2163 , n1823 );
nand ( n2165 , n2162 , n2164 );
not ( n2166 , n2146 );
not ( n2167 , n1707 );
nand ( n2168 , n2166 , n2167 );
and ( n2169 , n2168 , n1718 );
nor ( n2170 , n2169 , n2160 );
nor ( n2171 , n2165 , n2170 );
nand ( n2172 , n2158 , n2171 );
not ( n2173 , n1777 );
or ( n2174 , n2172 , n2173 );
or ( n2175 , n1772 , n1712 );
nand ( n2176 , n2174 , n2175 );
not ( n2177 , n2176 );
or ( n2178 , n2137 , n2177 );
or ( n2179 , n2176 , n2136 );
nand ( n2180 , n2178 , n2179 );
not ( n2181 , n2180 );
not ( n2182 , n2123 );
not ( n2183 , n1945 );
not ( n2184 , n2183 );
nor ( n2185 , n908 , n878 );
not ( n2186 , n2185 );
nand ( n2187 , n2184 , n2186 );
buf ( n2188 , n2187 );
or ( n2189 , n909 , n898 );
nand ( n2190 , n909 , n890 );
nand ( n2191 , n2189 , n2190 );
nor ( n2192 , n2188 , n2191 );
not ( n2193 , n2192 );
nor ( n2194 , n2182 , n2193 );
buf ( n2195 , n2194 );
not ( n2196 , n2195 );
or ( n2197 , n2181 , n2196 );
and ( n2198 , n2117 , n2121 , n2112 , n2115 );
nand ( n2199 , n2185 , n898 );
not ( n2200 , n2199 );
not ( n2201 , n2200 );
not ( n2202 , n2201 );
nand ( n2203 , n2198 , n2202 );
not ( n2204 , n2203 );
not ( n2205 , n1309 );
and ( n2206 , n2204 , n2205 );
nand ( n2207 , n2185 , n1950 );
nand ( n2208 , n2199 , n2207 );
not ( n2209 , n2208 );
buf ( n2210 , n2185 );
nand ( n2211 , n2209 , n2210 );
not ( n2212 , n2211 );
nand ( n2213 , n2118 , n2119 );
buf ( n2214 , n2213 );
not ( n2215 , n2214 );
nand ( n2216 , n2212 , n2215 );
or ( n2217 , n2216 , n1309 );
not ( n2218 , n61 );
nor ( n2219 , n2218 , n161 );
not ( n2220 , n2219 );
nand ( n2221 , n2217 , n2220 );
nor ( n2222 , n2206 , n2221 );
nand ( n2223 , n2197 , n2222 );
not ( n2224 , n2211 );
not ( n2225 , n2114 );
not ( n2226 , n2104 );
or ( n2227 , n2225 , n2226 );
nand ( n2228 , n2227 , n2097 );
nand ( n2229 , n2228 , n2116 );
not ( n2230 , n2104 );
not ( n2231 , n2111 );
or ( n2232 , n2230 , n2231 );
nand ( n2233 , n2232 , n2120 );
not ( n2234 , n2233 );
not ( n2235 , n2200 );
nand ( n2236 , n2235 , n2187 , n1952 );
nand ( n2237 , n2229 , n2234 , n2236 );
not ( n2238 , n2237 );
or ( n2239 , n2224 , n2238 );
nand ( n2240 , n2239 , n2215 );
nand ( n2241 , n2240 , n161 );
not ( n2242 , n2241 );
not ( n2243 , n2242 );
and ( n2244 , n47 , n39 );
and ( n2245 , n2244 , n51 );
and ( n2246 , n2245 , n35 );
nand ( n2247 , n2246 , n43 );
not ( n2248 , n2247 );
and ( n2249 , n59 , n2248 );
nand ( n2250 , n2249 , n55 );
not ( n2251 , n2250 );
not ( n2252 , n61 );
and ( n2253 , n2251 , n2252 );
and ( n2254 , n2250 , n61 );
nor ( n2255 , n2253 , n2254 );
nor ( n2256 , n2243 , n2255 );
nor ( n2257 , n2223 , n2256 );
and ( n2258 , n2083 , n1192 );
nand ( n2259 , n1706 , n2258 );
nand ( n2260 , n1212 , n1263 );
or ( n2261 , n1714 , n2260 );
or ( n2262 , n513 , n1196 );
not ( n2263 , n2262 );
nand ( n2264 , n1815 , n2263 );
and ( n2265 , n2259 , n2261 , n2264 );
not ( n2266 , n2265 );
not ( n2267 , n2262 );
not ( n2268 , n1815 );
not ( n2269 , n2268 );
or ( n2270 , n2267 , n2269 );
nand ( n2271 , n2080 , n1007 );
not ( n2272 , n2271 );
not ( n2273 , n2139 );
or ( n2274 , n2272 , n2273 );
not ( n2275 , n2271 );
nand ( n2276 , n2275 , n1822 );
nand ( n2277 , n2274 , n2276 );
not ( n2278 , n2277 );
not ( n2279 , n2278 );
not ( n2280 , n1146 );
nand ( n2281 , n1166 , n1763 , n2280 );
not ( n2282 , n2281 );
and ( n2283 , n1166 , n2280 );
nor ( n2284 , n2283 , n1763 );
nor ( n2285 , n2282 , n2284 );
not ( n2286 , n1112 );
not ( n2287 , n1120 );
or ( n2288 , n2286 , n2287 );
nor ( n2289 , n1078 , n1083 );
nand ( n2290 , n2288 , n2289 );
nand ( n2291 , n2290 , n1115 );
not ( n2292 , n2291 );
not ( n2293 , n1064 );
or ( n2294 , n2292 , n2293 );
not ( n2295 , n1061 );
nand ( n2296 , n2295 , n1062 );
nand ( n2297 , n2294 , n2296 );
and ( n2298 , n1167 , n2297 );
nand ( n2299 , n2285 , n2298 );
buf ( n2300 , n2281 );
nand ( n2301 , n2299 , n2300 );
not ( n2302 , n2301 );
or ( n2303 , n2279 , n2302 );
nand ( n2304 , n2303 , n2276 );
nand ( n2305 , n2270 , n2304 );
not ( n2306 , n2305 );
or ( n2307 , n2266 , n2306 );
not ( n2308 , n2260 );
not ( n2309 , n1714 );
or ( n2310 , n2308 , n2309 );
nand ( n2311 , n2310 , n2261 );
and ( n2312 , n2311 , n2261 );
or ( n2313 , n1706 , n2258 );
nand ( n2314 , n2313 , n2259 );
and ( n2315 , n2314 , n2259 , n2261 );
nor ( n2316 , n1233 , n1253 );
nor ( n2317 , n1772 , n2316 );
nor ( n2318 , n2312 , n2315 , n2317 );
nand ( n2319 , n2307 , n2318 );
nand ( n2320 , n1772 , n2316 );
nand ( n2321 , n1268 , n1287 );
nand ( n2322 , n2320 , n2321 );
not ( n2323 , n1801 );
and ( n2324 , n2322 , n2323 );
not ( n2325 , n2322 );
not ( n2326 , n1801 );
not ( n2327 , n2326 );
and ( n2328 , n2325 , n2327 );
or ( n2329 , n2324 , n2328 );
and ( n2330 , n2319 , n2329 );
not ( n2331 , n2319 );
not ( n2332 , n1801 );
and ( n2333 , n2321 , n2332 );
not ( n2334 , n2321 );
not ( n2335 , n2326 );
and ( n2336 , n2334 , n2335 );
or ( n2337 , n2333 , n2336 );
and ( n2338 , n2331 , n2337 );
or ( n2339 , n2330 , n2338 );
not ( n2340 , n2187 );
nand ( n2341 , n2340 , n2191 );
not ( n2342 , n2341 );
and ( n2343 , n2128 , n2342 );
nand ( n2344 , n2339 , n2343 );
buf ( n2345 , n2207 );
not ( n2346 , n2345 );
nand ( n2347 , n2122 , n2346 );
not ( n2348 , n2347 );
not ( n2349 , n1309 );
and ( n2350 , n1112 , n1083 );
and ( n2351 , n2350 , n1058 );
nand ( n2352 , n2351 , n1163 );
nor ( n2353 , n2352 , n1007 );
nand ( n2354 , n2353 , n1196 );
nor ( n2355 , n2354 , n1192 );
and ( n2356 , n2355 , n1230 );
nand ( n2357 , n2356 , n1253 );
nor ( n2358 , n2357 , n1287 );
not ( n2359 , n2358 );
not ( n2360 , n2359 );
or ( n2361 , n2349 , n2360 );
or ( n2362 , n2359 , n1309 );
nand ( n2363 , n2361 , n2362 );
nand ( n2364 , n2348 , n2363 );
nand ( n2365 , n2135 , n2257 , n2344 , n2364 );
not ( n2366 , n1177 );
nand ( n2367 , n2131 , n2366 );
or ( n2368 , n2246 , n43 );
nand ( n2369 , n2368 , n2247 , n2242 );
and ( n2370 , n1697 , n43 );
not ( n2371 , n2370 );
and ( n2372 , n2367 , n2369 , n2371 );
not ( n2373 , n2314 );
not ( n2374 , n2373 );
xor ( n2375 , n1815 , n2304 );
and ( n2376 , n2375 , n2263 );
and ( n2377 , n1815 , n2304 );
nor ( n2378 , n2376 , n2377 );
not ( n2379 , n2378 );
or ( n2380 , n2374 , n2379 );
or ( n2381 , n2378 , n2373 );
nand ( n2382 , n2380 , n2381 );
and ( n2383 , n2382 , n2343 );
or ( n2384 , n2355 , n1230 );
not ( n2385 , n2356 );
nand ( n2386 , n2384 , n2385 );
nor ( n2387 , n2347 , n2386 );
nor ( n2388 , n2383 , n2387 );
not ( n2389 , n2089 );
nand ( n2390 , n2088 , n1239 );
and ( n2391 , n2126 , n2389 , n2390 );
not ( n2392 , n2167 );
not ( n2393 , n1818 );
not ( n2394 , n2393 );
not ( n2395 , n1823 );
not ( n2396 , n2395 );
nand ( n2397 , n2156 , n2145 );
not ( n2398 , n2397 );
or ( n2399 , n2396 , n2398 );
nand ( n2400 , n2399 , n2140 );
not ( n2401 , n2400 );
or ( n2402 , n2394 , n2401 );
nand ( n2403 , n2402 , n2149 );
not ( n2404 , n2403 );
or ( n2405 , n2392 , n2404 );
or ( n2406 , n2403 , n2167 );
nand ( n2407 , n2405 , n2406 );
and ( n2408 , n2407 , n2195 );
nor ( n2409 , n2391 , n2408 );
not ( n2410 , n1230 );
nand ( n2411 , n2203 , n2216 );
buf ( n2412 , n2411 );
nand ( n2413 , n2410 , n2412 );
nand ( n2414 , n2372 , n2388 , n2409 , n2413 );
and ( n2415 , n118 , n1502 );
not ( n2416 , n118 );
not ( n2417 , n1502 );
and ( n2418 , n2416 , n2417 );
nor ( n2419 , n2415 , n2418 );
not ( n2420 , n2419 );
not ( n2421 , n121 );
not ( n2422 , n1487 );
or ( n2423 , n2421 , n2422 );
or ( n2424 , n1487 , n121 );
nand ( n2425 , n2423 , n2424 );
not ( n2426 , n2425 );
buf ( n2427 , n1542 );
not ( n2428 , n2427 );
not ( n2429 , n78 );
or ( n2430 , n2428 , n2429 );
or ( n2431 , n2427 , n78 );
nand ( n2432 , n2430 , n2431 );
not ( n2433 , n2432 );
not ( n2434 , n1570 );
not ( n2435 , n2434 );
not ( n2436 , n81 );
or ( n2437 , n2435 , n2436 );
or ( n2438 , n2434 , n81 );
nand ( n2439 , n2437 , n2438 );
not ( n2440 , n2439 );
not ( n2441 , n1395 );
not ( n2442 , n2441 );
not ( n2443 , n69 );
or ( n2444 , n2442 , n2443 );
or ( n2445 , n2441 , n69 );
nand ( n2446 , n2444 , n2445 );
not ( n2447 , n2446 );
not ( n2448 , n1359 );
not ( n2449 , n73 );
or ( n2450 , n2448 , n2449 );
or ( n2451 , n1359 , n73 );
nand ( n2452 , n2450 , n2451 );
not ( n2453 , n2452 );
nand ( n2454 , n62 , n1305 );
nand ( n2455 , n53 , n1283 );
nand ( n2456 , n2454 , n2455 );
not ( n2457 , n1225 );
nand ( n2458 , n2457 , n42 );
not ( n2459 , n1248 );
nand ( n2460 , n2459 , n57 );
nand ( n2461 , n2458 , n2460 );
nor ( n2462 , n2456 , n2461 );
not ( n2463 , n2462 );
and ( n2464 , n49 , n1024 );
not ( n2465 , n49 );
not ( n2466 , n1024 );
and ( n2467 , n2465 , n2466 );
nor ( n2468 , n2464 , n2467 );
not ( n2469 , n2468 );
and ( n2470 , n48 , n1005 );
not ( n2471 , n48 );
not ( n2472 , n1005 );
and ( n2473 , n2471 , n2472 );
nor ( n2474 , n2470 , n2473 );
not ( n2475 , n2474 );
xor ( n2476 , n1134 , n1159 );
not ( n2477 , n2476 );
nand ( n2478 , n6 , n147 );
not ( n2479 , n2478 );
not ( n2480 , n153 );
and ( n2481 , n2479 , n2480 );
and ( n2482 , n2478 , n153 );
nor ( n2483 , n2481 , n2482 );
or ( n2484 , n1107 , n2483 );
not ( n2485 , n153 );
or ( n2486 , n2478 , n2485 );
nand ( n2487 , n2484 , n2486 );
not ( n2488 , n2487 );
xnor ( n2489 , n1034 , n1054 );
not ( n2490 , n2489 );
or ( n2491 , n2488 , n2490 );
nand ( n2492 , n1054 , n155 );
nand ( n2493 , n2491 , n2492 );
not ( n2494 , n2493 );
or ( n2495 , n2477 , n2494 );
nand ( n2496 , n37 , n1160 );
nand ( n2497 , n2495 , n2496 );
not ( n2498 , n2497 );
or ( n2499 , n2475 , n2498 );
nand ( n2500 , n1005 , n48 );
nand ( n2501 , n2499 , n2500 );
not ( n2502 , n2501 );
or ( n2503 , n2469 , n2502 );
nand ( n2504 , n1024 , n49 );
nand ( n2505 , n2503 , n2504 );
and ( n2506 , n33 , n1187 );
not ( n2507 , n33 );
not ( n2508 , n1187 );
and ( n2509 , n2507 , n2508 );
nor ( n2510 , n2506 , n2509 );
and ( n2511 , n2505 , n2510 );
and ( n2512 , n1187 , n33 );
nor ( n2513 , n2511 , n2512 );
not ( n2514 , n2513 );
or ( n2515 , n2463 , n2514 );
not ( n2516 , n2462 );
and ( n2517 , n42 , n1225 );
not ( n2518 , n42 );
and ( n2519 , n2518 , n2457 );
nor ( n2520 , n2517 , n2519 );
not ( n2521 , n2520 );
or ( n2522 , n2516 , n2521 );
not ( n2523 , n2456 );
and ( n2524 , n57 , n2459 );
not ( n2525 , n57 );
and ( n2526 , n2525 , n1248 );
nor ( n2527 , n2524 , n2526 );
not ( n2528 , n2527 );
nand ( n2529 , n2528 , n2460 );
not ( n2530 , n2529 );
and ( n2531 , n2523 , n2530 );
and ( n2532 , n1305 , n705 );
not ( n2533 , n1305 );
and ( n2534 , n2533 , n62 );
nor ( n2535 , n2532 , n2534 );
buf ( n2536 , n2454 );
and ( n2537 , n2535 , n2536 );
nor ( n2538 , n2531 , n2537 );
nand ( n2539 , n2522 , n2538 );
and ( n2540 , n53 , n1283 );
not ( n2541 , n53 );
not ( n2542 , n1283 );
and ( n2543 , n2541 , n2542 );
nor ( n2544 , n2540 , n2543 );
or ( n2545 , n2456 , n2544 );
and ( n2546 , n65 , n1340 );
not ( n2547 , n65 );
and ( n2548 , n2547 , n1339 );
or ( n2549 , n2546 , n2548 );
nand ( n2550 , n2545 , n2549 );
nor ( n2551 , n2539 , n2550 );
nand ( n2552 , n2515 , n2551 );
nand ( n2553 , n65 , n1339 );
nand ( n2554 , n2552 , n2553 );
not ( n2555 , n2554 );
or ( n2556 , n2453 , n2555 );
not ( n2557 , n1359 );
nand ( n2558 , n2557 , n73 );
nand ( n2559 , n2556 , n2558 );
not ( n2560 , n2559 );
or ( n2561 , n2447 , n2560 );
nand ( n2562 , n69 , n1395 );
nand ( n2563 , n2561 , n2562 );
not ( n2564 , n2563 );
or ( n2565 , n2440 , n2564 );
nand ( n2566 , n81 , n1570 );
nand ( n2567 , n2565 , n2566 );
not ( n2568 , n2567 );
or ( n2569 , n2433 , n2568 );
not ( n2570 , n2427 );
nand ( n2571 , n2570 , n78 );
nand ( n2572 , n2569 , n2571 );
not ( n2573 , n2572 );
or ( n2574 , n2426 , n2573 );
not ( n2575 , n1487 );
nand ( n2576 , n2575 , n121 );
nand ( n2577 , n2574 , n2576 );
not ( n2578 , n2577 );
or ( n2579 , n2420 , n2578 );
nand ( n2580 , n118 , n1502 );
nand ( n2581 , n2579 , n2580 );
buf ( n2582 , n1452 );
not ( n2583 , n2582 );
xor ( n2584 , n112 , n2583 );
and ( n2585 , n2581 , n2584 );
and ( n2586 , n112 , n2583 );
nor ( n2587 , n2585 , n2586 );
not ( n2588 , n109 );
and ( n2589 , n2587 , n2588 );
not ( n2590 , n1959 );
not ( n2591 , n1946 );
nand ( n2592 , n2591 , n866 );
nand ( n2593 , n2590 , n2592 );
nor ( n2594 , n2593 , n1989 );
not ( n2595 , n782 );
nand ( n2596 , n2594 , n2595 );
not ( n2597 , n2596 );
not ( n2598 , n2597 );
nor ( n2599 , n2589 , n2598 );
not ( n2600 , n2587 );
nand ( n2601 , n2600 , n109 );
nand ( n2602 , n2599 , n2601 );
not ( n2603 , n2602 );
nand ( n2604 , n2603 , n890 );
xor ( n2605 , n1661 , n110 );
not ( n2606 , n2582 );
not ( n2607 , n113 );
not ( n2608 , n2607 );
and ( n2609 , n2606 , n2608 );
and ( n2610 , n117 , n2417 );
not ( n2611 , n117 );
and ( n2612 , n2611 , n1502 );
nor ( n2613 , n2610 , n2612 );
not ( n2614 , n2613 );
not ( n2615 , n2614 );
not ( n2616 , n122 );
not ( n2617 , n1487 );
or ( n2618 , n2616 , n2617 );
or ( n2619 , n1487 , n122 );
nand ( n2620 , n2618 , n2619 );
not ( n2621 , n2620 );
not ( n2622 , n79 );
not ( n2623 , n2427 );
or ( n2624 , n2622 , n2623 );
or ( n2625 , n2427 , n79 );
nand ( n2626 , n2624 , n2625 );
not ( n2627 , n2626 );
not ( n2628 , n82 );
not ( n2629 , n2434 );
or ( n2630 , n2628 , n2629 );
or ( n2631 , n82 , n2434 );
nand ( n2632 , n2630 , n2631 );
not ( n2633 , n2632 );
not ( n2634 , n70 );
not ( n2635 , n2441 );
or ( n2636 , n2634 , n2635 );
or ( n2637 , n2441 , n70 );
nand ( n2638 , n2636 , n2637 );
not ( n2639 , n2638 );
not ( n2640 , n74 );
not ( n2641 , n1359 );
or ( n2642 , n2640 , n2641 );
or ( n2643 , n1359 , n74 );
nand ( n2644 , n2642 , n2643 );
not ( n2645 , n2644 );
and ( n2646 , n58 , n2459 );
not ( n2647 , n2646 );
nand ( n2648 , n2457 , n41 );
nand ( n2649 , n2647 , n2648 );
nand ( n2650 , n1283 , n54 );
nand ( n2651 , n1305 , n63 );
nand ( n2652 , n2650 , n2651 );
nor ( n2653 , n2649 , n2652 );
nand ( n2654 , n1187 , n34 );
and ( n2655 , n2653 , n2654 );
not ( n2656 , n2655 );
and ( n2657 , n50 , n1024 );
not ( n2658 , n50 );
and ( n2659 , n2658 , n2466 );
nor ( n2660 , n2657 , n2659 );
not ( n2661 , n2660 );
and ( n2662 , n46 , n1005 );
not ( n2663 , n46 );
and ( n2664 , n2663 , n2472 );
nor ( n2665 , n2662 , n2664 );
not ( n2666 , n2665 );
and ( n2667 , n38 , n1160 );
not ( n2668 , n38 );
and ( n2669 , n2668 , n1159 );
nor ( n2670 , n2667 , n2669 );
not ( n2671 , n2670 );
nand ( n2672 , n6 , n148 );
and ( n2673 , n2672 , n152 );
not ( n2674 , n2672 );
not ( n2675 , n152 );
and ( n2676 , n2674 , n2675 );
nor ( n2677 , n2673 , n2676 );
or ( n2678 , n1107 , n2677 );
or ( n2679 , n2672 , n2675 );
nand ( n2680 , n2678 , n2679 );
not ( n2681 , n2680 );
not ( n2682 , n1054 );
and ( n2683 , n2682 , n1044 );
not ( n2684 , n2682 );
and ( n2685 , n2684 , n157 );
nor ( n2686 , n2683 , n2685 );
not ( n2687 , n2686 );
or ( n2688 , n2681 , n2687 );
nand ( n2689 , n1054 , n157 );
nand ( n2690 , n2688 , n2689 );
not ( n2691 , n2690 );
or ( n2692 , n2671 , n2691 );
nand ( n2693 , n1160 , n38 );
nand ( n2694 , n2692 , n2693 );
not ( n2695 , n2694 );
or ( n2696 , n2666 , n2695 );
nand ( n2697 , n1005 , n46 );
nand ( n2698 , n2696 , n2697 );
not ( n2699 , n2698 );
or ( n2700 , n2661 , n2699 );
nand ( n2701 , n1024 , n50 );
nand ( n2702 , n2700 , n2701 );
and ( n2703 , n34 , n1187 );
not ( n2704 , n34 );
and ( n2705 , n2704 , n2508 );
nor ( n2706 , n2703 , n2705 );
nand ( n2707 , n2702 , n2706 );
not ( n2708 , n2707 );
or ( n2709 , n2656 , n2708 );
and ( n2710 , n2457 , n41 );
not ( n2711 , n2457 );
not ( n2712 , n41 );
and ( n2713 , n2711 , n2712 );
nor ( n2714 , n2710 , n2713 );
not ( n2715 , n2714 );
not ( n2716 , n2715 );
not ( n2717 , n2653 );
or ( n2718 , n2716 , n2717 );
and ( n2719 , n63 , n1306 );
not ( n2720 , n63 );
and ( n2721 , n2720 , n1305 );
or ( n2722 , n2719 , n2721 );
not ( n2723 , n2722 );
not ( n2724 , n2651 );
not ( n2725 , n2724 );
and ( n2726 , n2723 , n2725 );
xor ( n2727 , n58 , n2459 );
or ( n2728 , n2646 , n2727 );
nor ( n2729 , n2652 , n2728 );
nor ( n2730 , n2726 , n2729 );
nand ( n2731 , n2718 , n2730 );
and ( n2732 , n54 , n2542 );
not ( n2733 , n54 );
and ( n2734 , n2733 , n1283 );
nor ( n2735 , n2732 , n2734 );
not ( n2736 , n2735 );
or ( n2737 , n2652 , n2736 );
and ( n2738 , n66 , n1340 );
not ( n2739 , n66 );
and ( n2740 , n2739 , n1339 );
or ( n2741 , n2738 , n2740 );
nand ( n2742 , n2737 , n2741 );
nor ( n2743 , n2731 , n2742 );
nand ( n2744 , n2709 , n2743 );
nand ( n2745 , n66 , n1339 );
nand ( n2746 , n2744 , n2745 );
not ( n2747 , n2746 );
or ( n2748 , n2645 , n2747 );
nand ( n2749 , n2557 , n74 );
nand ( n2750 , n2748 , n2749 );
not ( n2751 , n2750 );
or ( n2752 , n2639 , n2751 );
nand ( n2753 , n70 , n1395 );
nand ( n2754 , n2752 , n2753 );
not ( n2755 , n2754 );
or ( n2756 , n2633 , n2755 );
nand ( n2757 , n1570 , n82 );
nand ( n2758 , n2756 , n2757 );
not ( n2759 , n2758 );
or ( n2760 , n2627 , n2759 );
nand ( n2761 , n2570 , n79 );
nand ( n2762 , n2760 , n2761 );
not ( n2763 , n2762 );
or ( n2764 , n2621 , n2763 );
nand ( n2765 , n2575 , n122 );
nand ( n2766 , n2764 , n2765 );
not ( n2767 , n2766 );
or ( n2768 , n2615 , n2767 );
nand ( n2769 , n1502 , n117 );
nand ( n2770 , n2768 , n2769 );
and ( n2771 , n2582 , n2607 );
not ( n2772 , n2582 );
and ( n2773 , n2772 , n113 );
nor ( n2774 , n2771 , n2773 );
and ( n2775 , n2770 , n2774 );
nor ( n2776 , n2609 , n2775 );
xnor ( n2777 , n2605 , n2776 );
not ( n2778 , n2592 );
nand ( n2779 , n2595 , n1959 );
nor ( n2780 , n2778 , n2779 );
and ( n2781 , n1990 , n2780 );
buf ( n2782 , n2781 );
buf ( n2783 , n2782 );
nand ( n2784 , n2777 , n2783 );
not ( n2785 , n2594 );
nor ( n2786 , n2785 , n890 );
and ( n2787 , n2602 , n2786 );
not ( n2788 , n221 );
nand ( n2789 , n962 , n2592 );
and ( n2790 , n1990 , n2789 );
buf ( n2791 , n2790 );
not ( n2792 , n2791 );
or ( n2793 , n2788 , n2792 );
nand ( n2794 , n1697 , n111 );
nand ( n2795 , n2793 , n2794 );
nor ( n2796 , n2787 , n2795 );
nand ( n2797 , n2604 , n2784 , n2796 );
not ( n2798 , n2317 );
nand ( n2799 , n2798 , n2320 );
not ( n2800 , n2799 );
not ( n2801 , n2311 );
not ( n2802 , n2801 );
not ( n2803 , n2264 );
not ( n2804 , n2305 );
or ( n2805 , n2803 , n2804 );
nand ( n2806 , n2805 , n2373 );
nand ( n2807 , n2806 , n2259 );
not ( n2808 , n2807 );
or ( n2809 , n2802 , n2808 );
nand ( n2810 , n2809 , n2261 );
not ( n2811 , n2810 );
or ( n2812 , n2800 , n2811 );
or ( n2813 , n2810 , n2799 );
nand ( n2814 , n2812 , n2813 );
nand ( n2815 , n2814 , n2343 );
nand ( n2816 , n2412 , n1287 );
nand ( n2817 , n2090 , n1320 );
nand ( n2818 , n2817 , n2092 , n2126 );
not ( n2819 , n1777 );
not ( n2820 , n2172 );
or ( n2821 , n2819 , n2820 );
or ( n2822 , n2172 , n1777 );
nand ( n2823 , n2821 , n2822 );
nand ( n2824 , n2194 , n2823 );
and ( n2825 , n2357 , n1287 );
nor ( n2826 , n2825 , n2358 );
nand ( n2827 , n2348 , n2826 );
and ( n2828 , n2816 , n2818 , n2824 , n2827 );
not ( n2829 , n1290 );
not ( n2830 , n2131 );
or ( n2831 , n2829 , n2830 );
nand ( n2832 , n1697 , n55 );
nand ( n2833 , n2831 , n2832 );
or ( n2834 , n2249 , n55 );
nand ( n2835 , n2834 , n2250 );
nor ( n2836 , n2243 , n2835 );
nor ( n2837 , n2833 , n2836 );
nand ( n2838 , n2815 , n2828 , n2837 );
and ( n2839 , n2807 , n2311 );
not ( n2840 , n2807 );
and ( n2841 , n2840 , n2801 );
nor ( n2842 , n2839 , n2841 );
not ( n2843 , n2343 );
nor ( n2844 , n2842 , n2843 );
not ( n2845 , n2126 );
or ( n2846 , n2089 , n1274 );
nand ( n2847 , n2846 , n2090 );
nor ( n2848 , n2845 , n2847 );
xor ( n2849 , n59 , n2248 );
not ( n2850 , n2849 );
not ( n2851 , n2242 );
or ( n2852 , n2850 , n2851 );
nor ( n2853 , n2356 , n1254 );
nand ( n2854 , n2348 , n2853 );
nand ( n2855 , n2852 , n2854 );
nor ( n2856 , n2844 , n2848 , n2855 );
not ( n2857 , n1718 );
and ( n2858 , n2403 , n1707 );
not ( n2859 , n2147 );
nor ( n2860 , n2858 , n2859 );
not ( n2861 , n2860 );
or ( n2862 , n2857 , n2861 );
or ( n2863 , n2860 , n1718 );
nand ( n2864 , n2862 , n2863 );
nand ( n2865 , n2864 , n2195 );
nor ( n2866 , n2347 , n2385 );
or ( n2867 , n2866 , n2412 );
nand ( n2868 , n2867 , n1254 );
and ( n2869 , n2131 , n2087 );
and ( n2870 , n1697 , n59 );
nor ( n2871 , n2869 , n2870 );
nand ( n2872 , n2856 , n2865 , n2868 , n2871 );
not ( n2873 , n1195 );
not ( n2874 , n2130 );
or ( n2875 , n2873 , n2874 );
nand ( n2876 , n1697 , n35 );
nand ( n2877 , n2875 , n2876 );
or ( n2878 , n2245 , n35 );
not ( n2879 , n2246 );
nand ( n2880 , n2878 , n2879 );
nor ( n2881 , n2243 , n2880 );
nor ( n2882 , n2877 , n2881 );
nor ( n2883 , n2375 , n2262 );
not ( n2884 , n2883 );
nand ( n2885 , n2375 , n2262 );
nand ( n2886 , n2884 , n2885 );
and ( n2887 , n2886 , n2343 );
nand ( n2888 , n2084 , n2086 );
and ( n2889 , n2888 , n2088 );
and ( n2890 , n2126 , n2889 );
nor ( n2891 , n2887 , n2890 );
not ( n2892 , n1818 );
not ( n2893 , n2400 );
or ( n2894 , n2892 , n2893 );
or ( n2895 , n2400 , n1818 );
nand ( n2896 , n2894 , n2895 );
and ( n2897 , n2194 , n2896 );
and ( n2898 , n2354 , n1192 );
nor ( n2899 , n2898 , n2355 );
and ( n2900 , n2348 , n2899 );
nor ( n2901 , n2897 , n2900 );
not ( n2902 , n2411 );
not ( n2903 , n2902 );
nand ( n2904 , n2903 , n1192 );
nand ( n2905 , n2882 , n2891 , n2901 , n2904 );
not ( n2906 , n1029 );
not ( n2907 , n2353 );
or ( n2908 , n2906 , n2907 );
or ( n2909 , n2353 , n1029 );
nand ( n2910 , n2908 , n2909 );
and ( n2911 , n2346 , n2910 );
and ( n2912 , n2202 , n1029 );
nor ( n2913 , n2911 , n2912 );
not ( n2914 , n2913 );
and ( n2915 , n2397 , n2395 );
not ( n2916 , n2397 );
and ( n2917 , n2916 , n1823 );
nor ( n2918 , n2915 , n2917 );
nand ( n2919 , n2918 , n2192 );
and ( n2920 , n2301 , n2278 );
not ( n2921 , n2301 );
and ( n2922 , n2921 , n2277 );
nor ( n2923 , n2920 , n2922 );
nand ( n2924 , n2923 , n2342 );
not ( n2925 , n995 );
not ( n2926 , n2124 );
nor ( n2927 , n2926 , n1947 );
not ( n2928 , n2927 );
or ( n2929 , n2925 , n2928 );
not ( n2930 , n2082 );
not ( n2931 , n2930 );
or ( n2932 , n2931 , n2366 );
nor ( n2933 , n1946 , n2124 );
nand ( n2934 , n2932 , n2084 , n2933 );
nand ( n2935 , n2929 , n2934 );
nand ( n2936 , n2935 , n1999 );
nand ( n2937 , n2919 , n2924 , n2936 );
not ( n2938 , n2937 );
not ( n2939 , n2938 );
or ( n2940 , n2914 , n2939 );
nor ( n2941 , n2214 , n2233 );
not ( n2942 , n2229 );
nand ( n2943 , n2941 , n2942 );
not ( n2944 , n2943 );
nand ( n2945 , n2940 , n2944 );
not ( n2946 , n2212 );
not ( n2947 , n2946 );
not ( n2948 , n2943 );
or ( n2949 , n2947 , n2948 );
not ( n2950 , n1946 );
not ( n2951 , n1951 );
and ( n2952 , n2950 , n2951 );
nor ( n2953 , n2952 , n2213 );
nand ( n2954 , n2949 , n2953 );
nand ( n2955 , n2954 , n49 );
or ( n2956 , n2244 , n51 );
not ( n2957 , n2245 );
nand ( n2958 , n2956 , n2957 );
not ( n2959 , n2958 );
not ( n2960 , n2216 );
nand ( n2961 , n2959 , n2960 );
nand ( n2962 , n2945 , n2955 , n2961 );
and ( n2963 , n2937 , n2128 );
and ( n2964 , n1697 , n51 );
nor ( n2965 , n2963 , n2964 );
not ( n2966 , n2958 );
nand ( n2967 , n2966 , n2242 );
nand ( n2968 , n2348 , n2910 );
nand ( n2969 , n2412 , n1029 );
nand ( n2970 , n2965 , n2967 , n2968 , n2969 );
xor ( n2971 , n2774 , n2770 );
nand ( n2972 , n2971 , n2783 );
not ( n2973 , n2582 );
nand ( n2974 , n2594 , n2125 );
not ( n2975 , n2974 );
nand ( n2976 , n2973 , n2975 );
and ( n2977 , n2791 , n222 );
and ( n2978 , n1697 , n115 );
nor ( n2979 , n2977 , n2978 );
xor ( n2980 , n2584 , n2581 );
nand ( n2981 , n2597 , n2980 );
nand ( n2982 , n2972 , n2976 , n2979 , n2981 );
not ( n2983 , n2347 );
not ( n2984 , n2411 );
not ( n2985 , n2984 );
or ( n2986 , n2983 , n2985 );
nand ( n2987 , n2986 , n1084 );
nand ( n2988 , n2241 , n161 );
nand ( n2989 , n2988 , n146 );
nand ( n2990 , n1126 , n1085 );
not ( n2991 , n2990 );
not ( n2992 , n2188 );
not ( n2993 , n2992 );
or ( n2994 , n2991 , n2993 );
and ( n2995 , n2076 , n1120 );
nor ( n2996 , n2995 , n2077 );
and ( n2997 , n2933 , n2996 );
nand ( n2998 , n2997 , n1999 );
nand ( n2999 , n2994 , n2998 );
nand ( n3000 , n2128 , n2999 );
nand ( n3001 , n2987 , n2989 , n3000 );
not ( n3002 , n2933 );
nor ( n3003 , n3002 , n2079 );
not ( n3004 , n2078 );
not ( n3005 , n1147 );
nand ( n3006 , n3004 , n3005 );
and ( n3007 , n3003 , n3006 );
not ( n3008 , n1120 );
and ( n3009 , n2927 , n3008 );
nor ( n3010 , n3007 , n3009 );
and ( n3011 , n2291 , n1064 );
not ( n3012 , n2291 );
and ( n3013 , n3012 , n1065 );
nor ( n3014 , n3011 , n3013 );
and ( n3015 , n2342 , n3014 );
not ( n3016 , n2350 );
and ( n3017 , n3016 , n1062 );
nor ( n3018 , n3017 , n2351 );
not ( n3019 , n3018 );
nor ( n3020 , n3019 , n2345 );
nor ( n3021 , n3015 , n3020 );
nand ( n3022 , n3010 , n3021 );
not ( n3023 , n1999 );
nand ( n3024 , n3023 , n3021 );
and ( n3025 , n3022 , n3024 );
or ( n3026 , n1065 , n1129 );
nand ( n3027 , n3026 , n1130 );
nor ( n3028 , n2193 , n3027 );
nor ( n3029 , n3025 , n3028 );
not ( n3030 , n3029 );
nand ( n3031 , n3030 , n2128 );
not ( n3032 , n1058 );
nand ( n3033 , n3032 , n2411 );
nand ( n3034 , n2988 , n154 );
nand ( n3035 , n3031 , n3033 , n3034 );
and ( n3036 , n2352 , n1007 );
nor ( n3037 , n3036 , n2353 );
and ( n3038 , n2348 , n3037 );
xor ( n3039 , n47 , n39 );
and ( n3040 , n2242 , n3039 );
nor ( n3041 , n3038 , n3040 );
not ( n3042 , n1008 );
nand ( n3043 , n3042 , n2412 );
not ( n3044 , n2155 );
not ( n3045 , n1169 );
not ( n3046 , n3045 );
or ( n3047 , n3044 , n3046 );
or ( n3048 , n3045 , n2155 );
nand ( n3049 , n3047 , n3048 );
and ( n3050 , n2194 , n3049 );
not ( n3051 , n3005 );
not ( n3052 , n3051 );
not ( n3053 , n2927 );
or ( n3054 , n3052 , n3053 );
nand ( n3055 , n2081 , n1014 );
nand ( n3056 , n2930 , n3055 , n2933 );
nand ( n3057 , n3054 , n3056 );
nand ( n3058 , n3057 , n1999 );
nor ( n3059 , n2285 , n2298 );
not ( n3060 , n3059 );
nand ( n3061 , n3060 , n2342 , n2299 );
and ( n3062 , n3058 , n3061 );
or ( n3063 , n3062 , n2182 );
nand ( n3064 , n1697 , n47 );
nand ( n3065 , n3063 , n3064 );
nor ( n3066 , n3050 , n3065 );
nand ( n3067 , n3041 , n3043 , n3066 );
or ( n3068 , n2902 , n1163 );
or ( n3069 , n39 , n2243 );
and ( n3070 , n2351 , n1163 );
not ( n3071 , n2351 );
not ( n3072 , n1163 );
and ( n3073 , n3071 , n3072 );
nor ( n3074 , n3070 , n3073 );
and ( n3075 , n2348 , n3074 );
not ( n3076 , n2192 );
nor ( n3077 , n1132 , n1168 );
not ( n3078 , n3077 );
not ( n3079 , n1169 );
nand ( n3080 , n3078 , n3079 );
or ( n3081 , n3076 , n3080 );
not ( n3082 , n2079 );
and ( n3083 , n3082 , n994 );
nor ( n3084 , n3083 , n2595 );
buf ( n3085 , n2081 );
and ( n3086 , n3084 , n3085 );
and ( n3087 , n2295 , n2124 );
nor ( n3088 , n3086 , n3087 );
or ( n3089 , n3088 , n1954 );
nand ( n3090 , n3081 , n3089 );
not ( n3091 , n2297 );
nand ( n3092 , n3091 , n1168 );
not ( n3093 , n3092 );
nor ( n3094 , n3093 , n2298 );
and ( n3095 , n3094 , n2342 );
nor ( n3096 , n3090 , n3095 );
or ( n3097 , n3096 , n2182 );
nand ( n3098 , n1697 , n39 );
nand ( n3099 , n3097 , n3098 );
nor ( n3100 , n3075 , n3099 );
nand ( n3101 , n3068 , n3069 , n3100 );
nand ( n3102 , n2988 , n150 );
not ( n3103 , n1112 );
nand ( n3104 , n3103 , n2411 );
not ( n3105 , n1077 );
not ( n3106 , n2927 );
or ( n3107 , n3105 , n3106 );
not ( n3108 , n2077 );
not ( n3109 , n2295 );
and ( n3110 , n3108 , n3109 );
nor ( n3111 , n3110 , n2078 );
nand ( n3112 , n3111 , n2933 );
nand ( n3113 , n3107 , n3112 );
nand ( n3114 , n3113 , n1999 );
buf ( n3115 , n1116 );
xnor ( n3116 , n3115 , n1085 );
not ( n3117 , n3116 );
nand ( n3118 , n3117 , n2192 );
not ( n3119 , n2289 );
not ( n3120 , n3115 );
or ( n3121 , n3119 , n3120 );
or ( n3122 , n3115 , n2289 );
nand ( n3123 , n3121 , n3122 );
and ( n3124 , n2342 , n3123 );
and ( n3125 , n1113 , n1084 );
nor ( n3126 , n3125 , n2350 );
not ( n3127 , n3126 );
nor ( n3128 , n3127 , n2345 );
nor ( n3129 , n3124 , n3128 );
nand ( n3130 , n3114 , n3118 , n3129 );
nand ( n3131 , n2128 , n3130 );
nand ( n3132 , n3102 , n3104 , n3131 );
not ( n3133 , n52 );
and ( n3134 , n2953 , n2211 );
nor ( n3135 , n2229 , n2234 );
nand ( n3136 , n3134 , n3135 );
not ( n3137 , n3136 );
not ( n3138 , n3137 );
not ( n3139 , n3138 );
or ( n3140 , n3133 , n3139 );
not ( n3141 , n2918 );
not ( n3142 , n2191 );
nand ( n3143 , n3142 , n2199 );
buf ( n3144 , n3143 );
nor ( n3145 , n3141 , n3144 );
not ( n3146 , n2935 );
nand ( n3147 , n3146 , n2924 , n2913 );
nor ( n3148 , n3145 , n3147 );
or ( n3149 , n3148 , n3138 );
nand ( n3150 , n3140 , n3149 );
not ( n3151 , n50 );
nor ( n3152 , n2942 , n2234 );
nand ( n3153 , n3134 , n3152 );
not ( n3154 , n3153 );
or ( n3155 , n3151 , n3154 );
or ( n3156 , n3148 , n3153 );
nand ( n3157 , n3155 , n3156 );
not ( n3158 , n48 );
not ( n3159 , n2954 );
or ( n3160 , n3158 , n3159 );
and ( n3161 , n2960 , n3039 );
not ( n3162 , n2192 );
not ( n3163 , n3049 );
or ( n3164 , n3162 , n3163 );
nand ( n3165 , n3164 , n3058 );
and ( n3166 , n2346 , n3037 );
and ( n3167 , n2202 , n1007 );
nor ( n3168 , n3166 , n3167 );
nand ( n3169 , n3061 , n3168 );
nor ( n3170 , n3165 , n3169 );
nor ( n3171 , n3170 , n2943 );
nor ( n3172 , n3161 , n3171 );
nand ( n3173 , n3160 , n3172 );
not ( n3174 , n37 );
not ( n3175 , n2954 );
or ( n3176 , n3174 , n3175 );
not ( n3177 , n2216 );
not ( n3178 , n39 );
and ( n3179 , n3177 , n3178 );
nand ( n3180 , n2202 , n3072 );
not ( n3181 , n2345 );
nand ( n3182 , n3181 , n3074 );
and ( n3183 , n3180 , n3182 );
nand ( n3184 , n3096 , n3183 );
and ( n3185 , n3184 , n2944 );
nor ( n3186 , n3179 , n3185 );
nand ( n3187 , n3176 , n3186 );
not ( n3188 , n2613 );
not ( n3189 , n2766 );
or ( n3190 , n3188 , n3189 );
or ( n3191 , n2766 , n2613 );
nand ( n3192 , n3190 , n3191 );
and ( n3193 , n3192 , n2782 );
and ( n3194 , n1697 , n119 );
nor ( n3195 , n3193 , n3194 );
nand ( n3196 , n2975 , n1502 );
nand ( n3197 , n2791 , n223 );
xor ( n3198 , n2577 , n2419 );
nand ( n3199 , n3198 , n2597 );
nand ( n3200 , n3195 , n3196 , n3197 , n3199 );
not ( n3201 , n3136 );
not ( n3202 , n3144 );
nand ( n3203 , n3201 , n3202 );
not ( n3204 , n3203 );
not ( n3205 , n3204 );
not ( n3206 , n3049 );
or ( n3207 , n3205 , n3206 );
or ( n3208 , n3169 , n3057 );
and ( n3209 , n3137 , n3208 );
not ( n3210 , n3137 );
and ( n3211 , n3210 , n45 );
nor ( n3212 , n3209 , n3211 );
nand ( n3213 , n3207 , n3212 );
not ( n3214 , n155 );
not ( n3215 , n2954 );
or ( n3216 , n3214 , n3215 );
nand ( n3217 , n2202 , n1062 );
nand ( n3218 , n3029 , n3217 );
and ( n3219 , n3218 , n2944 );
not ( n3220 , n2216 );
and ( n3221 , n3220 , n154 );
nor ( n3222 , n3219 , n3221 );
nand ( n3223 , n3216 , n3222 );
or ( n3224 , n3203 , n3080 );
not ( n3225 , n3136 );
or ( n3226 , n3225 , n1138 );
not ( n3227 , n3095 );
not ( n3228 , n3088 );
nand ( n3229 , n3228 , n1948 );
nand ( n3230 , n3227 , n3183 , n3229 );
nand ( n3231 , n3225 , n3230 );
nand ( n3232 , n3224 , n3226 , n3231 );
or ( n3233 , n3203 , n3027 );
or ( n3234 , n3225 , n1037 );
not ( n3235 , n3022 );
nand ( n3236 , n3235 , n3217 );
nand ( n3237 , n3225 , n3236 );
nand ( n3238 , n3233 , n3234 , n3237 );
or ( n3239 , n3203 , n3116 );
not ( n3240 , n151 );
or ( n3241 , n3137 , n3240 );
not ( n3242 , n3113 );
nand ( n3243 , n2202 , n1113 );
nand ( n3244 , n3242 , n3129 , n3243 );
nand ( n3245 , n3244 , n3201 );
nand ( n3246 , n3239 , n3241 , n3245 );
not ( n3247 , n153 );
not ( n3248 , n2954 );
or ( n3249 , n3247 , n3248 );
not ( n3250 , n2216 );
not ( n3251 , n150 );
not ( n3252 , n3251 );
and ( n3253 , n3250 , n3252 );
not ( n3254 , n3130 );
nand ( n3255 , n3254 , n3243 );
and ( n3256 , n3255 , n2944 );
nor ( n3257 , n3253 , n3256 );
nand ( n3258 , n3249 , n3257 );
not ( n3259 , n2596 );
not ( n3260 , n2425 );
not ( n3261 , n2572 );
not ( n3262 , n3261 );
or ( n3263 , n3260 , n3262 );
or ( n3264 , n3261 , n2425 );
nand ( n3265 , n3263 , n3264 );
nand ( n3266 , n3259 , n3265 );
not ( n3267 , n1487 );
nand ( n3268 , n3267 , n2975 );
xor ( n3269 , n2620 , n2762 );
buf ( n3270 , n2781 );
and ( n3271 , n3269 , n3270 );
and ( n3272 , n1697 , n123 );
nor ( n3273 , n3271 , n3272 );
nand ( n3274 , n2791 , n224 );
nand ( n3275 , n3266 , n3268 , n3273 , n3274 );
not ( n3276 , n147 );
not ( n3277 , n2954 );
or ( n3278 , n3276 , n3277 );
and ( n3279 , n3220 , n146 );
nand ( n3280 , n2208 , n1084 );
not ( n3281 , n3280 );
nor ( n3282 , n2999 , n3281 );
nor ( n3283 , n3282 , n2943 );
nor ( n3284 , n3279 , n3283 );
nand ( n3285 , n3278 , n3284 );
not ( n3286 , n149 );
not ( n3287 , n3136 );
or ( n3288 , n3286 , n3287 );
not ( n3289 , n2342 );
nand ( n3290 , n3289 , n3143 );
nand ( n3291 , n3290 , n2990 );
not ( n3292 , n2997 );
and ( n3293 , n3291 , n3280 , n3292 );
or ( n3294 , n3293 , n3136 );
nand ( n3295 , n3288 , n3294 );
not ( n3296 , n2483 );
and ( n3297 , n2597 , n3296 );
not ( n3298 , n2677 );
and ( n3299 , n2782 , n3298 );
nor ( n3300 , n3297 , n3299 );
not ( n3301 , n1107 );
or ( n3302 , n3300 , n3301 );
nor ( n3303 , n2596 , n3296 );
not ( n3304 , n2677 );
not ( n3305 , n2781 );
or ( n3306 , n3304 , n3305 );
nand ( n3307 , n3306 , n2974 );
or ( n3308 , n3303 , n3307 );
nand ( n3309 , n3308 , n3301 );
not ( n3310 , n3251 );
not ( n3311 , n161 );
and ( n3312 , n3310 , n3311 );
buf ( n3313 , n2790 );
and ( n3314 , n3313 , n239 );
nor ( n3315 , n3312 , n3314 );
nand ( n3316 , n3302 , n3309 , n3315 );
or ( n3317 , n6 , n147 );
not ( n3318 , n2596 );
nand ( n3319 , n3317 , n2478 , n3318 );
nand ( n3320 , n2975 , n6 );
not ( n3321 , n6 );
and ( n3322 , n3321 , n1067 );
not ( n3323 , n2672 );
nor ( n3324 , n3322 , n3323 );
and ( n3325 , n3324 , n2782 );
not ( n3326 , n240 );
not ( n3327 , n2790 );
or ( n3328 , n3326 , n3327 );
nand ( n3329 , n1697 , n146 );
nand ( n3330 , n3328 , n3329 );
nor ( n3331 , n3325 , n3330 );
nand ( n3332 , n3319 , n3320 , n3331 );
and ( n3333 , n3153 , n1067 );
not ( n3334 , n3153 );
and ( n3335 , n3334 , n3293 );
nor ( n3336 , n3333 , n3335 );
buf ( n3337 , n2781 );
not ( n3338 , n2626 );
not ( n3339 , n2758 );
not ( n3340 , n3339 );
or ( n3341 , n3338 , n3340 );
or ( n3342 , n3339 , n2626 );
nand ( n3343 , n3341 , n3342 );
and ( n3344 , n3337 , n3343 );
and ( n3345 , n1697 , n77 );
nor ( n3346 , n3344 , n3345 );
nand ( n3347 , n2570 , n2975 );
nand ( n3348 , n2791 , n225 );
not ( n3349 , n2567 );
nand ( n3350 , n3349 , n2432 );
not ( n3351 , n3350 );
not ( n3352 , n2432 );
nand ( n3353 , n3352 , n2567 );
not ( n3354 , n3353 );
or ( n3355 , n3351 , n3354 );
not ( n3356 , n2596 );
nand ( n3357 , n3355 , n3356 );
nand ( n3358 , n3346 , n3347 , n3348 , n3357 );
nand ( n3359 , n2791 , n232 );
nand ( n3360 , n2975 , n2459 );
not ( n3361 , n2714 );
nand ( n3362 , n2707 , n2654 );
not ( n3363 , n3362 );
or ( n3364 , n3361 , n3363 );
nand ( n3365 , n3364 , n2648 );
xor ( n3366 , n3365 , n2727 );
and ( n3367 , n3337 , n3366 );
nor ( n3368 , n3367 , n2870 );
buf ( n3369 , n2513 );
or ( n3370 , n3369 , n2520 );
nand ( n3371 , n3370 , n2458 );
xor ( n3372 , n3371 , n2527 );
nand ( n3373 , n3318 , n3372 );
nand ( n3374 , n3359 , n3360 , n3368 , n3373 );
nand ( n3375 , n2791 , n226 );
not ( n3376 , n2434 );
nand ( n3377 , n3376 , n2975 );
not ( n3378 , n2632 );
not ( n3379 , n2754 );
not ( n3380 , n3379 );
or ( n3381 , n3378 , n3380 );
or ( n3382 , n3379 , n2632 );
nand ( n3383 , n3381 , n3382 );
and ( n3384 , n2782 , n3383 );
and ( n3385 , n1697 , n83 );
nor ( n3386 , n3384 , n3385 );
not ( n3387 , n2439 );
nand ( n3388 , n3387 , n2563 );
not ( n3389 , n3388 );
not ( n3390 , n2563 );
nand ( n3391 , n3390 , n2439 );
not ( n3392 , n3391 );
or ( n3393 , n3389 , n3392 );
nand ( n3394 , n3393 , n3356 );
nand ( n3395 , n3375 , n3377 , n3386 , n3394 );
not ( n3396 , n2638 );
not ( n3397 , n2750 );
not ( n3398 , n3397 );
or ( n3399 , n3396 , n3398 );
or ( n3400 , n3397 , n2638 );
nand ( n3401 , n3399 , n3400 );
and ( n3402 , n3401 , n3337 );
and ( n3403 , n1697 , n71 );
nor ( n3404 , n3402 , n3403 );
not ( n3405 , n2441 );
nand ( n3406 , n3405 , n2975 );
not ( n3407 , n2446 );
nand ( n3408 , n3407 , n2559 );
not ( n3409 , n3408 );
not ( n3410 , n2559 );
nand ( n3411 , n3410 , n2446 );
not ( n3412 , n3411 );
or ( n3413 , n3409 , n3412 );
nand ( n3414 , n3413 , n3356 );
nand ( n3415 , n2791 , n227 );
nand ( n3416 , n3404 , n3406 , n3414 , n3415 );
xor ( n3417 , n2746 , n2644 );
and ( n3418 , n3337 , n3417 );
and ( n3419 , n1697 , n75 );
nor ( n3420 , n3418 , n3419 );
not ( n3421 , n1359 );
nand ( n3422 , n3421 , n2975 );
nand ( n3423 , n2791 , n228 );
not ( n3424 , n2452 );
nand ( n3425 , n3424 , n2554 );
not ( n3426 , n3425 );
not ( n3427 , n2554 );
nand ( n3428 , n3427 , n2452 );
not ( n3429 , n3428 );
or ( n3430 , n3426 , n3429 );
not ( n3431 , n2596 );
nand ( n3432 , n3430 , n3431 );
nand ( n3433 , n3420 , n3422 , n3423 , n3432 );
not ( n3434 , n2741 );
and ( n3435 , n3365 , n2727 );
nor ( n3436 , n3435 , n2646 );
or ( n3437 , n3436 , n2735 );
nand ( n3438 , n3437 , n2650 );
and ( n3439 , n3438 , n2722 );
nor ( n3440 , n3439 , n2724 );
not ( n3441 , n3440 );
or ( n3442 , n3434 , n3441 );
or ( n3443 , n3440 , n2741 );
nand ( n3444 , n3442 , n3443 );
and ( n3445 , n3444 , n2782 );
and ( n3446 , n1697 , n67 );
nor ( n3447 , n3445 , n3446 );
not ( n3448 , n1340 );
nand ( n3449 , n3448 , n2975 );
and ( n3450 , n3371 , n2527 );
not ( n3451 , n2460 );
nor ( n3452 , n3450 , n3451 );
not ( n3453 , n2544 );
or ( n3454 , n3452 , n3453 );
nand ( n3455 , n3454 , n2455 );
not ( n3456 , n2535 );
and ( n3457 , n3455 , n3456 );
not ( n3458 , n2536 );
nor ( n3459 , n3457 , n3458 );
nand ( n3460 , n3459 , n2549 );
not ( n3461 , n3460 );
or ( n3462 , n3459 , n2549 );
not ( n3463 , n3462 );
or ( n3464 , n3461 , n3463 );
nand ( n3465 , n3464 , n3318 );
nand ( n3466 , n2791 , n229 );
nand ( n3467 , n3447 , n3449 , n3465 , n3466 );
nand ( n3468 , n2791 , n231 );
not ( n3469 , n2542 );
nand ( n3470 , n3469 , n2975 );
xor ( n3471 , n3436 , n2735 );
and ( n3472 , n3337 , n3471 );
not ( n3473 , n2832 );
nor ( n3474 , n3472 , n3473 );
xor ( n3475 , n3453 , n3452 );
nand ( n3476 , n3475 , n3318 );
nand ( n3477 , n3468 , n3470 , n3474 , n3476 );
xor ( n3478 , n3362 , n2714 );
and ( n3479 , n2782 , n3478 );
nor ( n3480 , n3479 , n2370 );
nand ( n3481 , n2975 , n2457 );
xor ( n3482 , n2520 , n3369 );
nand ( n3483 , n3482 , n3259 );
nand ( n3484 , n3313 , n233 );
nand ( n3485 , n3480 , n3481 , n3483 , n3484 );
nand ( n3486 , n2791 , n234 );
nand ( n3487 , n2975 , n1187 );
not ( n3488 , n2706 );
not ( n3489 , n2702 );
not ( n3490 , n3489 );
or ( n3491 , n3488 , n3490 );
or ( n3492 , n3489 , n2706 );
nand ( n3493 , n3491 , n3492 );
and ( n3494 , n3337 , n3493 );
not ( n3495 , n2876 );
nor ( n3496 , n3494 , n3495 );
not ( n3497 , n2505 );
nand ( n3498 , n3497 , n2510 );
not ( n3499 , n3498 );
not ( n3500 , n2510 );
nand ( n3501 , n3500 , n2505 );
not ( n3502 , n3501 );
or ( n3503 , n3499 , n3502 );
nand ( n3504 , n3503 , n3431 );
nand ( n3505 , n3486 , n3487 , n3496 , n3504 );
buf ( n3506 , n2119 );
buf ( n3507 , n1986 );
nand ( n3508 , n3506 , n3507 );
buf ( n3509 , n3508 );
not ( n3510 , n1959 );
or ( n3511 , n3510 , n148 );
or ( n3512 , n147 , n1959 );
nand ( n3513 , n3511 , n3512 , n2124 );
and ( n3514 , n3513 , n6 );
not ( n3515 , n3513 );
and ( n3516 , n3515 , n3321 );
nor ( n3517 , n3514 , n3516 );
nor ( n3518 , n3509 , n3517 );
not ( n3519 , n3064 );
nor ( n3520 , n3518 , n3519 );
nand ( n3521 , n1005 , n2975 );
not ( n3522 , n2665 );
not ( n3523 , n2694 );
not ( n3524 , n3523 );
or ( n3525 , n3522 , n3524 );
or ( n3526 , n3523 , n2665 );
nand ( n3527 , n3525 , n3526 );
and ( n3528 , n3270 , n3527 );
and ( n3529 , n2790 , n236 );
nor ( n3530 , n3528 , n3529 );
not ( n3531 , n2497 );
nand ( n3532 , n3531 , n2474 );
not ( n3533 , n3532 );
not ( n3534 , n2474 );
nand ( n3535 , n3534 , n2497 );
not ( n3536 , n3535 );
or ( n3537 , n3533 , n3536 );
nand ( n3538 , n3537 , n3259 );
nand ( n3539 , n3520 , n3521 , n3530 , n3538 );
nand ( n3540 , n2791 , n237 );
nand ( n3541 , n1160 , n2975 );
xor ( n3542 , n2690 , n2670 );
and ( n3543 , n3337 , n3542 );
not ( n3544 , n3098 );
nor ( n3545 , n3543 , n3544 );
not ( n3546 , n2476 );
nand ( n3547 , n3546 , n2493 );
not ( n3548 , n3547 );
not ( n3549 , n2493 );
nand ( n3550 , n3549 , n2476 );
not ( n3551 , n3550 );
or ( n3552 , n3548 , n3551 );
nand ( n3553 , n3552 , n3356 );
nand ( n3554 , n3540 , n3541 , n3545 , n3553 );
nand ( n3555 , n2791 , n230 );
not ( n3556 , n1306 );
nand ( n3557 , n3556 , n2975 );
xor ( n3558 , n3438 , n2722 );
and ( n3559 , n3337 , n3558 );
nor ( n3560 , n3559 , n2219 );
xor ( n3561 , n3455 , n3456 );
nand ( n3562 , n3561 , n3431 );
nand ( n3563 , n3555 , n3557 , n3560 , n3562 );
xor ( n3564 , n2698 , n2660 );
and ( n3565 , n2782 , n3564 );
nor ( n3566 , n3565 , n2964 );
nand ( n3567 , n2975 , n1024 );
xor ( n3568 , n2501 , n2468 );
nand ( n3569 , n3568 , n3431 );
nand ( n3570 , n3313 , n235 );
nand ( n3571 , n3566 , n3567 , n3569 , n3570 );
nor ( n3572 , n1041 , n161 );
nor ( n3573 , n3518 , n3572 );
not ( n3574 , n2682 );
nand ( n3575 , n3574 , n2975 );
xor ( n3576 , n2686 , n2680 );
and ( n3577 , n3270 , n3576 );
and ( n3578 , n2790 , n238 );
nor ( n3579 , n3577 , n3578 );
xor ( n3580 , n2489 , n2487 );
nand ( n3581 , n3580 , n3259 );
nand ( n3582 , n3573 , n3575 , n3579 , n3581 );
not ( n3583 , n177 );
and ( n3584 , n3509 , n3583 );
not ( n3585 , n3509 );
and ( n3586 , n3585 , n956 );
nor ( n3587 , n3584 , n3586 );
or ( n3588 , n961 , n3509 );
nand ( n3589 , n3509 , n178 );
nand ( n3590 , n3588 , n3589 );
not ( n3591 , n160 );
or ( n3592 , n2215 , n3591 );
not ( n3593 , n2941 );
nand ( n3594 , n3592 , n3593 );
buf ( n3595 , n3508 );
or ( n3596 , n3595 , n1435 );
nand ( n3597 , n3509 , n207 );
nand ( n3598 , n3596 , n3597 );
or ( n3599 , n3509 , n1559 );
nand ( n3600 , n3509 , n210 );
nand ( n3601 , n3599 , n3600 );
or ( n3602 , n3509 , n1495 );
nand ( n3603 , n3595 , n208 );
nand ( n3604 , n3602 , n3603 );
or ( n3605 , n3509 , n1521 );
nand ( n3606 , n3509 , n203 );
nand ( n3607 , n3605 , n3606 );
or ( n3608 , n3509 , n1602 );
nand ( n3609 , n3509 , n179 );
nand ( n3610 , n3608 , n3609 );
or ( n3611 , n3509 , n979 );
nand ( n3612 , n3509 , n176 );
nand ( n3613 , n3611 , n3612 );
or ( n3614 , n3595 , n1667 );
nand ( n3615 , n3595 , n173 );
nand ( n3616 , n3614 , n3615 );
or ( n3617 , n3595 , n1472 );
nand ( n3618 , n3509 , n204 );
nand ( n3619 , n3617 , n3618 );
or ( n3620 , n3595 , n1689 );
nand ( n3621 , n3595 , n205 );
nand ( n3622 , n3620 , n3621 );
or ( n3623 , n3595 , n994 );
nand ( n3624 , n3595 , n241 );
nand ( n3625 , n3623 , n3624 );
or ( n3626 , n3595 , n1120 );
nand ( n3627 , n3595 , n244 );
nand ( n3628 , n3626 , n3627 );
or ( n3629 , n3509 , n1516 );
nand ( n3630 , n3509 , n181 );
nand ( n3631 , n3629 , n3630 );
or ( n3632 , n3595 , n1481 );
nand ( n3633 , n3595 , n209 );
nand ( n3634 , n3632 , n3633 );
or ( n3635 , n3595 , n1385 );
nand ( n3636 , n3509 , n211 );
nand ( n3637 , n3635 , n3636 );
or ( n3638 , n3595 , n1375 );
nand ( n3639 , n3509 , n212 );
nand ( n3640 , n3638 , n3639 );
or ( n3641 , n3595 , n1329 );
nand ( n3642 , n3595 , n213 );
nand ( n3643 , n3641 , n3642 );
or ( n3644 , n3595 , n1320 );
nand ( n3645 , n3509 , n214 );
nand ( n3646 , n3644 , n3645 );
or ( n3647 , n3595 , n2133 );
nand ( n3648 , n3509 , n215 );
nand ( n3649 , n3647 , n3648 );
or ( n3650 , n3595 , n1239 );
nand ( n3651 , n3595 , n216 );
nand ( n3652 , n3650 , n3651 );
or ( n3653 , n3595 , n2086 );
nand ( n3654 , n3595 , n217 );
nand ( n3655 , n3653 , n3654 );
or ( n3656 , n3509 , n1574 );
nand ( n3657 , n3509 , n218 );
nand ( n3658 , n3656 , n3657 );
or ( n3659 , n3595 , n1177 );
nand ( n3660 , n3595 , n219 );
nand ( n3661 , n3659 , n3660 );
or ( n3662 , n3595 , n1014 );
nand ( n3663 , n3509 , n220 );
nand ( n3664 , n3662 , n3663 );
and ( n3665 , n3506 , n3507 );
nor ( n3666 , n2790 , n3665 );
or ( n3667 , n3005 , n3595 );
nand ( n3668 , n3595 , n242 );
nand ( n3669 , n3667 , n3668 );
or ( n3670 , n1061 , n3595 );
nand ( n3671 , n3595 , n243 );
nand ( n3672 , n3670 , n3671 );
or ( n3673 , n3509 , n1465 );
nand ( n3674 , n3509 , n180 );
nand ( n3675 , n3673 , n3674 );
or ( n3676 , n3595 , n1078 );
nand ( n3677 , n3595 , n245 );
nand ( n3678 , n3676 , n3677 );
or ( n3679 , n2101 , n1697 );
not ( n3680 , n193 );
or ( n3681 , n3680 , n161 );
nand ( n3682 , n3679 , n3681 );
not ( n3683 , n201 );
not ( n3684 , n1697 );
or ( n3685 , n3683 , n3684 );
or ( n3686 , n1452 , n1697 );
nand ( n3687 , n3685 , n3686 );
not ( n3688 , n198 );
not ( n3689 , n1697 );
or ( n3690 , n3688 , n3689 );
nand ( n3691 , n3690 , n899 );
not ( n3692 , n200 );
not ( n3693 , n1697 );
or ( n3694 , n3692 , n3693 );
or ( n3695 , n2417 , n1697 );
nand ( n3696 , n3694 , n3695 );
not ( n3697 , n182 );
not ( n3698 , n1697 );
or ( n3699 , n3697 , n3698 );
or ( n3700 , n2427 , n1697 );
nand ( n3701 , n3699 , n3700 );
not ( n3702 , n183 );
not ( n3703 , n1697 );
or ( n3704 , n3702 , n3703 );
or ( n3705 , n2434 , n1697 );
nand ( n3706 , n3704 , n3705 );
not ( n3707 , n184 );
not ( n3708 , n1697 );
or ( n3709 , n3707 , n3708 );
or ( n3710 , n2441 , n1697 );
nand ( n3711 , n3709 , n3710 );
not ( n3712 , n185 );
not ( n3713 , n1697 );
or ( n3714 , n3712 , n3713 );
or ( n3715 , n1359 , n1697 );
nand ( n3716 , n3714 , n3715 );
not ( n3717 , n162 );
not ( n3718 , n1697 );
or ( n3719 , n3717 , n3718 );
or ( n3720 , n1306 , n1697 );
nand ( n3721 , n3719 , n3720 );
not ( n3722 , n1140 );
and ( n3723 , n3722 , n161 );
and ( n3724 , n1697 , n187 );
nor ( n3725 , n3723 , n3724 );
not ( n3726 , n3725 );
and ( n3727 , n2457 , n161 );
and ( n3728 , n1697 , n165 );
nor ( n3729 , n3727 , n3728 );
not ( n3730 , n3729 );
not ( n3731 , n186 );
not ( n3732 , n1697 );
or ( n3733 , n3731 , n3732 );
or ( n3734 , n1340 , n1697 );
nand ( n3735 , n3733 , n3734 );
not ( n3736 , n189 );
not ( n3737 , n1697 );
or ( n3738 , n3736 , n3737 );
or ( n3739 , n410 , n1697 );
nand ( n3740 , n3738 , n3739 );
not ( n3741 , n163 );
not ( n3742 , n1697 );
or ( n3743 , n3741 , n3742 );
or ( n3744 , n2542 , n1697 );
nand ( n3745 , n3743 , n3744 );
not ( n3746 , n188 );
not ( n3747 , n1697 );
or ( n3748 , n3746 , n3747 );
or ( n3749 , n2125 , n1697 );
nand ( n3750 , n3748 , n3749 );
not ( n3751 , n192 );
not ( n3752 , n1697 );
or ( n3753 , n3751 , n3752 );
or ( n3754 , n1984 , n1697 );
nand ( n3755 , n3753 , n3754 );
not ( n3756 , n190 );
not ( n3757 , n1697 );
or ( n3758 , n3756 , n3757 );
not ( n3759 , n377 );
nand ( n3760 , n3759 , n378 , n1 , n161 );
nand ( n3761 , n3758 , n3760 );
not ( n3762 , n164 );
not ( n3763 , n1697 );
or ( n3764 , n3762 , n3763 );
or ( n3765 , n1248 , n1697 );
nand ( n3766 , n3764 , n3765 );
and ( n3767 , n3509 , n206 );
not ( n3768 , n3509 );
and ( n3769 , n3768 , n754 );
or ( n3770 , n3767 , n3769 );
and ( n3771 , n2215 , n2942 );
not ( n3772 , n2215 );
and ( n3773 , n3772 , n2114 );
nor ( n3774 , n3771 , n3773 );
and ( n3775 , n3509 , n174 );
not ( n3776 , n3509 );
and ( n3777 , n3776 , n800 );
or ( n3778 , n3775 , n3777 );
not ( n3779 , n3509 );
not ( n3780 , n175 );
or ( n3781 , n3779 , n3780 );
or ( n3782 , n970 , n3595 );
nand ( n3783 , n3781 , n3782 );
endmodule

