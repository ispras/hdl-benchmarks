// IWLS benchmark module "MinMax9b" printed on Wed May 29 22:12:32 2002
module MinMax9b(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \39 , \40 , \41 , \42 , \43 , \44 , \45 , \46 , \47 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ;
output
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ;
reg
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ;
wire
  \437 ,
  \438 ,
  \439 ,
  \[59] ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \462 ,
  \470 ,
  \478 ,
  \486 ,
  \494 ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \502 ,
  \510 ,
  \518 ,
  \[67] ,
  \526 ,
  \[68] ,
  \531 ,
  \536 ,
  \541 ,
  \546 ,
  \105 ,
  \107 ,
  \109 ,
  \551 ,
  \111 ,
  \113 ,
  \556 ,
  \115 ,
  \117 ,
  \561 ,
  \566 ,
  \571 ,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[76] ,
  \[78] ,
  \[35] ,
  \643 ,
  \[36] ,
  \651 ,
  \659 ,
  \[37] ,
  \667 ,
  \[38] ,
  \675 ,
  \[39] ,
  \683 ,
  \691 ,
  \699 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \710 ,
  \[87] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \83 ,
  \85 ,
  \87 ,
  \[50] ,
  \89 ,
  \91 ,
  \93 ,
  \95 ,
  \97 ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \409 ,
  \[56] ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \418 ,
  \419 ,
  \[57] ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \428 ,
  \[58] ,
  \430 ,
  \431 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ;
assign
  \437  = (\[74]  & \6 ) | (\[68]  & \425 ),
  \438  = (\437  & \436 ) | ((\437  & \435 ) | (\436  & \435 )),
  \439  = (\[72]  & \7 ) | (\[71]  & \414 ),
  \[59]  = \699 ,
  \440  = (\[74]  & \7 ) | (\[68]  & \424 ),
  \441  = (\440  & \439 ) | ((\440  & \438 ) | (\439  & \438 )),
  \442  = (\[72]  & \8 ) | (\[71]  & \413 ),
  \443  = (\[74]  & \8 ) | (\[68]  & \423 ),
  \444  = (\443  & \442 ) | ((\443  & \441 ) | (\442  & \441 )),
  \445  = (\[72]  & \9 ) | (\[71]  & \412 ),
  \446  = (\[74]  & \9 ) | (\[68]  & \422 ),
  \447  = (\446  & \445 ) | ((\446  & \444 ) | (\445  & \444 )),
  \448  = (\[72]  & \10 ) | (\[71]  & \411 ),
  \449  = (\[74]  & \10 ) | (\[68]  & \421 ),
  \450  = (\449  & \448 ) | ((\449  & \447 ) | (\448  & \447 )),
  \451  = (\[72]  & \11 ) | (\[71]  & \410 ),
  \452  = (\[74]  & \11 ) | (\[68]  & \420 ),
  \453  = (\452  & \451 ) | ((\452  & \450 ) | (\451  & \450 )),
  \454  = (\[72]  & \12 ) | (\[71]  & \409 ),
  \455  = (\[74]  & \12 ) | (\[68]  & \419 ),
  \462  = (\651  & (\431  & (\430  & \434 ))) | ((~\[62]  & (~\435  & \434 )) | ((\643  & (\431  & ~\435 )) | ((\[61]  & \531 ) | (\651  & ~\435 )))),
  \470  = (~\[62]  & (~\438  & \437 )) | ((\659  & (\437  & \435 )) | ((~\438  & (\435  & ~\59 )) | ((\[61]  & \536 ) | (\659  & ~\438 )))),
  \478  = (~\[62]  & (~\441  & \440 )) | ((\667  & (\440  & \438 )) | ((~\441  & (\438  & ~\60 )) | ((\[61]  & \541 ) | (\667  & ~\441 )))),
  \486  = (~\[62]  & (~\444  & \443 )) | ((\675  & (\443  & \441 )) | ((~\444  & (\441  & ~\61 )) | ((\[61]  & \546 ) | (\675  & ~\444 )))),
  \494  = (~\[62]  & (~\447  & \446 )) | ((\683  & (\446  & \444 )) | ((~\447  & (\444  & ~\62 )) | ((\[61]  & \551 ) | (\683  & ~\447 )))),
  \[60]  = \710 ,
  \[61]  = \3  | ~\2 ,
  \[62]  = \[61]  | \1 ,
  \[63]  = \83  | ~\30 ,
  \502  = (~\[62]  & (~\450  & \449 )) | ((\691  & (\449  & \447 )) | ((~\450  & (\447  & ~\63 )) | ((\[61]  & \556 ) | (\691  & ~\450 )))),
  \510  = (~\[62]  & (\452  & ~\453 )) | ((\699  & (\452  & \450 )) | ((\450  & (~\453  & ~\64 )) | ((\[61]  & \561 ) | (\699  & ~\453 )))),
  \518  = (~\[76]  & (~\[62]  & ~\455 )) | ((\[76]  & (~\[62]  & \455 )) | (\[61]  & \566 )),
  \[67]  = ~\[62]  & ~\83 ,
  \526  = (~\[62]  & (\455  & \453 )) | ((~\[62]  & (\454  & \453 )) | ((\710  & (\455  & \454 )) | (\[61]  & \710 ))),
  \[68]  = ~\[62]  & \428 ,
  \531  = (\[73]  & \13 ) | (\[70]  & \4 ),
  \536  = (\[73]  & \14 ) | (\[70]  & \5 ),
  \541  = (\[73]  & \15 ) | (\[70]  & \6 ),
  \546  = (\[73]  & \16 ) | (\[70]  & \7 ),
  \105  = (~\419  & \12 ) | (\419  & ~\12 ),
  \107  = (~\420  & \11 ) | (\420  & ~\11 ),
  \109  = (~\421  & \10 ) | (\421  & ~\10 ),
  \551  = (\[73]  & \17 ) | (\[70]  & \8 ),
  \111  = (~\422  & \9 ) | (\422  & ~\9 ),
  \113  = (~\423  & \8 ) | (\423  & ~\8 ),
  \556  = (\[73]  & \18 ) | (\[70]  & \9 ),
  \115  = (~\424  & \7 ) | (\424  & ~\7 ),
  \117  = (~\425  & \6 ) | (\425  & ~\6 ),
  \561  = (\[73]  & \19 ) | (\[70]  & \10 ),
  \566  = (\[73]  & \20 ) | (\[70]  & \11 ),
  \571  = (\[73]  & \21 ) | (\[70]  & \12 ),
  \[70]  = \2  & ~\1 ,
  \[71]  = ~\[62]  & ~\418 ,
  \[72]  = ~\[62]  & \418 ,
  \[73]  = ~\2  & ~\1 ,
  \[74]  = ~\[62]  & ~\428 ,
  \[76]  = (~\454  & ~\453 ) | (\454  & \453 ),
  \[78]  = ~\[62]  & \83 ,
  \[35]  = \531 ,
  \643  = ~\[62]  & \430 ,
  \[36]  = \536 ,
  \651  = ~\[62]  & \433 ,
  \659  = ~\[62]  & \436 ,
  \[37]  = \541 ,
  \667  = ~\[62]  & \439 ,
  \[38]  = \546 ,
  \675  = ~\[62]  & \442 ,
  \[39]  = \551 ,
  \683  = ~\[62]  & \445 ,
  \691  = ~\[62]  & \448 ,
  \699  = ~\[62]  & \451 ,
  \[40]  = \556 ,
  \[41]  = \561 ,
  \[42]  = \566 ,
  \710  = (~\[62]  & (~\571  & \454 )) | ((\[61]  & \571 ) | (\571  & \455 )),
  \[87]  = \38  | \21 ,
  \[43]  = \571 ,
  \[44]  = \57 ,
  \[45]  = \58 ,
  \[46]  = \59 ,
  \[47]  = \60 ,
  \[48]  = \61 ,
  \[49]  = \62 ,
  \39  = \462 ,
  \40  = \470 ,
  \41  = \478 ,
  \42  = \486 ,
  \43  = \494 ,
  \44  = \502 ,
  \45  = \510 ,
  \46  = \518 ,
  \47  = \526 ,
  \57  = \[62]  | \431 ,
  \58  = \[62]  | \434 ,
  \59  = \[62]  | \437 ,
  \60  = \[62]  | \440 ,
  \61  = \[62]  | \443 ,
  \62  = \[62]  | \446 ,
  \63  = \[62]  | \449 ,
  \64  = \[62]  | \452 ,
  \83  = (~\[62]  & (\38  & (~\37  & (~\36  & (~\35  & (~\34  & (~\33  & (~\32  & (~\31  & (~\30  & (\29  & (\28  & (\27  & (\26  & (\25  & (\24  & (\23  & (\22  & \21 )))))))))))))))))) | (~\[87]  & (~\[62]  & (~\37  & (~\36  & (~\35  & (~\34  & (~\33  & (~\32  & (~\31  & (~\30  & (\29  & (\28  & (\27  & (\26  & (\25  & (\24  & (\23  & \22 ))))))))))))))))),
  \85  = (~\409  & \12 ) | (\409  & ~\12 ),
  \87  = (~\410  & \11 ) | (\410  & ~\11 ),
  \[50]  = \63 ,
  \89  = (~\411  & \10 ) | (\411  & ~\10 ),
  \91  = (~\412  & \9 ) | (\412  & ~\9 ),
  \93  = (~\413  & \8 ) | (\413  & ~\8 ),
  \95  = (~\414  & \7 ) | (\414  & ~\7 ),
  \97  = (~\415  & \6 ) | (\415  & ~\6 ),
  \[51]  = \64 ,
  \[52]  = \643 ,
  \[53]  = \651 ,
  \[54]  = \659 ,
  \[55]  = \667 ,
  \409  = \[87]  & \[67] ,
  \[56]  = \675 ,
  \410  = \[67]  & \37 ,
  \411  = \[67]  & \36 ,
  \412  = \[67]  & \35 ,
  \413  = \[67]  & \34 ,
  \414  = \[67]  & \33 ,
  \415  = \[67]  & \32 ,
  \416  = \[67]  & \31 ,
  \418  = (\[63]  & (~\[62]  & (~\416  & (~\97  & (~\95  & (~\93  & (~\91  & (~\89  & (~\87  & (~\85  & \4 )))))))))) | ((\[63]  & (~\[62]  & (~\97  & (~\95  & (~\93  & (~\91  & (~\89  & (~\87  & (~\85  & (\5  & \4 )))))))))) | ((~\[62]  & (~\416  & (~\97  & (~\95  & (~\93  & (~\91  & (~\89  & (~\87  & (~\85  & \5 ))))))))) | ((~\[62]  & (\97  & (~\95  & (~\93  & (~\91  & (~\89  & (~\87  & (~\85  & \6 )))))))) | ((~\[62]  & (\95  & (~\93  & (~\91  & (~\89  & (~\87  & (~\85  & \7 ))))))) | ((~\[62]  & (\93  & (~\91  & (~\89  & (~\87  & (~\85  & \8 )))))) | ((~\[62]  & (\91  & (~\89  & (~\87  & (~\85  & \9 ))))) | ((~\[62]  & (\89  & (~\87  & (~\85  & \10 )))) | ((~\[62]  & (\87  & (~\85  & \11 ))) | (~\[62]  & (\85  & \12 )))))))))),
  \419  = (\409  & (\38  & \21 )) | \[78] ,
  \[57]  = \683 ,
  \420  = (~\[62]  & \29 ) | \[78] ,
  \421  = (~\[62]  & \28 ) | \[78] ,
  \422  = (~\[62]  & \27 ) | \[78] ,
  \423  = (~\[62]  & \26 ) | \[78] ,
  \424  = (~\[62]  & \25 ) | \[78] ,
  \425  = (~\[62]  & \24 ) | \[78] ,
  \426  = (~\[62]  & \23 ) | \[78] ,
  \428  = (\[67]  & (~\426  & (~\117  & (~\115  & (~\113  & (~\111  & (~\109  & (~\107  & (~\105  & (~\22  & \4 )))))))))) | ((\[67]  & (~\117  & (~\115  & (~\113  & (~\111  & (~\109  & (~\107  & (~\105  & (~\22  & (\5  & \4 )))))))))) | ((~\[62]  & (~\426  & (~\117  & (~\115  & (~\113  & (~\111  & (~\109  & (~\107  & (~\105  & \5 ))))))))) | ((~\[62]  & (\117  & (~\115  & (~\113  & (~\111  & (~\109  & (~\107  & (~\105  & \6 )))))))) | ((~\[62]  & (\115  & (~\113  & (~\111  & (~\109  & (~\107  & (~\105  & \7 ))))))) | ((~\[62]  & (\113  & (~\111  & (~\109  & (~\107  & (~\105  & \8 )))))) | ((~\[62]  & (\111  & (~\109  & (~\107  & (~\105  & \9 ))))) | ((~\[62]  & (\109  & (~\107  & (~\105  & \10 )))) | ((~\[62]  & (\107  & (~\105  & \11 ))) | (~\[62]  & (\105  & \12 )))))))))),
  \[58]  = \691 ,
  \430  = (\[72]  & \4 ) | (\[71]  & ~\[63] ),
  \431  = (\[74]  & \4 ) | ((\[68]  & \83 ) | (\[68]  & \22 )),
  \433  = (\[72]  & \5 ) | (\[71]  & \416 ),
  \434  = (\[74]  & \5 ) | (\[68]  & \426 ),
  \435  = (\431  & (\430  & \434 )) | ((\431  & (\430  & \433 )) | (\434  & \433 )),
  \436  = (\[72]  & \6 ) | (\[71]  & \415 );
always begin
  \13  = \[35] ;
  \14  = \[36] ;
  \15  = \[37] ;
  \16  = \[38] ;
  \17  = \[39] ;
  \18  = \[40] ;
  \19  = \[41] ;
  \20  = \[42] ;
  \21  = \[43] ;
  \22  = \[44] ;
  \23  = \[45] ;
  \24  = \[46] ;
  \25  = \[47] ;
  \26  = \[48] ;
  \27  = \[49] ;
  \28  = \[50] ;
  \29  = \[51] ;
  \30  = \[52] ;
  \31  = \[53] ;
  \32  = \[54] ;
  \33  = \[55] ;
  \34  = \[56] ;
  \35  = \[57] ;
  \36  = \[58] ;
  \37  = \[59] ;
  \38  = \[60] ;
end
initial begin
  \13  = 0;
  \14  = 0;
  \15  = 0;
  \16  = 0;
  \17  = 0;
  \18  = 0;
  \19  = 0;
  \20  = 0;
  \21  = 0;
  \22  = 1;
  \23  = 1;
  \24  = 1;
  \25  = 1;
  \26  = 1;
  \27  = 1;
  \28  = 1;
  \29  = 1;
  \30  = 0;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
end
endmodule

