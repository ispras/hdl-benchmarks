// IWLS benchmark module "pair" printed on Wed May 29 17:27:53 2002
module pair(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0, q0, r0, s0, t0, u0, v0, w0, x0, y0, z0, a1, b1, c1, d1, e1, f1, g1, h1, i1, j1, k1, l1, m1, n1, o1, p1, q1, r1, s1, t1, u1, v1, w1, x1, y1, z1, a2, b2, c2, d2, e2, f2, g2, h2, i2, j2, k2, l2, m2, n2, o2, p2, q2, r2, s2, t2, u2, v2, w2, x2, y2, z2, a3, b3, c3, d3, e3, f3, g3, h3, i3, j3, k3, l3, m3, n3, o3, p3, q3, r3, s3, t3, u3, v3, w3, x3, y3, z3, a4, b4, c4, d4, e4, f4, g4, h4, i4, j4, k4, l4, m4, n4, o4, p4, q4, r4, s4, t4, u4, v4, w4, x4, y4, z4, a5, b5, c5, d5, e5, f5, g5, h5, i5, j5, k5, l5, m5, n5, o5, p5, q5, r5, s5, t5, u5, v5, w5, x5, y5, z5, a6, b6, c6, d6, e6, f6, g6, h6, i6, j6, k6, l6, m6, n6, o6, p6, q6, r6, s6, t6, u6, v6, w6, x6, y6, z6, a7, b7, c7, d7, e7, f7, g7, h7, i7, j7, k7, l7, m7, n7, o7, p7, q7, r7, s7, t7, u7, v7, w7, x7, y7, z7, a8, b8, c8, d8, e8, f8, g8, h8, i8, j8, k8, l8, m8, n8, o8, p8, q8, r8, s8, t8, u8, v8, w8, x8, y8, z8, a9, b9, c9, d9, e9, f9, g9, h9, i9, j9, k9, l9, m9, n9, o9, p9, q9, r9, s9, t9, u9, v9, w9, x9, y9, z9, a10, b10, c10, d10, e10, f10, g10, h10, i10, j10, k10, l10, m10, n10, o10, p10, q10, r10, s10, t10, u10, v10, w10, x10, y10);
input
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  y,
  z,
  a0,
  a1,
  a2,
  a3,
  a4,
  a5,
  b0,
  b1,
  b2,
  b3,
  b4,
  b5,
  c0,
  c1,
  c2,
  c3,
  c4,
  c5,
  d0,
  d1,
  d2,
  d3,
  d4,
  d5,
  e0,
  e1,
  e2,
  e3,
  e4,
  e5,
  f0,
  f1,
  f2,
  f3,
  f4,
  f5,
  g0,
  g1,
  g2,
  g3,
  g4,
  g5,
  h0,
  h1,
  h2,
  h3,
  h4,
  h5,
  i0,
  i1,
  i2,
  i3,
  i4,
  i5,
  j0,
  j1,
  j2,
  j3,
  j4,
  j5,
  k0,
  k1,
  k2,
  k3,
  k4,
  k5,
  l0,
  l1,
  l2,
  l3,
  l4,
  l5,
  m0,
  m1,
  m2,
  m3,
  m4,
  m5,
  n0,
  n1,
  n2,
  n3,
  n4,
  n5,
  o0,
  o1,
  o2,
  o3,
  o4,
  o5,
  p0,
  p1,
  p2,
  p3,
  p4,
  p5,
  q0,
  q1,
  q2,
  q3,
  q4,
  q5,
  r0,
  r1,
  r2,
  r3,
  r4,
  r5,
  s0,
  s1,
  s2,
  s3,
  s4,
  t0,
  t1,
  t2,
  t3,
  t4,
  u0,
  u1,
  u2,
  u3,
  u4,
  v0,
  v1,
  v2,
  v3,
  v4,
  w0,
  w1,
  w2,
  w3,
  w4,
  x0,
  x1,
  x2,
  x3,
  x4,
  y0,
  y1,
  y2,
  y3,
  y4,
  z0,
  z1,
  z2,
  z3,
  z4;
output
  y10,
  a6,
  a7,
  a8,
  a9,
  b6,
  b7,
  b8,
  b9,
  c6,
  c7,
  c8,
  c9,
  d6,
  d7,
  d8,
  d9,
  e6,
  e7,
  e8,
  e9,
  f6,
  f7,
  f8,
  f9,
  g6,
  g7,
  g8,
  g9,
  h6,
  h7,
  h8,
  h9,
  i6,
  i7,
  i8,
  i9,
  j6,
  j7,
  j8,
  j9,
  k6,
  k7,
  k8,
  k9,
  l6,
  l7,
  l8,
  l9,
  m6,
  m7,
  m8,
  m9,
  n6,
  n7,
  n8,
  n9,
  o6,
  o7,
  o8,
  o9,
  p6,
  p7,
  p8,
  p9,
  q6,
  q7,
  q8,
  q9,
  a10,
  r6,
  r7,
  r8,
  r9,
  s5,
  s6,
  s7,
  s8,
  s9,
  t5,
  t6,
  t7,
  t8,
  t9,
  u5,
  u6,
  u7,
  u8,
  u9,
  v5,
  v6,
  v7,
  v8,
  v9,
  w5,
  w6,
  w7,
  w8,
  w9,
  x5,
  x6,
  x7,
  x8,
  x9,
  y5,
  y6,
  y7,
  y8,
  y9,
  z5,
  z6,
  z7,
  z8,
  z9,
  b10,
  c10,
  d10,
  e10,
  f10,
  g10,
  h10,
  i10,
  j10,
  k10,
  l10,
  m10,
  n10,
  o10,
  p10,
  q10,
  r10,
  s10,
  t10,
  u10,
  v10,
  w10,
  x10;
wire
  y17,
  y18,
  y19,
  y25,
  y26,
  y30,
  y31,
  y32,
  y33,
  y34,
  y35,
  y37,
  y40,
  y41,
  y42,
  y43,
  y45,
  y47,
  y48,
  y50,
  y52,
  y53,
  y54,
  y55,
  y56,
  z16,
  z19,
  z22,
  z23,
  z24,
  z26,
  z28,
  z29,
  \[0] ,
  z30,
  z31,
  z32,
  z33,
  z34,
  z35,
  z36,
  z38,
  \[1] ,
  z40,
  z41,
  z42,
  z44,
  z48,
  z49,
  \[2] ,
  z50,
  z51,
  z54,
  z55,
  z56,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  a21,
  a22,
  a24,
  a25,
  a26,
  a28,
  a30,
  a32,
  a33,
  a34,
  a35,
  a36,
  a37,
  a40,
  a42,
  a43,
  a45,
  a48,
  a50,
  a51,
  a53,
  a55,
  a56,
  a57,
  b16,
  b17,
  b18,
  b20,
  b21,
  b22,
  b24,
  b25,
  b30,
  b31,
  b32,
  b33,
  b34,
  b35,
  b36,
  b37,
  b39,
  b46,
  b48,
  b49,
  b51,
  b55,
  b56,
  b57,
  c18,
  c20,
  c21,
  c22,
  c23,
  c24,
  c25,
  c28,
  c29,
  c30,
  c31,
  c33,
  c34,
  c35,
  c36,
  c39,
  c41,
  c47,
  c48,
  c50,
  c52,
  c53,
  c54,
  c55,
  c56,
  c57,
  d17,
  d21,
  d22,
  d23,
  d27,
  d28,
  d29,
  d30,
  d31,
  d32,
  d34,
  d35,
  d36,
  d38,
  d39,
  d46,
  d47,
  d51,
  d55,
  d56,
  d57,
  e17,
  e18,
  e19,
  e20,
  e21,
  e23,
  e29,
  e32,
  e33,
  e34,
  e35,
  e36,
  e37,
  e38,
  e39,
  e40,
  e41,
  e42,
  e43,
  e44,
  e45,
  e46,
  e52,
  e55,
  e56,
  e57,
  f16,
  f17,
  f20,
  f21,
  f22,
  f26,
  f27,
  f28,
  f29,
  f30,
  f31,
  f32,
  f33,
  f34,
  f35,
  f36,
  f37,
  f38,
  f40,
  f48,
  f50,
  f51,
  f52,
  f53,
  f54,
  f55,
  f56,
  f57,
  g16,
  g19,
  g20,
  g23,
  g24,
  g25,
  g28,
  g29,
  g31,
  g32,
  g33,
  g34,
  g35,
  g36,
  g37,
  g38,
  g39,
  g40,
  g41,
  g42,
  g43,
  g44,
  g45,
  g46,
  g47,
  g48,
  g49,
  g51,
  g53,
  g54,
  g55,
  g56,
  h20,
  h22,
  h26,
  h27,
  h29,
  h31,
  h32,
  h33,
  h34,
  h35,
  h37,
  h38,
  h39,
  h40,
  h42,
  h43,
  h46,
  h53,
  h54,
  h55,
  h56,
  i17,
  i19,
  i20,
  i22,
  i23,
  i24,
  i25,
  i28,
  i33,
  i34,
  i35,
  i36,
  i38,
  i39,
  i40,
  i44,
  i45,
  i47,
  i48,
  i49,
  i51,
  i52,
  i53,
  i55,
  i56,
  j16,
  j17,
  j18,
  j22,
  j24,
  j25,
  j26,
  j27,
  j28,
  j34,
  j35,
  j37,
  j38,
  j39,
  j40,
  j42,
  j43,
  j44,
  j46,
  j47,
  j48,
  j49,
  j50,
  j51,
  j52,
  j54,
  j55,
  j56,
  k19,
  k20,
  k22,
  k26,
  k30,
  k33,
  k34,
  k35,
  k37,
  k38,
  k39,
  k40,
  k42,
  k43,
  k45,
  k46,
  k51,
  k52,
  k53,
  k54,
  k55,
  k56,
  l16,
  l17,
  l18,
  l22,
  l24,
  l25,
  l31,
  l32,
  l33,
  l34,
  l35,
  l37,
  l38,
  l40,
  l43,
  l44,
  l47,
  l48,
  l50,
  l51,
  l52,
  l54,
  l55,
  l56,
  m16,
  m17,
  m18,
  m19,
  m21,
  m22,
  m24,
  m25,
  m26,
  m27,
  m33,
  m34,
  m35,
  m38,
  m39,
  m40,
  m41,
  m42,
  m43,
  m49,
  m51,
  m52,
  m53,
  m54,
  m55,
  m56,
  n20,
  n21,
  n22,
  n25,
  n27,
  n29,
  n31,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n42,
  n43,
  n44,
  n45,
  n47,
  n49,
  n50,
  n53,
  n54,
  n55,
  n56,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  o16,
  o17,
  o19,
  o21,
  o23,
  o24,
  \[17] ,
  o25,
  o26,
  o27,
  o28,
  o31,
  o33,
  o34,
  \[18] ,
  o35,
  o36,
  o37,
  o39,
  o41,
  o42,
  o45,
  o47,
  o48,
  o49,
  o53,
  o54,
  o55,
  o56,
  \[21] ,
  \[22] ,
  \[23] ,
  \[24] ,
  \[26] ,
  p18,
  p21,
  p22,
  p24,
  \[27] ,
  p25,
  p28,
  p30,
  p31,
  p32,
  p33,
  p34,
  \[28] ,
  p35,
  p36,
  p37,
  p38,
  p39,
  p40,
  p41,
  p42,
  \[100] ,
  p43,
  \[29] ,
  p45,
  p46,
  p47,
  p49,
  p50,
  p51,
  \[101] ,
  p53,
  p54,
  p55,
  p56,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[30] ,
  \[108] ,
  \[31] ,
  \[109] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  q16,
  q18,
  q19,
  q20,
  q21,
  q22,
  q23,
  q24,
  \[37] ,
  q27,
  q28,
  q29,
  q30,
  q32,
  q33,
  q34,
  \[38] ,
  q35,
  q36,
  q37,
  q38,
  q39,
  q40,
  q42,
  \[110] ,
  q43,
  \[39] ,
  q48,
  q51,
  \[111] ,
  q53,
  q54,
  q55,
  q56,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[40] ,
  \[118] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  r16,
  r17,
  r18,
  r20,
  r21,
  r22,
  r23,
  r24,
  \[47] ,
  r25,
  r26,
  r27,
  r28,
  r29,
  r30,
  r31,
  r32,
  r33,
  r34,
  \[48] ,
  r35,
  r36,
  r37,
  r38,
  r40,
  r41,
  r43,
  r44,
  \[49] ,
  r45,
  r46,
  r47,
  r49,
  r50,
  \[121] ,
  r53,
  r54,
  r55,
  r56,
  \[122] ,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \[50] ,
  \[128] ,
  \[51] ,
  \[129] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  s16,
  s18,
  s22,
  s24,
  \[57] ,
  s25,
  s26,
  s28,
  s29,
  s30,
  s31,
  s32,
  s33,
  s34,
  \[58] ,
  s35,
  s36,
  s39,
  s40,
  s41,
  s42,
  \[130] ,
  s43,
  s44,
  \[59] ,
  s45,
  s46,
  s48,
  \[131] ,
  s53,
  s54,
  s55,
  s56,
  \[132] ,
  \[133] ,
  \[134] ,
  \[135] ,
  \[136] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  t17,
  t20,
  t21,
  t22,
  t23,
  \[67] ,
  t25,
  t26,
  t27,
  t28,
  t29,
  t30,
  t31,
  t32,
  t33,
  t34,
  \[68] ,
  t35,
  t37,
  t38,
  t39,
  t40,
  t41,
  t42,
  t44,
  \[69] ,
  t46,
  t47,
  t49,
  t50,
  t52,
  t54,
  t55,
  t56,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  u16,
  u18,
  u19,
  u22,
  u23,
  u24,
  \[77] ,
  u25,
  u26,
  u27,
  u28,
  u30,
  u31,
  u32,
  u33,
  u34,
  \[78] ,
  u35,
  u38,
  u39,
  u41,
  u42,
  u43,
  \[79] ,
  u45,
  u46,
  u49,
  u51,
  u52,
  u53,
  u54,
  u55,
  u56,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  v17,
  v19,
  v20,
  v21,
  v22,
  v23,
  v24,
  \[87] ,
  v26,
  v28,
  v29,
  v30,
  v31,
  v32,
  v33,
  v34,
  \[88] ,
  v35,
  v38,
  v39,
  v40,
  v41,
  v42,
  v43,
  v44,
  \[89] ,
  v45,
  v46,
  v48,
  v49,
  v50,
  v51,
  v52,
  v53,
  v54,
  v55,
  v56,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  w16,
  w18,
  w23,
  w24,
  \[97] ,
  w25,
  w29,
  w30,
  w32,
  w33,
  w34,
  \[98] ,
  w35,
  w39,
  w40,
  w43,
  w44,
  \[99] ,
  w46,
  w47,
  w51,
  w52,
  w53,
  w54,
  w55,
  w56,
  x18,
  x21,
  x23,
  x24,
  x25,
  x27,
  x29,
  x30,
  x31,
  x33,
  x34,
  x35,
  x40,
  x41,
  x42,
  x46,
  x49,
  x53,
  x54,
  x55,
  x56;
assign
  y10 = \[136] ,
  y17 = (~b17 & d1) | (b17 & ~d1),
  y18 = (~u18 & r18) | (u18 & ~r18),
  y19 = k1 | ~o1,
  y25 = (~x25 & k20) | ((~x25 & ~e3) | (~k20 & ~e3)),
  y26 = (~f2 & ~o26) | (f2 & o26),
  y30 = (~w2 & ~z30) | (w2 & z30),
  y31 = (~a3 & b32) | (a3 & ~b32),
  y32 = (~r32 & ~q32) | ((~r32 & ~e19) | (~q32 & e19)),
  y33 = ~s33 | (~r33 | (~q33 | ~p33)),
  y34 = ~y2 | ~n,
  y35 = ~u1 | ~r,
  y37 = ~o3 | (~n3 | (~m3 | ~l3)),
  y40 = j50 | e52,
  y41 = (~w3 & a42) | (w3 & ~a42),
  y42 = (~z3 & a43) | (z3 & ~a43),
  y43 = ~g41 & ~u43,
  y45 = n45 & (m4 & n4),
  y47 = ~b48 | ~a48,
  y48 = ~t50 | z,
  y50 = g49 | ~d47,
  y52 = (~t52 & (~m5 & h40)) | ((~t52 & (~m5 & ~o49)) | ((~t52 & (~m5 & m53)) | ((~t52 & (~n5 & h40)) | ((~t52 & (~n5 & ~o49)) | (~t52 & (~n5 & m53)))))),
  y53 = (~r5 & ~q5) | ((~r5 & ~p5) | (~q5 & ~p5)),
  y54 = ~k55 & (~m55 & ~l55),
  y55 = ~r3 | ~k0,
  y56 = ~z3 | ~o0,
  z16 = (~q16 & ~y0) | (q16 & y0),
  z19 = j1 | o1,
  z22 = (~b & (v22 & q1)) | ((~b & (v22 & r1)) | (~b & (v22 & p1))),
  z23 = (~q23 & ~o23) | ((~q23 & ~v19) | (~o23 & v19)),
  z24 = (~l24 & ~j24) | ((~l24 & ~v19) | (~j24 & v19)),
  z26 = (~y26 & ~q19) | ((~y26 & ~t1) | (q19 & ~t1)),
  z28 = (~q2 & ~r20) | (q2 & r20),
  z29 = (~g29 & ~e19) | (~e29 & e19),
  \[0]  = ~s35,
  z30 = r20 & ~x30,
  z31 = ~y31 | ~t20,
  z32 = (~d3 & c33) | (d3 & ~c33),
  z33 = ~l34 & (~n34 & ~m34),
  z34 = ~c3 | ~m,
  z35 = ~x1 | ~q,
  z36 = ~q5 | m53,
  z38 = (e38 & ~p3) | h0,
  \[1]  = ~d35,
  z40 = c52 & ~v40,
  z41 = (~l51 & ~n3) | ((l51 & ~y41) | (~y41 & ~n3)),
  z42 = (~l51 & ~q3) | ((l51 & ~y42) | (~y42 & ~q3)),
  z44 = (~h4 & ~n44) | (h4 & n44),
  z48 = (~y48 & o49) | (~y48 & ~d5),
  z49 = ~f5 & ~g5,
  \[2]  = ~o34,
  z50 = ~c47 & ~g0,
  z51 = (~u51 & ~k5) | (u51 & k5),
  z54 = ~r4 | ~u0,
  z55 = ~y55 | (~x55 | ~w55),
  z56 = ~c4 | ~n0,
  \[3]  = ~z33,
  \[4]  = ~k33,
  \[5]  = ~r56,
  \[6]  = ~c56,
  \[7]  = ~n55,
  \[8]  = ~y54,
  \[9]  = ~j54,
  a6 = \[8] ,
  a7 = \[34] ,
  a8 = \[60] ,
  a9 = \[86] ,
  b6 = \[9] ,
  b7 = \[35] ,
  b8 = \[61] ,
  b9 = \[87] ,
  c6 = \[10] ,
  c7 = \[36] ,
  c8 = \[62] ,
  c9 = \[88] ,
  d6 = \[11] ,
  d7 = \[37] ,
  d8 = \[63] ,
  d9 = \[89] ,
  e6 = \[12] ,
  e7 = \[38] ,
  e8 = \[64] ,
  e9 = \[90] ,
  f6 = \[13] ,
  f7 = \[39] ,
  f8 = \[65] ,
  f9 = \[91] ,
  g6 = \[14] ,
  g7 = \[40] ,
  g8 = \[66] ,
  g9 = \[92] ,
  h6 = \[15] ,
  h7 = \[41] ,
  h8 = \[67] ,
  h9 = \[93] ,
  i6 = \[16] ,
  i7 = \[42] ,
  i8 = \[68] ,
  i9 = \[94] ,
  j6 = \[17] ,
  j7 = \[43] ,
  j8 = \[69] ,
  j9 = \[95] ,
  k6 = \[18] ,
  k7 = \[44] ,
  k8 = \[70] ,
  k9 = \[96] ,
  l6 = a,
  l7 = \[45] ,
  l8 = \[71] ,
  l9 = \[97] ,
  m6 = e1,
  m7 = \[46] ,
  m8 = \[72] ,
  m9 = \[98] ,
  n6 = \[21] ,
  n7 = \[47] ,
  n8 = \[73] ,
  n9 = \[99] ,
  o6 = \[22] ,
  o7 = \[48] ,
  o8 = \[74] ,
  o9 = \[100] ,
  p6 = \[23] ,
  p7 = \[49] ,
  p8 = \[75] ,
  p9 = \[101] ,
  q6 = \[24] ,
  q7 = \[50] ,
  q8 = \[76] ,
  q9 = \[102] ,
  a10 = \[112] ,
  r6 = j1,
  r7 = \[51] ,
  r8 = \[77] ,
  r9 = \[103] ,
  a21 = p22 | (j18 | ~s18),
  a22 = f21 | p22,
  a24 = (~u1 & c24) | (u1 & ~c24),
  a25 = (~x1 & c25) | (x1 & ~c25),
  a26 = ~d21 & ~w25,
  a28 = m27 & k2,
  s5 = \[0] ,
  s6 = \[26] ,
  s7 = \[52] ,
  s8 = \[78] ,
  s9 = \[104] ,
  a30 = ~r20 | ~z29,
  a32 = e19 | t20,
  a33 = ~z32 | ~t20,
  a34 = ~v0 | ~w,
  a35 = ~z34 | (~y34 | ~x34),
  a36 = ~a2 | ~p,
  a37 = ~p5 | m53,
  t5 = \[1] ,
  t6 = \[27] ,
  t7 = \[53] ,
  t8 = \[79] ,
  t9 = \[105] ,
  a40 = p3 | (o3 | ~n3),
  a42 = ~g41 & ~x41,
  a43 = ~g41 & ~x42,
  a45 = (~v50 & ~z44) | ((v50 & ~v3) | (~z44 & ~v3)),
  a48 = ~c48 & ~g47,
  u5 = \[2] ,
  u6 = \[28] ,
  u7 = \[54] ,
  u8 = \[80] ,
  u9 = \[106] ,
  a50 = (~z49 & (~x49 & ~z)) | ((~z49 & (~f5 & ~z)) | (x49 & (~f5 & ~z))),
  a51 = i5 | ~o5,
  a53 = ~y52 | ~i53,
  a55 = ~w4 | ~t0,
  a56 = ~r55 | (~q55 | (~p55 | ~o55)),
  a57 = ~i3 | ~m0,
  v5 = \[3] ,
  v6 = \[29] ,
  v7 = \[55] ,
  v8 = \[81] ,
  v9 = \[107] ,
  w5 = \[4] ,
  w6 = \[30] ,
  w7 = \[56] ,
  w8 = \[82] ,
  w9 = \[108] ,
  x5 = \[5] ,
  x6 = \[31] ,
  x7 = \[57] ,
  x8 = \[83] ,
  x9 = \[109] ,
  y5 = \[6] ,
  y6 = \[32] ,
  y7 = \[58] ,
  y8 = \[84] ,
  y9 = \[110] ,
  z5 = \[7] ,
  z6 = \[33] ,
  z7 = \[59] ,
  z8 = \[85] ,
  z9 = \[111] ,
  b10 = \[113] ,
  b16 = ~j1 | o28,
  b17 = ~e17 | ~d17,
  b18 = b | ~o19,
  b20 = (~o28 & j1) | ((o28 & ~j1) | b),
  b21 = ~v0 | (h22 | ~r1),
  b22 = ~p21 | h22,
  b24 = (~a24 & k20) | ((~a24 & ~y2) | (~k20 & ~y2)),
  b25 = (~a25 & k20) | ((~a25 & ~b3) | (~k20 & ~b3)),
  b30 = (~t2 & ~a30) | (t2 & a30),
  b31 = (~r30 & ~p30) | ((~r30 & ~e19) | (~p30 & e19)),
  b32 = r20 & ~x31,
  b33 = e19 | t20,
  b34 = ~a1 | ~v,
  b35 = ~s34 | (~r34 | (~q34 | ~p34)),
  b36 = ~t2 | ~o,
  b37 = (~p36 & ~i3) | h0,
  b39 = q3 | ~z38,
  b46 = n45 & m4,
  b48 = y50 & y4,
  b49 = (~y48 & ~e5) | (~y48 & r49),
  b51 = g5 | o5,
  b55 = ~d4 | ~s0,
  b56 = ~v55 | (~u55 | (~t55 | ~s55)),
  b57 = ~p3 | ~l0,
  c10 = \[114] ,
  c18 = (~b18 & r18) | (~b18 & ~h1),
  c20 = o19 & ~h20,
  c21 = ~q20 & ~p22,
  c22 = ~b22 | ~a22,
  c23 = (~u22 & (t22 & ~q1)) | ((~u22 & (~r1 & ~q1)) | ((u22 & (~t22 & ~r1)) | ((u22 & (t22 & ~p1)) | ((u22 & (~r1 & ~p1)) | ((~t22 & (~r1 & ~q1)) | ((t22 & (~q1 & ~p1)) | (~r1 & (~q1 & ~p1)))))))),
  c24 = ~d21 & ~z23,
  c25 = ~d21 & ~z24,
  c28 = (~k2 & m27) | (k2 & ~m27),
  c29 = (~q2 & ~r2) | h29,
  c30 = ~b30 | ~t20,
  c31 = (~x2 & ~d31) | (x2 & d31),
  c33 = r20 & ~y32,
  c34 = ~b2 | ~u,
  c35 = ~w34 | (~v34 | (~u34 | ~t34)),
  c36 = ~a3 | ~n,
  c39 = (g38 & p3) | h0,
  c41 = (~u3 & ~g41) | (u3 & g41),
  c47 = \[121]  | c5,
  c48 = ~x4 | (~w4 | ~v4),
  c50 = (f50 & (~x49 & ~f5)) | ((f50 & (x49 & ~g5)) | (f50 & (~g5 & ~f5))),
  c52 = d0 | ~p51,
  c53 = ~u52 | ~w52,
  c54 = (~z & (y53 & q5)) | ((~z & (y53 & r5)) | (~z & (y53 & p5))),
  c55 = ~h4 | ~r0,
  c56 = ~o56 & (~q56 & ~p56),
  c57 = ~t3 | ~k0,
  d10 = \[115] ,
  d17 = ~f17 & ~j16,
  d21 = ~h & ~c21,
  d22 = ~q21 & (~e21 & ~c22),
  d23 = (~u22 & (t22 & ~r1)) | ((~u22 & (~r1 & ~p1)) | ((u22 & (~t22 & ~p1)) | ((u22 & (t22 & ~q1)) | ((u22 & (~q1 & ~p1)) | ((~t22 & (~r1 & ~p1)) | ((t22 & (~r1 & ~q1)) | (~r1 & (~q1 & ~p1)))))))),
  d27 = (~g2 & ~j26) | (g2 & j26),
  d28 = (~c28 & ~q19) | ((~c28 & ~x1) | (q19 & ~x1)),
  d29 = ~j & ~r22,
  d30 = e19 | t20,
  d31 = r20 & ~b31,
  d32 = (~o31 & ~l31) | ((~o31 & ~e19) | (~l31 & e19)),
  d34 = ~f2 | ~t,
  d35 = ~p35 & (~r35 & ~q35),
  d36 = ~e3 | ~m,
  d38 = ~l3 & b37,
  d39 = ~c39 | ~q3,
  d46 = (~m4 & n45) | (m4 & ~n45),
  d47 = (~c47 & ~r5) | (~c47 & m53),
  d51 = (~p46 & h5) | ((p46 & ~h5) | z),
  d55 = ~m4 | ~q0,
  d56 = ~t4 | ~u0,
  d57 = ~c57 | (~b57 | ~a57),
  e10 = \[116] ,
  e17 = u19 & c1,
  e18 = (~b18 & ~i1) | (~b18 & u18),
  e19 = ~g20 & ~g,
  e20 = w0 & ~v0,
  e21 = ~b & (~n1 & (m1 & ~l1)),
  e23 = (~u22 & (t22 & ~p1)) | ((~u22 & (~q1 & ~p1)) | ((u22 & (~t22 & ~q1)) | ((u22 & (t22 & ~r1)) | ((u22 & (~r1 & ~q1)) | ((~t22 & (~q1 & ~p1)) | ((t22 & (~r1 & ~p1)) | (~r1 & (~q1 & ~p1)))))))),
  e29 = (~d29 & ~c29) | (~d29 & s2),
  e32 = (~b3 & h32) | (b3 & ~h32),
  e33 = (~t32 & ~s32) | ((~t32 & ~e19) | (~s32 & e19)),
  e34 = ~k2 | ~s,
  e35 = ~x0 | ~w,
  e36 = ~d36 | (~c36 | ~b36),
  e37 = (~r36 & i3) | h0,
  e38 = j3 & b37,
  e39 = ~p3 | ~q3,
  e40 = t3 | (s3 | (r3 | q3)),
  e41 = (~l51 & ~l3) | ((l51 & ~c41) | (~c41 & ~l3)),
  e42 = ~x3 & p41,
  e43 = ~a4 & k42,
  e44 = j0 | ~q5,
  e45 = (~i4 & ~i44) | (i4 & i44),
  e46 = (~v50 & ~d46) | ((v50 & ~z3) | (~d46 & ~z3)),
  e52 = ~l52 & ~z,
  e55 = ~m5 | ~p0,
  e56 = ~y4 | ~t0,
  e57 = ~v56 | (~u56 | (~t56 | ~s56)),
  f10 = \[117] ,
  f16 = \[21]  | g1,
  f17 = ~b1 | (~a1 | ~z0),
  f20 = g19 & v0,
  f21 = (v17 & (r1 & ~c)) | ((v17 & (~d1 & ~c)) | (~r1 & (~d1 & ~c))),
  f22 = ~i22 | (h20 | ~k22),
  f26 = l | ~q1,
  f27 = ~o26 & (f2 & h2),
  f28 = (~l2 & a28) | (l2 & ~a28),
  f29 = (q2 & r2) | h29,
  f30 = z2 | (y2 | (x2 | w2)),
  f31 = (~u30 & ~t30) | ((~u30 & ~e19) | (~t30 & e19)),
  f32 = ~e32 | ~t20,
  f33 = (~e3 & i33) | (e3 & ~i33),
  f34 = ~m1 | ~r,
  f35 = ~c1 | ~v,
  f36 = ~w35 | (~v35 | (~u35 | ~t35)),
  f37 = (~j50 & ~f3) | (j50 & f3),
  f38 = e37 & l3,
  f40 = ~r3 & ~b39,
  f48 = y50 & (v4 & ~g47),
  f50 = t50 & ~j51,
  f51 = s4 & ~r4,
  f52 = (~c47 & ~g49) | ~k51,
  f53 = m52 | u53,
  f54 = (~x53 & (w53 & ~q5)) | ((~x53 & (~r5 & ~q5)) | ((x53 & (~w53 & ~r5)) | ((x53 & (w53 & ~p5)) | ((x53 & (~r5 & ~p5)) | ((~w53 & (~r5 & ~q5)) | ((w53 & (~q5 & ~p5)) | (~r5 & (~q5 & ~p5)))))))),
  f55 = ~r5 | ~o0,
  f56 = ~f4 | ~s0,
  f57 = ~z56 | (~y56 | (~x56 | ~w56)),
  g10 = \[118] ,
  g16 = (~f16 & ~r1) | (~f16 & h22),
  g19 = ~d1 & (~w0 & i19),
  g20 = ~s18 & ~p22,
  g23 = (~s1 & ~d21) | (s1 & d21),
  g24 = ~v1 & r23,
  g25 = ~y1 & m24,
  g28 = (~f28 & ~q19) | ((~f28 & ~y1) | (q19 & ~y1)),
  g29 = (~d29 & ~f29) | (~d29 & ~s2),
  g31 = (~y2 & ~h31) | (y2 & h31),
  g32 = e19 | t20,
  g33 = ~f33 | ~t20,
  g34 = ~r1 | ~q,
  g35 = ~d2 | ~u,
  g36 = ~a36 | (~z35 | (~y35 | ~x35)),
  g37 = (~g3 & ~h37) | (g3 & h37),
  g38 = k3 & e37,
  g39 = (~j50 & ~k38) | ((j50 & ~j38) | (~k38 & ~j38)),
  g40 = ~d39 & r3,
  g41 = ~f0 & ~k52,
  g42 = r41 & x3,
  g43 = m42 & a4,
  g44 = d4 & e4,
  g45 = ~n44 & (h4 & j4),
  g46 = (~n4 & b46) | (n4 & ~b46),
  g47 = ~u4 | (~t4 | (~s4 | ~r4)),
  g48 = y50 & (~c48 & ~g47),
  g49 = d5 | ~i49,
  g51 = l50 & r4,
  g53 = ~h40 | m53,
  g54 = (~x53 & (w53 & ~r5)) | ((~x53 & (~r5 & ~p5)) | ((x53 & (~w53 & ~p5)) | ((x53 & (w53 & ~q5)) | ((x53 & (~q5 & ~p5)) | ((~w53 & (~r5 & ~p5)) | ((w53 & (~r5 & ~q5)) | (~r5 & (~q5 & ~p5)))))))),
  g55 = ~p5 | ~n0,
  g56 = ~k4 | ~r0,
  h10 = y,
  h20 = ~b & (~n1 & (~m1 & l1)),
  h22 = ~m22 | ~l22,
  h26 = b2 & c2,
  h27 = ~o26 & f2,
  h29 = ~j & ~s22,
  h31 = r20 & ~f31,
  h32 = r20 & ~d32,
  h33 = e19 | t20,
  h34 = ~p1 | ~p,
  h35 = ~i2 | ~t,
  h37 = c52 & ~f37,
  h38 = ~m3 & (~l3 & b37),
  h39 = (~o3 & k39) | (o3 & ~k39),
  h40 = ~e40 & ~a40,
  h42 = ~y3 & (~x3 & p41),
  h43 = ~b4 & (~a4 & k42),
  h46 = (~v50 & ~g46) | ((v50 & ~a4) | (~g46 & ~a4)),
  h53 = ~g53 | ~f53,
  h54 = (~x53 & (w53 & ~p5)) | ((~x53 & (~q5 & ~p5)) | ((x53 & (~w53 & ~q5)) | ((x53 & (w53 & ~r5)) | ((x53 & (~r5 & ~q5)) | ((~w53 & (~q5 & ~p5)) | ((w53 & (~r5 & ~p5)) | (~r5 & (~q5 & ~p5)))))))),
  h55 = ~f3 | ~m0,
  h56 = ~o4 | ~q0,
  i10 = a5,
  i17 = u19 & (z0 & ~j16),
  i19 = ~c1 & (~b1 & (~a1 & m19)),
  i20 = ~v0 & g19,
  i22 = r18 | ~e21,
  i23 = (~g23 & k20) | ((~g23 & ~w2) | (~k20 & ~w2)),
  i24 = t23 & v1,
  i25 = o24 & y1,
  i28 = (~m2 & x27) | (m2 & ~x27),
  i33 = r20 & ~e33,
  i34 = ~q2 | ~o,
  i35 = ~m2 | ~s,
  i36 = (~f3 & ~c52) | (f3 & c52),
  i38 = e37 & (l3 & m3),
  i39 = ~h39 | ~e52,
  i40 = ~s3 & (~r3 & ~b39),
  i44 = (d4 & (e4 & f4)) | ~e44,
  i45 = ~n44 & h4,
  i47 = y50 & r4,
  i48 = y50 & (w4 & (v4 & ~g47)),
  i49 = r49 | (~v49 | ~u49),
  i51 = ~p49 & ~u53,
  i52 = u53 | (g49 | ~p49),
  i53 = ~v52 & (~l52 & ~h53),
  i55 = ~m3 | ~l0,
  i56 = ~v3 | ~p0,
  j10 = \[121] ,
  j16 = ~y0 | (~x0 | (~w0 | ~v0)),
  j17 = u19 & (~f17 & ~j16),
  j18 = h1 | ~l18,
  j22 = ~m21 | (r18 | p21),
  j24 = ~w1 & (~v1 & r23),
  j25 = ~z1 & (~y1 & m24),
  j26 = (b2 & (c2 & d2)) | ~f26,
  j27 = f27 & i2,
  j28 = (~i28 & ~q19) | ((~i28 & ~z1) | (q19 & ~z1)),
  j34 = ~x2 | ~n,
  j35 = ~t1 | ~r,
  j37 = (~j50 & ~q36) | ((j50 & ~n36) | (~q36 & ~n36)),
  j38 = ~n3 & (~m3 & (~l3 & b37)),
  j39 = j50 | e52,
  j40 = ~d39 & (r3 & s3),
  j42 = r41 & (x3 & y3),
  j43 = m42 & (a4 & b4),
  j44 = (~e4 & ~d4) | (e4 & d4),
  j46 = (~o4 & y45) | (o4 & ~y45),
  j47 = y50 & ~g47,
  j48 = (~j47 & ~v4) | (j47 & v4),
  j49 = ~d5 | ~z48,
  j50 = ~i51 & ~e0,
  j51 = ~z & (~n5 & (~m5 & l5)),
  j52 = ~r4 | (m53 | ~r5),
  j54 = ~v54 & (~x54 & ~w54),
  j55 = ~q3 | ~k0,
  j56 = ~y3 | ~o0,
  k10 = \[122] ,
  k19 = ~y0 & ~x0,
  k20 = (~h20 & p22) | (~h20 & ~f20),
  k22 = h22 | ~j22,
  k26 = (~c2 & ~b2) | (c2 & b2),
  k30 = ~z2 | (~y2 | (~x2 | ~w2)),
  k33 = ~w33 & (~y33 & ~x33),
  k34 = ~b3 | ~m,
  k35 = ~w1 | ~q,
  k37 = (~h3 & ~l37) | (h3 & l37),
  k38 = e37 & (l3 & (m3 & n3)),
  k39 = c52 & ~g39,
  k40 = ~e39 & (r3 & (s3 & t3)),
  k42 = (p41 & (~x3 & (~y3 & ~z3))) | i0,
  k43 = (~z50 & ~m42) | ((z50 & ~k42) | (~m42 & ~k42)),
  k45 = g45 & k4,
  k46 = (~v50 & ~j46) | ((v50 & ~b4) | (~j46 & ~b4)),
  k51 = ~r4 & l50,
  k52 = ~q51 & ~u53,
  k53 = ~n53 | (j51 | ~p53),
  k54 = ~l5 | ~u0,
  k55 = ~j55 | (~i55 | ~h55),
  k56 = ~b4 | ~n0,
  l10 = \[123] ,
  l16 = u19 & v0,
  l17 = u19 & (a1 & (z0 & ~j16)),
  l18 = u18 | (~y18 | ~x18),
  l22 = m1 & l1,
  l24 = t23 & (v1 & w1),
  l25 = o24 & (y1 & z1),
  l31 = (q30 & ~a3) | j,
  l32 = a3 | (z2 | ~y2),
  l33 = ~l1 | ~w,
  l34 = ~k34 | (~j34 | ~i34),
  l35 = ~z1 | ~p,
  l37 = c52 & ~j37,
  l38 = (~j50 & ~e37) | ((j50 & ~b37) | (~e37 & ~b37)),
  l40 = (~j50 & d39) | ((j50 & b39) | (d39 & b39)),
  l43 = (~a4 & n43) | (a4 & ~n43),
  l44 = (~f4 & ~g44) | (f4 & g44),
  l47 = y50 & (s4 & r4),
  l48 = (~f48 & ~w4) | (f48 & w4),
  l50 = ~z4 & (~s4 & n50),
  l51 = (~j51 & u53) | (~j51 & ~g51),
  l52 = ~z & (~n5 & (m5 & ~l5)),
  l54 = ~v4 | ~t0,
  l55 = ~c55 | (~b55 | (~a55 | ~z54)),
  l56 = ~h3 | ~m0,
  m10 = \[124] ,
  m16 = u19 & ~j16,
  m17 = (~m16 & ~z0) | (m16 & z0),
  m18 = ~h1 | ~c18,
  m19 = ~z0 & k19,
  m21 = c3 & (d3 & e3),
  m22 = ~b & ~n1,
  m24 = (r23 & (~v1 & (~w1 & ~x1))) | k,
  m25 = (~o24 & ~m24) | ((~o24 & ~v19) | (~m24 & v19)),
  m26 = (~d2 & ~h26) | (d2 & h26),
  m27 = (f27 & (i2 & j2)) | l,
  m33 = ~z0 | ~v,
  m34 = ~d34 | (~c34 | (~b34 | ~a34)),
  m35 = ~s2 | ~o,
  m38 = (~l3 & ~n38) | (l3 & n38),
  m39 = (~j50 & ~g38) | ((j50 & ~e38) | (~g38 & ~e38)),
  m40 = (~r3 & ~n40) | (r3 & n40),
  m41 = ~v3 & ~u3,
  m42 = (r41 & (x3 & (y3 & z3))) | i0,
  m43 = (~l51 & ~r3) | ((l51 & ~l43) | (~l43 & ~r3)),
  m49 = ~u49 | (~v49 | o49),
  m51 = ~j5 & k5,
  m52 = (s48 & (r5 & ~a0)) | ((s48 & (~z4 & ~a0)) | (~r5 & (~z4 & ~a0))),
  m53 = ~r53 | ~q53,
  m54 = c52 | ~s0,
  m55 = ~g55 | (~f55 | (~e55 | ~d55)),
  m56 = ~o3 | ~l0,
  n10 = \[125] ,
  n20 = (p22 & (r1 & ~v0)) | ((v20 & (r1 & ~v0)) | ((p22 & h22) | (h22 & v20))),
  n21 = ~b & (n1 & (m1 & l1)),
  n22 = n1 | ~q22,
  n25 = (~y1 & p25) | (y1 & ~p25),
  n27 = (~h2 & h27) | (h2 & ~h27),
  n29 = (~e29 & ~t2) | j,
  n31 = b3 | ~l31,
  n33 = r20 | ~u,
  n34 = ~h34 | (~g34 | (~f34 | ~e34)),
  n35 = ~z2 | ~n,
  n36 = (~f3 & ~g3) | s36,
  n37 = (~j50 & ~r36) | (j50 & ~p36),
  n38 = c52 & ~l38,
  n39 = (~p3 & q39) | (p3 & ~q39),
  n40 = c52 & ~l40,
  n42 = (~z50 & ~r41) | ((z50 & ~p41) | (~r41 & ~p41)),
  n43 = ~g41 & ~k43,
  n44 = ~t44 | ~g4,
  n45 = (g45 & (k4 & l4)) | j0,
  n47 = y50 & (t4 & (s4 & r4)),
  n49 = ~e5 | ~b49,
  n50 = ~y4 & (~x4 & (~w4 & r50)),
  n53 = o49 | ~l52,
  n54 = ~g4 | ~r0,
  n55 = ~z55 & (~b56 & ~a56),
  n56 = ~s3 | ~k0,
  \[10]  = ~s16 & ~r16,
  \[11]  = ~s16 & ~u16,
  \[12]  = ~s16 & ~w16,
  \[13]  = ~s16 & ~z16,
  \[14]  = ~s16 & ~m17,
  \[15]  = ~s16 & ~o17,
  o10 = \[126] ,
  \[16]  = ~s16 & ~r17,
  o16 = u19 & (w0 & v0),
  o17 = (~i17 & ~a1) | (i17 & a1),
  o19 = b | (~l1 | (m1 | ~n1)),
  o21 = (~n21 & ~m21) | ((~n21 & p21) | ((~n21 & r18) | (~n21 & h22))),
  o23 = ~t1 & ~s1,
  o24 = (t23 & (v1 & (w1 & x1))) | k,
  \[17]  = ~s16 & ~t17,
  o25 = (~n25 & k20) | ((~n25 & ~c3) | (~k20 & ~c3)),
  o26 = ~t26 | ~e2,
  o27 = (~n27 & ~q19) | ((~n27 & ~u1) | (q19 & ~u1)),
  o28 = ~n2 | (~e2 | ~t26),
  o31 = (s30 & a3) | j,
  o33 = ~e2 | ~t,
  o34 = ~a35 & (~c35 & ~b35),
  \[18]  = ~s16 & ~y17,
  o35 = ~d3 | ~m,
  o36 = ~h0 & ~a37,
  o37 = ~c52 | ~n37,
  o39 = ~n39 | ~e52,
  o41 = u3 & v3,
  o42 = (~x3 & q42) | (x3 & ~q42),
  o45 = (~j4 & i45) | (j4 & ~i45),
  o47 = (~y50 & ~r4) | (y50 & r4),
  o48 = (~i48 & ~x4) | (i48 & x4),
  o49 = b5 | ~a5,
  o53 = ~k40 | (o49 | h40),
  o54 = p46 | ~q0,
  o55 = ~s4 | ~u0,
  o56 = ~n56 | (~m56 | ~l56),
  \[21]  = i1 | ~p18,
  \[22]  = ~m18 | ~l18,
  \[23]  = ~q18 | ~p18,
  \[24]  = ~c20 | ~b20,
  p10 = g5,
  \[26]  = ~b & f22,
  p18 = ~x18 | (~y18 | r18),
  p21 = ~p32 & ~l32,
  p22 = ~b & n22,
  p24 = (~t23 & ~r23) | ((~t23 & ~v19) | (~r23 & v19)),
  \[27]  = ~b & v21,
  p25 = ~d21 & ~m25,
  p28 = ~f2 | ~h2,
  p30 = ~w2 & n29,
  p31 = ~o31 | ~b3,
  p32 = e3 | (d3 | (c3 | b3)),
  p33 = o28 | ~s,
  p34 = ~w0 | ~w,
  \[28]  = ~b & x21,
  p35 = ~o35 | (~n35 | ~m35),
  p36 = (~o36 & ~n36) | (~o36 & h3),
  p37 = (~i3 & ~o37) | (i3 & o37),
  p38 = (~j50 & ~f38) | ((j50 & ~d38) | (~f38 & ~d38)),
  p39 = j50 | e52,
  p40 = (~j50 & ~g40) | ((j50 & ~f40) | (~g40 & ~f40)),
  p41 = (~u3 & (~v3 & ~w3)) | i0,
  p42 = (~l51 & ~o3) | ((l51 & ~o42) | (~o42 & ~o3)),
  \[100]  = z | ~a45,
  p43 = (~z50 & ~g43) | ((z50 & ~e43) | (~g43 & ~e43)),
  \[29]  = ~p22,
  p45 = (~v50 & ~o45) | ((v50 & ~w3) | (~o45 & ~w3)),
  p46 = ~p4 | (~g4 | ~t44),
  p47 = ~t50 | (z | (~j52 | ~i52)),
  p49 = ~c5 & ~\[121] ,
  p50 = ~u4 & ~t4,
  p51 = (u53 & (r5 & ~r4)) | ((f52 & (r5 & ~r4)) | ((u53 & ~m51) | (f52 & ~m51))),
  \[101]  = z | ~e45,
  p53 = m53 | ~o53,
  p54 = ~n5 | ~p0,
  p55 = ~x4 | ~t0,
  p56 = ~g56 | (~f56 | (~e56 | ~d56)),
  \[102]  = z | ~p45,
  \[103]  = z | ~s45,
  \[104]  = z | ~v45,
  \[105]  = z | ~e46,
  \[106]  = z | ~h46,
  \[107]  = z | ~k46,
  \[30]  = ~c23 | ~z22,
  \[108]  = ~v46 & (~r46 & (~s46 & ~t46)),
  \[31]  = ~d23 & z22,
  \[109]  = z | ~x46,
  \[32]  = ~e23 & z22,
  \[33]  = ~b & ~i23,
  \[34]  = ~b & ~w23,
  \[35]  = ~b & ~b24,
  q10 = \[128] ,
  \[36]  = b | ~r24,
  q16 = u19 & (x0 & (w0 & v0)),
  q18 = ~i1 | ~e18,
  q19 = ~o19 | ~o28,
  q20 = (~q1 & (~p1 & ~i19)) | ((~q1 & (~p1 & ~r1)) | ((~q1 & (~k19 & ~i19)) | ((~q1 & (~k19 & ~r1)) | ((~p1 & (~m19 & ~i19)) | ((~p1 & (~m19 & ~r1)) | ((~m19 & (~k19 & ~i19)) | ((~m19 & (~k19 & ~r1)) | ~e20))))))),
  q21 = ~b & (n1 & (~m1 & ~l1)),
  q22 = ~m1 & ~l1,
  q23 = s1 & t1,
  q24 = (~v1 & s24) | (v1 & ~s24),
  \[37]  = b | ~w24,
  q27 = (~i2 & f27) | (i2 & ~f27),
  q28 = ~i2 | (~j2 | ~k2),
  q29 = (~g29 & t2) | j,
  q30 = u2 & n29,
  q32 = ~c3 & ~n31,
  q33 = ~n1 | ~r,
  q34 = ~b1 | ~v,
  \[38]  = b | ~b25,
  q35 = ~h35 | (~g35 | (~f35 | ~e35)),
  q36 = (f3 & g3) | s36,
  q37 = ~p37 | ~e52,
  q38 = (~m3 & ~r38) | (m3 & r38),
  q39 = c52 & ~m39,
  q40 = (~s3 & t40) | (s3 & ~t40),
  q42 = ~g41 & ~n42,
  \[110]  = ~p47 & ~o47,
  q43 = (~b4 & s43) | (b4 & ~s43),
  \[39]  = ~b & ~o25,
  q48 = (~g48 & ~y4) | (g48 & y4),
  q51 = (~r50 & (~p50 & ~n50)) | ((~r50 & (~p50 & ~r5)) | ((~r50 & (~n50 & ~p5)) | ((~r50 & (~r5 & ~p5)) | ((~p50 & (~n50 & ~q5)) | ((~p50 & (~r5 & ~q5)) | ((~n50 & (~p5 & ~q5)) | ((~r5 & (~p5 & ~q5)) | ~f51))))))),
  \[111]  = ~p47 & ~r47,
  q53 = m5 & l5,
  q54 = e52 | ~o0,
  q55 = ~e4 | ~s0,
  q56 = ~k56 | (~j56 | (~i56 | ~h56)),
  \[112]  = ~p47 & ~t47,
  \[113]  = ~p47 & ~w47,
  \[114]  = ~p47 & ~j48,
  \[115]  = ~p47 & ~l48,
  \[116]  = ~p47 & ~o48,
  \[117]  = ~p47 & ~q48,
  \[40]  = b | ~t25,
  \[118]  = ~p47 & ~v48,
  \[41]  = b | ~y25,
  \[42]  = b | ~b2,
  \[43]  = b | ~k26,
  \[44]  = b | ~m26,
  \[45]  = b | ~v26,
  r10 = \[129] ,
  \[46]  = b | ~z26,
  r16 = (~u19 & ~v0) | (u19 & v0),
  r17 = (~l17 & ~b1) | (l17 & b1),
  r18 = f1 | ~e1,
  r20 = f | ~n20,
  r21 = (~q21 & (~h20 & ~p21)) | (~q21 & (~h20 & h22)),
  r22 = ~p1 | h22,
  r23 = (~s1 & (~t1 & ~u1)) | k,
  r24 = (~q24 & k20) | ((~q24 & ~z2) | (~k20 & ~z2)),
  \[47]  = b | ~d27,
  r25 = (~i25 & ~g25) | ((~i25 & ~v19) | (~g25 & v19)),
  r26 = ~j26 | ~g2,
  r27 = (~q27 & ~q19) | ((~q27 & ~v1) | (q19 & ~v1)),
  r28 = ~l2 | (~m2 | ~o2),
  r29 = (~e19 & ~q2) | (e19 & q2),
  r30 = q29 & w2,
  r31 = (~w30 & ~v30) | ((~w30 & ~e19) | (~v30 & e19)),
  r32 = ~p31 & c3,
  r33 = t20 | ~q,
  r34 = ~c2 | ~u,
  \[48]  = b | ~o27,
  r35 = ~l35 | (~k35 | (~j35 | ~i35)),
  r36 = (~o36 & ~q36) | (~o36 & ~h3),
  r37 = j50 | e52,
  r38 = c52 & ~p38,
  r40 = ~q40 | ~e52,
  r41 = (u3 & (v3 & w3)) | i0,
  r43 = (~l51 & ~s3) | ((l51 & ~q43) | (~q43 & ~s3)),
  r44 = ~i44 | ~i4,
  \[49]  = b | ~r27,
  r45 = (~k4 & g45) | (k4 & ~g45),
  r46 = ~h4 | ~j4,
  r47 = (~i47 & ~s4) | (i47 & s4),
  r49 = ~t49 | ~g5,
  r50 = ~v4 & p50,
  \[121]  = e5 | ~m49,
  r53 = ~z & ~n5,
  r54 = ~q5 | ~n0,
  r55 = ~j4 | ~r0,
  r56 = ~d57 & (~f57 & ~e57),
  \[122]  = ~j49 | ~i49,
  \[123]  = ~n49 | ~m49,
  \[124]  = f50 & ~a50,
  \[125]  = ~z & ~c50,
  \[126]  = ~f50 | ~d51,
  \[50]  = b | ~u27,
  \[128]  = ~w51 & ~v51,
  \[51]  = b | ~d28,
  \[129]  = ~w51 & ~z51,
  \[52]  = b | ~g28,
  \[53]  = b | ~j28,
  \[54]  = ~t28 & (~p28 & (~q28 & ~r28)),
  \[55]  = b | ~v28,
  s10 = \[130] ,
  \[56]  = (~b16 & ~a) | ((b16 & p2) | (p2 & ~a)),
  s16 = ~o19 | (b | (~b21 | ~a21)),
  s18 = ~g1 & ~\[21] ,
  s22 = ~q1 | h22,
  s24 = ~d21 & ~p24,
  \[57]  = t20 & ~z28,
  s25 = (~z1 & u25) | (z1 & ~u25),
  s26 = ~p1 & ~l,
  s28 = x27 & m2,
  s29 = (~r2 & ~t29) | (r2 & t29),
  s30 = v2 & q29,
  s31 = (~z2 & v31) | (z2 & ~v31),
  s32 = ~d3 & (~c3 & ~n31),
  s33 = ~q1 | ~p,
  s34 = ~h2 | ~t,
  \[58]  = t20 & ~s29,
  s35 = ~e36 & (~g36 & ~f36),
  s36 = ~h0 & ~z36,
  s39 = (~j50 & ~c39) | ((j50 & ~z38) | (~c39 & ~z38)),
  s40 = j50 | e52,
  s41 = (~z50 & ~u3) | (z50 & u3),
  s42 = (~z50 & ~g42) | ((z50 & ~e42) | (~g42 & ~e42)),
  \[130]  = ~z & k53,
  s43 = ~g41 & ~p43,
  s44 = ~p5 & ~j0,
  \[59]  = t20 & ~w29,
  s45 = (~v50 & ~r45) | ((v50 & ~x3) | (~r45 & ~x3)),
  s46 = ~k4 | (~l4 | ~m4),
  s48 = ~z4 | y47,
  \[131]  = ~z & a53,
  s53 = n5 | ~v53,
  s54 = ~k40 | ~m0,
  s55 = ~n4 | ~q0,
  s56 = ~u4 | ~u0,
  \[132]  = ~z & c53,
  \[133]  = ~u53,
  \[134]  = ~f54 | ~c54,
  \[135]  = ~g54 & c54,
  \[136]  = ~h54 & c54,
  \[60]  = ~d30 | ~c30,
  \[61]  = (~f30 & t20) | ((~f30 & e19) | (~t20 & e19)),
  \[62]  = ~k30 & t20,
  \[63]  = t20 & ~y30,
  \[64]  = t20 & ~c31,
  \[65]  = t20 & ~g31,
  t10 = \[131] ,
  \[66]  = ~u31 | ~t31,
  t17 = (~j17 & ~c1) | (j17 & c1),
  t20 = ~e21 & ~b,
  t21 = (~n21 & (~m1 & p21)) | ((~n21 & (~m1 & ~r18)) | ((~n21 & (~m1 & h22)) | ((~n21 & (~n1 & p21)) | ((~n21 & (~n1 & ~r18)) | (~n21 & (~n1 & h22)))))),
  t22 = ~n21 & ~e,
  t23 = (s1 & (t1 & u1)) | k,
  \[67]  = ~a32 | ~z31,
  t25 = (~s25 & k20) | ((~s25 & ~d3) | (~k20 & ~d3)),
  t26 = ~s26 | ~r26,
  t27 = (~j2 & j27) | (j2 & ~j27),
  t28 = ~b & q19,
  t29 = r20 & ~r29,
  t30 = ~x2 & (~w2 & n29),
  t31 = ~s31 | ~t20,
  t32 = ~p31 & (c3 & d3),
  t33 = ~m21 | ~o,
  t34 = ~l2 | ~s,
  \[68]  = ~g32 | ~f32,
  t35 = ~y0 | ~w,
  t37 = o3 | (n3 | (m3 | l3)),
  t38 = (~j50 & ~i38) | ((j50 & ~h38) | (~i38 & ~h38)),
  t39 = (~q3 & w39) | (q3 & ~w39),
  t40 = c52 & ~p40,
  t41 = (~v3 & v41) | (v3 & ~v41),
  t42 = (~y3 & v42) | (y3 & ~v42),
  t44 = ~s44 | ~r44,
  \[69]  = t20 & ~v32,
  t46 = ~n4 | (~o4 | ~q4),
  t47 = (~l47 & ~t4) | (l47 & t4),
  t49 = ~b51 | ~a51,
  t50 = z | (~l5 | (m5 | ~n5)),
  t52 = ~z & (n5 & (m5 & l5)),
  t54 = ~l3 | ~l0,
  t55 = ~u3 | ~p0,
  t56 = ~z4 | ~t0,
  \[70]  = ~b33 | ~a33,
  \[71]  = ~h33 | ~g33,
  \[72]  = e52 & ~i36,
  \[73]  = e52 & ~g37,
  \[74]  = e52 & ~k37,
  \[75]  = ~r37 | ~q37,
  u10 = \[132] ,
  \[76]  = (~e52 & j50) | ((e52 & ~t37) | (~t37 & j50)),
  u16 = (~l16 & ~w0) | (l16 & w0),
  u18 = ~w18 | ~j1,
  u19 = j18 | ~g16,
  u22 = ~q21 & ~d,
  u23 = (~v19 & ~s1) | (v19 & s1),
  u24 = (~i24 & ~g24) | ((~i24 & ~v19) | (~g24 & v19)),
  \[77]  = ~y37 & e52,
  u25 = ~d21 & ~r25,
  u26 = (~e2 & t26) | (e2 & ~t26),
  u27 = (~t27 & ~q19) | ((~t27 & ~w1) | (q19 & ~w1)),
  u28 = (~o2 & s28) | (o2 & ~s28),
  u30 = q29 & (w2 & x2),
  u31 = e19 | t20,
  u32 = (p31 & n31) | ((p31 & ~e19) | (n31 & e19)),
  u33 = ~w2 | ~n,
  u34 = ~s1 | ~r,
  \[78]  = e52 & ~m38,
  u35 = ~d1 | ~v,
  u38 = (~n3 & ~v38) | (n3 & v38),
  u39 = ~t39 | ~e52,
  u41 = (~l51 & ~m3) | ((l51 & ~t41) | (~t41 & ~m3)),
  u42 = (~l51 & ~p3) | ((l51 & ~t42) | (~t42 & ~p3)),
  u43 = (~z50 & ~j43) | ((z50 & ~h43) | (~j43 & ~h43)),
  \[79]  = e52 & ~q38,
  u45 = (~l4 & k45) | (l4 & ~k45),
  u46 = y45 & o4,
  u49 = ~d5 & ~e5,
  u51 = j5 & ~m53,
  u52 = (~t52 & ~k40) | ((~t52 & h40) | ((~t52 & o49) | (~t52 & m53))),
  u53 = ~z & s53,
  u54 = ~h40 | ~k0,
  u55 = ~x3 | ~o0,
  u56 = ~i4 | ~s0,
  \[80]  = e52 & ~u38,
  \[81]  = ~j39 | ~i39,
  \[82]  = ~p39 | ~o39,
  \[83]  = ~v39 | ~u39,
  \[84]  = e52 & ~m40,
  \[85]  = ~s40 | ~r40,
  v10 = \[133] ,
  \[86]  = ~y40 | ~x40,
  v17 = ~d1 | b17,
  v19 = ~f16 & ~i,
  v20 = (~f16 & ~j18) | ~i20,
  v21 = ~t21 | ~d22,
  v22 = (~r1 & ~q1) | ((~r1 & ~p1) | (~q1 & ~p1)),
  v23 = (~t1 & x23) | (t1 & ~x23),
  v24 = (~w1 & x24) | (w1 & ~x24),
  \[87]  = ~z & ~e41,
  v26 = (~u26 & ~q19) | ((~u26 & ~s1) | (q19 & ~s1)),
  v28 = (~u28 & ~q19) | ((~u28 & ~a2) | (q19 & ~a2)),
  v29 = (~f29 & ~c29) | ((~f29 & ~e19) | (~c29 & e19)),
  v30 = ~y2 & (~x2 & (~w2 & n29)),
  v31 = r20 & ~r31,
  v32 = (~c3 & ~w32) | (c3 & w32),
  v33 = ~p21 | ~m,
  v34 = ~v1 | ~q,
  \[88]  = ~z & ~u41,
  v35 = ~g2 | ~u,
  v38 = c52 & ~t38,
  v39 = j50 | e52,
  v40 = (~j50 & ~j40) | ((j50 & ~i40) | (~j40 & ~i40)),
  v41 = ~g41 & ~s41,
  v42 = ~g41 & ~s42,
  v43 = (~c4 & y43) | (c4 & ~y43),
  v44 = (~g4 & t44) | (g4 & ~t44),
  \[89]  = ~z & ~z41,
  v45 = (~v50 & ~u45) | ((v50 & ~y3) | (~u45 & ~y3)),
  v46 = ~z & v50,
  v48 = (~y47 & z4) | (y47 & ~z4),
  v49 = (~r49 & o49) | (r49 & ~o49),
  v50 = ~t50 | ~p46,
  v51 = (~m53 & j5) | (m53 & ~j5),
  v52 = ~z & (n5 & (~m5 & ~l5)),
  v53 = ~m5 & ~l5,
  v54 = ~u54 | (~t54 | ~s54),
  v55 = ~a4 | ~n0,
  v56 = ~l4 | ~r0,
  \[90]  = z | ~p42,
  \[91]  = z | ~u42,
  \[92]  = z | ~z42,
  \[93]  = ~z & ~m43,
  \[94]  = z | ~r43,
  \[95]  = z | ~w43,
  w10 = \[134] ,
  \[96]  = z | ~d4,
  w16 = (~o16 & ~x0) | (o16 & x0),
  w18 = ~z19 | ~y19,
  w23 = (~v23 & k20) | ((~v23 & ~x2) | (~k20 & ~x2)),
  w24 = (~v24 & k20) | ((~v24 & ~a3) | (~k20 & ~a3)),
  \[97]  = z | ~j44,
  w25 = (~l25 & ~j25) | ((~l25 & ~v19) | (~j25 & v19)),
  w29 = (~s2 & ~x29) | (s2 & x29),
  w30 = q29 & (w2 & (x2 & y2)),
  w32 = r20 & ~u32,
  w33 = ~v33 | (~u33 | ~t33),
  w34 = ~y1 | ~p,
  \[98]  = z | ~l44,
  w35 = ~j2 | ~t,
  w39 = c52 & ~s39,
  w40 = (~t3 & z40) | (t3 & ~z40),
  w43 = (~l51 & ~t3) | ((l51 & ~v43) | (~v43 & ~t3)),
  w44 = (~v50 & ~v44) | ((v50 & ~u3) | (~v44 & ~u3)),
  \[99]  = z | ~w44,
  w46 = (~q4 & u46) | (q4 & ~u46),
  w47 = (~n47 & ~u4) | (n47 & u4),
  w51 = m51 | z,
  w52 = (~v52 & (~j51 & ~h40)) | (~v52 & (~j51 & m53)),
  w53 = ~t52 & ~c0,
  w54 = ~n54 | (~m54 | (~l54 | ~k54)),
  w55 = ~g3 | ~m0,
  w56 = ~q4 | ~q0,
  x10 = \[135] ,
  x18 = ~h1 & ~i1,
  x21 = ~o21 | ~r21,
  x23 = ~d21 & ~u23,
  x24 = ~d21 & ~u24,
  x25 = (~a2 & a26) | (a2 & ~a26),
  x27 = m27 & (k2 & l2),
  x29 = r20 & ~v29,
  x30 = (~q29 & ~n29) | ((~q29 & ~e19) | (~n29 & e19)),
  x31 = (~s30 & ~q30) | ((~s30 & ~e19) | (~q30 & e19)),
  x33 = ~o33 | (~n33 | (~m33 | ~l33)),
  x34 = ~r2 | ~o,
  x35 = ~o2 | ~s,
  x40 = ~w40 | ~e52,
  x41 = (~z50 & ~o41) | ((z50 & ~m41) | (~o41 & ~m41)),
  x42 = (~z50 & ~j42) | ((z50 & ~h42) | (~j42 & ~h42)),
  x46 = (~v50 & ~w46) | ((v50 & ~c4) | (~w46 & ~c4)),
  x49 = h5 | ~\[126] ,
  x53 = ~v52 & ~b0,
  x54 = ~r54 | (~q54 | (~p54 | ~o54)),
  x55 = ~n3 | ~l0,
  x56 = ~w3 | ~p0;
endmodule

