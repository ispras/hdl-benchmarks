//NOTE: no-implementation module stub

module lmi_dcache (
    input wire CLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire DISABLEC,
    input wire INVALIDATE,
    input wire MEMSEQUENTIAL,
    input wire MEMZEROFIRST,
    input wire MEMFULLWORD,
    input wire EXT_DCREQRAM_R,
    input wire DC_GNTRAM_R,
    input wire DATAIN,
    output wire DC_DATAOUT,
    output wire DC_DATAOE,
    output wire DC_LBCOE,
    input wire NEXTADDR,
    input wire NEXTRDOP,
    input wire NEXTWROP,
    input wire NEXTBE,
    input wire NEXTSX,
    input wire DWORD_E,
    output wire EXCP,
    output wire DS_VAL,
    output wire DC_VAL,
    output wire LACK,
    output wire X_HALT_R,
    output wire DC_MISS_P,
    output wire DC_MISS_R,
    output wire DC_BAREMISS_R,
    output wire DC_HALT_W_R,
    output wire DC_HALT_M_R,
    output wire DC_CSTWBUS,
    output wire DC_RPQUIETIFNBA,
    output wire DC_RPQUIETIFB,
    output wire DC_RPALGNIFNBNA,
    output wire DC_RPALGNIFB,
    input wire DC_TAGINDEX,
    input wire DCR_TAGRD,
    input wire DC_TAGWR,
    input wire DC_TAGWE,
    input wire DC_TAGWEN,
    input wire DC_TAGRE,
    input wire DC_TAGREN,
    input wire DC_TAGCS,
    input wire DC_TAGCSN,
    input wire DCC_TAGMASK,
    input wire DC_DATAINDEX,
    input wire DCR_DATARD,
    input wire DC_DATAWR,
    input wire DC_DATAWE,
    input wire DC_DATAWEN,
    input wire DC_DATARE,
    input wire DC_DATAREN,
    input wire DC_DATACS,
    input wire DC_DATACSN,
    input wire DC_USEPROCIN
);

endmodule
