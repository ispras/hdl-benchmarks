//NOTE: no-implementation module stub

module GtCLK_FJK3 (
    output Q,
    output QN,
    input CP,
    input CD,
    input SD,
    input J,
    input K
);

endmodule
