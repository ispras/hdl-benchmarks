// IWLS benchmark module "too_large" printed on Wed May 29 17:29:21 2002
module too_large(a, b, c, d, e, f, g, h, i, j, k, l, m, n, o, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0, g0, h0, i0, j0, k0, l0, m0, n0, o0, p0);
input
  g0,
  h0,
  i0,
  j0,
  k0,
  l0,
  a,
  b,
  c,
  d,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m0,
  m,
  n,
  o,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0,
  d0,
  e0,
  f0;
output
  n0,
  o0,
  p0;
wire
  g1,
  g2,
  h1,
  h2,
  i1,
  i2,
  j1,
  j2,
  k1,
  l1,
  m1,
  n1,
  o1,
  p1,
  \[0] ,
  q1,
  \[1] ,
  r1,
  \[2] ,
  s1,
  t1,
  u1,
  v1,
  w0,
  w1,
  x0,
  x1,
  y0,
  y1,
  z0,
  z1,
  a1,
  a2,
  b1,
  b2,
  c1,
  c2,
  d1,
  d2,
  e1,
  e2,
  f1,
  f2;
assign
  g1 = j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (w & (~q & (~o & ~m)))))))),
  g2 = ~i0 & (~g0 & (~f0 & (~e0 & (d0 & (~c0 & (~a0 & (~y & w))))))),
  h1 = j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (w & (~r & (~q & ~o)))))))),
  h2 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (w & (~q & (~n & ~m)))))))),
  i1 = j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (w & (~q & (~n & ~m)))))))),
  i2 = i0 & (~g0 & (~f0 & (~e0 & (d0 & (~c0 & (~y & (~\x  & w))))))),
  j1 = i0 & (h0 & (~d0 & (~c0 & (~b0 & (z & (~y & (~\x  & (~q & (~o & ~m))))))))),
  j2 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (w & (~r & (~q & ~n)))))))),
  k1 = j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (w & (~r & (~q & ~n)))))))),
  l1 = i0 & (h0 & (~d0 & (~c0 & (~b0 & (z & (~y & (~\x  & (~r & (~q & ~o))))))))),
  m1 = j0 & (~i0 & (h0 & (~g0 & (~f0 & (~e0 & (~d0 & (~c0 & z))))))),
  n0 = \[0] ,
  n1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (v & (~q & (~o & ~m))))))))),
  o0 = \[1] ,
  o1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (v & (~r & (~q & ~o))))))))),
  p0 = \[2] ,
  p1 = ~i0 & (h0 & (~g0 & (~f0 & (~e0 & (~d0 & (~c0 & (~a0 & (z & ~y)))))))),
  \[0]  = (~a0 & (~y & (~v & (~g0 & (~s & (d & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (~g0 & (~s & (d & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (~g0 & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (~s & (d & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (~s & (d & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~v & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~a0 & (~y & (~g0 & (~s & (d & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~a0 & (~y & (~s & (d & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~g0 & (~s & (d & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~g0 & (~s & (d & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~s & (d & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (~s & (d & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~g0 & (~s & (d & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~s & (d & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))))) | ((~f0 & (~b & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~o & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~o & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~o & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~o & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~o & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~g & (~f & (~e & ~c))))))))))))))))) | ((~f0 & (~b & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e))))))))))))))))) | ((~k & (~a0 & (~y & (~v & (~g0 & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (~a0 & (~y & (~v & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((~k & (~a0 & (~y & (~v & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~k & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~g & (~f & ~e))))))))))))))))) | ((~o & (~a0 & (~y & (~v & (~g0 & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((~o & (~a0 & (~y & (~v & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((~o & (~a0 & (~y & (~v & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~o & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~o & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))))) | ((~m & (~f0 & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~g & (~f & ~e)))))))))))))))) | ((~m & (~f0 & (~o & (~a0 & (~y & (~v & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~g & (~f & ~e)))))))))))))))) | ((~m & (~f0 & (~o & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~o & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~o & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~o & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~g & (~f & ~e)))))))))))))))) | ((~m & (~f0 & (~a0 & (~y & (~v & (k0 & (~j0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~g & (~f & ~e)))))))))))))))) | ((~m & (~f0 & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~f0 & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~o & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~b & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c)))))))))))))))) | ((~m & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~o & (~a0 & (~y & (~v & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~o & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~o & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~o & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~o & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~o & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~o & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~a0 & (~y & (~v & (~g0 & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~a0 & (~y & (~v & (k0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~m & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~c))))))))))))))) | ((~e0 & (~f0 & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~c)))))))))))))) | ((~e0 & (~f0 & (~o & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & ~c)))))))))))))) | ((~e0 & (~f0 & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~c)))))))))))))) | ((~e0 & (~f0 & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & ~c)))))))))))))) | ((~e0 & (~m & (~f0 & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & ~q))))))))))))) | ((~e0 & (~m & (~f0 & (~o & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~q & ~i))))))))))))) | ((~e0 & (~m & (~f0 & (~o & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~i))))))))))))) | ((~e0 & (~m & (~f0 & (~o & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~i))))))))))))) | ((~e0 & (~m & (~f0 & (~a0 & (~y & (~v & (~g0 & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~q & ~n))))))))))))) | ((~e0 & (~m & (~f0 & (~a0 & (~y & (~v & (k0 & (~j0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~i))))))))))))) | ((~e0 & (~m & (~f0 & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~i))))))))))))) | ((~e0 & (~m & (~f0 & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~i))))))))))))) | ((~e0 & (~f0 & (~o & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~i))))))))))))) | ((~e0 & (~f0 & (~o & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~i))))))))))))) | ((~e0 & (~f0 & (~a0 & (~y & (k0 & (~j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~i))))))))))))) | ((~e0 & (~f0 & (~y & (k0 & (~j0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~i))))))))))))) | ((~e0 & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & ~c))))))))))))) | ((~e0 & (~o & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & ~c))))))))))))) | ((~e0 & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & ~c))))))))))))) | ((~e0 & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & ~c))))))))))))) | ((~m & (f0 & (k & (~y & (v & (~s & (d & (i0 & (~c0 & (~b0 & (~\x  & (~q & (~n & h))))))))))))) | ((~m & (f0 & (k & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~t & (~q & (~n & (~l & h))))))))))))) | ((~m & (f0 & (k & (~y & (~s & (d & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & h))))))))))))) | ((~m & (f0 & (k & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~q & (~n & (~l & h))))))))))))) | ((~m & (f0 & (k & (v & (~s & (d & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~q & (~n & h))))))))))))) | ((~m & (f0 & (k & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~t & (~q & (~n & (~l & h))))))))))))) | ((~m & (f0 & (k & (~s & (d & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & h))))))))))))) | ((~m & (f0 & (k & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~q & (~n & (~l & h))))))))))))) | ((f0 & (k & (~y & (v & (~s & (d & (i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h))))))))))))) | ((f0 & (k & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & h))))))))))))) | ((f0 & (k & (~y & (~s & (d & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h))))))))))))) | ((f0 & (k & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & h))))))))))))) | ((f0 & (k & (v & (~s & (d & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h))))))))))))) | ((f0 & (k & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & h))))))))))))) | ((f0 & (k & (~s & (d & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h))))))))))))) | ((f0 & (k & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & h))))))))))))) | ((~a0 & (~y & (~v & (~s & (d & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & c))))))))))))) | ((~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & c))))))))))))) | ((~e0 & (~m & (~o & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~q & ~h)))))))))))) | ((~e0 & (~m & (~o & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (~o & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~h)))))))))))) | ((~e0 & (~m & (~o & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (~o & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~h)))))))))))) | ((~e0 & (~m & (~o & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (~o & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~h)))))))))))) | ((~e0 & (~m & (~o & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (~a0 & (~y & (~v & (~g0 & (k0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~h)))))))))))) | ((~e0 & (~m & (~a0 & (~y & (~v & (k0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~m & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~h)))))))))))) | ((~e0 & (~m & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~m & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~h)))))))))))) | ((~e0 & (~m & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~m & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & ~h)))))))))))) | ((~e0 & (~m & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~o & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~h)))))))))))) | ((~e0 & (~o & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & ~h)))))))))))) | ((~e0 & (~o & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~h)))))))))))) | ((~e0 & (~o & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & ~h)))))))))))) | ((~e0 & (~o & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~h)))))))))))) | ((~e0 & (~o & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & ~h)))))))))))) | ((~e0 & (~a0 & (~y & (~g0 & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~h)))))))))))) | ((~e0 & (~a0 & (~y & (k0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~h)))))))))))) | ((~e0 & (~y & (k0 & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & ~h)))))))))))) | ((~e0 & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & ~h)))))))))))) | ((~e0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & ~h)))))))))))) | ((~m & (f0 & (k & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~q & (n & h)))))))))))) | ((~m & (f0 & (k & (~o & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (n & h)))))))))))) | ((~m & (f0 & (k & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~q & (n & h)))))))))))) | ((~m & (f0 & (k & (~o & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (n & h)))))))))))) | ((~m & (f0 & (k & (~a0 & (~y & (~s & (d & (~c0 & (~b0 & (~\x  & (~q & (~n & h)))))))))))) | ((~m & (f0 & (k & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~t & (~q & (~n & (~l & h)))))))))))) | ((f0 & (k & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & h)))))))))))) | ((f0 & (k & (~o & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & h)))))))))))) | ((f0 & (k & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & h)))))))))))) | ((f0 & (k & (~o & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & h)))))))))))) | ((f0 & (k & (~a0 & (~y & (~s & (d & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h)))))))))))) | ((f0 & (k & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & h)))))))))))) | ((~k & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & c)))))))))))) | ((~o & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & c)))))))))))) | ((~m & (f0 & (k & (~o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~q & (n & h))))))))))) | ((~m & (f0 & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~q & (~j & h))))))))))) | ((~m & (f0 & (~o & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~j & h))))))))))) | ((~m & (f0 & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~q & (~j & h))))))))))) | ((~m & (f0 & (~o & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~j & h))))))))))) | ((~m & (f0 & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~j & h))))))))))) | ((~m & (f0 & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~j & h))))))))))) | ((~m & (f0 & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~j & h))))))))))) | ((~m & (f0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~j & h))))))))))) | ((f0 & (k & (~o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & h))))))))))) | ((f0 & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & h))))))))))) | ((f0 & (~o & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & h))))))))))) | ((f0 & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & h))))))))))) | ((f0 & (~o & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & h))))))))))) | ((f0 & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & h))))))))))) | ((f0 & (~y & (i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & h))))))))))) | ((f0 & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & h))))))))))) | ((f0 & (j0 & (~i0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & h))))))))))) | ((a & (~m & (~o & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & ~q)))))))))) | ((a & (~m & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((a & (~o & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))) | ((a & (~a0 & (~y & (~v & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((z & (h0 & (~m & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & ~q)))))))))) | ((z & (h0 & (~m & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & ~q)))))))))) | ((z & (h0 & (~o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))) | ((z & (h0 & (~o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))) | ((h0 & (~m & (o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((h0 & (~m & (o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((h0 & (o & (~y & (v & (i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((h0 & (o & (v & (j0 & (~i0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((u & (~m & (~o & (~y & (~v & (i0 & (d0 & (~c0 & (~b0 & (~\x  & ~q)))))))))) | ((u & (~m & (~o & (~v & (j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & ~q)))))))))) | ((u & (~m & (~y & (~v & (i0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((u & (~m & (~v & (j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((u & (~o & (~y & (~v & (i0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))) | ((u & (~o & (~v & (j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))) | ((u & (~y & (~v & (i0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((u & (~v & (j0 & (~i0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((~m & (f0 & (~o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~q & (~j & h)))))))))) | ((~m & (f0 & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~q & (~n & (~j & h)))))))))) | ((f0 & (~o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & h)))))))))) | ((f0 & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & h)))))))))) | ((z & (h0 & (~e0 & (~f0 & (~a0 & (~y & (v & (~g0 & (~i0 & ~c0))))))))) | ((z & (h0 & (~e0 & (~f0 & (~y & (v & (~g0 & (i0 & (~c0 & ~\x ))))))))) | ((h0 & (~e0 & (~f0 & (o & (~a0 & (~y & (v & (~g0 & (~i0 & ~c0))))))))) | ((h0 & (~e0 & (~f0 & (o & (~a0 & (~y & (~g0 & (~i0 & (~d0 & ~c0))))))))) | ((h0 & (~e0 & (~f0 & (o & (~y & (v & (~g0 & (i0 & (~c0 & ~\x ))))))))) | ((h0 & (~m & (o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~q & ~n))))))))) | ((h0 & (o & (~a0 & (~y & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n))))))))) | ((u & (~e0 & (~f0 & (~a0 & (~y & (~v & (~g0 & (~i0 & (d0 & ~c0))))))))) | ((u & (~e0 & (~f0 & (~y & (~v & (~g0 & (i0 & (d0 & (~c0 & ~\x ))))))))) | ((~e0 & (~f0 & (~a0 & (~y & (~g0 & (k0 & (~j0 & (~i0 & (~d0 & ~c0))))))))) | ((~e0 & (~f0 & (~y & (~g0 & (k0 & (~j0 & (i0 & (~d0 & (~c0 & ~\x ))))))))) | ((~e0 & (~f0 & (~y & (~g0 & (k0 & (i0 & (~d0 & (~c0 & (~\x  & ~h))))))))) | ((z & (h0 & (~e0 & (~f0 & (v & (~g0 & (j0 & (~i0 & ~c0)))))))) | ((h0 & (~e0 & (~f0 & (o & (v & (~g0 & (j0 & (~i0 & ~c0)))))))) | ((u & (~e0 & (~f0 & (~v & (~g0 & (j0 & (~i0 & (d0 & ~c0)))))))) | ((~e0 & (~f0 & (~g0 & (k0 & (j0 & (~i0 & (~d0 & (~c0 & ~h)))))))) | (j2 | (i2 | (h2 | (g2 | (f2 | (e2 | (d2 | (c2 | (b2 | (a2 | (z1 | (y1 | (x1 | (w1 | (v1 | (t1 | (s1 | (q1 | (p1 | (m1 | (l1 | (k1 | (j1 | (i1 | (h1 | (g1 | (f1 | (e1 | (d1 | (c1 | (b1 | (a1 | (z0 | (y0 | (x0 | w0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  q1 = i0 & (h0 & (~g0 & (~f0 & (~e0 & (~d0 & (~c0 & (z & (~y & ~\x )))))))),
  \[1]  = (~j0 & (~g0 & (~s & (d & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~j0 & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~j0 & (~s & (d & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~j0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~g0 & (~s & (d & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~s & (d & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))))))) | ((~k & (~j0 & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~k & (~j0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~i & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~k & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~k & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~i0 & (~c & (j0 & (~g0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e))))))))))))))))))) | ((~i0 & (~c & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & ~e))))))))))))))))))) | ((~i0 & (~c & (j0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))))) | ((~i0 & (~c & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~j0 & (~g0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~j0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~g0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~h & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))))) | ((i0 & (~c & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))))) | ((~c & (~j0 & (~g0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e))))))))))))))))))) | ((~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~g & (~f & ~e))))))))))))))))))) | ((~c & (~j0 & (~s & (d & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e))))))))))))))))))) | ((~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~t & (~r & (~q & (~n & (~l & (~j & (~i & (~g & (~f & ~e))))))))))))))))))) | ((~o & (~j0 & (~g0 & (~s & (d & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~j0 & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~l & (~j & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~j0 & (~s & (d & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~i & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~j0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~l & (~j & (~i & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~g0 & (~s & (d & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~l & (~j & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (~s & (d & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~i & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~o & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~t & (~r & (~q & (~l & (~j & (~i & (~h & (~g & (~f & (~e & ~a))))))))))))))))))) | ((~b & (~j0 & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~b & (~j0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~i & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~b & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~b & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~k & (~i0 & (~c & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~k & (~i0 & (~c & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~k & (i0 & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~k & (i0 & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~k & (i0 & (~c & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~k & (i0 & (~c & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~k & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~k & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~k & (~o & (~j0 & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~k & (~o & (~j0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~i & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~k & (~o & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~k & (~o & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~j & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (~g0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~l & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~t & (~r & (~q & (~l & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (~g0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~g0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~h & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((i0 & (~c & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~i & (~h & (~g & (~f & ~e)))))))))))))))))) | ((~c & (~o & (~j0 & (~g0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~g & (~f & ~e)))))))))))))))))) | ((~c & (~o & (~j0 & (~s & (d & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~t & (~r & (~q & (~l & (~j & (~i & (~g & (~f & ~e)))))))))))))))))) | ((~o & (~j0 & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (n & (~j & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~o & (~j0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (n & (~j & (~i & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~o & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (n & (~j & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~o & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))))) | ((~m & (~j0 & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~g & (~f & (~e & ~a))))))))))))))))) | ((~m & (~j0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~i & (~g & (~f & (~e & ~a))))))))))))))))) | ((~m & (~g0 & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~h & (~g & (~f & (~e & ~a))))))))))))))))) | ((~m & (l0 & (~h0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~i & (~h & (~g & (~f & (~e & ~a))))))))))))))))) | ((~b & (~i0 & (~c & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & ~e))))))))))))))))) | ((~b & (~i0 & (~c & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~b & (i0 & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~g & (~f & ~e))))))))))))))))) | ((~b & (i0 & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~i & (~g & (~f & ~e))))))))))))))))) | ((~b & (i0 & (~c & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~h & (~g & (~f & ~e))))))))))))))))) | ((~b & (i0 & (~c & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~b & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~g & (~f & ~e))))))))))))))))) | ((~b & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & (~i & (~g & (~f & ~e))))))))))))))))) | ((~b & (~o & (~j0 & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~g & (~f & (~e & ~a))))))))))))))))) | ((~b & (~o & (~j0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~i & (~g & (~f & (~e & ~a))))))))))))))))) | ((~b & (~o & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~h & (~g & (~f & (~e & ~a))))))))))))))))) | ((~b & (~o & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~i & (~h & (~g & (~f & (~e & ~a))))))))))))))))) | ((~k & (~i0 & (~c & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (~i0 & (~c & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (i0 & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~g & (~f & ~e))))))))))))))))) | ((~k & (i0 & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((~k & (i0 & (~c & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (i0 & (~c & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~k & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~j & (~g & (~f & ~e))))))))))))))))) | ((~k & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((~i0 & (~c & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~g & (~f & ~e))))))))))))))))) | ((i0 & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((i0 & (~c & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~h & (~g & (~f & ~e))))))))))))))))) | ((i0 & (~c & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~i & (~h & (~g & (~f & ~e))))))))))))))))) | ((~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~g & (~f & ~e))))))))))))))))) | ((~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (n & (~j & (~i & (~g & (~f & ~e))))))))))))))))) | ((~m & (~i0 & (~c & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~h & (~g & (~f & ~e)))))))))))))))) | ((~m & (~i0 & (~c & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & ~e)))))))))))))))) | ((~m & (i0 & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & (~g & (~f & ~e)))))))))))))))) | ((~m & (i0 & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & (~i & (~g & (~f & ~e)))))))))))))))) | ((~m & (i0 & (~c & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & (~h & (~g & (~f & ~e)))))))))))))))) | ((~m & (i0 & (~c & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & (~i & (~h & (~g & (~f & ~e)))))))))))))))) | ((~m & (~c & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~n & (~g & (~f & ~e)))))))))))))))) | ((~m & (~c & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~n & (~i & (~g & (~f & ~e)))))))))))))))) | ((~m & (~o & (~j0 & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~g & (~f & (~e & ~a)))))))))))))))) | ((~m & (~o & (~j0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~i & (~g & (~f & (~e & ~a)))))))))))))))) | ((~m & (~o & (~g0 & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~h & (~g & (~f & (~e & ~a)))))))))))))))) | ((~m & (~o & (l0 & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~i & (~h & (~g & (~f & (~e & ~a)))))))))))))))) | ((~b & (~i0 & (~c & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~h & (~g & (~f & ~e)))))))))))))))) | ((~b & (~i0 & (~c & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & ~e)))))))))))))))) | ((~b & (i0 & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~g & (~f & ~e)))))))))))))))) | ((~b & (i0 & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~i & (~g & (~f & ~e)))))))))))))))) | ((~b & (i0 & (~c & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~h & (~g & (~f & ~e)))))))))))))))) | ((~b & (i0 & (~c & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~i & (~h & (~g & (~f & ~e)))))))))))))))) | ((~b & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~g & (~f & ~e)))))))))))))))) | ((~b & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~i & (~g & (~f & ~e)))))))))))))))) | ((~m & (~i0 & (~c & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~i0 & (~c & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (i0 & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~g & (~f & ~e))))))))))))))) | ((~m & (i0 & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~i & (~g & (~f & ~e))))))))))))))) | ((~m & (i0 & (~c & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (i0 & (~c & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~i & (~h & (~g & (~f & ~e))))))))))))))) | ((~m & (~c & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~g & (~f & ~e))))))))))))))) | ((~m & (~c & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~i & (~g & (~f & ~e))))))))))))))) | ((~e0 & (~m & (~j0 & (~g0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & ~a)))))))))))))) | ((~e0 & (~m & (~j0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~i & ~a)))))))))))))) | ((~e0 & (~m & (~g0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~h & ~a)))))))))))))) | ((~e0 & (~m & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~n & (~i & (~h & ~a)))))))))))))) | ((~e0 & (~j0 & (~g0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & ~a)))))))))))))) | ((~e0 & (~j0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~i & ~a)))))))))))))) | ((~e0 & (~g0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~h & ~a)))))))))))))) | ((~e0 & (l0 & (~h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~n & (~i & (~h & ~a)))))))))))))) | ((f0 & (~e0 & (~m & (~i0 & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~n))))))))))))) | ((f0 & (~e0 & (~m & (i0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & ~n))))))))))))) | ((f0 & (~e0 & (~m & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & ~n))))))))))))) | ((f0 & (~e0 & (~i0 & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n))))))))))))) | ((f0 & (~e0 & (i0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & ~n))))))))))))) | ((f0 & (~e0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & ~n))))))))))))) | ((~e0 & (~m & (~i0 & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & (~i & ~h))))))))))))) | ((~e0 & (~m & (i0 & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & ~i))))))))))))) | ((~e0 & (~m & (i0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & (~i & ~h))))))))))))) | ((~e0 & (~m & (~o & (~j0 & (~g0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & ~a))))))))))))) | ((~e0 & (~m & (~o & (~j0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~i & ~a))))))))))))) | ((~e0 & (~m & (~o & (~g0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~h & ~a))))))))))))) | ((~e0 & (~m & (~o & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~q & (~i & (~h & ~a))))))))))))) | ((~e0 & (~m & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~n & ~i))))))))))))) | ((~e0 & (~i0 & (j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & (~i & ~h))))))))))))) | ((~e0 & (i0 & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & ~i))))))))))))) | ((~e0 & (i0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & (~i & ~h))))))))))))) | ((~e0 & (~o & (~j0 & (~g0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & ~a))))))))))))) | ((~e0 & (~o & (~j0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~i & ~a))))))))))))) | ((~e0 & (~o & (~g0 & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~h & ~a))))))))))))) | ((~e0 & (~o & (l0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & (~i & (~h & ~a))))))))))))) | ((~e0 & (~j0 & (l0 & (~h0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & ~i))))))))))))) | ((f0 & (~e0 & (~m & (~i0 & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & ~q)))))))))))) | ((f0 & (~e0 & (~m & (i0 & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & ~q)))))))))))) | ((f0 & (~e0 & (~m & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & ~q)))))))))))) | ((f0 & (~e0 & (~i0 & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & ~q)))))))))))) | ((f0 & (~e0 & (i0 & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & ~q)))))))))))) | ((f0 & (~e0 & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & ~q)))))))))))) | ((~e0 & (~m & (~i0 & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (i0 & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & ~i)))))))))))) | ((~e0 & (~m & (i0 & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~i & ~h)))))))))))) | ((~e0 & (~m & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & ~i)))))))))))) | ((~e0 & (~i0 & (~o & (j0 & (l0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~i & ~h)))))))))))) | ((~e0 & (i0 & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & ~i)))))))))))) | ((~e0 & (i0 & (~o & (l0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~i & ~h)))))))))))) | ((~e0 & (~o & (~j0 & (l0 & (~d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & ~i)))))))))))) | ((z & (~m & (~i0 & (~o & (j0 & (h0 & (~c0 & (~b0 & (~\x  & (u & ~q)))))))))) | ((z & (~m & (~i0 & (j0 & (h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & ~n)))))))))) | ((z & (~m & (~i0 & (j0 & (h0 & (~c0 & (~b0 & (~\x  & (u & (~q & ~n)))))))))) | ((z & (~m & (i0 & (~o & (h0 & (~c0 & (~b0 & (~y & (~\x  & (u & ~q)))))))))) | ((z & (~m & (i0 & (h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & ~n)))))))))) | ((z & (~m & (i0 & (h0 & (~c0 & (~b0 & (~y & (~\x  & (u & (~q & ~n)))))))))) | ((z & (~i0 & (~o & (j0 & (h0 & (~c0 & (~b0 & (~\x  & (u & (~r & ~q)))))))))) | ((z & (~i0 & (j0 & (h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n)))))))))) | ((z & (~i0 & (j0 & (h0 & (~c0 & (~b0 & (~\x  & (u & (~r & (~q & ~n)))))))))) | ((z & (i0 & (~o & (h0 & (~c0 & (~b0 & (~y & (~\x  & (u & (~r & ~q)))))))))) | ((z & (i0 & (h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & ~n)))))))))) | ((z & (i0 & (h0 & (~c0 & (~b0 & (~y & (~\x  & (u & (~r & (~q & ~n)))))))))) | ((~f0 & (~e0 & (~i0 & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~a0 & ~y)))))))))) | ((~f0 & (~e0 & (~i0 & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~a0 & ~y)))))))))) | ((~f0 & (~e0 & (i0 & (~o & (~j0 & (~g0 & (l0 & (~d0 & (~c0 & (~y & ~\x )))))))))) | ((~f0 & (~e0 & (i0 & (~o & (~g0 & (l0 & (~d0 & (~c0 & (~y & (~\x  & ~h)))))))))) | ((~f0 & (~e0 & (i0 & (~j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~y & ~\x )))))))))) | ((~f0 & (~e0 & (i0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & (~y & (~\x  & ~h)))))))))) | ((f0 & (~m & (~i0 & (~o & (j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & h)))))))))) | ((f0 & (~m & (~i0 & (~o & (j0 & (~c0 & (~b0 & (~\x  & (u & (~q & h)))))))))) | ((f0 & (~m & (~i0 & (j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (~n & h)))))))))) | ((f0 & (~m & (~i0 & (j0 & (~c0 & (~b0 & (~\x  & (u & (~q & (~n & h)))))))))) | ((f0 & (~m & (i0 & (~o & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & h)))))))))) | ((f0 & (~m & (i0 & (~o & (~c0 & (~b0 & (~y & (~\x  & (u & (~q & h)))))))))) | ((f0 & (~m & (i0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (~n & h)))))))))) | ((f0 & (~m & (i0 & (~c0 & (~b0 & (~y & (~\x  & (u & (~q & (~n & h)))))))))) | ((f0 & (~i0 & (~o & (j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & h)))))))))) | ((f0 & (~i0 & (~o & (j0 & (~c0 & (~b0 & (~\x  & (u & (~r & (~q & h)))))))))) | ((f0 & (~i0 & (j0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (~n & h)))))))))) | ((f0 & (~i0 & (j0 & (~c0 & (~b0 & (~\x  & (u & (~r & (~q & (~n & h)))))))))) | ((f0 & (i0 & (~o & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & h)))))))))) | ((f0 & (i0 & (~o & (~c0 & (~b0 & (~y & (~\x  & (u & (~r & (~q & h)))))))))) | ((f0 & (i0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (~n & h)))))))))) | ((f0 & (i0 & (~c0 & (~b0 & (~y & (~\x  & (u & (~r & (~q & (~n & h)))))))))) | ((c & (~o & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & ~q)))))))))) | ((c & (d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~u & (~r & (~q & ~n)))))))))) | ((v & (~m & (~i0 & (~o & (j0 & (d0 & (~c0 & (~b0 & (~\x  & ~q))))))))) | ((v & (~m & (~i0 & (j0 & (d0 & (~c0 & (~b0 & (~\x  & (~q & ~n))))))))) | ((v & (~m & (i0 & (~o & (d0 & (~c0 & (~b0 & (~y & (~\x  & ~q))))))))) | ((v & (~m & (i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & ~n))))))))) | ((v & (~i0 & (~o & (j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & ~q))))))))) | ((v & (~i0 & (j0 & (d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & ~n))))))))) | ((v & (i0 & (~o & (d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & ~q))))))))) | ((v & (i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & ~n))))))))) | ((z & (~f0 & (~e0 & (~i0 & (~g0 & (h0 & (~c0 & (~a0 & (~y & u))))))))) | ((z & (~f0 & (~e0 & (i0 & (~g0 & (h0 & (~c0 & (~y & (~\x  & u))))))))) | ((z & (~m & (h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & ~n))))))))) | ((z & (h0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & ~n))))))))) | ((~f0 & (~e0 & (~i0 & (~o & (j0 & (~g0 & (l0 & (~d0 & (~c0 & ~h))))))))) | ((~f0 & (~e0 & (~i0 & (j0 & (~g0 & (l0 & (~h0 & (~d0 & (~c0 & ~h))))))))) | ((f0 & (~m & (~o & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & h))))))))) | ((f0 & (~m & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~q & (~n & h))))))))) | ((f0 & (~o & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & h))))))))) | ((f0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~r & (~q & (~n & h))))))))) | ((v & (~f0 & (~e0 & (~i0 & (~g0 & (d0 & (~c0 & (~a0 & ~y)))))))) | ((v & (~f0 & (~e0 & (i0 & (~g0 & (d0 & (~c0 & (~y & ~\x )))))))) | ((z & (~f0 & (~e0 & (~i0 & (j0 & (~g0 & (h0 & (~c0 & u)))))))) | ((v & (~f0 & (~e0 & (~i0 & (j0 & (~g0 & (d0 & ~c0))))))) | (j2 | (i2 | (h2 | (g2 | (f2 | (e2 | (d2 | (c2 | (b2 | (a2 | (y1 | (x1 | (w1 | (u1 | (r1 | (q1 | (p1 | (o1 | (n1 | (m1 | (l1 | (k1 | (j1 | (i1 | (h1 | (g1 | (z0 | (y0 | (x0 | w0)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  r1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (v & (~q & (~n & ~m))))))))),
  \[2]  = (~m & (~d & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~m & (~d & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~m & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~m & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c)))))))))))))))) | ((~d & (~b & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~d & (~b & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~d0 & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (~d0 & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (~d0 & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (~d0 & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (t & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (t & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (t & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (t & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c)))))))))))))))) | ((~b & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((~b & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c)))))))))))))))) | ((d & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (i0 & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~s & (~j & ~c))))))))))))))) | ((d & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~s & (~j & ~c))))))))))))))) | ((d & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~s & (~j & ~c))))))))))))))) | ((d & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~s & (~j & ~c))))))))))))))) | ((d & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~s & (~j & ~c))))))))))))))) | ((i0 & (~d0 & (~t & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & (~l & (~j & ~c))))))))))))))) | ((i0 & (~d0 & (~t & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & (~l & (~j & ~c))))))))))))))) | ((i0 & (~d0 & (~t & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~l & (~j & ~c))))))))))))))) | ((i0 & (~d0 & (~t & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~l & (~j & ~c))))))))))))))) | ((~d0 & (~t & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~l & (~j & ~c))))))))))))))) | ((~d0 & (~t & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~l & (~j & ~c))))))))))))))) | ((~d0 & (~t & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~l & (~j & ~c))))))))))))))) | ((~d0 & (~t & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~l & (~j & ~c))))))))))))))) | ((~t & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~l & (~j & ~c))))))))))))))) | ((~t & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~l & (~j & ~c))))))))))))))) | ((~t & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~l & (~j & ~c))))))))))))))) | ((~t & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~l & (~j & ~c))))))))))))))) | ((~k & (~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~m & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~m & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~m & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~m & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (i0 & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (~d0 & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (~d0 & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (~d0 & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (j & ~c)))))))))))))) | ((~k & (~b & (~i & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~b & (~i & (~g & (~f & (~e & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~b & (~g & (~f & (~e & (~h0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (~b & (~g & (~f & (~e & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c)))))))))))))) | ((~k & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & (~j & ~c)))))))))))))) | ((~k & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & (~j & ~c)))))))))))))) | ((~k & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (~j & ~c)))))))))))))) | ((~k & (i0 & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (~j & ~c)))))))))))))) | ((~k & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~j & ~c)))))))))))))) | ((~k & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~j & ~c)))))))))))))) | ((~k & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~j & ~c)))))))))))))) | ((~k & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~j & ~c)))))))))))))) | ((~k & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (~j & ~c)))))))))))))) | ((~k & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (~j & ~c)))))))))))))) | ((~k & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~j & ~c)))))))))))))) | ((~k & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~j & ~c)))))))))))))) | ((k & (m & (~d & (t & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~n)))))))))))))) | ((k & (m & (~d & (t & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~n)))))))))))))) | ((k & (m & (~d & (t & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~n)))))))))))))) | ((k & (m & (~d & (t & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~n)))))))))))))) | ((k & (m & (~d & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & l)))))))))))))) | ((k & (m & (~d & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & l)))))))))))))) | ((k & (m & (~d & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & l)))))))))))))) | ((k & (m & (~d & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & l)))))))))))))) | ((k & (m & (t & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & ~n)))))))))))))) | ((k & (m & (t & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & ~n)))))))))))))) | ((k & (m & (t & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & ~n)))))))))))))) | ((k & (m & (t & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & ~n)))))))))))))) | ((k & (m & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & l)))))))))))))) | ((k & (m & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & l)))))))))))))) | ((k & (m & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & l)))))))))))))) | ((k & (m & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & l)))))))))))))) | ((d & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & (~s & (~j & ~c)))))))))))))) | ((d & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & (~s & (~j & ~c)))))))))))))) | ((d & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & (~s & (~j & ~c)))))))))))))) | ((d & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & (~s & (~j & ~c)))))))))))))) | ((d & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~s & (~j & ~c)))))))))))))) | ((d & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & (~s & (~j & ~c)))))))))))))) | ((d & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & (~s & (~j & ~c)))))))))))))) | ((d & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~s & (~j & ~c)))))))))))))) | ((d & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~s & (~j & ~c)))))))))))))) | ((~i0 & (~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & (~l & (~j & ~c)))))))))))))) | ((~i0 & (~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & (~l & (~j & ~c)))))))))))))) | ((~i0 & (~d0 & (~t & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & (~l & (~j & ~c)))))))))))))) | ((~i0 & (~d0 & (~t & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & (~l & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & (~l & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & (~l & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~t & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & (~l & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~t & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & (~l & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & (n & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & (n & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & (n & (~j & ~c)))))))))))))) | ((i0 & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & (n & (~j & ~c)))))))))))))) | ((~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~l & (~j & ~c)))))))))))))) | ((~d0 & (~t & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~l & (~j & ~c)))))))))))))) | ((~d0 & (~t & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~l & (~j & ~c)))))))))))))) | ((~d0 & (~t & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~l & (~j & ~c)))))))))))))) | ((~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (n & (~j & ~c)))))))))))))) | ((~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (n & (~j & ~c)))))))))))))) | ((~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (n & (~j & ~c)))))))))))))) | ((~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (n & (~j & ~c)))))))))))))) | ((~t & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & (~l & (~j & ~c)))))))))))))) | ((~t & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & (~l & (~j & ~c)))))))))))))) | ((~t & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~l & (~j & ~c)))))))))))))) | ((~t & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~l & (~j & ~c)))))))))))))) | ((~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & (n & (~j & ~c)))))))))))))) | ((~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & (n & (~j & ~c)))))))))))))) | ((~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (n & (~j & ~c)))))))))))))) | ((~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (n & (~j & ~c)))))))))))))) | ((~k & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & (~j & ~c))))))))))))) | ((~k & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & (~j & ~c))))))))))))) | ((~k & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & (~j & ~c))))))))))))) | ((~k & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & (~j & ~c))))))))))))) | ((~k & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & (~j & ~c))))))))))))) | ((~k & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & (~j & ~c))))))))))))) | ((~k & (i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & (~j & ~c))))))))))))) | ((~k & (i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & (~j & ~c))))))))))))) | ((~k & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~j & ~c))))))))))))) | ((~k & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~j & ~c))))))))))))) | ((~k & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~j & ~c))))))))))))) | ((~k & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~j & ~c))))))))))))) | ((~k & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & (~j & ~c))))))))))))) | ((~k & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & (~j & ~c))))))))))))) | ((~k & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (~j & ~c))))))))))))) | ((~k & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (~j & ~c))))))))))))) | ((k & (m & (~d & (t & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~n))))))))))))) | ((k & (m & (~d & (t & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~n))))))))))))) | ((k & (m & (~d & (t & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~n))))))))))))) | ((k & (m & (~d & (t & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~n))))))))))))) | ((k & (m & (~d & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & l))))))))))))) | ((k & (m & (~d & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & l))))))))))))) | ((k & (m & (~d & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & l))))))))))))) | ((k & (m & (~d & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & l))))))))))))) | ((k & (m & (t & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & ~n))))))))))))) | ((k & (m & (t & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & ~n))))))))))))) | ((k & (m & (t & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & ~n))))))))))))) | ((k & (m & (t & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & ~n))))))))))))) | ((k & (m & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & l))))))))))))) | ((k & (m & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & l))))))))))))) | ((k & (m & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & l))))))))))))) | ((k & (m & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & l))))))))))))) | ((~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & ~c))))))))))))) | ((~m & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & ~c))))))))))))) | ((~m & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & ~c))))))))))))) | ((~m & (i0 & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & ~c))))))))))))) | ((~m & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & ~c))))))))))))) | ((~m & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & ~c))))))))))))) | ((~m & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & ~c))))))))))))) | ((~m & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & ~c))))))))))))) | ((~m & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))))))) | ((~m & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))))))) | ((~m & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))))))) | ((~m & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))))))) | ((m & (~d & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & j))))))))))))) | ((m & (~d & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & j))))))))))))) | ((m & (~d & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & j))))))))))))) | ((m & (~d & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & j))))))))))))) | ((m & (~d & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & j))))))))))))) | ((m & (~d & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & j))))))))))))) | ((m & (~d & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & j))))))))))))) | ((m & (~d & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & j))))))))))))) | ((m & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & j))))))))))))) | ((m & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & j))))))))))))) | ((m & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & j))))))))))))) | ((m & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & j))))))))))))) | ((m & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & j))))))))))))) | ((m & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & j))))))))))))) | ((m & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & j))))))))))))) | ((m & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & j))))))))))))) | ((~d & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c))))))))))))) | ((~d & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c))))))))))))) | ((~d & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (j & ~c))))))))))))) | ((~d & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (j & ~c))))))))))))) | ((~d & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c))))))))))))) | ((~d & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c))))))))))))) | ((~d & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (~n & (l & (j & ~c))))))))))))) | ((~d & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (~n & (l & (j & ~c))))))))))))) | ((~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~y & ~c))))))))))))) | ((~b & (i0 & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~z & (~y & ~c))))))))))))) | ((~b & (i0 & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~y & ~c))))))))))))) | ((~b & (i0 & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~z & (~y & ~c))))))))))))) | ((~b & (~d0 & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & ~c))))))))))))) | ((~b & (~d0 & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & ~c))))))))))))) | ((~b & (~d0 & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & ~c))))))))))))) | ((~b & (~d0 & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & ~c))))))))))))) | ((~b & (~i & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))))))) | ((~b & (~i & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))))))) | ((~b & (~g & (~f & (~e & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))))))) | ((~b & (~g & (~f & (~e & (~f0 & (m0 & (~j0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))))))) | ((~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & (n & (~j & ~c))))))))))))) | ((~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & (n & (~j & ~c))))))))))))) | ((~i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & (n & (~j & ~c))))))))))))) | ((~i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & (n & (~j & ~c))))))))))))) | ((i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & (n & (~j & ~c))))))))))))) | ((i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & (n & (~j & ~c))))))))))))) | ((i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & (n & (~j & ~c))))))))))))) | ((i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & (n & (~j & ~c))))))))))))) | ((~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (n & (~j & ~c))))))))))))) | ((~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (n & (~j & ~c))))))))))))) | ((~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (n & (~j & ~c))))))))))))) | ((~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (n & (~j & ~c))))))))))))) | ((t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c))))))))))))) | ((t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c))))))))))))) | ((t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (j & ~c))))))))))))) | ((t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (j & ~c))))))))))))) | ((~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & (n & (~j & ~c))))))))))))) | ((~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & (n & (~j & ~c))))))))))))) | ((~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c))))))))))))) | ((~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c))))))))))))) | ((~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & (n & (~j & ~c))))))))))))) | ((~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & (n & (~j & ~c))))))))))))) | ((~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (s & (~n & (l & (j & ~c))))))))))))) | ((m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (s & (~n & (l & (j & ~c))))))))))))) | ((~m & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & ~c)))))))))))) | ((~m & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & ~c)))))))))))) | ((~m & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & ~c)))))))))))) | ((~m & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & ~c)))))))))))) | ((~m & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & ~c)))))))))))) | ((~m & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & ~c)))))))))))) | ((~m & (i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & ~c)))))))))))) | ((~m & (i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & ~c)))))))))))) | ((~m & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & ~c)))))))))))) | ((~m & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & ~c)))))))))))) | ((~m & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & ~c)))))))))))) | ((~m & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & ~c)))))))))))) | ((~m & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))))) | ((~m & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))))) | ((~m & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))))) | ((~m & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))))) | ((~d & (i0 & (~d0 & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~y & (~n & j)))))))))))) | ((~d & (i0 & (~d0 & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~z & (~y & (~n & j)))))))))))) | ((~d & (i0 & (~d0 & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~y & (~n & j)))))))))))) | ((~d & (i0 & (~d0 & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & (~y & (~n & j)))))))))))) | ((~d & (i0 & (~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~y & (~n & (l & j)))))))))))) | ((~d & (i0 & (~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~z & (~y & (~n & (l & j)))))))))))) | ((~d & (i0 & (~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~y & (~n & (l & j)))))))))))) | ((~d & (i0 & (~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & (~y & (~n & (l & j)))))))))))) | ((~d & (~d0 & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~n & j)))))))))))) | ((~d & (~d0 & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~n & j)))))))))))) | ((~d & (~d0 & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~n & j)))))))))))) | ((~d & (~d0 & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~n & j)))))))))))) | ((~d & (~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~n & (l & j)))))))))))) | ((~d & (~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & j)))))))))))) | ((~d & (~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~n & (l & j)))))))))))) | ((~d & (~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~n & (l & j)))))))))))) | ((~b & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~c0 & ~c)))))))))))) | ((~b & (~i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (j0 & (~c0 & (~z & ~c)))))))))))) | ((~b & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (j0 & (~g0 & (~c0 & ~c)))))))))))) | ((~b & (~i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (j0 & (~g0 & (~c0 & (~z & ~c)))))))))))) | ((~b & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~y & ~c)))))))))))) | ((~b & (i0 & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~z & (~y & ~c)))))))))))) | ((~b & (i0 & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~y & ~c)))))))))))) | ((~b & (i0 & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~z & (~y & ~c)))))))))))) | ((~b & (~d0 & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & ~c)))))))))))) | ((~b & (~d0 & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & ~c)))))))))))) | ((~b & (~d0 & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & ~c)))))))))))) | ((~b & (~d0 & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & ~c)))))))))))) | ((~b & (~i & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))))) | ((~b & (~i & (~h & (~g & (~f & (~e & (m0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))))) | ((~b & (~h & (~g & (~f & (~e & (~h0 & (m0 & (~g0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))))) | ((~b & (~h & (~g & (~f & (~e & (m0 & (~g0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))))) | ((i0 & (~d0 & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~y & (s & (~n & j)))))))))))) | ((i0 & (~d0 & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~z & (~y & (s & (~n & j)))))))))))) | ((i0 & (~d0 & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~y & (s & (~n & j)))))))))))) | ((i0 & (~d0 & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & (~y & (s & (~n & j)))))))))))) | ((i0 & (~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~y & (s & (~n & (l & j)))))))))))) | ((i0 & (~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~z & (~y & (s & (~n & (l & j)))))))))))) | ((i0 & (~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~y & (s & (~n & (l & j)))))))))))) | ((i0 & (~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & (~y & (s & (~n & (l & j)))))))))))) | ((~d0 & (t & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (s & (~n & j)))))))))))) | ((~d0 & (t & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & j)))))))))))) | ((~d0 & (t & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (s & (~n & j)))))))))))) | ((~d0 & (t & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & j)))))))))))) | ((~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (s & (~n & (l & j)))))))))))) | ((~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & j)))))))))))) | ((~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (s & (~n & (l & j)))))))))))) | ((~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (s & (~n & (l & j)))))))))))) | ((~k & (m & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j))))))))))) | ((~k & (m & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j))))))))))) | ((~k & (m & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j))))))))))) | ((~k & (m & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j))))))))))) | ((~k & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (j & ~c))))))))))) | ((~k & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c))))))))))) | ((~k & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & (j & ~c))))))))))) | ((~k & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & (j & ~c))))))))))) | ((m & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j))))))))))) | ((m & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j))))))))))) | ((m & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j))))))))))) | ((m & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j))))))))))) | ((~k & (i0 & (~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~y & j)))))))))) | ((~k & (i0 & (~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~z & (~y & j)))))))))) | ((~k & (i0 & (~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~y & j)))))))))) | ((~k & (i0 & (~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & (~y & j)))))))))) | ((~k & (~d0 & (~i & (~h0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & j)))))))))) | ((~k & (~d0 & (~i & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & j)))))))))) | ((~k & (~d0 & (~h0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & j)))))))))) | ((~k & (~d0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & j)))))))))) | ((m & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j)))))))))) | ((m & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j)))))))))) | ((m & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & j)))))))))) | ((m & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & j)))))))))) | ((~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))) | ((~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))) | ((~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~c)))))))))) | ((~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c)))))))))) | ((i0 & (~d0 & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & ~y))))))))) | ((i0 & (~d0 & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~z & ~y))))))))) | ((i0 & (~d0 & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & ~y))))))))) | ((i0 & (~d0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~z & ~y))))))))) | ((~d0 & (~i & (~h0 & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & ~y))))))))) | ((~d0 & (~i & (~f0 & (m0 & (~j0 & (~e0 & (~c0 & (~a0 & (~z & ~y))))))))) | ((~d0 & (~h0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & ~y))))))))) | ((~d0 & (~f0 & (m0 & (~j0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & ~y))))))))) | ((~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))) | ((~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))) | ((~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~y & (~w & ~c))))))))) | ((~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & (~y & (~w & ~c))))))))) | ((~i0 & (~d0 & (~i & (~h & (~h0 & (m0 & (j0 & (~e0 & ~c0)))))))) | ((~i0 & (~d0 & (~i & (~h & (m0 & (j0 & (~e0 & (~c0 & ~z)))))))) | ((~i0 & (~d0 & (~h & (~h0 & (m0 & (j0 & (~g0 & (~e0 & ~c0)))))))) | ((~i0 & (~d0 & (~h & (m0 & (j0 & (~g0 & (~e0 & (~c0 & ~z)))))))) | ((i0 & (~d0 & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & ~y)))))))) | ((i0 & (~d0 & (~i & (~h & (m0 & (~e0 & (~c0 & (~z & ~y)))))))) | ((i0 & (~d0 & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & ~y)))))))) | ((i0 & (~d0 & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~z & ~y)))))))) | ((~d0 & (~i & (~h & (~h0 & (m0 & (~e0 & (~c0 & (~a0 & ~y)))))))) | ((~d0 & (~i & (~h & (m0 & (~e0 & (~c0 & (~a0 & (~z & ~y)))))))) | ((~d0 & (~h & (~h0 & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & ~y)))))))) | ((~d0 & (~h & (m0 & (~g0 & (~e0 & (~c0 & (~a0 & (~z & ~y)))))))) | ((r & (m & (~i0 & (~d0 & (f0 & (j0 & ~c0)))))) | ((r & (m & (~i0 & (~d0 & (j0 & (g0 & ~c0)))))) | ((r & (m & (~i0 & (~d0 & (j0 & (e0 & ~c0)))))) | ((r & (m & (~i0 & (f0 & (j0 & (~c0 & w)))))) | ((r & (m & (~i0 & (j0 & (g0 & (~c0 & w)))))) | ((r & (m & (~i0 & (j0 & (e0 & (~c0 & w)))))) | ((r & (m & (i0 & (~d0 & (f0 & (~c0 & ~y)))))) | ((r & (m & (i0 & (~d0 & (g0 & (~c0 & ~y)))))) | ((r & (m & (i0 & (~d0 & (e0 & (~c0 & ~y)))))) | ((r & (m & (i0 & (f0 & (~c0 & (~y & w)))))) | ((r & (m & (i0 & (g0 & (~c0 & (~y & w)))))) | ((r & (m & (i0 & (e0 & (~c0 & (~y & w)))))) | ((r & (m & (d0 & (~c0 & (~a0 & (~y & ~w)))))) | ((~i0 & (~d0 & (o & (f0 & (j0 & (~c0 & n)))))) | ((~i0 & (~d0 & (o & (j0 & (g0 & (~c0 & n)))))) | ((~i0 & (~d0 & (o & (j0 & (e0 & (~c0 & n)))))) | ((~i0 & (o & (f0 & (j0 & (~c0 & (w & n)))))) | ((~i0 & (o & (j0 & (g0 & (~c0 & (w & n)))))) | ((~i0 & (o & (j0 & (e0 & (~c0 & (w & n)))))) | ((i0 & (~d0 & (o & (f0 & (~c0 & (~y & n)))))) | ((i0 & (~d0 & (o & (g0 & (~c0 & (~y & n)))))) | ((i0 & (~d0 & (o & (e0 & (~c0 & (~y & n)))))) | ((i0 & (o & (f0 & (~c0 & (~y & (w & n)))))) | ((i0 & (o & (g0 & (~c0 & (~y & (w & n)))))) | ((i0 & (o & (e0 & (~c0 & (~y & (w & n)))))) | ((d0 & (o & (~c0 & (~a0 & (~y & (~w & n)))))) | ((v & (~i0 & (d0 & (j0 & (~c0 & ~w))))) | ((v & (i0 & (d0 & (~c0 & (~y & ~w))))) | ((u & (~i0 & (d0 & (j0 & (~c0 & ~w))))) | ((u & (i0 & (d0 & (~c0 & (~y & ~w))))) | ((r & (m & (f0 & (~c0 & (~a0 & ~y))))) | ((r & (m & (g0 & (~c0 & (~a0 & ~y))))) | ((r & (m & (e0 & (~c0 & (~a0 & ~y))))) | ((b0 & (~i0 & (~d0 & (f0 & (j0 & ~c0))))) | ((b0 & (~i0 & (~d0 & (j0 & (g0 & ~c0))))) | ((b0 & (~i0 & (~d0 & (j0 & (e0 & ~c0))))) | ((b0 & (~i0 & (f0 & (j0 & (~c0 & w))))) | ((b0 & (~i0 & (j0 & (g0 & (~c0 & w))))) | ((b0 & (~i0 & (j0 & (e0 & (~c0 & w))))) | ((b0 & (i0 & (~d0 & (f0 & (~c0 & ~y))))) | ((b0 & (i0 & (~d0 & (g0 & (~c0 & ~y))))) | ((b0 & (i0 & (~d0 & (e0 & (~c0 & ~y))))) | ((b0 & (i0 & (f0 & (~c0 & (~y & w))))) | ((b0 & (i0 & (g0 & (~c0 & (~y & w))))) | ((b0 & (i0 & (e0 & (~c0 & (~y & w))))) | ((b0 & (d0 & (~c0 & (~a0 & (~y & ~w))))) | ((q & (~i0 & (~d0 & (f0 & (j0 & ~c0))))) | ((q & (~i0 & (~d0 & (j0 & (g0 & ~c0))))) | ((q & (~i0 & (~d0 & (j0 & (e0 & ~c0))))) | ((q & (~i0 & (f0 & (j0 & (~c0 & w))))) | ((q & (~i0 & (j0 & (g0 & (~c0 & w))))) | ((q & (~i0 & (j0 & (e0 & (~c0 & w))))) | ((q & (i0 & (~d0 & (f0 & (~c0 & ~y))))) | ((q & (i0 & (~d0 & (g0 & (~c0 & ~y))))) | ((q & (i0 & (~d0 & (e0 & (~c0 & ~y))))) | ((q & (i0 & (f0 & (~c0 & (~y & w))))) | ((q & (i0 & (g0 & (~c0 & (~y & w))))) | ((q & (i0 & (e0 & (~c0 & (~y & w))))) | ((q & (d0 & (~c0 & (~a0 & (~y & ~w))))) | ((~i0 & (~d0 & (f0 & (\x  & (j0 & ~c0))))) | ((~i0 & (~d0 & (\x  & (j0 & (g0 & ~c0))))) | ((~i0 & (~d0 & (\x  & (j0 & (e0 & ~c0))))) | ((~i0 & (h0 & (o & (j0 & (~c0 & w))))) | ((~i0 & (f0 & (\x  & (j0 & (~c0 & w))))) | ((~i0 & (\x  & (j0 & (g0 & (~c0 & w))))) | ((~i0 & (\x  & (j0 & (e0 & (~c0 & w))))) | ((i0 & (h0 & (o & (~c0 & (~y & w))))) | ((d0 & (\x  & (~c0 & (~a0 & (~y & ~w))))) | ((o & (f0 & (~c0 & (~a0 & (~y & n))))) | ((o & (g0 & (~c0 & (~a0 & (~y & n))))) | ((o & (e0 & (~c0 & (~a0 & (~y & n))))) | ((b0 & (f0 & (~c0 & (~a0 & ~y)))) | ((b0 & (g0 & (~c0 & (~a0 & ~y)))) | ((b0 & (e0 & (~c0 & (~a0 & ~y)))) | ((q & (f0 & (~c0 & (~a0 & ~y)))) | ((q & (g0 & (~c0 & (~a0 & ~y)))) | ((q & (e0 & (~c0 & (~a0 & ~y)))) | ((i0 & (~d0 & (\x  & (~c0 & ~y)))) | ((i0 & (\x  & (~c0 & (~y & w)))) | ((h0 & (o & (~c0 & (~a0 & ~y)))) | ((f0 & (\x  & (~c0 & (~a0 & ~y)))) | ((\x  & (g0 & (~c0 & (~a0 & ~y)))) | ((\x  & (e0 & (~c0 & (~a0 & ~y)))) | (z1 | (v1 | (u1 | (t1 | (s1 | (r1 | (o1 | (n1 | (f1 | (e1 | (d1 | (c1 | (b1 | a1))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))),
  s1 = j0 & (~i0 & (h0 & (~g0 & (~f0 & (~e0 & (~d0 & (~c0 & o))))))),
  t1 = i0 & (h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~q & (o & (~n & ~m))))))))),
  u1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (v & (~r & (~q & ~n))))))))),
  v1 = i0 & (h0 & (~d0 & (~c0 & (~b0 & (~y & (~\x  & (~r & (~q & (o & ~n))))))))),
  w0 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~v & (~u & (~q & (~o & (~m & c)))))))))),
  w1 = i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (w & (~q & (~o & ~m)))))))),
  x0 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~v & (~u & (~q & (~n & (~m & c)))))))))),
  x1 = i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (w & (~r & (~q & ~o)))))))),
  y0 = j0 & (~i0 & (h0 & (~d0 & (~c0 & (~b0 & (z & (~\x  & (~q & (~o & ~m))))))))),
  y1 = h0 & (~c0 & (~b0 & (~a0 & (z & (~y & (~\x  & (~q & (~o & ~m)))))))),
  z0 = j0 & (~i0 & (h0 & (~d0 & (~c0 & (~b0 & (z & (~\x  & (~r & (~q & ~o))))))))),
  z1 = i0 & (h0 & (~g0 & (~f0 & (~e0 & (~d0 & (~c0 & (~y & (~\x  & o)))))))),
  a1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (~v & (u & (~q & (~o & ~m)))))))))),
  a2 = h0 & (~c0 & (~b0 & (~a0 & (z & (~y & (~\x  & (~r & (~q & ~o)))))))),
  b1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (~v & (u & (~r & (~q & ~o)))))))))),
  b2 = j0 & (~i0 & (~g0 & (~f0 & (~e0 & (d0 & (~c0 & w)))))),
  c1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (~v & (u & (~q & (~n & ~m)))))))))),
  c2 = i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (w & (~q & (~n & ~m)))))))),
  d1 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (~w & (~v & (u & (~r & (~q & ~n)))))))))),
  d2 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (w & (~q & (~o & ~m)))))))),
  e1 = j0 & (~i0 & (h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~q & (o & (~n & ~m))))))))),
  e2 = i0 & (d0 & (~c0 & (~b0 & (~y & (~\x  & (w & (~r & (~q & ~n)))))))),
  f1 = j0 & (~i0 & (h0 & (~d0 & (~c0 & (~b0 & (~\x  & (~r & (~q & (o & ~n))))))))),
  f2 = d0 & (~c0 & (~b0 & (~a0 & (~y & (~\x  & (w & (~r & (~q & ~o))))))));
endmodule

