// IWLS benchmark module "Min_Max9_4" printed on Wed May 29 22:12:22 2002
module Min_Max9_4(\1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \40 , \41 , \42 , \43 , \44 , \45 , \46 , \47 , \48 );
input
  \1 ,
  \2 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ;
output
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ;
reg
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ,
  \34 ,
  \35 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ;
wire
  \[60] ,
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \375 ,
  \376 ,
  \377 ,
  \378 ,
  \379 ,
  \[61] ,
  \380 ,
  \381 ,
  \383 ,
  \384 ,
  \385 ,
  \386 ,
  \387 ,
  \388 ,
  \389 ,
  \[62] ,
  \391 ,
  \392 ,
  \393 ,
  \394 ,
  \395 ,
  \396 ,
  \397 ,
  \399 ,
  \400 ,
  \401 ,
  \402 ,
  \403 ,
  \404 ,
  \405 ,
  \407 ,
  \408 ,
  \409 ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \420 ,
  \421 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \428 ,
  \429 ,
  \430 ,
  \431 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \438 ,
  \439 ,
  \440 ,
  \441 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \463 ,
  \464 ,
  \465 ,
  \466 ,
  \468 ,
  \470 ,
  \471 ,
  \473 ,
  \474 ,
  \476 ,
  \478 ,
  \479 ,
  \481 ,
  \482 ,
  \484 ,
  \486 ,
  \487 ,
  \489 ,
  \490 ,
  \492 ,
  \494 ,
  \495 ,
  \497 ,
  \498 ,
  \500 ,
  \502 ,
  \503 ,
  \505 ,
  \506 ,
  \508 ,
  \510 ,
  \511 ,
  \513 ,
  \514 ,
  \516 ,
  \518 ,
  \519 ,
  \521 ,
  \522 ,
  \524 ,
  \526 ,
  \527 ,
  \529 ,
  \530 ,
  \532 ,
  \534 ,
  \535 ,
  \537 ,
  \538 ,
  \540 ,
  \543 ,
  \546 ,
  \548 ,
  \551 ,
  \554 ,
  \556 ,
  \559 ,
  \562 ,
  \564 ,
  \567 ,
  \570 ,
  \572 ,
  \575 ,
  \578 ,
  \580 ,
  \583 ,
  \586 ,
  \588 ,
  \591 ,
  \594 ,
  \596 ,
  \599 ,
  \602 ,
  \604 ,
  \607 ,
  \610 ,
  \612 ,
  \613 ,
  \614 ,
  \615 ,
  \616 ,
  \617 ,
  \618 ,
  \619 ,
  \620 ,
  \621 ,
  \622 ,
  \623 ,
  \624 ,
  \625 ,
  \626 ,
  \627 ,
  \628 ,
  \629 ,
  \630 ,
  \631 ,
  \632 ,
  \633 ,
  \634 ,
  \635 ,
  \636 ,
  \637 ,
  \638 ,
  \639 ,
  \640 ,
  \641 ,
  \642 ,
  \643 ,
  \644 ,
  \645 ,
  \646 ,
  \647 ,
  \648 ,
  \649 ,
  \650 ,
  \651 ,
  \652 ,
  \653 ,
  \654 ,
  \655 ,
  \656 ,
  \657 ,
  \658 ,
  \659 ,
  \660 ,
  \661 ,
  \662 ,
  \663 ,
  \664 ,
  \665 ,
  \666 ,
  \667 ,
  \668 ,
  \669 ,
  \670 ,
  \671 ,
  \672 ,
  \673 ,
  \674 ,
  \675 ,
  \676 ,
  \677 ,
  \678 ,
  \679 ,
  \680 ,
  \681 ,
  \682 ,
  \683 ,
  \684 ,
  \685 ,
  \686 ,
  \687 ,
  \688 ,
  \689 ,
  \690 ,
  \691 ,
  \692 ,
  \693 ,
  \694 ,
  \695 ,
  \696 ,
  \697 ,
  \698 ,
  \699 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \700 ,
  \66 ,
  \701 ,
  \703 ,
  \705 ,
  \706 ,
  \707 ,
  \708 ,
  \709 ,
  \710 ,
  \711 ,
  \712 ,
  \713 ,
  \714 ,
  \715 ,
  \716 ,
  \717 ,
  \718 ,
  \719 ,
  \83 ,
  \85 ,
  \720 ,
  \721 ,
  \87 ,
  \722 ,
  \723 ,
  \89 ,
  \724 ,
  \725 ,
  \726 ,
  \727 ,
  \728 ,
  \729 ,
  \91 ,
  \93 ,
  \95 ,
  \730 ,
  \97 ,
  \732 ,
  \99 ,
  \734 ,
  \735 ,
  \736 ,
  \737 ,
  \738 ,
  \739 ,
  \740 ,
  \741 ,
  \742 ,
  \743 ,
  \744 ,
  \745 ,
  \746 ,
  \747 ,
  \748 ,
  \749 ,
  \750 ,
  \751 ,
  \752 ,
  \753 ,
  \754 ,
  \755 ,
  \756 ,
  \757 ,
  \758 ,
  \759 ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \103 ,
  \105 ,
  \107 ,
  \109 ,
  \111 ,
  \113 ,
  \115 ,
  \117 ,
  \119 ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \[52] ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ,
  \322 ,
  \323 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \367 ,
  \368 ,
  \369 ;
assign
  \[60]  = \594 ,
  \370  = \369  & \2 ,
  \371  = \15  & ~\2 ,
  \372  = \371  | \370 ,
  \373  = \372  & ~\1 ,
  \375  = \290  & ~\3 ,
  \376  = \7  & \3 ,
  \377  = \376  | \375 ,
  \378  = \377  & \2 ,
  \379  = \16  & ~\2 ,
  \[61]  = \602 ,
  \380  = \379  | \378 ,
  \381  = \380  & ~\1 ,
  \383  = \291  & ~\3 ,
  \384  = \8  & \3 ,
  \385  = \384  | \383 ,
  \386  = \385  & \2 ,
  \387  = \17  & ~\2 ,
  \388  = \387  | \386 ,
  \389  = \388  & ~\1 ,
  \[62]  = \610 ,
  \391  = \292  & ~\3 ,
  \392  = \9  & \3 ,
  \393  = \392  | \391 ,
  \394  = \393  & \2 ,
  \395  = \18  & ~\2 ,
  \396  = \395  | \394 ,
  \397  = \396  & ~\1 ,
  \399  = \293  & ~\3 ,
  \400  = \10  & \3 ,
  \401  = \400  | \399 ,
  \402  = \401  & \2 ,
  \403  = \19  & ~\2 ,
  \404  = \403  | \402 ,
  \405  = \404  & ~\1 ,
  \407  = \294  & ~\3 ,
  \408  = \11  & \3 ,
  \409  = \408  | \407 ,
  \410  = \409  & \2 ,
  \411  = \20  & ~\2 ,
  \412  = \411  | \410 ,
  \413  = \412  & ~\1 ,
  \415  = \286  & ~\3 ,
  \416  = \12  & \3 ,
  \417  = \416  | \415 ,
  \418  = \417  & \2 ,
  \419  = \21  & ~\2 ,
  \420  = \419  | \418 ,
  \421  = \420  & ~\1 ,
  \423  = \4  & \2 ,
  \424  = \13  & ~\2 ,
  \425  = \424  | \423 ,
  \426  = \425  & ~\1 ,
  \428  = \5  & \2 ,
  \429  = \14  & ~\2 ,
  \430  = \429  | \428 ,
  \431  = \430  & ~\1 ,
  \433  = \6  & \2 ,
  \434  = \15  & ~\2 ,
  \435  = \434  | \433 ,
  \436  = \435  & ~\1 ,
  \438  = \7  & \2 ,
  \439  = \16  & ~\2 ,
  \440  = \439  | \438 ,
  \441  = \440  & ~\1 ,
  \443  = \8  & \2 ,
  \444  = \17  & ~\2 ,
  \445  = \444  | \443 ,
  \446  = \445  & ~\1 ,
  \448  = \9  & \2 ,
  \449  = \18  & ~\2 ,
  \450  = \449  | \448 ,
  \451  = \450  & ~\1 ,
  \453  = \10  & \2 ,
  \454  = \19  & ~\2 ,
  \455  = \454  | \453 ,
  \456  = \455  & ~\1 ,
  \458  = \11  & \2 ,
  \459  = \20  & ~\2 ,
  \460  = \459  | \458 ,
  \461  = \460  & ~\1 ,
  \463  = \12  & \2 ,
  \464  = \21  & ~\2 ,
  \465  = \464  | \463 ,
  \466  = \465  & ~\1 ,
  \468  = \326  & ~\3 ,
  \470  = \468  | \3 ,
  \471  = \470  & \2 ,
  \473  = \471  | ~\2 ,
  \474  = \473  & ~\1 ,
  \476  = \329  & ~\3 ,
  \478  = \476  | \3 ,
  \479  = \478  & \2 ,
  \481  = \479  | ~\2 ,
  \482  = \481  & ~\1 ,
  \484  = \332  & ~\3 ,
  \486  = \484  | \3 ,
  \487  = \486  & \2 ,
  \489  = \487  | ~\2 ,
  \490  = \489  & ~\1 ,
  \492  = \335  & ~\3 ,
  \494  = \492  | \3 ,
  \495  = \494  & \2 ,
  \497  = \495  | ~\2 ,
  \498  = \497  & ~\1 ,
  \500  = \338  & ~\3 ,
  \502  = \500  | \3 ,
  \503  = \502  & \2 ,
  \505  = \503  | ~\2 ,
  \506  = \505  & ~\1 ,
  \508  = \341  & ~\3 ,
  \510  = \508  | \3 ,
  \511  = \510  & \2 ,
  \513  = \511  | ~\2 ,
  \514  = \513  & ~\1 ,
  \516  = \344  & ~\3 ,
  \518  = \516  | \3 ,
  \519  = \518  & \2 ,
  \521  = \519  | ~\2 ,
  \522  = \521  & ~\1 ,
  \524  = \347  & ~\3 ,
  \526  = \524  | \3 ,
  \527  = \526  & \2 ,
  \529  = \527  | ~\2 ,
  \530  = \529  & ~\1 ,
  \532  = \350  & ~\3 ,
  \534  = \532  | \3 ,
  \535  = \534  & \2 ,
  \537  = \535  | ~\2 ,
  \538  = \537  & ~\1 ,
  \540  = \325  & ~\3 ,
  \543  = \540  & \2 ,
  \546  = \543  & ~\1 ,
  \548  = \328  & ~\3 ,
  \551  = \548  & \2 ,
  \554  = \551  & ~\1 ,
  \556  = \331  & ~\3 ,
  \559  = \556  & \2 ,
  \562  = \559  & ~\1 ,
  \564  = \334  & ~\3 ,
  \567  = \564  & \2 ,
  \570  = \567  & ~\1 ,
  \572  = \337  & ~\3 ,
  \575  = \572  & \2 ,
  \578  = \575  & ~\1 ,
  \580  = \340  & ~\3 ,
  \583  = \580  & \2 ,
  \586  = \583  & ~\1 ,
  \588  = \343  & ~\3 ,
  \591  = \588  & \2 ,
  \594  = \591  & ~\1 ,
  \596  = \346  & ~\3 ,
  \599  = \596  & \2 ,
  \602  = \599  & ~\1 ,
  \604  = \349  & ~\3 ,
  \607  = \604  & \2 ,
  \610  = \607  & ~\1 ,
  \612  = \323  & \30 ,
  \613  = ~\323  & \12 ,
  \614  = \613  | \612 ,
  \615  = ~\3  & \2 ,
  \616  = \615  & ~\1 ,
  \617  = ~\322  & \39 ,
  \618  = \322  & \12 ,
  \619  = \618  | \617 ,
  \620  = ~\3  & \2 ,
  \621  = \620  & ~\1 ,
  \622  = \323  & \29 ,
  \623  = ~\323  & \11 ,
  \624  = \623  | \622 ,
  \625  = ~\3  & \2 ,
  \626  = \625  & ~\1 ,
  \627  = ~\322  & \38 ,
  \628  = \322  & \11 ,
  \629  = \628  | \627 ,
  \630  = ~\3  & \2 ,
  \631  = \630  & ~\1 ,
  \632  = \323  & \28 ,
  \633  = ~\323  & \10 ,
  \634  = \633  | \632 ,
  \635  = ~\3  & \2 ,
  \636  = \635  & ~\1 ,
  \637  = ~\322  & \37 ,
  \638  = \322  & \10 ,
  \639  = \638  | \637 ,
  \640  = ~\3  & \2 ,
  \641  = \640  & ~\1 ,
  \642  = \323  & \27 ,
  \643  = ~\323  & \9 ,
  \644  = \643  | \642 ,
  \645  = ~\3  & \2 ,
  \646  = \645  & ~\1 ,
  \647  = ~\322  & \36 ,
  \648  = \322  & \9 ,
  \649  = \648  | \647 ,
  \650  = ~\3  & \2 ,
  \651  = \650  & ~\1 ,
  \652  = \323  & \26 ,
  \653  = ~\323  & \8 ,
  \654  = \653  | \652 ,
  \655  = ~\3  & \2 ,
  \656  = \655  & ~\1 ,
  \657  = ~\322  & \35 ,
  \658  = \322  & \8 ,
  \659  = \658  | \657 ,
  \660  = ~\3  & \2 ,
  \661  = \660  & ~\1 ,
  \662  = \323  & \25 ,
  \663  = ~\323  & \7 ,
  \664  = \663  | \662 ,
  \665  = ~\3  & \2 ,
  \666  = \665  & ~\1 ,
  \667  = ~\322  & \34 ,
  \668  = \322  & \7 ,
  \669  = \668  | \667 ,
  \670  = ~\3  & \2 ,
  \671  = \670  & ~\1 ,
  \672  = \323  & \24 ,
  \673  = ~\323  & \6 ,
  \674  = \673  | \672 ,
  \675  = ~\3  & \2 ,
  \676  = \675  & ~\1 ,
  \677  = ~\322  & \33 ,
  \678  = \322  & \6 ,
  \679  = \678  | \677 ,
  \680  = ~\3  & \2 ,
  \681  = \680  & ~\1 ,
  \682  = \323  & \23 ,
  \683  = ~\323  & \5 ,
  \684  = \683  | \682 ,
  \685  = ~\3  & \2 ,
  \686  = \685  & ~\1 ,
  \687  = ~\322  & \32 ,
  \688  = \322  & \5 ,
  \689  = \688  | \687 ,
  \690  = ~\3  & \2 ,
  \691  = \690  & ~\1 ,
  \692  = \323  & \22 ,
  \693  = ~\323  & \4 ,
  \694  = \693  | \692 ,
  \695  = ~\3  & \2 ,
  \696  = \695  & ~\1 ,
  \697  = ~\322  & \31 ,
  \698  = \322  & \4 ,
  \699  = \698  | \697 ,
  \40  = \357 ,
  \41  = \365 ,
  \42  = \373 ,
  \43  = \381 ,
  \44  = \389 ,
  \45  = \397 ,
  \46  = \405 ,
  \47  = \413 ,
  \48  = \421 ,
  \58  = \474  | \1 ,
  \59  = \482  | \1 ,
  \60  = \490  | \1 ,
  \61  = \498  | \1 ,
  \62  = \506  | \1 ,
  \63  = \514  | \1 ,
  \64  = \522  | \1 ,
  \65  = \530  | \1 ,
  \700  = ~\3  & \2 ,
  \66  = \538  | \1 ,
  \701  = \700  & ~\1 ,
  \703  = \119  & \4 ,
  \705  = \703  & ~\117 ,
  \706  = \117  & \5 ,
  \707  = \706  | \705 ,
  \708  = \707  & ~\115 ,
  \709  = \115  & \6 ,
  \710  = \709  | \708 ,
  \711  = \710  & ~\113 ,
  \712  = \113  & \7 ,
  \713  = \712  | \711 ,
  \714  = \713  & ~\111 ,
  \715  = \111  & \8 ,
  \716  = \715  | \714 ,
  \717  = \716  & ~\109 ,
  \718  = \109  & \9 ,
  \719  = \718  | \717 ,
  \83  = (~\12  & \39 ) | (\12  & ~\39 ),
  \85  = (~\11  & \38 ) | (\11  & ~\38 ),
  \720  = \719  & ~\107 ,
  \721  = \107  & \10 ,
  \87  = (~\10  & \37 ) | (\10  & ~\37 ),
  \722  = \721  | \720 ,
  \723  = \722  & ~\105 ,
  \89  = (~\9  & \36 ) | (\9  & ~\36 ),
  \724  = \105  & \11 ,
  \725  = \724  | \723 ,
  \726  = \725  & ~\103 ,
  \727  = \103  & \12 ,
  \728  = \727  | \726 ,
  \729  = ~\3  & \2 ,
  \91  = (~\8  & \35 ) | (\8  & ~\35 ),
  \93  = (~\7  & \34 ) | (\7  & ~\34 ),
  \95  = (~\6  & \33 ) | (\6  & ~\33 ),
  \730  = \729  & ~\1 ,
  \97  = (~\5  & \32 ) | (\5  & ~\32 ),
  \732  = \99  & \4 ,
  \99  = (~\4  & \31 ) | (\4  & ~\31 ),
  \734  = \732  & ~\97 ,
  \735  = \97  & \5 ,
  \736  = \735  | \734 ,
  \737  = \736  & ~\95 ,
  \738  = \95  & \6 ,
  \739  = \738  | \737 ,
  \740  = \739  & ~\93 ,
  \741  = \93  & \7 ,
  \742  = \741  | \740 ,
  \743  = \742  & ~\91 ,
  \744  = \91  & \8 ,
  \745  = \744  | \743 ,
  \746  = \745  & ~\89 ,
  \747  = \89  & \9 ,
  \748  = \747  | \746 ,
  \749  = \748  & ~\87 ,
  \750  = \87  & \10 ,
  \751  = \750  | \749 ,
  \752  = \751  & ~\85 ,
  \753  = \85  & \11 ,
  \754  = \753  | \752 ,
  \755  = \754  & ~\83 ,
  \756  = \83  & \12 ,
  \757  = \756  | \755 ,
  \758  = ~\3  & \2 ,
  \759  = \758  & ~\1 ,
  \[36]  = \426 ,
  \[37]  = \431 ,
  \[38]  = \436 ,
  \[39]  = \441 ,
  \103  = (~\12  & \30 ) | (\12  & ~\30 ),
  \105  = (~\11  & \29 ) | (\11  & ~\29 ),
  \107  = (~\10  & \28 ) | (\10  & ~\28 ),
  \109  = (~\9  & \27 ) | (\9  & ~\27 ),
  \111  = (~\8  & \26 ) | (\8  & ~\26 ),
  \113  = (~\7  & \25 ) | (\7  & ~\25 ),
  \115  = (~\6  & \24 ) | (\6  & ~\24 ),
  \117  = (~\5  & \23 ) | (\5  & ~\23 ),
  \119  = (~\4  & \22 ) | (\4  & ~\22 ),
  \[40]  = \446 ,
  \[41]  = \451 ,
  \[42]  = \456 ,
  \[43]  = \461 ,
  \[44]  = \466 ,
  \[45]  = \58 ,
  \[46]  = \59 ,
  \[47]  = \60 ,
  \[48]  = \61 ,
  \[49]  = \62 ,
  \[50]  = \63 ,
  \[51]  = \64 ,
  \286  = (\350  & \349 ) | ((\350  & \348 ) | (\349  & \348 )),
  \287  = (~\329  & (~\328  & \327 )) | ((~\329  & (\328  & ~\327 )) | ((\329  & (~\328  & ~\327 )) | (\329  & (\328  & \327 )))),
  \288  = (~\332  & (~\331  & \330 )) | ((~\332  & (\331  & ~\330 )) | ((\332  & (~\331  & ~\330 )) | (\332  & (\331  & \330 )))),
  \289  = (~\335  & (~\334  & \333 )) | ((~\335  & (\334  & ~\333 )) | ((\335  & (~\334  & ~\333 )) | (\335  & (\334  & \333 )))),
  \[52]  = \65 ,
  \290  = (~\338  & (~\337  & \336 )) | ((~\338  & (\337  & ~\336 )) | ((\338  & (~\337  & ~\336 )) | (\338  & (\337  & \336 )))),
  \291  = (~\341  & (~\340  & \339 )) | ((~\341  & (\340  & ~\339 )) | ((\341  & (~\340  & ~\339 )) | (\341  & (\340  & \339 )))),
  \292  = (~\344  & (~\343  & \342 )) | ((~\344  & (\343  & ~\342 )) | ((\344  & (~\343  & ~\342 )) | (\344  & (\343  & \342 )))),
  \293  = (~\347  & (~\346  & \345 )) | ((~\347  & (\346  & ~\345 )) | ((\347  & (~\346  & ~\345 )) | (\347  & (\346  & \345 )))),
  \294  = (~\350  & (~\349  & \348 )) | ((~\350  & (\349  & ~\348 )) | ((\350  & (~\349  & ~\348 )) | (\350  & (\349  & \348 )))),
  \[53]  = \66 ,
  \[54]  = \546 ,
  \[55]  = \554 ,
  \[56]  = \562 ,
  \[57]  = \570 ,
  \[58]  = \578 ,
  \[59]  = \586 ,
  \322  = \759  & \757 ,
  \323  = \730  & \728 ,
  \325  = \701  & \699 ,
  \326  = \696  & \694 ,
  \327  = \326  & \325 ,
  \328  = \691  & \689 ,
  \329  = \686  & \684 ,
  \330  = (\329  & \328 ) | ((\329  & \327 ) | (\328  & \327 )),
  \331  = \681  & \679 ,
  \332  = \676  & \674 ,
  \333  = (\332  & \331 ) | ((\332  & \330 ) | (\331  & \330 )),
  \334  = \671  & \669 ,
  \335  = \666  & \664 ,
  \336  = (\335  & \334 ) | ((\335  & \333 ) | (\334  & \333 )),
  \337  = \661  & \659 ,
  \338  = \656  & \654 ,
  \339  = (\338  & \337 ) | ((\338  & \336 ) | (\337  & \336 )),
  \340  = \651  & \649 ,
  \341  = \646  & \644 ,
  \342  = (\341  & \340 ) | ((\341  & \339 ) | (\340  & \339 )),
  \343  = \641  & \639 ,
  \344  = \636  & \634 ,
  \345  = (\344  & \343 ) | ((\344  & \342 ) | (\343  & \342 )),
  \346  = \631  & \629 ,
  \347  = \626  & \624 ,
  \348  = (\347  & \346 ) | ((\347  & \345 ) | (\346  & \345 )),
  \349  = \621  & \619 ,
  \350  = \616  & \614 ,
  \351  = \287  & ~\3 ,
  \352  = \4  & \3 ,
  \353  = \352  | \351 ,
  \354  = \353  & \2 ,
  \355  = \13  & ~\2 ,
  \356  = \355  | \354 ,
  \357  = \356  & ~\1 ,
  \359  = \288  & ~\3 ,
  \360  = \5  & \3 ,
  \361  = \360  | \359 ,
  \362  = \361  & \2 ,
  \363  = \14  & ~\2 ,
  \364  = \363  | \362 ,
  \365  = \364  & ~\1 ,
  \367  = \289  & ~\3 ,
  \368  = \6  & \3 ,
  \369  = \368  | \367 ;
always begin
  \13  = \[36] ;
  \14  = \[37] ;
  \15  = \[38] ;
  \16  = \[39] ;
  \17  = \[40] ;
  \18  = \[41] ;
  \19  = \[42] ;
  \20  = \[43] ;
  \21  = \[44] ;
  \22  = \[45] ;
  \23  = \[46] ;
  \24  = \[47] ;
  \25  = \[48] ;
  \26  = \[49] ;
  \27  = \[50] ;
  \28  = \[51] ;
  \29  = \[52] ;
  \30  = \[53] ;
  \31  = \[54] ;
  \32  = \[55] ;
  \33  = \[56] ;
  \34  = \[57] ;
  \35  = \[58] ;
  \36  = \[59] ;
  \37  = \[60] ;
  \38  = \[61] ;
  \39  = \[62] ;
end
initial begin
  \22  = 1;
  \23  = 1;
  \24  = 1;
  \25  = 1;
  \26  = 1;
  \27  = 1;
  \28  = 1;
  \29  = 1;
  \30  = 1;
  \31  = 0;
  \32  = 0;
  \33  = 0;
  \34  = 0;
  \35  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
end
endmodule

