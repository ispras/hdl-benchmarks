//NOTE: no-implementation module stub

module EREG15LC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire WSCR_we,
    input wire [14:0] DMD,
    output reg [14:0] WSCR,
    input wire RST
);

endmodule
