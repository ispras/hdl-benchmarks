// IWLS benchmark module "frg1" printed on Wed May 29 16:34:07 2002
module frg1(a, b, c, e, f, g, h, i, j, k, l, m, n, o, p, q, r, s, t, u, v, w, \x , y, z, a0, b0, c0, d0, e0, f0);
input
  a,
  b,
  c,
  e,
  f,
  g,
  h,
  i,
  j,
  k,
  l,
  m,
  n,
  o,
  p,
  q,
  r,
  s,
  t,
  u,
  v,
  w,
  \x ,
  y,
  z,
  a0,
  b0,
  c0;
output
  d0,
  e0,
  f0;
wire
  \[25] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[30] ,
  \[4] ,
  \[31] ,
  \[6] ,
  \[8] ,
  \[10] ,
  \[9] ,
  \[12] ;
assign
  \[25]  = (\[4]  & ~w) | \[8] ,
  \[27]  = (\[4]  & ~z) | \[12] ,
  \[28]  = (~\x  & (~w & ~o)) | ((~\x  & ~h) | ((~o & ~m) | (~m & ~h))),
  \[29]  = (\[25]  & (~y & ~o)) | ((\[4]  & (~o & ~m)) | ((\[8]  & ~y) | (\[8]  & ~m))),
  \[0]  = (\[30]  & (\[9]  & (\[4]  & (~v & (~r & (~p & ~h)))))) | ((\[10]  & (\[6]  & (\[4]  & (~r & (~q & (~p & ~o)))))) | ((\[8]  & (~z & (~y & (~v & (~u & (~r & ~q)))))) | ((\[9]  & (\[4]  & (~r & (~p & (~k & ~h))))) | ((\[8]  & (~z & (~y & (~r & (~q & ~k))))) | ((\[8]  & (~v & (~u & (~r & (~q & ~m))))) | ((\[30]  & (\[4]  & (~v & (~l & ~h)))) | ((\[8]  & (~z & (~v & (~r & ~h)))) | ((\[8]  & (~z & (~r & (~k & ~h)))) | ((\[8]  & (~v & (~r & (~m & ~h)))) | ((\[8]  & (~r & (~q & (~m & ~k)))) | ((\[8]  & (~r & (~m & (~k & ~h)))) | ((\[30]  & (\[28]  & (\[12]  & ~p))) | ((\[29]  & (~u & (~q & ~g))) | ((\[29]  & (~q & (~k & ~g))) | ((\[28]  & (\[12]  & (~p & ~k))) | ((\[27]  & (~\x  & (~n & ~h))) | ((\[25]  & (~y & (~n & ~g))) | ((\[12]  & (~\x  & (~w & ~n))) | ((\[12]  & (~w & (~o & ~g))) | ((\[12]  & (~w & (~n & ~g))) | ((\[12]  & (~o & (~m & ~g))) | ((\[8]  & (~z & (~y & ~n))) | ((\[8]  & (~z & (~n & ~h))) | ((\[8]  & (~v & (~u & ~l))) | ((\[8]  & (~v & (~l & ~h))) | ((\[4]  & (~u & (~l & ~g))) | ((\[30]  & (\[12]  & ~l)) | ((\[12]  & (~l & ~g)) | ((\[10]  & (\[4]  & ~n)) | ((\[6]  & (\[4]  & ~l)) | ((\[4]  & (~n & ~l)) | ((\[4]  & (~h & ~g)) | ((~\[3]  & (~c0 & ~c)) | ((\[8]  & ~i) | (c & ~b))))))))))))))))))))))))))))))))))),
  \[1]  = (~a0 & f) | ((f & e) | \[31] ),
  \[2]  = (\[31]  & ~e) | (~b0 & ~e),
  \[3]  = e | a,
  d0 = \[0] ,
  \[30]  = ~t & ~s,
  \[4]  = \[3]  & ~c,
  e0 = \[1] ,
  \[31]  = c | a,
  f0 = \[2] ,
  \[6]  = (\[30]  & (~v & ~u)) | ~k,
  \[8]  = \[4]  & ~j,
  \[10]  = (\[9]  & (~y & ~w)) | ~m,
  \[9]  = (~z & ~\x ) | ~m,
  \[12]  = \[4]  & ~i;
endmodule

