module carry_sum (sin, cin, sout, cout);
  input sin;
  input cin;
  output sout;
  output cout;
endmodule
