// IWLS benchmark module "bigkey" printed on Wed May 29 21:51:26 2002
module bigkey(\key<255> , \key<254> , \key<253> , \key<252> , \key<251> , \key<250> , \key<249> , \key<248> , \key<247> , \key<246> , \key<245> , \key<244> , \key<243> , \key<242> , \key<241> , \key<240> , \key<239> , \key<238> , \key<237> , \key<236> , \key<235> , \key<234> , \key<233> , \key<232> , \key<231> , \key<230> , \key<229> , \key<228> , \key<227> , \key<226> , \key<225> , \key<224> , \key<223> , \key<222> , \key<221> , \key<220> , \key<219> , \key<218> , \key<217> , \key<216> , \key<215> , \key<214> , \key<213> , \key<212> , \key<211> , \key<210> , \key<209> , \key<208> , \key<207> , \key<206> , \key<205> , \key<204> , \key<203> , \key<202> , \key<201> , \key<200> , \key<199> , \key<198> , \key<197> , \key<196> , \key<195> , \key<194> , \key<193> , \key<192> , \key<191> , \key<190> , \key<189> , \key<188> , \key<187> , \key<186> , \key<185> , \key<184> , \key<183> , \key<182> , \key<181> , \key<180> , \key<179> , \key<178> , \key<177> , \key<176> , \key<175> , \key<174> , \key<173> , \key<172> , \key<171> , \key<170> , \key<169> , \key<168> , \key<167> , \key<166> , \key<165> , \key<164> , \key<163> , \key<162> , \key<161> , \key<160> , \key<159> , \key<158> , \key<157> , \key<156> , \key<155> , \key<154> , \key<153> , \key<152> , \key<151> , \key<150> , \key<149> , \key<148> , \key<147> , \key<146> , \key<145> , \key<144> , \key<143> , \key<142> , \key<141> , \key<140> , \key<139> , \key<138> , \key<137> , \key<136> , \key<135> , \key<134> , \key<133> , \key<132> , \key<131> , \key<130> , \key<129> , \key<128> , \key<127> , \key<126> , \key<125> , \key<124> , \key<123> , \key<122> , \key<121> , \key<120> , \key<119> , \key<118> , \key<117> , \key<116> , \key<115> , \key<114> , \key<113> , \key<112> , \key<111> , \key<110> , \key<109> , \key<108> , \key<107> , \key<106> , \key<105> , \key<104> , \key<103> , \key<102> , \key<101> , \key<100> , \key<99> , \key<98> , \key<97> , \key<96> , \key<95> , \key<94> , \key<93> , \key<92> , \key<91> , \key<90> , \key<89> , \key<88> , \key<87> , \key<86> , \key<85> , \key<84> , \key<83> , \key<82> , \key<81> , \key<80> , \key<79> , \key<78> , \key<77> , \key<76> , \key<75> , \key<74> , \key<73> , \key<72> , \key<71> , \key<70> , \key<69> , \key<68> , \key<67> , \key<66> , \key<65> , \key<64> , \key<63> , \key<62> , \key<61> , \key<60> , \key<59> , \key<58> , \key<57> , \key<56> , \key<55> , \key<54> , \key<53> , \key<52> , \key<51> , \key<50> , \key<49> , \key<48> , \key<47> , \key<46> , \key<45> , \key<44> , \key<43> , \key<42> , \key<41> , \key<40> , \key<39> , \key<38> , \key<37> , \key<36> , \key<35> , \key<34> , \key<33> , \key<32> , \key<31> , \key<30> , \key<29> , \key<28> , \key<27> , \key<26> , \key<25> , \key<24> , \key<23> , \key<22> , \key<21> , \key<20> , \key<19> , \key<18> , \key<17> , \key<16> , \key<15> , \key<14> , \key<13> , \key<12> , \key<11> , \key<10> , \key<9> , \key<8> , \key<7> , \key<6> , \key<5> , \key<4> , \key<3> , \key<2> , \key<1> , \key<0> , \encrypt<0> , \start<0> , \count<3> , \count<2> , \count<1> , \count<0> , \new_count<3> , \new_count<2> , \new_count<1> , \new_count<0> , \data_ready<0> , \KSi<191> , \KSi<190> , \KSi<189> , \KSi<188> , \KSi<187> , \KSi<186> , \KSi<185> , \KSi<184> , \KSi<183> , \KSi<182> , \KSi<181> , \KSi<180> , \KSi<179> , \KSi<178> , \KSi<177> , \KSi<176> , \KSi<175> , \KSi<174> , \KSi<173> , \KSi<172> , \KSi<171> , \KSi<170> , \KSi<169> , \KSi<168> , \KSi<167> , \KSi<166> , \KSi<165> , \KSi<164> , \KSi<163> , \KSi<162> , \KSi<161> , \KSi<160> , \KSi<159> , \KSi<158> , \KSi<157> , \KSi<156> , \KSi<155> , \KSi<154> , \KSi<153> , \KSi<152> , \KSi<151> , \KSi<150> , \KSi<149> , \KSi<148> , \KSi<147> , \KSi<146> , \KSi<145> , \KSi<144> , \KSi<143> , \KSi<142> , \KSi<141> , \KSi<140> , \KSi<139> , \KSi<138> , \KSi<137> , \KSi<136> , \KSi<135> , \KSi<134> , \KSi<133> , \KSi<132> , \KSi<131> , \KSi<130> , \KSi<129> , \KSi<128> , \KSi<127> , \KSi<126> , \KSi<125> , \KSi<124> , \KSi<123> , \KSi<122> , \KSi<121> , \KSi<120> , \KSi<119> , \KSi<118> , \KSi<117> , \KSi<116> , \KSi<115> , \KSi<114> , \KSi<113> , \KSi<112> , \KSi<111> , \KSi<110> , \KSi<109> , \KSi<108> , \KSi<107> , \KSi<106> , \KSi<105> , \KSi<104> , \KSi<103> , \KSi<102> , \KSi<101> , \KSi<100> , \KSi<99> , \KSi<98> , \KSi<97> , \KSi<96> , \KSi<95> , \KSi<94> , \KSi<93> , \KSi<92> , \KSi<91> , \KSi<90> , \KSi<89> , \KSi<88> , \KSi<87> , \KSi<86> , \KSi<85> , \KSi<84> , \KSi<83> , \KSi<82> , \KSi<81> , \KSi<80> , \KSi<79> , \KSi<78> , \KSi<77> , \KSi<76> , \KSi<75> , \KSi<74> , \KSi<73> , \KSi<72> , \KSi<71> , \KSi<70> , \KSi<69> , \KSi<68> , \KSi<67> , \KSi<66> , \KSi<65> , \KSi<64> , \KSi<63> , \KSi<62> , \KSi<61> , \KSi<60> , \KSi<59> , \KSi<58> , \KSi<57> , \KSi<56> , \KSi<55> , \KSi<54> , \KSi<53> , \KSi<52> , \KSi<51> , \KSi<50> , \KSi<49> , \KSi<48> , \KSi<47> , \KSi<46> , \KSi<45> , \KSi<44> , \KSi<43> , \KSi<42> , \KSi<41> , \KSi<40> , \KSi<39> , \KSi<38> , \KSi<37> , \KSi<36> , \KSi<35> , \KSi<34> , \KSi<33> , \KSi<32> , \KSi<31> , \KSi<30> , \KSi<29> , \KSi<28> , \KSi<27> , \KSi<26> , \KSi<25> , \KSi<24> , \KSi<23> , \KSi<22> , \KSi<21> , \KSi<20> , \KSi<19> , \KSi<18> , \KSi<17> , \KSi<16> , \KSi<15> , \KSi<14> , \KSi<13> , \KSi<12> , \KSi<11> , \KSi<10> , \KSi<9> , \KSi<8> , \KSi<7> , \KSi<6> , \KSi<5> , \KSi<4> , \KSi<3> , \KSi<2> , \KSi<1> , \KSi<0> );
input
  \key<156> ,
  \key<155> ,
  \key<158> ,
  \key<157> ,
  \key<159> ,
  \key<240> ,
  \key<14> ,
  \key<13> ,
  \key<242> ,
  \key<12> ,
  \key<241> ,
  \key<11> ,
  \key<244> ,
  \key<10> ,
  \key<243> ,
  \key<246> ,
  \key<245> ,
  \key<248> ,
  \key<247> ,
  \key<249> ,
  \key<19> ,
  \key<18> ,
  \key<17> ,
  \key<0> ,
  \key<16> ,
  \key<1> ,
  \key<15> ,
  \key<2> ,
  \key<230> ,
  \key<24> ,
  \key<3> ,
  \key<23> ,
  \key<4> ,
  \key<232> ,
  \key<22> ,
  \key<5> ,
  \key<231> ,
  \key<21> ,
  \key<6> ,
  \key<234> ,
  \key<20> ,
  \key<7> ,
  \key<233> ,
  \key<8> ,
  \key<236> ,
  \key<9> ,
  \key<235> ,
  \key<238> ,
  \key<237> ,
  \key<239> ,
  \key<29> ,
  \key<28> ,
  \key<27> ,
  \key<26> ,
  \key<25> ,
  \key<220> ,
  \key<34> ,
  \key<33> ,
  \key<222> ,
  \key<32> ,
  \key<221> ,
  \key<31> ,
  \key<224> ,
  \key<30> ,
  \key<223> ,
  \key<226> ,
  \key<225> ,
  \key<228> ,
  \key<227> ,
  \key<229> ,
  \key<39> ,
  \key<38> ,
  \key<37> ,
  \key<36> ,
  \key<35> ,
  \key<210> ,
  \key<44> ,
  \key<43> ,
  \key<212> ,
  \key<42> ,
  \key<211> ,
  \key<41> ,
  \key<214> ,
  \key<40> ,
  \key<213> ,
  \key<216> ,
  \key<215> ,
  \key<218> ,
  \key<217> ,
  \key<219> ,
  \key<49> ,
  \key<48> ,
  \key<47> ,
  \key<46> ,
  \key<45> ,
  \key<200> ,
  \key<54> ,
  \key<53> ,
  \key<202> ,
  \key<52> ,
  \key<201> ,
  \key<51> ,
  \key<204> ,
  \key<50> ,
  \key<203> ,
  \key<206> ,
  \key<205> ,
  \key<208> ,
  \key<207> ,
  \key<209> ,
  \key<59> ,
  \key<58> ,
  \key<57> ,
  \key<56> ,
  \key<55> ,
  \key<64> ,
  \key<63> ,
  \key<62> ,
  \key<61> ,
  \key<60> ,
  \key<69> ,
  \key<68> ,
  \key<67> ,
  \key<66> ,
  \key<65> ,
  \key<74> ,
  \key<73> ,
  \key<72> ,
  \key<71> ,
  \key<70> ,
  \key<79> ,
  \key<78> ,
  \key<77> ,
  \key<76> ,
  \key<75> ,
  \key<84> ,
  \key<83> ,
  \key<82> ,
  \key<81> ,
  \key<80> ,
  \key<89> ,
  \key<88> ,
  \key<87> ,
  \key<86> ,
  \key<85> ,
  \key<94> ,
  \key<93> ,
  \key<92> ,
  \key<91> ,
  \key<90> ,
  \key<99> ,
  \key<98> ,
  \key<97> ,
  \key<96> ,
  \key<95> ,
  \start<0> ,
  \key<140> ,
  \key<250> ,
  \key<142> ,
  \key<252> ,
  \key<141> ,
  \key<251> ,
  \key<144> ,
  \key<254> ,
  \key<143> ,
  \key<253> ,
  \key<146> ,
  \key<145> ,
  \key<255> ,
  \key<148> ,
  \key<147> ,
  \key<149> ,
  \key<130> ,
  \key<132> ,
  \key<131> ,
  \key<134> ,
  \key<133> ,
  \key<136> ,
  \key<135> ,
  \key<138> ,
  \key<137> ,
  \key<139> ,
  \count<0> ,
  \count<3> ,
  \key<120> ,
  \count<1> ,
  \key<122> ,
  \count<2> ,
  \key<121> ,
  \key<124> ,
  \key<123> ,
  \key<126> ,
  \key<125> ,
  \key<128> ,
  \key<127> ,
  \key<129> ,
  \key<110> ,
  \key<112> ,
  \key<111> ,
  \key<114> ,
  \key<113> ,
  \key<116> ,
  \key<115> ,
  \key<118> ,
  \key<117> ,
  \key<119> ,
  \key<100> ,
  \key<102> ,
  \key<101> ,
  \key<104> ,
  \key<103> ,
  \key<106> ,
  \key<105> ,
  \key<108> ,
  \key<107> ,
  \key<109> ,
  \key<190> ,
  \key<192> ,
  \key<191> ,
  \key<194> ,
  \key<193> ,
  \key<196> ,
  \key<195> ,
  \key<198> ,
  \key<197> ,
  \key<199> ,
  \key<180> ,
  \key<182> ,
  \key<181> ,
  \key<184> ,
  \key<183> ,
  \key<186> ,
  \key<185> ,
  \key<188> ,
  \key<187> ,
  \key<189> ,
  \key<170> ,
  \key<172> ,
  \key<171> ,
  \key<174> ,
  \key<173> ,
  \key<176> ,
  \key<175> ,
  \key<178> ,
  \key<177> ,
  \key<179> ,
  \encrypt<0> ,
  \key<160> ,
  \key<162> ,
  \key<161> ,
  \key<164> ,
  \key<163> ,
  \key<166> ,
  \key<165> ,
  \key<168> ,
  \key<167> ,
  \key<169> ,
  \key<150> ,
  \key<152> ,
  \key<151> ,
  \key<154> ,
  \key<153> ;
output
  \KSi<130> ,
  \KSi<131> ,
  \KSi<132> ,
  \KSi<133> ,
  \KSi<134> ,
  \KSi<135> ,
  \KSi<136> ,
  \KSi<137> ,
  \KSi<138> ,
  \KSi<139> ,
  \KSi<100> ,
  \KSi<101> ,
  \KSi<102> ,
  \KSi<103> ,
  \KSi<104> ,
  \KSi<105> ,
  \KSi<106> ,
  \KSi<107> ,
  \KSi<108> ,
  \KSi<109> ,
  \KSi<190> ,
  \KSi<191> ,
  \KSi<160> ,
  \KSi<161> ,
  \KSi<162> ,
  \KSi<163> ,
  \KSi<164> ,
  \KSi<165> ,
  \KSi<166> ,
  \KSi<167> ,
  \KSi<168> ,
  \KSi<169> ,
  \KSi<150> ,
  \KSi<151> ,
  \KSi<152> ,
  \KSi<153> ,
  \KSi<154> ,
  \KSi<155> ,
  \KSi<156> ,
  \KSi<157> ,
  \KSi<158> ,
  \KSi<159> ,
  \KSi<0> ,
  \KSi<1> ,
  \KSi<2> ,
  \KSi<3> ,
  \KSi<4> ,
  \KSi<180> ,
  \KSi<5> ,
  \KSi<181> ,
  \KSi<6> ,
  \KSi<182> ,
  \KSi<7> ,
  \KSi<183> ,
  \KSi<8> ,
  \KSi<184> ,
  \KSi<9> ,
  \KSi<185> ,
  \KSi<186> ,
  \KSi<187> ,
  \KSi<188> ,
  \KSi<189> ,
  \KSi<170> ,
  \KSi<171> ,
  \KSi<172> ,
  \KSi<173> ,
  \KSi<174> ,
  \KSi<175> ,
  \KSi<176> ,
  \KSi<177> ,
  \KSi<178> ,
  \KSi<179> ,
  \new_count<0> ,
  \new_count<3> ,
  \new_count<1> ,
  \new_count<2> ,
  \KSi<12> ,
  \KSi<11> ,
  \KSi<14> ,
  \KSi<13> ,
  \KSi<10> ,
  \KSi<19> ,
  \KSi<16> ,
  \KSi<15> ,
  \KSi<18> ,
  \KSi<17> ,
  \KSi<22> ,
  \KSi<21> ,
  \KSi<24> ,
  \KSi<23> ,
  \KSi<20> ,
  \KSi<29> ,
  \KSi<26> ,
  \KSi<25> ,
  \KSi<28> ,
  \KSi<27> ,
  \KSi<32> ,
  \KSi<31> ,
  \KSi<34> ,
  \KSi<33> ,
  \KSi<30> ,
  \KSi<39> ,
  \KSi<36> ,
  \KSi<35> ,
  \KSi<38> ,
  \KSi<37> ,
  \KSi<42> ,
  \KSi<41> ,
  \KSi<44> ,
  \KSi<43> ,
  \KSi<40> ,
  \KSi<49> ,
  \KSi<46> ,
  \KSi<45> ,
  \KSi<48> ,
  \KSi<47> ,
  \KSi<52> ,
  \KSi<51> ,
  \KSi<54> ,
  \KSi<53> ,
  \KSi<50> ,
  \KSi<59> ,
  \KSi<56> ,
  \KSi<55> ,
  \KSi<58> ,
  \KSi<57> ,
  \KSi<62> ,
  \KSi<61> ,
  \KSi<64> ,
  \KSi<63> ,
  \KSi<60> ,
  \KSi<69> ,
  \KSi<66> ,
  \data_ready<0> ,
  \KSi<65> ,
  \KSi<68> ,
  \KSi<67> ,
  \KSi<72> ,
  \KSi<71> ,
  \KSi<74> ,
  \KSi<73> ,
  \KSi<70> ,
  \KSi<79> ,
  \KSi<76> ,
  \KSi<75> ,
  \KSi<78> ,
  \KSi<77> ,
  \KSi<82> ,
  \KSi<81> ,
  \KSi<84> ,
  \KSi<83> ,
  \KSi<80> ,
  \KSi<89> ,
  \KSi<86> ,
  \KSi<85> ,
  \KSi<88> ,
  \KSi<87> ,
  \KSi<92> ,
  \KSi<91> ,
  \KSi<94> ,
  \KSi<93> ,
  \KSi<90> ,
  \KSi<99> ,
  \KSi<96> ,
  \KSi<95> ,
  \KSi<98> ,
  \KSi<97> ,
  \KSi<120> ,
  \KSi<121> ,
  \KSi<122> ,
  \KSi<123> ,
  \KSi<124> ,
  \KSi<125> ,
  \KSi<126> ,
  \KSi<127> ,
  \KSi<128> ,
  \KSi<129> ,
  \KSi<110> ,
  \KSi<111> ,
  \KSi<112> ,
  \KSi<113> ,
  \KSi<114> ,
  \KSi<115> ,
  \KSi<116> ,
  \KSi<117> ,
  \KSi<118> ,
  \KSi<119> ,
  \KSi<140> ,
  \KSi<141> ,
  \KSi<142> ,
  \KSi<143> ,
  \KSi<144> ,
  \KSi<145> ,
  \KSi<146> ,
  \KSi<147> ,
  \KSi<148> ,
  \KSi<149> ;
reg
  \D<0> ,
  \D<1> ,
  \D<2> ,
  \D<3> ,
  \D<4> ,
  \D<5> ,
  \D<6> ,
  \C<10> ,
  \D<7> ,
  \C<11> ,
  \D<8> ,
  \C<12> ,
  \D<9> ,
  \C<13> ,
  \C<14> ,
  \C<15> ,
  \C<16> ,
  \C<17> ,
  \C<18> ,
  \C<19> ,
  \C<20> ,
  \C<21> ,
  \C<22> ,
  \C<23> ,
  \C<24> ,
  \C<25> ,
  \C<26> ,
  \C<27> ,
  \C<28> ,
  \C<29> ,
  \C<30> ,
  \C<31> ,
  \C<32> ,
  \C<33> ,
  \C<34> ,
  \C<35> ,
  \C<36> ,
  \C<37> ,
  \C<38> ,
  \C<39> ,
  \C<40> ,
  \C<41> ,
  \C<42> ,
  \C<43> ,
  \C<44> ,
  \C<45> ,
  \C<46> ,
  \C<47> ,
  \C<48> ,
  \C<49> ,
  \C<50> ,
  \C<51> ,
  \C<52> ,
  \C<53> ,
  \C<54> ,
  \C<55> ,
  \C<56> ,
  \C<57> ,
  \C<58> ,
  \C<59> ,
  \C<60> ,
  \C<61> ,
  \C<62> ,
  \C<63> ,
  \C<64> ,
  \C<65> ,
  \C<66> ,
  \C<67> ,
  \C<68> ,
  \C<69> ,
  \C<70> ,
  \C<71> ,
  \C<72> ,
  \C<73> ,
  \C<74> ,
  \C<75> ,
  \C<76> ,
  \C<77> ,
  \C<78> ,
  \C<79> ,
  \C<80> ,
  \C<81> ,
  \C<82> ,
  \C<83> ,
  \C<84> ,
  \C<85> ,
  \C<86> ,
  \C<87> ,
  \C<88> ,
  \C<89> ,
  \C<90> ,
  \C<91> ,
  \D<10> ,
  \C<92> ,
  \D<11> ,
  \C<93> ,
  \D<12> ,
  \C<94> ,
  \D<13> ,
  \C<95> ,
  \D<14> ,
  \C<96> ,
  \D<15> ,
  \C<97> ,
  \D<16> ,
  \C<98> ,
  \D<17> ,
  \C<99> ,
  \D<18> ,
  \D<19> ,
  \D<20> ,
  \D<21> ,
  \D<22> ,
  \D<23> ,
  \D<24> ,
  \D<25> ,
  \D<26> ,
  \D<27> ,
  \D<28> ,
  \D<29> ,
  \D<30> ,
  \D<31> ,
  \D<32> ,
  \D<33> ,
  \D<34> ,
  \D<35> ,
  \D<36> ,
  \D<37> ,
  \D<38> ,
  \D<39> ,
  \D<40> ,
  \D<41> ,
  \D<42> ,
  \D<43> ,
  \D<44> ,
  \D<45> ,
  \D<46> ,
  \D<47> ,
  \D<48> ,
  \D<49> ,
  \D<50> ,
  \D<51> ,
  \D<52> ,
  \D<53> ,
  \D<54> ,
  \D<55> ,
  \D<56> ,
  \D<57> ,
  \D<58> ,
  \D<59> ,
  \D<60> ,
  \D<61> ,
  \D<62> ,
  \D<63> ,
  \D<64> ,
  \D<65> ,
  \D<66> ,
  \D<67> ,
  \D<68> ,
  \D<69> ,
  \C<100> ,
  \D<70> ,
  \C<101> ,
  \D<71> ,
  \C<102> ,
  \D<72> ,
  \C<103> ,
  \D<73> ,
  \C<104> ,
  \D<74> ,
  \C<105> ,
  \D<75> ,
  \C<106> ,
  \D<76> ,
  \C<107> ,
  \D<77> ,
  \C<108> ,
  \C<0> ,
  \D<78> ,
  \C<109> ,
  \C<1> ,
  \D<79> ,
  \C<2> ,
  \C<3> ,
  \C<4> ,
  \C<5> ,
  \C<6> ,
  \C<7> ,
  \C<110> ,
  \C<8> ,
  \D<80> ,
  \C<111> ,
  \C<9> ,
  \D<81> ,
  \D<82> ,
  \D<83> ,
  \D<84> ,
  \D<85> ,
  \D<86> ,
  \D<87> ,
  \D<88> ,
  \D<89> ,
  \D<90> ,
  \D<91> ,
  \D<92> ,
  \D<93> ,
  \D<94> ,
  \D<95> ,
  \D<96> ,
  \D<97> ,
  \D<98> ,
  \D<99> ,
  \D<100> ,
  \D<101> ,
  \D<102> ,
  \D<103> ,
  \D<104> ,
  \D<105> ,
  \D<106> ,
  \D<107> ,
  \D<108> ,
  \D<109> ,
  \D<110> ,
  \D<111> ;
wire
  \[568] ,
  \[758] ,
  \new_D<98> ,
  \[569] ,
  \[759] ,
  \new_D<91> ,
  \new_D<92> ,
  \new_D<93> ,
  \new_D<94> ,
  \[570] ,
  \[760] ,
  \new_D<90> ,
  \[571] ,
  \[761] ,
  \[572] ,
  \[762] ,
  \[573] ,
  \[763] ,
  \[574] ,
  \[764] ,
  \[575] ,
  \[765] ,
  \[576] ,
  \[766] ,
  \[577] ,
  \[767] ,
  \[578] ,
  \[768] ,
  \new_C<111> ,
  \[579] ,
  \[769] ,
  \new_C<110> ,
  \[580] ,
  \[770] ,
  \[581] ,
  \[771] ,
  \[582] ,
  \[772] ,
  \[583] ,
  \[773] ,
  \[584] ,
  \[774] ,
  \[585] ,
  \[775] ,
  \[586] ,
  \[776] ,
  \[587] ,
  \[777] ,
  \[588] ,
  \[778] ,
  \[589] ,
  \[779] ,
  \[590] ,
  \[780] ,
  \[591] ,
  \[781] ,
  \[592] ,
  \[782] ,
  \[593] ,
  \[783] ,
  \[594] ,
  \[784] ,
  \[595] ,
  \[785] ,
  \[596] ,
  \[786] ,
  \[597] ,
  \[787] ,
  \[598] ,
  \[788] ,
  \[599] ,
  \[789] ,
  \[790] ,
  \[791] ,
  \new_D<59> ,
  \[792] ,
  \[793] ,
  \[794] ,
  \[795] ,
  \new_D<55> ,
  \[796] ,
  \new_D<56> ,
  \[797] ,
  \new_D<57> ,
  \[798] ,
  \new_D<58> ,
  \[799] ,
  \new_D<51> ,
  \new_D<52> ,
  \new_D<53> ,
  \new_D<54> ,
  \new_D<50> ,
  \new_D<69> ,
  \new_D<65> ,
  \new_D<66> ,
  \new_D<67> ,
  \new_D<68> ,
  \new_D<61> ,
  \new_D<62> ,
  \new_D<63> ,
  \new_D<64> ,
  \new_D<60> ,
  \new_D<79> ,
  \new_D<75> ,
  \new_D<76> ,
  \new_D<77> ,
  \new_D<78> ,
  \new_D<71> ,
  \new_D<72> ,
  \new_D<73> ,
  \new_D<74> ,
  \new_D<70> ,
  \new_D<111> ,
  \new_D<89> ,
  \new_D<85> ,
  \new_D<110> ,
  \new_D<86> ,
  \new_D<87> ,
  \new_D<88> ,
  \new_D<81> ,
  \new_D<82> ,
  \new_D<83> ,
  \new_D<84> ,
  \new_C<109> ,
  \new_D<80> ,
  \new_C<106> ,
  \new_C<105> ,
  \new_C<108> ,
  \new_C<107> ,
  \new_C<102> ,
  \new_C<101> ,
  \new_C<104> ,
  \new_C<103> ,
  \new_C<100> ,
  \[600] ,
  \[601] ,
  \[602] ,
  \[603] ,
  \[224] ,
  \[604] ,
  \[225] ,
  \[605] ,
  \[226] ,
  \[606] ,
  \[227] ,
  \[607] ,
  \[228] ,
  \[608] ,
  \[609] ,
  \[610] ,
  \[800] ,
  \[421] ,
  \[611] ,
  \[801] ,
  \[422] ,
  \[612] ,
  \[802] ,
  \[423] ,
  \[613] ,
  \[803] ,
  \[424] ,
  \[614] ,
  \[804] ,
  \[425] ,
  \[615] ,
  \[805] ,
  \[426] ,
  \[616] ,
  \[806] ,
  \new_D<1> ,
  \[427] ,
  \[617] ,
  \[807] ,
  \new_D<2> ,
  \[428] ,
  \[618] ,
  \[808] ,
  \new_D<3> ,
  \[429] ,
  \[619] ,
  \[809] ,
  \new_D<4> ,
  \new_D<0> ,
  \new_D<9> ,
  \[430] ,
  \[620] ,
  \[810] ,
  \[431] ,
  \[621] ,
  \[811] ,
  \[432] ,
  \[622] ,
  \[812] ,
  \new_D<5> ,
  \[433] ,
  \[623] ,
  \[813] ,
  \new_D<6> ,
  \[434] ,
  \[624] ,
  \[814] ,
  \new_D<7> ,
  \[435] ,
  \[625] ,
  \[815] ,
  \new_D<8> ,
  \[436] ,
  \[626] ,
  \[816] ,
  \[437] ,
  \[627] ,
  \[817] ,
  \[438] ,
  \[628] ,
  \[818] ,
  \[439] ,
  \[629] ,
  \[819] ,
  \[440] ,
  \[630] ,
  \[820] ,
  \[441] ,
  \[631] ,
  \[821] ,
  \[442] ,
  \[632] ,
  \[822] ,
  \[443] ,
  \[633] ,
  \[823] ,
  \[444] ,
  \[634] ,
  \[824] ,
  \[445] ,
  \[635] ,
  \[825] ,
  \[446] ,
  \[636] ,
  \[826] ,
  \[447] ,
  \[637] ,
  \[827] ,
  \[448] ,
  \[638] ,
  \[828] ,
  \[449] ,
  \[639] ,
  \new_D<109> ,
  \[829] ,
  \new_D<106> ,
  \new_D<105> ,
  \new_D<108> ,
  \new_D<107> ,
  \[450] ,
  \[640] ,
  \new_D<102> ,
  \[830] ,
  \[451] ,
  \[641] ,
  \new_D<101> ,
  \[831] ,
  \[452] ,
  \[642] ,
  \new_D<104> ,
  \[832] ,
  \[453] ,
  \[643] ,
  \new_D<103> ,
  \[833] ,
  \[454] ,
  \[644] ,
  \[834] ,
  \[455] ,
  \[645] ,
  \[835] ,
  \[456] ,
  \[646] ,
  \new_D<100> ,
  \[836] ,
  \[457] ,
  \[647] ,
  \[837] ,
  \[458] ,
  \[648] ,
  \[838] ,
  \[459] ,
  \[649] ,
  \[839] ,
  \[460] ,
  \new_C<19> ,
  \[650] ,
  \[840] ,
  \[461] ,
  \[651] ,
  \[841] ,
  \[462] ,
  \[652] ,
  \[842] ,
  \[463] ,
  \[653] ,
  \[843] ,
  \[464] ,
  \new_C<15> ,
  \[654] ,
  \[844] ,
  \[465] ,
  \new_C<16> ,
  \[655] ,
  \[845] ,
  \[466] ,
  \new_C<17> ,
  \[656] ,
  \[846] ,
  \[467] ,
  \new_C<18> ,
  \[657] ,
  \[847] ,
  \[468] ,
  \new_C<11> ,
  \[658] ,
  \[848] ,
  \[469] ,
  \new_C<12> ,
  \[659] ,
  \[849] ,
  \new_C<13> ,
  \new_C<14> ,
  \$$COND0<0>5.1 ,
  \new_C<10> ,
  \[470] ,
  \new_C<29> ,
  \[660] ,
  \[850] ,
  \[471] ,
  \[661] ,
  \[851] ,
  \[472] ,
  \[662] ,
  \[852] ,
  \[473] ,
  \[663] ,
  \[853] ,
  \[474] ,
  \new_C<25> ,
  \[664] ,
  \[854] ,
  \[475] ,
  \new_C<26> ,
  \[665] ,
  \[855] ,
  \[476] ,
  \new_C<27> ,
  \[666] ,
  \[856] ,
  \[477] ,
  \new_C<28> ,
  \[667] ,
  \[857] ,
  \[478] ,
  \new_C<21> ,
  \[668] ,
  \[858] ,
  \[479] ,
  \new_C<22> ,
  \[669] ,
  \[859] ,
  \new_C<23> ,
  \new_C<24> ,
  \new_C<20> ,
  \[480] ,
  \new_C<39> ,
  \[670] ,
  \[860] ,
  \[481] ,
  \[671] ,
  \[861] ,
  \[482] ,
  \[672] ,
  \[862] ,
  \[483] ,
  \[673] ,
  \[863] ,
  \[484] ,
  \new_C<35> ,
  \[674] ,
  \[864] ,
  \[485] ,
  \new_C<36> ,
  \[675] ,
  \[865] ,
  \[486] ,
  \new_C<37> ,
  \[676] ,
  \[866] ,
  \[487] ,
  \new_C<38> ,
  \[677] ,
  \[867] ,
  \[488] ,
  \new_C<31> ,
  \[678] ,
  \[868] ,
  \[489] ,
  \new_C<32> ,
  \[679] ,
  \[869] ,
  \new_C<33> ,
  \new_C<34> ,
  \new_C<30> ,
  \[490] ,
  \new_C<49> ,
  \[680] ,
  \[870] ,
  \[491] ,
  \[681] ,
  \[871] ,
  \[492] ,
  \[682] ,
  \[872] ,
  \[493] ,
  \[683] ,
  \[873] ,
  \[494] ,
  \new_C<45> ,
  \[684] ,
  \[874] ,
  \[495] ,
  \new_C<46> ,
  \[685] ,
  \[875] ,
  \[496] ,
  \new_C<47> ,
  \[686] ,
  \[876] ,
  \[497] ,
  \new_C<48> ,
  \[687] ,
  \[877] ,
  \[498] ,
  \new_C<41> ,
  \[688] ,
  \[878] ,
  \[499] ,
  \new_C<42> ,
  \[689] ,
  \[879] ,
  \new_C<43> ,
  \new_C<44> ,
  \new_C<40> ,
  \[690] ,
  \[880] ,
  \[691] ,
  \[692] ,
  \[882] ,
  \[693] ,
  \[694] ,
  \[695] ,
  \[696] ,
  \[697] ,
  \[698] ,
  \[699] ,
  \new_C<99> ,
  \new_D<19> ,
  \new_C<95> ,
  \new_C<96> ,
  \new_D<15> ,
  \new_C<97> ,
  \new_D<16> ,
  \new_C<98> ,
  \new_D<17> ,
  \new_C<91> ,
  \new_D<18> ,
  \new_C<92> ,
  \new_D<11> ,
  \new_C<93> ,
  \new_D<12> ,
  \new_C<94> ,
  \new_D<13> ,
  \new_D<14> ,
  \new_C<90> ,
  \new_D<10> ,
  \new_D<29> ,
  \new_D<25> ,
  \new_D<26> ,
  \new_D<27> ,
  \new_D<28> ,
  \new_D<21> ,
  \new_D<22> ,
  \new_D<23> ,
  \new_D<24> ,
  \[500] ,
  \new_D<20> ,
  \[501] ,
  \new_D<39> ,
  \[502] ,
  \[503] ,
  \[504] ,
  \[505] ,
  \new_D<35> ,
  \[506] ,
  \new_D<36> ,
  \[507] ,
  \new_D<37> ,
  \[508] ,
  \new_D<38> ,
  \[509] ,
  \new_D<31> ,
  \new_D<32> ,
  \new_D<33> ,
  \new_D<34> ,
  \[510] ,
  \[700] ,
  \new_D<30> ,
  \[511] ,
  \[701] ,
  \new_D<49> ,
  \[512] ,
  \[702] ,
  \[513] ,
  \[703] ,
  \[514] ,
  \[704] ,
  \[515] ,
  \[705] ,
  \new_D<45> ,
  \[516] ,
  \[706] ,
  \new_C<1> ,
  \new_D<46> ,
  \[517] ,
  \[707] ,
  \new_C<2> ,
  \new_D<47> ,
  \[518] ,
  \[708] ,
  \new_C<3> ,
  \new_D<48> ,
  \[519] ,
  \[709] ,
  \new_C<4> ,
  \new_D<41> ,
  \new_D<42> ,
  \new_D<43> ,
  \new_D<44> ,
  \new_C<0> ,
  \new_C<9> ,
  \[520] ,
  \new_C<59> ,
  \[710] ,
  \new_D<40> ,
  \[521] ,
  \[711] ,
  \[522] ,
  \[712] ,
  \new_C<5> ,
  \[523] ,
  \[713] ,
  \new_C<6> ,
  \[524] ,
  \new_C<55> ,
  \[714] ,
  \new_C<7> ,
  \[525] ,
  \new_C<56> ,
  \[715] ,
  \new_C<8> ,
  \[526] ,
  \new_C<57> ,
  \[716] ,
  \[527] ,
  \new_C<58> ,
  \[717] ,
  \[528] ,
  \new_C<51> ,
  \[718] ,
  \[529] ,
  \new_C<52> ,
  \[719] ,
  \new_C<53> ,
  \new_C<54> ,
  \new_C<50> ,
  \[530] ,
  \new_C<69> ,
  \[720] ,
  \[531] ,
  \[721] ,
  \[532] ,
  \[722] ,
  \[533] ,
  \[723] ,
  \[534] ,
  \new_C<65> ,
  \[724] ,
  \[535] ,
  \new_C<66> ,
  \[725] ,
  \[536] ,
  \new_C<67> ,
  \[726] ,
  \[537] ,
  \new_C<68> ,
  \[727] ,
  \[538] ,
  \new_C<61> ,
  \[728] ,
  \[539] ,
  \new_C<62> ,
  \[729] ,
  \new_C<63> ,
  \new_C<64> ,
  \new_C<60> ,
  \[540] ,
  \new_C<79> ,
  \[730] ,
  \[541] ,
  \[731] ,
  \[542] ,
  \[732] ,
  \[543] ,
  \[733] ,
  \[544] ,
  \new_C<75> ,
  \[734] ,
  \[545] ,
  \new_C<76> ,
  \[735] ,
  \[546] ,
  \new_C<77> ,
  \[736] ,
  \[547] ,
  \new_C<78> ,
  \[737] ,
  \[548] ,
  \new_C<71> ,
  \[738] ,
  \[549] ,
  \new_C<72> ,
  \[739] ,
  \new_C<73> ,
  \new_C<74> ,
  \new_C<70> ,
  \[550] ,
  \new_C<89> ,
  \[740] ,
  \[551] ,
  \[741] ,
  \[552] ,
  \[742] ,
  \[553] ,
  \[743] ,
  \[554] ,
  \new_C<85> ,
  \[744] ,
  \[555] ,
  \new_C<86> ,
  \[745] ,
  \[556] ,
  \new_C<87> ,
  \[746] ,
  \[557] ,
  \new_C<88> ,
  \[747] ,
  \[558] ,
  \new_C<81> ,
  \[748] ,
  \[559] ,
  \new_C<82> ,
  \[749] ,
  \new_C<83> ,
  \new_C<84> ,
  \new_C<80> ,
  \[560] ,
  \[750] ,
  \[561] ,
  \[751] ,
  \new_D<99> ,
  \[562] ,
  \[752] ,
  \[563] ,
  \[753] ,
  \[564] ,
  \[754] ,
  \[565] ,
  \[755] ,
  \$$COND1<0>8.1 ,
  \new_D<95> ,
  \[566] ,
  \[756] ,
  \new_D<96> ,
  \[567] ,
  \[757] ,
  \new_D<97> ;
assign
  \[568]  = \new_D<76> ,
  \[758]  = (~\D<60>  & \C<60> ) | (\D<60>  & ~\C<60> ),
  \new_D<98>  = (\[648]  & (\D<98>  & \C<98> )) | ((\[682]  & \[652] ) | ((~\[681]  & \[650] ) | ((\[681]  & \[649] ) | ((\[654]  & \key<197> ) | (\[651]  & \key<205> ))))),
  \[569]  = \new_D<75> ,
  \[759]  = \D<59>  | \C<59> ,
  \new_D<91>  = (\[648]  & (\D<91>  & \C<91> )) | ((\[696]  & \[652] ) | ((~\[695]  & \[650] ) | ((\[695]  & \[649] ) | ((\[654]  & \key<253> ) | (\[651]  & \key<198> ))))),
  \new_D<92>  = (\[648]  & (\D<92>  & \C<92> )) | ((\[694]  & \[652] ) | ((~\[693]  & \[650] ) | ((\[693]  & \[649] ) | ((\[654]  & \key<245> ) | (\[651]  & \key<253> ))))),
  \new_D<93>  = (\[648]  & (\D<93>  & \C<93> )) | ((\[692]  & \[652] ) | ((~\[691]  & \[650] ) | ((\[691]  & \[649] ) | ((\[654]  & \key<237> ) | (\[651]  & \key<245> ))))),
  \new_D<94>  = (\[648]  & (\D<94>  & \C<94> )) | ((\[690]  & \[652] ) | ((~\[689]  & \[650] ) | ((\[689]  & \[649] ) | ((\[654]  & \key<229> ) | (\[651]  & \key<237> ))))),
  \KSi<130>  = \D<32> ,
  \KSi<131>  = \D<47> ,
  \KSi<132>  = \D<43> ,
  \[570]  = \new_D<74> ,
  \[760]  = (~\D<59>  & \C<59> ) | (\D<59>  & ~\C<59> ),
  \KSi<133>  = \D<48> ,
  \new_D<90>  = (\[648]  & (\D<90>  & \C<90> )) | ((\[698]  & \[652] ) | ((~\[697]  & \[650] ) | ((\[697]  & \[649] ) | ((\[654]  & \key<198> ) | (\[651]  & \key<206> ))))),
  \[571]  = \new_D<73> ,
  \[761]  = \D<58>  | \C<58> ,
  \KSi<134>  = \D<38> ,
  \[572]  = \new_D<72> ,
  \[762]  = (~\D<58>  & \C<58> ) | (\D<58>  & ~\C<58> ),
  \KSi<135>  = \D<55> ,
  \[573]  = \new_D<71> ,
  \[763]  = \D<57>  | \C<57> ,
  \KSi<136>  = \D<33> ,
  \[574]  = \new_D<70> ,
  \[764]  = (~\D<57>  & \C<57> ) | (\D<57>  & ~\C<57> ),
  \KSi<137>  = \D<52> ,
  \[575]  = \new_D<69> ,
  \[765]  = \D<56>  | \C<56> ,
  \KSi<138>  = \D<45> ,
  \[576]  = \new_D<68> ,
  \[766]  = (~\D<56>  & \C<56> ) | (\D<56>  & ~\C<56> ),
  \KSi<139>  = \D<31> ,
  \[577]  = \new_D<67> ,
  \[767]  = \D<55>  | \C<55> ,
  \[578]  = \new_D<66> ,
  \[768]  = (~\D<55>  & \C<55> ) | (\D<55>  & ~\C<55> ),
  \new_C<111>  = (\[647]  & (\D<111>  & \C<111> )) | ((\[656]  & \[653] ) | ((~\[655]  & \[649] ) | ((\[655]  & \[650] ) | ((\[654]  & \key<56> ) | (\[651]  & \key<227> ))))),
  \[579]  = \new_D<65> ,
  \[769]  = \D<54>  | \C<54> ,
  \new_C<110>  = (\[647]  & (\D<110>  & \C<110> )) | ((\[658]  & \[653] ) | ((~\[657]  & \[649] ) | ((\[657]  & \[650] ) | ((\[654]  & \key<227> ) | (\[651]  & \key<235> ))))),
  \[580]  = \new_D<64> ,
  \[770]  = (~\D<54>  & \C<54> ) | (\D<54>  & ~\C<54> ),
  \[581]  = \new_D<63> ,
  \[771]  = \D<53>  | \C<53> ,
  \[582]  = \new_D<62> ,
  \[772]  = (~\D<53>  & \C<53> ) | (\D<53>  & ~\C<53> ),
  \[583]  = \new_D<61> ,
  \[773]  = \D<52>  | \C<52> ,
  \[584]  = \new_D<60> ,
  \[774]  = (~\D<52>  & \C<52> ) | (\D<52>  & ~\C<52> ),
  \[585]  = \new_D<59> ,
  \[775]  = \D<51>  | \C<51> ,
  \[586]  = \new_D<58> ,
  \[776]  = (~\D<51>  & \C<51> ) | (\D<51>  & ~\C<51> ),
  \[587]  = \new_D<57> ,
  \[777]  = \D<50>  | \C<50> ,
  \[588]  = \new_D<56> ,
  \[778]  = (~\D<50>  & \C<50> ) | (\D<50>  & ~\C<50> ),
  \[589]  = \new_D<55> ,
  \[779]  = \D<49>  | \C<49> ,
  \[590]  = \new_D<54> ,
  \[780]  = (~\D<49>  & \C<49> ) | (\D<49>  & ~\C<49> ),
  \[591]  = \new_D<53> ,
  \[781]  = \D<48>  | \C<48> ,
  \[592]  = \new_D<52> ,
  \[782]  = (~\D<48>  & \C<48> ) | (\D<48>  & ~\C<48> ),
  \[593]  = \new_D<51> ,
  \[783]  = \D<47>  | \C<47> ,
  \[594]  = \new_D<50> ,
  \[784]  = (~\D<47>  & \C<47> ) | (\D<47>  & ~\C<47> ),
  \[595]  = \new_D<49> ,
  \[785]  = \D<46>  | \C<46> ,
  \[596]  = \new_D<48> ,
  \[786]  = (~\D<46>  & \C<46> ) | (\D<46>  & ~\C<46> ),
  \[597]  = \new_D<47> ,
  \[787]  = \D<45>  | \C<45> ,
  \[598]  = \new_D<46> ,
  \[788]  = (~\D<45>  & \C<45> ) | (\D<45>  & ~\C<45> ),
  \[599]  = \new_D<45> ,
  \[789]  = \D<44>  | \C<44> ,
  \KSi<100>  = \D<18> ,
  \KSi<101>  = \D<26> ,
  \KSi<102>  = \D<1> ,
  \[790]  = (~\D<44>  & \C<44> ) | (\D<44>  & ~\C<44> ),
  \KSi<103>  = \D<11> ,
  \[791]  = \D<43>  | \C<43> ,
  \KSi<104>  = \D<22> ,
  \new_D<59>  = (\[648]  & (\D<59>  & \C<59> )) | ((\[760]  & \[652] ) | ((~\[759]  & \[650] ) | ((\[759]  & \[649] ) | ((\[654]  & \key<158> ) | (\[651]  & \key<166> ))))),
  \[792]  = (~\D<43>  & \C<43> ) | (\D<43>  & ~\C<43> ),
  \KSi<105>  = \D<16> ,
  \[793]  = \D<42>  | \C<42> ,
  \KSi<106>  = \D<4> ,
  \[794]  = (~\D<42>  & \C<42> ) | (\D<42>  & ~\C<42> ),
  \KSi<107>  = \D<19> ,
  \[795]  = \D<41>  | \C<41> ,
  \KSi<108>  = \D<15> ,
  \new_D<55>  = (\[648]  & (\D<55>  & \C<55> )) | ((\[768]  & \[652] ) | ((~\[767]  & \[650] ) | ((\[767]  & \[649] ) | ((\[654]  & \key<190> ) | (\[651]  & \key<67> ))))),
  \[796]  = (~\D<41>  & \C<41> ) | (\D<41>  & ~\C<41> ),
  \KSi<109>  = \D<20> ,
  \new_D<56>  = (\[648]  & (\D<56>  & \C<56> )) | ((\[766]  & \[652] ) | ((~\[765]  & \[650] ) | ((\[765]  & \[649] ) | ((\[654]  & \key<182> ) | (\[651]  & \key<190> ))))),
  \[797]  = \D<40>  | \C<40> ,
  \new_D<57>  = (\[648]  & (\D<57>  & \C<57> )) | ((\[764]  & \[652] ) | ((~\[763]  & \[650] ) | ((\[763]  & \[649] ) | ((\[654]  & \key<174> ) | (\[651]  & \key<182> ))))),
  \[798]  = (~\D<40>  & \C<40> ) | (\D<40>  & ~\C<40> ),
  \new_D<58>  = (\[648]  & (\D<58>  & \C<58> )) | ((\[762]  & \[652] ) | ((~\[761]  & \[650] ) | ((\[761]  & \[649] ) | ((\[654]  & \key<166> ) | (\[651]  & \key<174> ))))),
  \[799]  = \D<39>  | \C<39> ,
  \new_D<51>  = (\[648]  & (\D<51>  & \C<51> )) | ((\[776]  & \[652] ) | ((~\[775]  & \[650] ) | ((\[775]  & \[649] ) | ((\[654]  & \key<91> ) | (\[651]  & \key<68> ))))),
  \new_D<52>  = (\[648]  & (\D<52>  & \C<52> )) | ((\[774]  & \[652] ) | ((~\[773]  & \[650] ) | ((\[773]  & \[649] ) | ((\[654]  & \key<83> ) | (\[651]  & \key<91> ))))),
  \new_D<53>  = (\[648]  & (\D<53>  & \C<53> )) | ((\[772]  & \[652] ) | ((~\[771]  & \[650] ) | ((\[771]  & \[649] ) | ((\[654]  & \key<75> ) | (\[651]  & \key<83> ))))),
  \new_D<54>  = (\[648]  & (\D<54>  & \C<54> )) | ((\[770]  & \[652] ) | ((~\[769]  & \[650] ) | ((\[769]  & \[649] ) | ((\[654]  & \key<67> ) | (\[651]  & \key<75> ))))),
  \new_D<50>  = (\[648]  & (\D<50>  & \C<50> )) | ((\[778]  & \[652] ) | ((~\[777]  & \[650] ) | ((\[777]  & \[649] ) | ((\[654]  & \key<68> ) | (\[651]  & \key<76> ))))),
  \new_D<69>  = (\[648]  & (\D<69>  & \C<69> )) | ((\[740]  & \[652] ) | ((~\[739]  & \[650] ) | ((\[739]  & \[649] ) | ((\[654]  & \key<141> ) | (\[651]  & \key<149> ))))),
  \new_D<65>  = (\[648]  & (\D<65>  & \C<65> )) | ((\[748]  & \[652] ) | ((~\[747]  & \[650] ) | ((\[747]  & \[649] ) | ((\[654]  & \key<173> ) | (\[651]  & \key<181> ))))),
  \new_D<66>  = (\[648]  & (\D<66>  & \C<66> )) | ((\[746]  & \[652] ) | ((~\[745]  & \[650] ) | ((\[745]  & \[649] ) | ((\[654]  & \key<165> ) | (\[651]  & \key<173> ))))),
  \new_D<67>  = (\[648]  & (\D<67>  & \C<67> )) | ((\[744]  & \[652] ) | ((~\[743]  & \[650] ) | ((\[743]  & \[649] ) | ((\[654]  & \key<157> ) | (\[651]  & \key<165> ))))),
  \new_D<68>  = (\[648]  & (\D<68>  & \C<68> )) | ((\[742]  & \[652] ) | ((~\[741]  & \[650] ) | ((\[741]  & \[649] ) | ((\[654]  & \key<149> ) | (\[651]  & \key<157> ))))),
  \new_D<61>  = (\[648]  & (\D<61>  & \C<61> )) | ((\[756]  & \[652] ) | ((~\[755]  & \[650] ) | ((\[755]  & \[649] ) | ((\[654]  & \key<142> ) | (\[651]  & \key<150> ))))),
  \new_D<62>  = (\[648]  & (\D<62>  & \C<62> )) | ((\[754]  & \[652] ) | ((~\[753]  & \[650] ) | ((\[753]  & \[649] ) | ((\[654]  & \key<134> ) | (\[651]  & \key<142> ))))),
  \new_D<63>  = (\[648]  & (\D<63>  & \C<63> )) | ((\[752]  & \[652] ) | ((~\[751]  & \[650] ) | ((\[751]  & \[649] ) | ((\[654]  & \key<189> ) | (\[651]  & \key<134> ))))),
  \new_D<64>  = (\[648]  & (\D<64>  & \C<64> )) | ((\[750]  & \[652] ) | ((~\[749]  & \[650] ) | ((\[749]  & \[649] ) | ((\[654]  & \key<181> ) | (\[651]  & \key<189> ))))),
  \new_D<60>  = (\[648]  & (\D<60>  & \C<60> )) | ((\[758]  & \[652] ) | ((~\[757]  & \[650] ) | ((\[757]  & \[649] ) | ((\[654]  & \key<150> ) | (\[651]  & \key<158> ))))),
  \new_D<79>  = (\[648]  & (\D<79>  & \C<79> )) | ((\[720]  & \[652] ) | ((~\[719]  & \[650] ) | ((\[719]  & \[649] ) | ((\[654]  & \key<155> ) | (\[651]  & \key<132> ))))),
  \new_D<75>  = (\[648]  & (\D<75>  & \C<75> )) | ((\[728]  & \[652] ) | ((~\[727]  & \[650] ) | ((\[727]  & \[649] ) | ((\[654]  & \key<156> ) | (\[651]  & \key<164> ))))),
  \new_D<76>  = (\[648]  & (\D<76>  & \C<76> )) | ((\[726]  & \[652] ) | ((~\[725]  & \[650] ) | ((\[725]  & \[649] ) | ((\[654]  & \key<148> ) | (\[651]  & \key<156> ))))),
  \new_D<77>  = (\[648]  & (\D<77>  & \C<77> )) | ((\[724]  & \[652] ) | ((~\[723]  & \[650] ) | ((\[723]  & \[649] ) | ((\[654]  & \key<140> ) | (\[651]  & \key<148> ))))),
  \new_D<78>  = (\[648]  & (\D<78>  & \C<78> )) | ((\[722]  & \[652] ) | ((~\[721]  & \[650] ) | ((\[721]  & \[649] ) | ((\[654]  & \key<132> ) | (\[651]  & \key<140> ))))),
  \new_D<71>  = (\[648]  & (\D<71>  & \C<71> )) | ((\[736]  & \[652] ) | ((~\[735]  & \[650] ) | ((\[735]  & \[649] ) | ((\[654]  & \key<188> ) | (\[651]  & \key<133> ))))),
  \new_D<72>  = (\[648]  & (\D<72>  & \C<72> )) | ((\[734]  & \[652] ) | ((~\[733]  & \[650] ) | ((\[733]  & \[649] ) | ((\[654]  & \key<180> ) | (\[651]  & \key<188> ))))),
  \new_D<73>  = (\[648]  & (\D<73>  & \C<73> )) | ((\[732]  & \[652] ) | ((~\[731]  & \[650] ) | ((\[731]  & \[649] ) | ((\[654]  & \key<172> ) | (\[651]  & \key<180> ))))),
  \new_D<74>  = (\[648]  & (\D<74>  & \C<74> )) | ((\[730]  & \[652] ) | ((~\[729]  & \[650] ) | ((\[729]  & \[649] ) | ((\[654]  & \key<164> ) | (\[651]  & \key<172> ))))),
  \KSi<190>  = \D<84> ,
  \KSi<191>  = \D<87> ,
  \new_D<70>  = (\[648]  & (\D<70>  & \C<70> )) | ((\[738]  & \[652] ) | ((~\[737]  & \[650] ) | ((\[737]  & \[649] ) | ((\[654]  & \key<133> ) | (\[651]  & \key<141> ))))),
  \new_D<111>  = (\[648]  & (\D<111>  & \C<111> )) | ((\[656]  & \[652] ) | ((~\[655]  & \[650] ) | ((\[655]  & \[649] ) | ((\[654]  & \key<62> ) | (\[651]  & \key<195> ))))),
  \new_D<89>  = (\[648]  & (\D<89>  & \C<89> )) | ((\[700]  & \[652] ) | ((~\[699]  & \[650] ) | ((\[699]  & \[649] ) | ((\[654]  & \key<206> ) | (\[651]  & \key<214> ))))),
  \new_D<85>  = (\[648]  & (\D<85>  & \C<85> )) | ((\[708]  & \[652] ) | ((~\[707]  & \[650] ) | ((\[707]  & \[649] ) | ((\[654]  & \key<238> ) | (\[651]  & \key<246> ))))),
  \new_D<110>  = (\[648]  & (\D<110>  & \C<110> )) | ((\[658]  & \[652] ) | ((~\[657]  & \[650] ) | ((\[657]  & \[649] ) | ((\[654]  & \key<195> ) | (\[651]  & \key<203> ))))),
  \new_D<86>  = (\[648]  & (\D<86>  & \C<86> )) | ((\[706]  & \[652] ) | ((~\[705]  & \[650] ) | ((\[705]  & \[649] ) | ((\[654]  & \key<230> ) | (\[651]  & \key<238> ))))),
  \new_D<87>  = (\[648]  & (\D<87>  & \C<87> )) | ((\[704]  & \[652] ) | ((~\[703]  & \[650] ) | ((\[703]  & \[649] ) | ((\[654]  & \key<222> ) | (\[651]  & \key<230> ))))),
  \new_D<88>  = (\[648]  & (\D<88>  & \C<88> )) | ((\[702]  & \[652] ) | ((~\[701]  & \[650] ) | ((\[701]  & \[649] ) | ((\[654]  & \key<214> ) | (\[651]  & \key<222> ))))),
  \new_D<81>  = (\[648]  & (\D<81>  & \C<81> )) | ((\[716]  & \[652] ) | ((~\[715]  & \[650] ) | ((\[715]  & \[649] ) | ((\[654]  & \key<139> ) | (\[651]  & \key<147> ))))),
  \new_D<82>  = (\[648]  & (\D<82>  & \C<82> )) | ((\[714]  & \[652] ) | ((~\[713]  & \[650] ) | ((\[713]  & \[649] ) | ((\[654]  & \key<131> ) | (\[651]  & \key<139> ))))),
  \new_D<83>  = (\[648]  & (\D<83>  & \C<83> )) | ((\[712]  & \[652] ) | ((~\[711]  & \[650] ) | ((\[711]  & \[649] ) | ((\[654]  & \key<254> ) | (\[651]  & \key<131> ))))),
  \new_D<84>  = (\[648]  & (\D<84>  & \C<84> )) | ((\[710]  & \[652] ) | ((~\[709]  & \[650] ) | ((\[709]  & \[649] ) | ((\[654]  & \key<246> ) | (\[651]  & \key<254> ))))),
  \new_C<109>  = (\[647]  & (\D<109>  & \C<109> )) | ((\[660]  & \[653] ) | ((~\[659]  & \[649] ) | ((\[659]  & \[650] ) | ((\[654]  & \key<235> ) | (\[651]  & \key<243> ))))),
  \new_D<80>  = (\[648]  & (\D<80>  & \C<80> )) | ((\[718]  & \[652] ) | ((~\[717]  & \[650] ) | ((\[717]  & \[649] ) | ((\[654]  & \key<147> ) | (\[651]  & \key<155> ))))),
  \new_C<106>  = (\[647]  & (\D<106>  & \C<106> )) | ((\[666]  & \[653] ) | ((~\[665]  & \[649] ) | ((\[665]  & \[650] ) | ((\[654]  & \key<194> ) | (\[651]  & \key<202> ))))),
  \new_C<105>  = (\[647]  & (\D<105>  & \C<105> )) | ((\[668]  & \[653] ) | ((~\[667]  & \[649] ) | ((\[667]  & \[650] ) | ((\[654]  & \key<202> ) | (\[651]  & \key<210> ))))),
  \new_C<108>  = (\[647]  & (\D<108>  & \C<108> )) | ((\[662]  & \[653] ) | ((~\[661]  & \[649] ) | ((\[661]  & \[650] ) | ((\[654]  & \key<243> ) | (\[651]  & \key<251> ))))),
  \new_C<107>  = (\[647]  & (\D<107>  & \C<107> )) | ((\[664]  & \[653] ) | ((~\[663]  & \[649] ) | ((\[663]  & \[650] ) | ((\[654]  & \key<251> ) | (\[651]  & \key<194> ))))),
  \new_C<102>  = (\[647]  & (\D<102>  & \C<102> )) | ((\[674]  & \[653] ) | ((~\[673]  & \[649] ) | ((\[673]  & \[650] ) | ((\[654]  & \key<226> ) | (\[651]  & \key<234> ))))),
  \new_C<101>  = (\[647]  & (\D<101>  & \C<101> )) | ((\[676]  & \[653] ) | ((~\[675]  & \[649] ) | ((\[675]  & \[650] ) | ((\[654]  & \key<234> ) | (\[651]  & \key<242> ))))),
  \new_C<104>  = (\[647]  & (\D<104>  & \C<104> )) | ((\[670]  & \[653] ) | ((~\[669]  & \[649] ) | ((\[669]  & \[650] ) | ((\[654]  & \key<210> ) | (\[651]  & \key<218> ))))),
  \new_C<103>  = (\[647]  & (\D<103>  & \C<103> )) | ((\[672]  & \[653] ) | ((~\[671]  & \[649] ) | ((\[671]  & \[650] ) | ((\[654]  & \key<218> ) | (\[651]  & \key<226> ))))),
  \new_C<100>  = (\[647]  & (\D<100>  & \C<100> )) | ((\[678]  & \[653] ) | ((~\[677]  & \[649] ) | ((\[677]  & \[650] ) | ((\[654]  & \key<242> ) | (\[651]  & \key<250> ))))),
  \KSi<160>  = \D<61> ,
  \KSi<161>  = \D<80> ,
  \KSi<162>  = \D<73> ,
  \[600]  = \new_D<44> ,
  \KSi<163>  = \D<69> ,
  \[601]  = \new_D<43> ,
  \KSi<164>  = \D<77> ,
  \[602]  = \new_D<42> ,
  \KSi<165>  = \D<63> ,
  \[603]  = \new_D<41> ,
  \KSi<166>  = \D<56> ,
  \[224]  = (\[880]  & (~\$$COND1<0>8.1  & (~\[225]  & ~\start<0> ))) | ((\[880]  & (\$$COND1<0>8.1  & \[225] )) | ((~\$$COND1<0>8.1  & (\count<3>  & ~\start<0> )) | ((\$$COND1<0>8.1  & (\[225]  & ~\count<3> )) | ((\[227]  & (~\[225]  & \count<3> )) | \[882] )))),
  \[604]  = \new_D<40> ,
  \KSi<167>  = \D<59> ,
  \[225]  = (\[646]  & (~\[227]  & (\count<1>  & ~\count<2> ))) | ((\[227]  & (~\count<1>  & (~\count<2>  & ~\encrypt<0> ))) | ((\[646]  & (~\count<1>  & \count<2> )) | ((~\[227]  & (\count<2>  & ~\encrypt<0> )) | ((\[880]  & \[227] ) | \[882] )))),
  \[605]  = \new_D<39> ,
  \KSi<168>  = \D<104> ,
  \[226]  = (\[646]  & (~\[227]  & ~\count<1> )) | ((~\[227]  & (\count<1>  & ~\encrypt<0> )) | ((\[227]  & (~\count<1>  & ~\encrypt<0> )) | ((\[227]  & (\count<1>  & \encrypt<0> )) | \[882] ))),
  \[606]  = \new_D<38> ,
  \KSi<169>  = \D<107> ,
  \[227]  = (~\count<0>  & ~\start<0> ) | \[651] ,
  \[607]  = \new_D<37> ,
  \[228]  = (\[653]  & (\$$COND1<0>8.1  & \count<1> )) | (\[649]  & \$$COND0<0>5.1 ),
  \[608]  = \new_D<36> ,
  \[609]  = \new_D<35> ,
  \KSi<150>  = \D<57> ,
  \KSi<151>  = \D<67> ,
  \KSi<152>  = \D<78> ,
  \[610]  = \new_D<34> ,
  \[800]  = (~\D<39>  & \C<39> ) | (\D<39>  & ~\C<39> ),
  \KSi<153>  = \D<70> ,
  \[421]  = \new_C<111> ,
  \[611]  = \new_D<33> ,
  \[801]  = \D<38>  | \C<38> ,
  \KSi<154>  = \D<60> ,
  \[422]  = \new_C<110> ,
  \[612]  = \new_D<32> ,
  \[802]  = (~\D<38>  & \C<38> ) | (\D<38>  & ~\C<38> ),
  \KSi<155>  = \D<75> ,
  \[423]  = \new_C<109> ,
  \[613]  = \new_D<31> ,
  \[803]  = \D<37>  | \C<37> ,
  \KSi<156>  = \D<71> ,
  \[424]  = \new_C<108> ,
  \[614]  = \new_D<30> ,
  \[804]  = (~\D<37>  & \C<37> ) | (\D<37>  & ~\C<37> ),
  \KSi<157>  = \D<76> ,
  \[425]  = \new_C<107> ,
  \[615]  = \new_D<29> ,
  \[805]  = \D<36>  | \C<36> ,
  \KSi<158>  = \D<66> ,
  \[426]  = \new_C<106> ,
  \[616]  = \new_D<28> ,
  \[806]  = (~\D<36>  & \C<36> ) | (\D<36>  & ~\C<36> ),
  \KSi<159>  = \D<83> ,
  \new_D<1>  = (\[648]  & (\D<1>  & \C<1> )) | ((\[876]  & \[652] ) | ((~\[875]  & \[650] ) | ((\[875]  & \[649] ) | ((\[654]  & \key<46> ) | (\[651]  & \key<54> ))))),
  \[427]  = \new_C<105> ,
  \[617]  = \new_D<27> ,
  \[807]  = \D<35>  | \C<35> ,
  \new_D<2>  = (\[648]  & (\D<2>  & \C<2> )) | ((\[874]  & \[652] ) | ((~\[873]  & \[650] ) | ((\[873]  & \[649] ) | ((\[654]  & \key<38> ) | (\[651]  & \key<46> ))))),
  \[428]  = \new_C<104> ,
  \[618]  = \new_D<26> ,
  \[808]  = (~\D<35>  & \C<35> ) | (\D<35>  & ~\C<35> ),
  \new_D<3>  = (\[648]  & (\D<3>  & \C<3> )) | ((\[872]  & \[652] ) | ((~\[871]  & \[650] ) | ((\[871]  & \[649] ) | ((\[654]  & \key<30> ) | (\[651]  & \key<38> ))))),
  \[429]  = \new_C<103> ,
  \[619]  = \new_D<25> ,
  \[809]  = \D<34>  | \C<34> ,
  \KSi<0>  = \C<13> ,
  \new_D<4>  = (\[648]  & (\D<4>  & \C<4> )) | ((\[870]  & \[652] ) | ((~\[869]  & \[650] ) | ((\[869]  & \[649] ) | ((\[654]  & \key<22> ) | (\[651]  & \key<30> ))))),
  \KSi<1>  = \C<16> ,
  \KSi<2>  = \C<10> ,
  \KSi<3>  = \C<23> ,
  \KSi<4>  = \C<0> ,
  \KSi<180>  = \D<99> ,
  \new_D<0>  = (\[648]  & (\D<0>  & \C<0> )) | ((\[878]  & \[652] ) | ((~\[877]  & \[650] ) | ((\[877]  & \[649] ) | ((\[654]  & \key<54> ) | (\[651]  & \key<62> ))))),
  \KSi<5>  = \C<4> ,
  \KSi<181>  = \D<104> ,
  \new_D<9>  = (\[648]  & (\D<9>  & \C<9> )) | ((\[860]  & \[652] ) | ((~\[859]  & \[650] ) | ((\[859]  & \[649] ) | ((\[654]  & \key<45> ) | (\[651]  & \key<53> ))))),
  \KSi<6>  = \C<2> ,
  \KSi<182>  = \D<94> ,
  \[430]  = \new_C<102> ,
  \[620]  = \new_D<24> ,
  \[810]  = (~\D<34>  & \C<34> ) | (\D<34>  & ~\C<34> ),
  \KSi<7>  = \C<27> ,
  \KSi<183>  = \D<111> ,
  \[431]  = \new_C<101> ,
  \[621]  = \new_D<23> ,
  \[811]  = \D<33>  | \C<33> ,
  \KSi<8>  = \C<14> ,
  \KSi<184>  = \D<89> ,
  \[432]  = \new_C<100> ,
  \[622]  = \new_D<22> ,
  \[812]  = (~\D<33>  & \C<33> ) | (\D<33>  & ~\C<33> ),
  \KSi<9>  = \C<5> ,
  \KSi<185>  = \D<108> ,
  \new_D<5>  = (\[648]  & (\D<5>  & \C<5> )) | ((\[868]  & \[652] ) | ((~\[867]  & \[650] ) | ((\[867]  & \[649] ) | ((\[654]  & \key<14> ) | (\[651]  & \key<22> ))))),
  \[433]  = \new_C<99> ,
  \[623]  = \new_D<21> ,
  \[813]  = \D<32>  | \C<32> ,
  \KSi<186>  = \D<101> ,
  \new_D<6>  = (\[648]  & (\D<6>  & \C<6> )) | ((\[866]  & \[652] ) | ((~\[865]  & \[650] ) | ((\[865]  & \[649] ) | ((\[654]  & \key<6> ) | (\[651]  & \key<14> ))))),
  \[434]  = \new_C<98> ,
  \[624]  = \new_D<20> ,
  \[814]  = (~\D<32>  & \C<32> ) | (\D<32>  & ~\C<32> ),
  \KSi<187>  = \D<87> ,
  \new_D<7>  = (\[648]  & (\D<7>  & \C<7> )) | ((\[864]  & \[652] ) | ((~\[863]  & \[650] ) | ((\[863]  & \[649] ) | ((\[654]  & \key<61> ) | (\[651]  & \key<6> ))))),
  \[435]  = \new_C<97> ,
  \[625]  = \new_D<19> ,
  \[815]  = \D<31>  | \C<31> ,
  \KSi<188>  = \D<105> ,
  \new_D<8>  = (\[648]  & (\D<8>  & \C<8> )) | ((\[862]  & \[652] ) | ((~\[861]  & \[650] ) | ((\[861]  & \[649] ) | ((\[654]  & \key<53> ) | (\[651]  & \key<61> ))))),
  \[436]  = \new_C<96> ,
  \[626]  = \new_D<18> ,
  \[816]  = (~\D<31>  & \C<31> ) | (\D<31>  & ~\C<31> ),
  \KSi<189>  = \D<91> ,
  \[437]  = \new_C<95> ,
  \[627]  = \new_D<17> ,
  \[817]  = \D<30>  | \C<30> ,
  \[438]  = \new_C<94> ,
  \[628]  = \new_D<16> ,
  \[818]  = (~\D<30>  & \C<30> ) | (\D<30>  & ~\C<30> ),
  \[439]  = \new_C<93> ,
  \[629]  = \new_D<15> ,
  \[819]  = \D<29>  | \C<29> ,
  \KSi<170>  = \D<86> ,
  \KSi<171>  = \D<92> ,
  \KSi<172>  = \D<102> ,
  \[440]  = \new_C<92> ,
  \[630]  = \new_D<14> ,
  \[820]  = (~\D<29>  & \C<29> ) | (\D<29>  & ~\C<29> ),
  \KSi<173>  = \D<110> ,
  \[441]  = \new_C<91> ,
  \[631]  = \new_D<13> ,
  \[821]  = \D<28>  | \C<28> ,
  \KSi<174>  = \D<85> ,
  \[442]  = \new_C<90> ,
  \[632]  = \new_D<12> ,
  \[822]  = (~\D<28>  & \C<28> ) | (\D<28>  & ~\C<28> ),
  \KSi<175>  = \D<95> ,
  \[443]  = \new_C<89> ,
  \[633]  = \new_D<11> ,
  \[823]  = \D<27>  | \C<27> ,
  \KSi<176>  = \D<106> ,
  \[444]  = \new_C<88> ,
  \[634]  = \new_D<10> ,
  \[824]  = (~\D<27>  & \C<27> ) | (\D<27>  & ~\C<27> ),
  \KSi<177>  = \D<100> ,
  \[445]  = \new_C<87> ,
  \[635]  = \new_D<9> ,
  \[825]  = \D<26>  | \C<26> ,
  \KSi<178>  = \D<88> ,
  \[446]  = \new_C<86> ,
  \[636]  = \new_D<8> ,
  \[826]  = (~\D<26>  & \C<26> ) | (\D<26>  & ~\C<26> ),
  \KSi<179>  = \D<103> ,
  \[447]  = \new_C<85> ,
  \[637]  = \new_D<7> ,
  \[827]  = \D<25>  | \C<25> ,
  \[448]  = \new_C<84> ,
  \[638]  = \new_D<6> ,
  \[828]  = (~\D<25>  & \C<25> ) | (\D<25>  & ~\C<25> ),
  \[449]  = \new_C<83> ,
  \[639]  = \new_D<5> ,
  \new_D<109>  = (\[648]  & (\D<109>  & \C<109> )) | ((\[660]  & \[652] ) | ((~\[659]  & \[650] ) | ((\[659]  & \[649] ) | ((\[654]  & \key<203> ) | (\[651]  & \key<211> ))))),
  \[829]  = \D<24>  | \C<24> ,
  \new_D<106>  = (\[648]  & (\D<106>  & \C<106> )) | ((\[666]  & \[652] ) | ((~\[665]  & \[650] ) | ((\[665]  & \[649] ) | ((\[654]  & \key<196> ) | (\[651]  & \key<204> ))))),
  \new_D<105>  = (\[648]  & (\D<105>  & \C<105> )) | ((\[668]  & \[652] ) | ((~\[667]  & \[650] ) | ((\[667]  & \[649] ) | ((\[654]  & \key<204> ) | (\[651]  & \key<212> ))))),
  \new_D<108>  = (\[648]  & (\D<108>  & \C<108> )) | ((\[662]  & \[652] ) | ((~\[661]  & \[650] ) | ((\[661]  & \[649] ) | ((\[654]  & \key<211> ) | (\[651]  & \key<219> ))))),
  \new_D<107>  = (\[648]  & (\D<107>  & \C<107> )) | ((\[664]  & \[652] ) | ((~\[663]  & \[650] ) | ((\[663]  & \[649] ) | ((\[654]  & \key<219> ) | (\[651]  & \key<196> ))))),
  \[450]  = \new_C<82> ,
  \[640]  = \new_D<4> ,
  \new_D<102>  = (\[648]  & (\D<102>  & \C<102> )) | ((\[674]  & \[652] ) | ((~\[673]  & \[650] ) | ((\[673]  & \[649] ) | ((\[654]  & \key<228> ) | (\[651]  & \key<172> ))))),
  \[830]  = (~\D<24>  & \C<24> ) | (\D<24>  & ~\C<24> ),
  \[451]  = \new_C<81> ,
  \[641]  = \new_D<3> ,
  \new_D<101>  = (\[648]  & (\D<101>  & \C<101> )) | ((\[676]  & \[652] ) | ((~\[675]  & \[650] ) | ((\[675]  & \[649] ) | ((\[654]  & \key<172> ) | (\[651]  & \key<244> ))))),
  \[831]  = \D<23>  | \C<23> ,
  \[452]  = \new_C<80> ,
  \[642]  = \new_D<2> ,
  \new_D<104>  = (\[648]  & (\D<104>  & \C<104> )) | ((\[670]  & \[652] ) | ((~\[669]  & \[650] ) | ((\[669]  & \[649] ) | ((\[654]  & \key<212> ) | (\[651]  & \key<220> ))))),
  \[832]  = (~\D<23>  & \C<23> ) | (\D<23>  & ~\C<23> ),
  \[453]  = \new_C<79> ,
  \[643]  = \new_D<1> ,
  \new_D<103>  = (\[648]  & (\D<103>  & \C<103> )) | ((\[672]  & \[652] ) | ((~\[671]  & \[650] ) | ((\[671]  & \[649] ) | ((\[654]  & \key<220> ) | (\[651]  & \key<228> ))))),
  \[833]  = \D<22>  | \C<22> ,
  \[454]  = \new_C<78> ,
  \[644]  = \new_D<0> ,
  \[834]  = (~\D<22>  & \C<22> ) | (\D<22>  & ~\C<22> ),
  \[455]  = \new_C<77> ,
  \[645]  = ~\start<0>  & ~\encrypt<0> ,
  \[835]  = \D<21>  | \C<21> ,
  \[456]  = \new_C<76> ,
  \[646]  = ~\start<0>  & \encrypt<0> ,
  \new_D<100>  = (\[648]  & (\D<100>  & \C<100> )) | ((\[678]  & \[652] ) | ((~\[677]  & \[650] ) | ((\[677]  & \[649] ) | ((\[654]  & \key<244> ) | (\[651]  & \key<252> ))))),
  \[836]  = (~\D<21>  & \C<21> ) | (\D<21>  & ~\C<21> ),
  \[457]  = \new_C<75> ,
  \[647]  = (\$$COND0<0>5.1  & ~\start<0> ) | \[645] ,
  \[837]  = \D<20>  | \C<20> ,
  \[458]  = \new_C<74> ,
  \[648]  = (~\$$COND0<0>5.1  & ~\start<0> ) | \[645] ,
  \[838]  = (~\D<20>  & \C<20> ) | (\D<20>  & ~\C<20> ),
  \[459]  = \new_C<73> ,
  \[649]  = \[645]  & \$$COND1<0>8.1 ,
  \[839]  = \D<19>  | \C<19> ,
  \[460]  = \new_C<72> ,
  \new_C<19>  = (\[647]  & (\D<19>  & \C<19> )) | ((\[840]  & \[653] ) | ((~\[839]  & \[649] ) | ((\[839]  & \[650] ) | ((\[654]  & \key<26> ) | (\[651]  & \key<34> ))))),
  \[650]  = \[645]  & ~\$$COND1<0>8.1 ,
  \[840]  = (~\D<19>  & \C<19> ) | (\D<19>  & ~\C<19> ),
  \[461]  = \new_C<71> ,
  \[651]  = \start<0>  & ~\encrypt<0> ,
  \[841]  = \D<18>  | \C<18> ,
  \[462]  = \new_C<70> ,
  \[652]  = \[646]  & \$$COND0<0>5.1 ,
  \[842]  = (~\D<18>  & \C<18> ) | (\D<18>  & ~\C<18> ),
  \[463]  = \new_C<69> ,
  \[653]  = \[646]  & ~\$$COND0<0>5.1 ,
  \[843]  = \D<17>  | \C<17> ,
  \[464]  = \new_C<68> ,
  \new_C<15>  = (\[647]  & (\D<15>  & \C<15> )) | ((\[848]  & \[653] ) | ((~\[847]  & \[649] ) | ((\[847]  & \[650] ) | ((\[654]  & \key<58> ) | (\[651]  & \key<1> ))))),
  \[654]  = \start<0>  & \encrypt<0> ,
  \[844]  = (~\D<17>  & \C<17> ) | (\D<17>  & ~\C<17> ),
  \[465]  = \new_C<67> ,
  \new_C<16>  = (\[647]  & (\D<16>  & \C<16> )) | ((\[846]  & \[653] ) | ((~\[845]  & \[649] ) | ((\[845]  & \[650] ) | ((\[654]  & \key<50> ) | (\[651]  & \key<58> ))))),
  \[655]  = \D<111>  | \C<111> ,
  \[845]  = \D<16>  | \C<16> ,
  \[466]  = \new_C<66> ,
  \new_C<17>  = (\[647]  & (\D<17>  & \C<17> )) | ((\[844]  & \[653] ) | ((~\[843]  & \[649] ) | ((\[843]  & \[650] ) | ((\[654]  & \key<42> ) | (\[651]  & \key<50> ))))),
  \[656]  = (~\D<111>  & \C<111> ) | (\D<111>  & ~\C<111> ),
  \[846]  = (~\D<16>  & \C<16> ) | (\D<16>  & ~\C<16> ),
  \[467]  = \new_C<65> ,
  \new_C<18>  = (\[647]  & (\D<18>  & \C<18> )) | ((\[842]  & \[653] ) | ((~\[841]  & \[649] ) | ((\[841]  & \[650] ) | ((\[654]  & \key<34> ) | (\[651]  & \key<42> ))))),
  \[657]  = \D<110>  | \C<110> ,
  \[847]  = \D<15>  | \C<15> ,
  \[468]  = \new_C<64> ,
  \new_C<11>  = (\[647]  & (\D<11>  & \C<11> )) | ((\[856]  & \[653] ) | ((~\[855]  & \[649] ) | ((\[855]  & \[650] ) | ((\[654]  & \key<25> ) | (\[651]  & \key<33> ))))),
  \[658]  = (~\D<110>  & \C<110> ) | (\D<110>  & ~\C<110> ),
  \[848]  = (~\D<15>  & \C<15> ) | (\D<15>  & ~\C<15> ),
  \[469]  = \new_C<63> ,
  \new_C<12>  = (\[647]  & (\D<12>  & \C<12> )) | ((\[854]  & \[653] ) | ((~\[853]  & \[649] ) | ((\[853]  & \[650] ) | ((\[654]  & \key<17> ) | (\[651]  & \key<25> ))))),
  \[659]  = \D<109>  | \C<109> ,
  \[849]  = \D<14>  | \C<14> ,
  \new_C<13>  = (\[647]  & (\D<13>  & \C<13> )) | ((\[852]  & \[653] ) | ((~\[851]  & \[649] ) | ((\[851]  & \[650] ) | ((\[654]  & \key<9> ) | (\[651]  & \key<17> ))))),
  \new_C<14>  = (\[647]  & (\D<14>  & \C<14> )) | ((\[850]  & \[653] ) | ((~\[849]  & \[649] ) | ((\[849]  & \[650] ) | ((\[654]  & \key<1> ) | (\[651]  & \key<9> ))))),
  \$$COND0<0>5.1  = (\[880]  & (~\count<0>  & \count<3> )) | ((\[880]  & (\count<0>  & ~\count<3> )) | (\$$COND1<0>8.1  & (~\count<0>  & ~\count<3> ))),
  \new_C<10>  = (\[647]  & (\D<10>  & \C<10> )) | ((\[858]  & \[653] ) | ((~\[857]  & \[649] ) | ((\[857]  & \[650] ) | ((\[654]  & \key<33> ) | (\[651]  & \key<41> ))))),
  \[470]  = \new_C<62> ,
  \new_C<29>  = (\[647]  & (\D<29>  & \C<29> )) | ((\[820]  & \[653] ) | ((~\[819]  & \[649] ) | ((\[819]  & \[650] ) | ((\[654]  & \key<104> ) | (\[651]  & \key<112> ))))),
  \[660]  = (~\D<109>  & \C<109> ) | (\D<109>  & ~\C<109> ),
  \[850]  = (~\D<14>  & \C<14> ) | (\D<14>  & ~\C<14> ),
  \[471]  = \new_C<61> ,
  \[661]  = \D<108>  | \C<108> ,
  \[851]  = \D<13>  | \C<13> ,
  \[472]  = \new_C<60> ,
  \[662]  = (~\D<108>  & \C<108> ) | (\D<108>  & ~\C<108> ),
  \[852]  = (~\D<13>  & \C<13> ) | (\D<13>  & ~\C<13> ),
  \[473]  = \new_C<59> ,
  \[663]  = \D<107>  | \C<107> ,
  \[853]  = \D<12>  | \C<12> ,
  \[474]  = \new_C<58> ,
  \new_C<25>  = (\[647]  & (\D<25>  & \C<25> )) | ((\[828]  & \[653] ) | ((~\[827]  & \[649] ) | ((\[827]  & \[650] ) | ((\[654]  & \key<43> ) | (\[651]  & \key<51> ))))),
  \[664]  = (~\D<107>  & \C<107> ) | (\D<107>  & ~\C<107> ),
  \[854]  = (~\D<12>  & \C<12> ) | (\D<12>  & ~\C<12> ),
  \[475]  = \new_C<57> ,
  \new_C<26>  = (\[647]  & (\D<26>  & \C<26> )) | ((\[826]  & \[653] ) | ((~\[825]  & \[649] ) | ((\[825]  & \[650] ) | ((\[654]  & \key<35> ) | (\[651]  & \key<43> ))))),
  \[665]  = \D<106>  | \C<106> ,
  \[855]  = \D<11>  | \C<11> ,
  \[476]  = \new_C<56> ,
  \new_C<27>  = (\[647]  & (\D<27>  & \C<27> )) | ((\[824]  & \[653] ) | ((~\[823]  & \[649] ) | ((\[823]  & \[650] ) | ((\[654]  & \key<120> ) | (\[651]  & \key<35> ))))),
  \[666]  = (~\D<106>  & \C<106> ) | (\D<106>  & ~\C<106> ),
  \[856]  = (~\D<11>  & \C<11> ) | (\D<11>  & ~\C<11> ),
  \[477]  = \new_C<55> ,
  \new_C<28>  = (\[647]  & (\D<28>  & \C<28> )) | ((\[822]  & \[653] ) | ((~\[821]  & \[649] ) | ((\[821]  & \[650] ) | ((\[654]  & \key<112> ) | (\[651]  & \key<120> ))))),
  \[667]  = \D<105>  | \C<105> ,
  \[857]  = \D<10>  | \C<10> ,
  \[478]  = \new_C<54> ,
  \new_C<21>  = (\[647]  & (\D<21>  & \C<21> )) | ((\[836]  & \[653] ) | ((~\[835]  & \[649] ) | ((\[835]  & \[650] ) | ((\[654]  & \key<10> ) | (\[651]  & \key<18> ))))),
  \[668]  = (~\D<105>  & \C<105> ) | (\D<105>  & ~\C<105> ),
  \[858]  = (~\D<10>  & \C<10> ) | (\D<10>  & ~\C<10> ),
  \[479]  = \new_C<53> ,
  \new_C<22>  = (\[647]  & (\D<22>  & \C<22> )) | ((\[834]  & \[653] ) | ((~\[833]  & \[649] ) | ((\[833]  & \[650] ) | ((\[654]  & \key<2> ) | (\[651]  & \key<10> ))))),
  \[669]  = \D<104>  | \C<104> ,
  \[859]  = \D<9>  | \C<9> ,
  \new_C<23>  = (\[647]  & (\D<23>  & \C<23> )) | ((\[832]  & \[653] ) | ((~\[831]  & \[649] ) | ((\[831]  & \[650] ) | ((\[654]  & \key<59> ) | (\[651]  & \key<2> ))))),
  \new_C<24>  = (\[647]  & (\D<24>  & \C<24> )) | ((\[830]  & \[653] ) | ((~\[829]  & \[649] ) | ((\[829]  & \[650] ) | ((\[654]  & \key<51> ) | (\[651]  & \key<59> ))))),
  \new_C<20>  = (\[647]  & (\D<20>  & \C<20> )) | ((\[838]  & \[653] ) | ((~\[837]  & \[649] ) | ((\[837]  & \[650] ) | ((\[654]  & \key<18> ) | (\[651]  & \key<26> ))))),
  \[480]  = \new_C<52> ,
  \new_C<39>  = (\[647]  & (\D<39>  & \C<39> )) | ((\[800]  & \[653] ) | ((~\[799]  & \[649] ) | ((\[799]  & \[650] ) | ((\[654]  & \key<89> ) | (\[651]  & \key<97> ))))),
  \[670]  = (~\D<104>  & \C<104> ) | (\D<104>  & ~\C<104> ),
  \[860]  = (~\D<9>  & \C<9> ) | (\D<9>  & ~\C<9> ),
  \[481]  = \new_C<51> ,
  \[671]  = \D<103>  | \C<103> ,
  \[861]  = \D<8>  | \C<8> ,
  \[482]  = \new_C<50> ,
  \[672]  = (~\D<103>  & \C<103> ) | (\D<103>  & ~\C<103> ),
  \[862]  = (~\D<8>  & \C<8> ) | (\D<8>  & ~\C<8> ),
  \[483]  = \new_C<49> ,
  \[673]  = \D<102>  | \C<102> ,
  \[863]  = \D<7>  | \C<7> ,
  \[484]  = \new_C<48> ,
  \new_C<35>  = (\[647]  & (\D<35>  & \C<35> )) | ((\[808]  & \[653] ) | ((~\[807]  & \[649] ) | ((\[807]  & \[650] ) | ((\[654]  & \key<121> ) | (\[651]  & \key<64> ))))),
  \[674]  = (~\D<102>  & \C<102> ) | (\D<102>  & ~\C<102> ),
  \[864]  = (~\D<7>  & \C<7> ) | (\D<7>  & ~\C<7> ),
  \[485]  = \new_C<47> ,
  \new_C<36>  = (\[647]  & (\D<36>  & \C<36> )) | ((\[806]  & \[653] ) | ((~\[805]  & \[649] ) | ((\[805]  & \[650] ) | ((\[654]  & \key<113> ) | (\[651]  & \key<121> ))))),
  \[675]  = \D<101>  | \C<101> ,
  \[865]  = \D<6>  | \C<6> ,
  \[486]  = \new_C<46> ,
  \new_C<37>  = (\[647]  & (\D<37>  & \C<37> )) | ((\[804]  & \[653] ) | ((~\[803]  & \[649] ) | ((\[803]  & \[650] ) | ((\[654]  & \key<105> ) | (\[651]  & \key<113> ))))),
  \[676]  = (~\D<101>  & \C<101> ) | (\D<101>  & ~\C<101> ),
  \[866]  = (~\D<6>  & \C<6> ) | (\D<6>  & ~\C<6> ),
  \[487]  = \new_C<45> ,
  \new_C<38>  = (\[647]  & (\D<38>  & \C<38> )) | ((\[802]  & \[653] ) | ((~\[801]  & \[649] ) | ((\[801]  & \[650] ) | ((\[654]  & \key<97> ) | (\[651]  & \key<105> ))))),
  \[677]  = \D<100>  | \C<100> ,
  \[867]  = \D<5>  | \C<5> ,
  \[488]  = \new_C<44> ,
  \new_C<31>  = (\[647]  & (\D<31>  & \C<31> )) | ((\[816]  & \[653] ) | ((~\[815]  & \[649] ) | ((\[815]  & \[650] ) | ((\[654]  & \key<88> ) | (\[651]  & \key<96> ))))),
  \[678]  = (~\D<100>  & \C<100> ) | (\D<100>  & ~\C<100> ),
  \[868]  = (~\D<5>  & \C<5> ) | (\D<5>  & ~\C<5> ),
  \[489]  = \new_C<43> ,
  \new_C<32>  = (\[647]  & (\D<32>  & \C<32> )) | ((\[814]  & \[653] ) | ((~\[813]  & \[649] ) | ((\[813]  & \[650] ) | ((\[654]  & \key<80> ) | (\[651]  & \key<88> ))))),
  \[679]  = \D<99>  | \C<99> ,
  \[869]  = \D<4>  | \C<4> ,
  \new_C<33>  = (\[647]  & (\D<33>  & \C<33> )) | ((\[812]  & \[653] ) | ((~\[811]  & \[649] ) | ((\[811]  & \[650] ) | ((\[654]  & \key<72> ) | (\[651]  & \key<80> ))))),
  \new_C<34>  = (\[647]  & (\D<34>  & \C<34> )) | ((\[810]  & \[653] ) | ((~\[809]  & \[649] ) | ((\[809]  & \[650] ) | ((\[654]  & \key<64> ) | (\[651]  & \key<72> ))))),
  \new_C<30>  = (\[647]  & (\D<30>  & \C<30> )) | ((\[818]  & \[653] ) | ((~\[817]  & \[649] ) | ((\[817]  & \[650] ) | ((\[654]  & \key<96> ) | (\[651]  & \key<104> ))))),
  \[490]  = \new_C<42> ,
  \new_C<49>  = (\[647]  & (\D<49>  & \C<49> )) | ((\[780]  & \[653] ) | ((~\[779]  & \[649] ) | ((\[779]  & \[650] ) | ((\[654]  & \key<74> ) | (\[651]  & \key<82> ))))),
  \[680]  = (~\D<99>  & \C<99> ) | (\D<99>  & ~\C<99> ),
  \[870]  = (~\D<4>  & \C<4> ) | (\D<4>  & ~\C<4> ),
  \[491]  = \new_C<41> ,
  \[681]  = \D<98>  | \C<98> ,
  \[871]  = \D<3>  | \C<3> ,
  \[492]  = \new_C<40> ,
  \[682]  = (~\D<98>  & \C<98> ) | (\D<98>  & ~\C<98> ),
  \[872]  = (~\D<3>  & \C<3> ) | (\D<3>  & ~\C<3> ),
  \[493]  = \new_C<39> ,
  \[683]  = \D<97>  | \C<97> ,
  \[873]  = \D<2>  | \C<2> ,
  \[494]  = \new_C<38> ,
  \new_C<45>  = (\[647]  & (\D<45>  & \C<45> )) | ((\[788]  & \[653] ) | ((~\[787]  & \[649] ) | ((\[787]  & \[650] ) | ((\[654]  & \key<106> ) | (\[651]  & \key<114> ))))),
  \[684]  = (~\D<97>  & \C<97> ) | (\D<97>  & ~\C<97> ),
  \[874]  = (~\D<2>  & \C<2> ) | (\D<2>  & ~\C<2> ),
  \[495]  = \new_C<37> ,
  \new_C<46>  = (\[647]  & (\D<46>  & \C<46> )) | ((\[786]  & \[653] ) | ((~\[785]  & \[649] ) | ((\[785]  & \[650] ) | ((\[654]  & \key<98> ) | (\[651]  & \key<106> ))))),
  \[685]  = \D<96>  | \C<96> ,
  \[875]  = \D<1>  | \C<1> ,
  \[496]  = \new_C<36> ,
  \new_C<47>  = (\[647]  & (\D<47>  & \C<47> )) | ((\[784]  & \[653] ) | ((~\[783]  & \[649] ) | ((\[783]  & \[650] ) | ((\[654]  & \key<90> ) | (\[651]  & \key<98> ))))),
  \[686]  = (~\D<96>  & \C<96> ) | (\D<96>  & ~\C<96> ),
  \[876]  = (~\D<1>  & \C<1> ) | (\D<1>  & ~\C<1> ),
  \[497]  = \new_C<35> ,
  \new_C<48>  = (\[647]  & (\D<48>  & \C<48> )) | ((\[782]  & \[653] ) | ((~\[781]  & \[649] ) | ((\[781]  & \[650] ) | ((\[654]  & \key<82> ) | (\[651]  & \key<90> ))))),
  \[687]  = \D<95>  | \C<95> ,
  \[877]  = \D<0>  | \C<0> ,
  \[498]  = \new_C<34> ,
  \new_C<41>  = (\[647]  & (\D<41>  & \C<41> )) | ((\[796]  & \[653] ) | ((~\[795]  & \[649] ) | ((\[795]  & \[650] ) | ((\[654]  & \key<73> ) | (\[651]  & \key<81> ))))),
  \[688]  = (~\D<95>  & \C<95> ) | (\D<95>  & ~\C<95> ),
  \[878]  = (~\D<0>  & \C<0> ) | (\D<0>  & ~\C<0> ),
  \[499]  = \new_C<33> ,
  \new_C<42>  = (\[647]  & (\D<42>  & \C<42> )) | ((\[794]  & \[653] ) | ((~\[793]  & \[649] ) | ((\[793]  & \[650] ) | ((\[654]  & \key<65> ) | (\[651]  & \key<73> ))))),
  \[689]  = \D<94>  | \C<94> ,
  \[879]  = ~\count<0>  | ~\count<3> ,
  \new_count<0>  = \[227] ,
  \new_C<43>  = (\[647]  & (\D<43>  & \C<43> )) | ((\[792]  & \[653] ) | ((~\[791]  & \[649] ) | ((\[791]  & \[650] ) | ((\[654]  & \key<122> ) | (\[651]  & \key<65> ))))),
  \new_C<44>  = (\[647]  & (\D<44>  & \C<44> )) | ((\[790]  & \[653] ) | ((~\[789]  & \[649] ) | ((\[789]  & \[650] ) | ((\[654]  & \key<114> ) | (\[651]  & \key<122> ))))),
  \new_count<3>  = \[224] ,
  \new_count<1>  = \[226] ,
  \new_C<40>  = (\[647]  & (\D<40>  & \C<40> )) | ((\[798]  & \[653] ) | ((~\[797]  & \[649] ) | ((\[797]  & \[650] ) | ((\[654]  & \key<81> ) | (\[651]  & \key<89> ))))),
  \new_count<2>  = \[225] ,
  \[690]  = (~\D<94>  & \C<94> ) | (\D<94>  & ~\C<94> ),
  \[880]  = \count<1>  & \count<2> ,
  \[691]  = \D<93>  | \C<93> ,
  \[692]  = (~\D<93>  & \C<93> ) | (\D<93>  & ~\C<93> ),
  \[882]  = \[227]  & \start<0> ,
  \[693]  = \D<92>  | \C<92> ,
  \[694]  = (~\D<92>  & \C<92> ) | (\D<92>  & ~\C<92> ),
  \[695]  = \D<91>  | \C<91> ,
  \[696]  = (~\D<91>  & \C<91> ) | (\D<91>  & ~\C<91> ),
  \[697]  = \D<90>  | \C<90> ,
  \[698]  = (~\D<90>  & \C<90> ) | (\D<90>  & ~\C<90> ),
  \[699]  = \D<89>  | \C<89> ,
  \KSi<12>  = \C<22> ,
  \KSi<11>  = \C<9> ,
  \KSi<14>  = \C<11> ,
  \KSi<13>  = \C<18> ,
  \KSi<10>  = \C<20> ,
  \KSi<19>  = \C<6> ,
  \KSi<16>  = \C<25> ,
  \KSi<15>  = \C<3> ,
  \KSi<18>  = \C<15> ,
  \KSi<17>  = \C<7> ,
  \KSi<22>  = \C<12> ,
  \KSi<21>  = \C<19> ,
  \KSi<24>  = \C<41> ,
  \KSi<23>  = \C<1> ,
  \KSi<20>  = \C<26> ,
  \KSi<29>  = \C<32> ,
  \KSi<26>  = \C<38> ,
  \KSi<25>  = \C<44> ,
  \KSi<28>  = \C<28> ,
  \KSi<27>  = \C<51> ,
  \KSi<32>  = \C<42> ,
  \KSi<31>  = \C<55> ,
  \KSi<34>  = \C<48> ,
  \KSi<33>  = \C<33> ,
  \KSi<30>  = \C<30> ,
  \KSi<39>  = \C<31> ,
  \KSi<36>  = \C<50> ,
  \KSi<35>  = \C<37> ,
  \KSi<38>  = \C<39> ,
  \KSi<37>  = \C<46> ,
  \KSi<42>  = \C<43> ,
  \KSi<41>  = \C<35> ,
  \KSi<44>  = \C<54> ,
  \KSi<43>  = \C<34> ,
  \new_C<99>  = (\[647]  & (\D<99>  & \C<99> )) | ((\[680]  & \[653] ) | ((~\[679]  & \[649] ) | ((\[679]  & \[650] ) | ((\[654]  & \key<250> ) | (\[651]  & \key<193> ))))),
  \new_D<19>  = (\[648]  & (\D<19>  & \C<19> )) | ((\[840]  & \[652] ) | ((~\[839]  & \[650] ) | ((\[839]  & \[649] ) | ((\[654]  & \key<28> ) | (\[651]  & \key<36> ))))),
  \KSi<40>  = \C<53> ,
  \new_C<95>  = (\[647]  & (\D<95>  & \C<95> )) | ((\[688]  & \[653] ) | ((~\[687]  & \[649] ) | ((\[687]  & \[650] ) | ((\[654]  & \key<217> ) | (\[651]  & \key<225> ))))),
  \KSi<49>  = \C<72> ,
  \new_C<96>  = (\[647]  & (\D<96>  & \C<96> )) | ((\[686]  & \[653] ) | ((~\[685]  & \[649] ) | ((\[685]  & \[650] ) | ((\[654]  & \key<209> ) | (\[651]  & \key<217> ))))),
  \new_D<15>  = (\[648]  & (\D<15>  & \C<15> )) | ((\[848]  & \[652] ) | ((~\[847]  & \[650] ) | ((\[847]  & \[649] ) | ((\[654]  & \key<60> ) | (\[651]  & \key<5> ))))),
  \new_C<97>  = (\[647]  & (\D<97>  & \C<97> )) | ((\[684]  & \[653] ) | ((~\[683]  & \[649] ) | ((\[683]  & \[650] ) | ((\[654]  & \key<201> ) | (\[651]  & \key<209> ))))),
  \new_D<16>  = (\[648]  & (\D<16>  & \C<16> )) | ((\[846]  & \[652] ) | ((~\[845]  & \[650] ) | ((\[845]  & \[649] ) | ((\[654]  & \key<52> ) | (\[651]  & \key<60> ))))),
  \new_C<98>  = (\[647]  & (\D<98>  & \C<98> )) | ((\[682]  & \[653] ) | ((~\[681]  & \[649] ) | ((\[681]  & \[650] ) | ((\[654]  & \key<193> ) | (\[651]  & \key<201> ))))),
  \new_D<17>  = (\[648]  & (\D<17>  & \C<17> )) | ((\[844]  & \[652] ) | ((~\[843]  & \[650] ) | ((\[843]  & \[649] ) | ((\[654]  & \key<44> ) | (\[651]  & \key<52> ))))),
  \KSi<46>  = \C<40> ,
  \new_C<91>  = (\[647]  & (\D<91>  & \C<91> )) | ((\[696]  & \[653] ) | ((~\[695]  & \[649] ) | ((\[695]  & \[650] ) | ((\[654]  & \key<249> ) | (\[651]  & \key<192> ))))),
  \new_D<18>  = (\[648]  & (\D<18>  & \C<18> )) | ((\[842]  & \[652] ) | ((~\[841]  & \[650] ) | ((\[841]  & \[649] ) | ((\[654]  & \key<36> ) | (\[651]  & \key<44> ))))),
  \KSi<45>  = \C<47> ,
  \new_C<92>  = (\[647]  & (\D<92>  & \C<92> )) | ((\[694]  & \[653] ) | ((~\[693]  & \[649] ) | ((\[693]  & \[650] ) | ((\[654]  & \key<241> ) | (\[651]  & \key<249> ))))),
  \new_D<11>  = (\[648]  & (\D<11>  & \C<11> )) | ((\[856]  & \[652] ) | ((~\[855]  & \[650] ) | ((\[855]  & \[649] ) | ((\[654]  & \key<29> ) | (\[651]  & \key<37> ))))),
  \KSi<48>  = \C<69> ,
  \new_C<93>  = (\[647]  & (\D<93>  & \C<93> )) | ((\[692]  & \[653] ) | ((~\[691]  & \[649] ) | ((\[691]  & \[650] ) | ((\[654]  & \key<233> ) | (\[651]  & \key<241> ))))),
  \new_D<12>  = (\[648]  & (\D<12>  & \C<12> )) | ((\[854]  & \[652] ) | ((~\[853]  & \[650] ) | ((\[853]  & \[649] ) | ((\[654]  & \key<21> ) | (\[651]  & \key<29> ))))),
  \KSi<47>  = \C<29> ,
  \new_C<94>  = (\[647]  & (\D<94>  & \C<94> )) | ((\[690]  & \[653] ) | ((~\[689]  & \[649] ) | ((\[689]  & \[650] ) | ((\[654]  & \key<225> ) | (\[651]  & \key<233> ))))),
  \new_D<13>  = (\[648]  & (\D<13>  & \C<13> )) | ((\[852]  & \[652] ) | ((~\[851]  & \[650] ) | ((\[851]  & \[649] ) | ((\[654]  & \key<13> ) | (\[651]  & \key<21> ))))),
  \KSi<52>  = \C<56> ,
  \new_D<14>  = (\[648]  & (\D<14>  & \C<14> )) | ((\[850]  & \[652] ) | ((~\[849]  & \[650] ) | ((\[849]  & \[649] ) | ((\[654]  & \key<5> ) | (\[651]  & \key<13> ))))),
  \KSi<51>  = \C<79> ,
  \KSi<54>  = \C<58> ,
  \KSi<53>  = \C<60> ,
  \new_C<90>  = (\[647]  & (\D<90>  & \C<90> )) | ((\[698]  & \[653] ) | ((~\[697]  & \[649] ) | ((\[697]  & \[650] ) | ((\[654]  & \key<192> ) | (\[651]  & \key<200> ))))),
  \new_D<10>  = (\[648]  & (\D<10>  & \C<10> )) | ((\[858]  & \[652] ) | ((~\[857]  & \[650] ) | ((\[857]  & \[649] ) | ((\[654]  & \key<37> ) | (\[651]  & \key<45> ))))),
  \new_D<29>  = (\[648]  & (\D<29>  & \C<29> )) | ((\[820]  & \[652] ) | ((~\[819]  & \[650] ) | ((\[819]  & \[649] ) | ((\[654]  & \key<110> ) | (\[651]  & \key<118> ))))),
  \KSi<50>  = \C<66> ,
  \KSi<59>  = \C<65> ,
  \new_D<25>  = (\[648]  & (\D<25>  & \C<25> )) | ((\[828]  & \[652] ) | ((~\[827]  & \[650] ) | ((\[827]  & \[649] ) | ((\[654]  & \key<11> ) | (\[651]  & \key<19> ))))),
  \new_D<26>  = (\[648]  & (\D<26>  & \C<26> )) | ((\[826]  & \[652] ) | ((~\[825]  & \[650] ) | ((\[825]  & \[649] ) | ((\[654]  & \key<3> ) | (\[651]  & \key<11> ))))),
  \new_D<27>  = (\[648]  & (\D<27>  & \C<27> )) | ((\[824]  & \[652] ) | ((~\[823]  & \[650] ) | ((\[823]  & \[649] ) | ((\[654]  & \key<126> ) | (\[651]  & \key<3> ))))),
  \KSi<56>  = \C<70> ,
  \new_D<28>  = (\[648]  & (\D<28>  & \C<28> )) | ((\[822]  & \[652] ) | ((~\[821]  & \[650] ) | ((\[821]  & \[649] ) | ((\[654]  & \key<118> ) | (\[651]  & \key<126> ))))),
  \KSi<55>  = \C<83> ,
  \new_D<21>  = (\[648]  & (\D<21>  & \C<21> )) | ((\[836]  & \[652] ) | ((~\[835]  & \[650] ) | ((\[835]  & \[649] ) | ((\[654]  & \key<12> ) | (\[651]  & \key<20> ))))),
  \KSi<58>  = \C<76> ,
  \new_D<22>  = (\[648]  & (\D<22>  & \C<22> )) | ((\[834]  & \[652] ) | ((~\[833]  & \[650] ) | ((\[833]  & \[649] ) | ((\[654]  & \key<4> ) | (\[651]  & \key<12> ))))),
  \KSi<57>  = \C<61> ,
  \new_D<23>  = (\[648]  & (\D<23>  & \C<23> )) | ((\[832]  & \[652] ) | ((~\[831]  & \[650] ) | ((\[831]  & \[649] ) | ((\[654]  & \key<27> ) | (\[651]  & \key<4> ))))),
  \KSi<62>  = \C<67> ,
  \new_D<24>  = (\[648]  & (\D<24>  & \C<24> )) | ((\[830]  & \[652] ) | ((~\[829]  & \[650] ) | ((\[829]  & \[649] ) | ((\[654]  & \key<19> ) | (\[651]  & \key<27> ))))),
  \KSi<61>  = \C<74> ,
  \KSi<64>  = \C<81> ,
  \KSi<63>  = \C<59> ,
  \[500]  = \new_C<32> ,
  \new_D<20>  = (\[648]  & (\D<20>  & \C<20> )) | ((\[838]  & \[652] ) | ((~\[837]  & \[650] ) | ((\[837]  & \[649] ) | ((\[654]  & \key<20> ) | (\[651]  & \key<28> ))))),
  \[501]  = \new_C<31> ,
  \new_D<39>  = (\[648]  & (\D<39>  & \C<39> )) | ((\[800]  & \[652] ) | ((~\[799]  & \[650] ) | ((\[799]  & \[649] ) | ((\[654]  & \key<93> ) | (\[651]  & \key<101> ))))),
  \KSi<60>  = \C<78> ,
  \[502]  = \new_C<30> ,
  \[503]  = \new_C<29> ,
  \[504]  = \new_C<28> ,
  \KSi<69>  = \C<75> ,
  \[505]  = \new_C<27> ,
  \new_D<35>  = (\[648]  & (\D<35>  & \C<35> )) | ((\[808]  & \[652] ) | ((~\[807]  & \[650] ) | ((\[807]  & \[649] ) | ((\[654]  & \key<125> ) | (\[651]  & \key<70> ))))),
  \[506]  = \new_C<26> ,
  \new_D<36>  = (\[648]  & (\D<36>  & \C<36> )) | ((\[806]  & \[652] ) | ((~\[805]  & \[650] ) | ((\[805]  & \[649] ) | ((\[654]  & \key<117> ) | (\[651]  & \key<125> ))))),
  \[507]  = \new_C<25> ,
  \new_D<37>  = (\[648]  & (\D<37>  & \C<37> )) | ((\[804]  & \[652] ) | ((~\[803]  & \[650] ) | ((\[803]  & \[649] ) | ((\[654]  & \key<109> ) | (\[651]  & \key<117> ))))),
  \KSi<66>  = \C<71> ,
  \[508]  = \new_C<24> ,
  \data_ready<0>  = \[228] ,
  \new_D<38>  = (\[648]  & (\D<38>  & \C<38> )) | ((\[802]  & \[652] ) | ((~\[801]  & \[650] ) | ((\[801]  & \[649] ) | ((\[654]  & \key<101> ) | (\[651]  & \key<109> ))))),
  \KSi<65>  = \C<63> ,
  \[509]  = \new_C<23> ,
  \new_D<31>  = (\[648]  & (\D<31>  & \C<31> )) | ((\[816]  & \[652] ) | ((~\[815]  & \[650] ) | ((\[815]  & \[649] ) | ((\[654]  & \key<94> ) | (\[651]  & \key<102> ))))),
  \KSi<68>  = \C<82> ,
  \new_D<32>  = (\[648]  & (\D<32>  & \C<32> )) | ((\[814]  & \[652] ) | ((~\[813]  & \[650] ) | ((\[813]  & \[649] ) | ((\[654]  & \key<86> ) | (\[651]  & \key<94> ))))),
  \KSi<67>  = \C<62> ,
  \new_D<33>  = (\[648]  & (\D<33>  & \C<33> )) | ((\[812]  & \[652] ) | ((~\[811]  & \[650] ) | ((\[811]  & \[649] ) | ((\[654]  & \key<78> ) | (\[651]  & \key<86> ))))),
  \KSi<72>  = \C<97> ,
  \new_D<34>  = (\[648]  & (\D<34>  & \C<34> )) | ((\[810]  & \[652] ) | ((~\[809]  & \[650] ) | ((\[809]  & \[649] ) | ((\[654]  & \key<70> ) | (\[651]  & \key<78> ))))),
  \KSi<71>  = \C<57> ,
  \KSi<74>  = \C<94> ,
  \KSi<73>  = \C<100> ,
  \[510]  = \new_C<22> ,
  \[700]  = (~\D<89>  & \C<89> ) | (\D<89>  & ~\C<89> ),
  \new_D<30>  = (\[648]  & (\D<30>  & \C<30> )) | ((\[818]  & \[652] ) | ((~\[817]  & \[650] ) | ((\[817]  & \[649] ) | ((\[654]  & \key<102> ) | (\[651]  & \key<110> ))))),
  \[511]  = \new_C<21> ,
  \[701]  = \D<88>  | \C<88> ,
  \new_D<49>  = (\[648]  & (\D<49>  & \C<49> )) | ((\[780]  & \[652] ) | ((~\[779]  & \[650] ) | ((\[779]  & \[649] ) | ((\[654]  & \key<76> ) | (\[651]  & \key<84> ))))),
  \KSi<70>  = \C<68> ,
  \[512]  = \new_C<20> ,
  \[702]  = (~\D<88>  & \C<88> ) | (\D<88>  & ~\C<88> ),
  \[513]  = \new_C<19> ,
  \[703]  = \D<87>  | \C<87> ,
  \[514]  = \new_C<18> ,
  \[704]  = (~\D<87>  & \C<87> ) | (\D<87>  & ~\C<87> ),
  \KSi<79>  = \C<111> ,
  \[515]  = \new_C<17> ,
  \[705]  = \D<86>  | \C<86> ,
  \new_D<45>  = (\[648]  & (\D<45>  & \C<45> )) | ((\[788]  & \[652] ) | ((~\[787]  & \[650] ) | ((\[787]  & \[649] ) | ((\[654]  & \key<44> ) | (\[651]  & \key<116> ))))),
  \[516]  = \new_C<16> ,
  \[706]  = (~\D<86>  & \C<86> ) | (\D<86>  & ~\C<86> ),
  \new_C<1>  = (\[647]  & (\D<1>  & \C<1> )) | ((\[876]  & \[653] ) | ((~\[875]  & \[649] ) | ((\[875]  & \[650] ) | ((\[654]  & \key<40> ) | (\[651]  & \key<48> ))))),
  \new_D<46>  = (\[648]  & (\D<46>  & \C<46> )) | ((\[786]  & \[652] ) | ((~\[785]  & \[650] ) | ((\[785]  & \[649] ) | ((\[654]  & \key<100> ) | (\[651]  & \key<44> ))))),
  \[517]  = \new_C<15> ,
  \[707]  = \D<85>  | \C<85> ,
  \new_C<2>  = (\[647]  & (\D<2>  & \C<2> )) | ((\[874]  & \[653] ) | ((~\[873]  & \[649] ) | ((\[873]  & \[650] ) | ((\[654]  & \key<32> ) | (\[651]  & \key<40> ))))),
  \new_D<47>  = (\[648]  & (\D<47>  & \C<47> )) | ((\[784]  & \[652] ) | ((~\[783]  & \[650] ) | ((\[783]  & \[649] ) | ((\[654]  & \key<92> ) | (\[651]  & \key<100> ))))),
  \KSi<76>  = \C<84> ,
  \[518]  = \new_C<14> ,
  \[708]  = (~\D<85>  & \C<85> ) | (\D<85>  & ~\C<85> ),
  \new_C<3>  = (\[647]  & (\D<3>  & \C<3> )) | ((\[872]  & \[653] ) | ((~\[871]  & \[649] ) | ((\[871]  & \[650] ) | ((\[654]  & \key<24> ) | (\[651]  & \key<32> ))))),
  \new_D<48>  = (\[648]  & (\D<48>  & \C<48> )) | ((\[782]  & \[652] ) | ((~\[781]  & \[650] ) | ((\[781]  & \[649] ) | ((\[654]  & \key<84> ) | (\[651]  & \key<92> ))))),
  \KSi<75>  = \C<107> ,
  \[519]  = \new_C<13> ,
  \[709]  = \D<84>  | \C<84> ,
  \new_C<4>  = (\[647]  & (\D<4>  & \C<4> )) | ((\[870]  & \[653] ) | ((~\[869]  & \[649] ) | ((\[869]  & \[650] ) | ((\[654]  & \key<16> ) | (\[651]  & \key<24> ))))),
  \new_D<41>  = (\[648]  & (\D<41>  & \C<41> )) | ((\[796]  & \[652] ) | ((~\[795]  & \[650] ) | ((\[795]  & \[649] ) | ((\[654]  & \key<77> ) | (\[651]  & \key<85> ))))),
  \KSi<78>  = \C<86> ,
  \new_D<42>  = (\[648]  & (\D<42>  & \C<42> )) | ((\[794]  & \[652] ) | ((~\[793]  & \[650] ) | ((\[793]  & \[649] ) | ((\[654]  & \key<69> ) | (\[651]  & \key<77> ))))),
  \KSi<77>  = \C<88> ,
  \new_D<43>  = (\[648]  & (\D<43>  & \C<43> )) | ((\[792]  & \[652] ) | ((~\[791]  & \[650] ) | ((\[791]  & \[649] ) | ((\[654]  & \key<124> ) | (\[651]  & \key<69> ))))),
  \KSi<82>  = \C<104> ,
  \new_D<44>  = (\[648]  & (\D<44>  & \C<44> )) | ((\[790]  & \[652] ) | ((~\[789]  & \[650] ) | ((\[789]  & \[649] ) | ((\[654]  & \key<116> ) | (\[651]  & \key<124> ))))),
  \KSi<81>  = \C<89> ,
  \new_C<0>  = (\[647]  & (\D<0>  & \C<0> )) | ((\[878]  & \[653] ) | ((~\[877]  & \[649] ) | ((\[877]  & \[650] ) | ((\[654]  & \key<48> ) | (\[651]  & \key<56> ))))),
  \KSi<84>  = \C<106> ,
  \new_C<9>  = (\[647]  & (\D<9>  & \C<9> )) | ((\[860]  & \[653] ) | ((~\[859]  & \[649] ) | ((\[859]  & \[650] ) | ((\[654]  & \key<41> ) | (\[651]  & \key<49> ))))),
  \KSi<83>  = \C<93> ,
  \[520]  = \new_C<12> ,
  \new_C<59>  = (\[647]  & (\D<59>  & \C<59> )) | ((\[760]  & \[653] ) | ((~\[759]  & \[649] ) | ((\[759]  & \[650] ) | ((\[654]  & \key<152> ) | (\[651]  & \key<160> ))))),
  \[710]  = (~\D<84>  & \C<84> ) | (\D<84>  & ~\C<84> ),
  \new_D<40>  = (\[648]  & (\D<40>  & \C<40> )) | ((\[798]  & \[652] ) | ((~\[797]  & \[650] ) | ((\[797]  & \[649] ) | ((\[654]  & \key<85> ) | (\[651]  & \key<93> ))))),
  \[521]  = \new_C<11> ,
  \[711]  = \D<83>  | \C<83> ,
  \KSi<80>  = \C<98> ,
  \[522]  = \new_C<10> ,
  \[712]  = (~\D<83>  & \C<83> ) | (\D<83>  & ~\C<83> ),
  \new_C<5>  = (\[647]  & (\D<5>  & \C<5> )) | ((\[868]  & \[653] ) | ((~\[867]  & \[649] ) | ((\[867]  & \[650] ) | ((\[654]  & \key<8> ) | (\[651]  & \key<16> ))))),
  \[523]  = \new_C<9> ,
  \[713]  = \D<82>  | \C<82> ,
  \new_C<6>  = (\[647]  & (\D<6>  & \C<6> )) | ((\[866]  & \[653] ) | ((~\[865]  & \[649] ) | ((\[865]  & \[650] ) | ((\[654]  & \key<0> ) | (\[651]  & \key<8> ))))),
  \[524]  = \new_C<8> ,
  \new_C<55>  = (\[647]  & (\D<55>  & \C<55> )) | ((\[768]  & \[653] ) | ((~\[767]  & \[649] ) | ((\[767]  & \[650] ) | ((\[654]  & \key<184> ) | (\[651]  & \key<99> ))))),
  \[714]  = (~\D<82>  & \C<82> ) | (\D<82>  & ~\C<82> ),
  \new_C<7>  = (\[647]  & (\D<7>  & \C<7> )) | ((\[864]  & \[653] ) | ((~\[863]  & \[649] ) | ((\[863]  & \[650] ) | ((\[654]  & \key<57> ) | (\[651]  & \key<0> ))))),
  \KSi<89>  = \C<91> ,
  \[525]  = \new_C<7> ,
  \new_C<56>  = (\[647]  & (\D<56>  & \C<56> )) | ((\[766]  & \[653] ) | ((~\[765]  & \[649] ) | ((\[765]  & \[650] ) | ((\[654]  & \key<176> ) | (\[651]  & \key<184> ))))),
  \[715]  = \D<81>  | \C<81> ,
  \new_C<8>  = (\[647]  & (\D<8>  & \C<8> )) | ((\[862]  & \[653] ) | ((~\[861]  & \[649] ) | ((\[861]  & \[650] ) | ((\[654]  & \key<49> ) | (\[651]  & \key<57> ))))),
  \[526]  = \new_C<6> ,
  \new_C<57>  = (\[647]  & (\D<57>  & \C<57> )) | ((\[764]  & \[653] ) | ((~\[763]  & \[649] ) | ((\[763]  & \[650] ) | ((\[654]  & \key<168> ) | (\[651]  & \key<176> ))))),
  \[716]  = (~\D<81>  & \C<81> ) | (\D<81>  & ~\C<81> ),
  \[527]  = \new_C<5> ,
  \new_C<58>  = (\[647]  & (\D<58>  & \C<58> )) | ((\[762]  & \[653] ) | ((~\[761]  & \[649] ) | ((\[761]  & \[650] ) | ((\[654]  & \key<160> ) | (\[651]  & \key<168> ))))),
  \[717]  = \D<80>  | \C<80> ,
  \KSi<86>  = \C<95> ,
  \[528]  = \new_C<4> ,
  \new_C<51>  = (\[647]  & (\D<51>  & \C<51> )) | ((\[776]  & \[653] ) | ((~\[775]  & \[649] ) | ((\[775]  & \[650] ) | ((\[654]  & \key<123> ) | (\[651]  & \key<66> ))))),
  \[718]  = (~\D<80>  & \C<80> ) | (\D<80>  & ~\C<80> ),
  \KSi<85>  = \C<102> ,
  \[529]  = \new_C<3> ,
  \new_C<52>  = (\[647]  & (\D<52>  & \C<52> )) | ((\[774]  & \[653] ) | ((~\[773]  & \[649] ) | ((\[773]  & \[650] ) | ((\[654]  & \key<115> ) | (\[651]  & \key<123> ))))),
  \[719]  = \D<79>  | \C<79> ,
  \KSi<88>  = \C<109> ,
  \new_C<53>  = (\[647]  & (\D<53>  & \C<53> )) | ((\[772]  & \[653] ) | ((~\[771]  & \[649] ) | ((\[771]  & \[650] ) | ((\[654]  & \key<107> ) | (\[651]  & \key<115> ))))),
  \KSi<87>  = \C<87> ,
  \new_C<54>  = (\[647]  & (\D<54>  & \C<54> )) | ((\[770]  & \[653] ) | ((~\[769]  & \[649] ) | ((\[769]  & \[650] ) | ((\[654]  & \key<99> ) | (\[651]  & \key<107> ))))),
  \KSi<92>  = \C<110> ,
  \KSi<91>  = \C<90> ,
  \KSi<94>  = \C<96> ,
  \KSi<93>  = \C<103> ,
  \new_C<50>  = (\[647]  & (\D<50>  & \C<50> )) | ((\[778]  & \[653] ) | ((~\[777]  & \[649] ) | ((\[777]  & \[650] ) | ((\[654]  & \key<66> ) | (\[651]  & \key<74> ))))),
  \[530]  = \new_C<2> ,
  \new_C<69>  = (\[647]  & (\D<69>  & \C<69> )) | ((\[740]  & \[653] ) | ((~\[739]  & \[649] ) | ((\[739]  & \[650] ) | ((\[654]  & \key<137> ) | (\[651]  & \key<145> ))))),
  \[720]  = (~\D<79>  & \C<79> ) | (\D<79>  & ~\C<79> ),
  \[531]  = \new_C<1> ,
  \[721]  = \D<78>  | \C<78> ,
  \KSi<90>  = \C<109> ,
  \[532]  = \new_C<0> ,
  \[722]  = (~\D<78>  & \C<78> ) | (\D<78>  & ~\C<78> ),
  \[533]  = \new_D<111> ,
  \[723]  = \D<77>  | \C<77> ,
  \[534]  = \new_D<110> ,
  \new_C<65>  = (\[647]  & (\D<65>  & \C<65> )) | ((\[748]  & \[653] ) | ((~\[747]  & \[649] ) | ((\[747]  & \[650] ) | ((\[654]  & \key<169> ) | (\[651]  & \key<177> ))))),
  \[724]  = (~\D<77>  & \C<77> ) | (\D<77>  & ~\C<77> ),
  \KSi<99>  = \D<8> ,
  \[535]  = \new_D<109> ,
  \new_C<66>  = (\[647]  & (\D<66>  & \C<66> )) | ((\[746]  & \[653] ) | ((~\[745]  & \[649] ) | ((\[745]  & \[650] ) | ((\[654]  & \key<161> ) | (\[651]  & \key<169> ))))),
  \[725]  = \D<76>  | \C<76> ,
  \[536]  = \new_D<108> ,
  \new_C<67>  = (\[647]  & (\D<67>  & \C<67> )) | ((\[744]  & \[653] ) | ((~\[743]  & \[649] ) | ((\[743]  & \[650] ) | ((\[654]  & \key<153> ) | (\[651]  & \key<161> ))))),
  \[726]  = (~\D<76>  & \C<76> ) | (\D<76>  & ~\C<76> ),
  \[537]  = \new_D<107> ,
  \new_C<68>  = (\[647]  & (\D<68>  & \C<68> )) | ((\[742]  & \[653] ) | ((~\[741]  & \[649] ) | ((\[741]  & \[650] ) | ((\[654]  & \key<145> ) | (\[651]  & \key<153> ))))),
  \[727]  = \D<75>  | \C<75> ,
  \KSi<96>  = \D<12> ,
  \[538]  = \new_D<106> ,
  \new_C<61>  = (\[647]  & (\D<61>  & \C<61> )) | ((\[756]  & \[653] ) | ((~\[755]  & \[649] ) | ((\[755]  & \[650] ) | ((\[654]  & \key<136> ) | (\[651]  & \key<144> ))))),
  \[728]  = (~\D<75>  & \C<75> ) | (\D<75>  & ~\C<75> ),
  \KSi<95>  = \C<85> ,
  \[539]  = \new_D<105> ,
  \new_C<62>  = (\[647]  & (\D<62>  & \C<62> )) | ((\[754]  & \[653] ) | ((~\[753]  & \[649] ) | ((\[753]  & \[650] ) | ((\[654]  & \key<128> ) | (\[651]  & \key<136> ))))),
  \[729]  = \D<74>  | \C<74> ,
  \KSi<98>  = \D<2> ,
  \new_C<63>  = (\[647]  & (\D<63>  & \C<63> )) | ((\[752]  & \[653] ) | ((~\[751]  & \[649] ) | ((\[751]  & \[650] ) | ((\[654]  & \key<185> ) | (\[651]  & \key<128> ))))),
  \KSi<97>  = \D<23> ,
  \new_C<64>  = (\[647]  & (\D<64>  & \C<64> )) | ((\[750]  & \[653] ) | ((~\[749]  & \[649] ) | ((\[749]  & \[650] ) | ((\[654]  & \key<177> ) | (\[651]  & \key<185> ))))),
  \KSi<120>  = \D<40> ,
  \KSi<121>  = \D<51> ,
  \new_C<60>  = (\[647]  & (\D<60>  & \C<60> )) | ((\[758]  & \[653] ) | ((~\[757]  & \[649] ) | ((\[757]  & \[650] ) | ((\[654]  & \key<144> ) | (\[651]  & \key<152> ))))),
  \KSi<122>  = \D<30> ,
  \[540]  = \new_D<104> ,
  \new_C<79>  = (\[647]  & (\D<79>  & \C<79> )) | ((\[720]  & \[653] ) | ((~\[719]  & \[649] ) | ((\[719]  & \[650] ) | ((\[654]  & \key<187> ) | (\[651]  & \key<130> ))))),
  \[730]  = (~\D<74>  & \C<74> ) | (\D<74>  & ~\C<74> ),
  \KSi<123>  = \D<36> ,
  \[541]  = \new_D<103> ,
  \[731]  = \D<73>  | \C<73> ,
  \KSi<124>  = \D<46> ,
  \[542]  = \new_D<102> ,
  \[732]  = (~\D<73>  & \C<73> ) | (\D<73>  & ~\C<73> ),
  \KSi<125>  = \D<54> ,
  \[543]  = \new_D<101> ,
  \[733]  = \D<72>  | \C<72> ,
  \KSi<126>  = \D<29> ,
  \[544]  = \new_D<100> ,
  \new_C<75>  = (\[647]  & (\D<75>  & \C<75> )) | ((\[728]  & \[653] ) | ((~\[727]  & \[649] ) | ((\[727]  & \[650] ) | ((\[654]  & \key<154> ) | (\[651]  & \key<162> ))))),
  \[734]  = (~\D<72>  & \C<72> ) | (\D<72>  & ~\C<72> ),
  \KSi<127>  = \D<39> ,
  \[545]  = \new_D<99> ,
  \new_C<76>  = (\[647]  & (\D<76>  & \C<76> )) | ((\[726]  & \[653] ) | ((~\[725]  & \[649] ) | ((\[725]  & \[650] ) | ((\[654]  & \key<146> ) | (\[651]  & \key<154> ))))),
  \[735]  = \D<71>  | \C<71> ,
  \KSi<128>  = \D<50> ,
  \[546]  = \new_D<98> ,
  \new_C<77>  = (\[647]  & (\D<77>  & \C<77> )) | ((\[724]  & \[653] ) | ((~\[723]  & \[649] ) | ((\[723]  & \[650] ) | ((\[654]  & \key<138> ) | (\[651]  & \key<146> ))))),
  \[736]  = (~\D<71>  & \C<71> ) | (\D<71>  & ~\C<71> ),
  \KSi<129>  = \D<44> ,
  \[547]  = \new_D<97> ,
  \new_C<78>  = (\[647]  & (\D<78>  & \C<78> )) | ((\[722]  & \[653] ) | ((~\[721]  & \[649] ) | ((\[721]  & \[650] ) | ((\[654]  & \key<130> ) | (\[651]  & \key<138> ))))),
  \[737]  = \D<70>  | \C<70> ,
  \[548]  = \new_D<96> ,
  \new_C<71>  = (\[647]  & (\D<71>  & \C<71> )) | ((\[736]  & \[653] ) | ((~\[735]  & \[649] ) | ((\[735]  & \[650] ) | ((\[654]  & \key<186> ) | (\[651]  & \key<129> ))))),
  \[738]  = (~\D<70>  & \C<70> ) | (\D<70>  & ~\C<70> ),
  \[549]  = \new_D<95> ,
  \new_C<72>  = (\[647]  & (\D<72>  & \C<72> )) | ((\[734]  & \[653] ) | ((~\[733]  & \[649] ) | ((\[733]  & \[650] ) | ((\[654]  & \key<178> ) | (\[651]  & \key<186> ))))),
  \[739]  = \D<69>  | \C<69> ,
  \new_C<73>  = (\[647]  & (\D<73>  & \C<73> )) | ((\[732]  & \[653] ) | ((~\[731]  & \[649] ) | ((\[731]  & \[650] ) | ((\[654]  & \key<170> ) | (\[651]  & \key<178> ))))),
  \new_C<74>  = (\[647]  & (\D<74>  & \C<74> )) | ((\[730]  & \[653] ) | ((~\[729]  & \[649] ) | ((\[729]  & \[650] ) | ((\[654]  & \key<162> ) | (\[651]  & \key<170> ))))),
  \KSi<110>  = \D<10> ,
  \KSi<111>  = \D<27> ,
  \new_C<70>  = (\[647]  & (\D<70>  & \C<70> )) | ((\[738]  & \[653] ) | ((~\[737]  & \[649] ) | ((\[737]  & \[650] ) | ((\[654]  & \key<129> ) | (\[651]  & \key<137> ))))),
  \KSi<112>  = \D<5> ,
  \[550]  = \new_D<94> ,
  \new_C<89>  = (\[647]  & (\D<89>  & \C<89> )) | ((\[700]  & \[653] ) | ((~\[699]  & \[649] ) | ((\[699]  & \[650] ) | ((\[654]  & \key<200> ) | (\[651]  & \key<208> ))))),
  \[740]  = (~\D<69>  & \C<69> ) | (\D<69>  & ~\C<69> ),
  \KSi<113>  = \D<24> ,
  \[551]  = \new_D<93> ,
  \[741]  = \D<68>  | \C<68> ,
  \KSi<114>  = \D<17> ,
  \[552]  = \new_D<92> ,
  \[742]  = (~\D<68>  & \C<68> ) | (\D<68>  & ~\C<68> ),
  \KSi<115>  = \D<13> ,
  \[553]  = \new_D<91> ,
  \[743]  = \D<67>  | \C<67> ,
  \KSi<116>  = \D<21> ,
  \[554]  = \new_D<90> ,
  \new_C<85>  = (\[647]  & (\D<85>  & \C<85> )) | ((\[708]  & \[653] ) | ((~\[707]  & \[649] ) | ((\[707]  & \[650] ) | ((\[654]  & \key<232> ) | (\[651]  & \key<240> ))))),
  \[744]  = (~\D<67>  & \C<67> ) | (\D<67>  & ~\C<67> ),
  \KSi<117>  = \D<7> ,
  \[555]  = \new_D<89> ,
  \new_C<86>  = (\[647]  & (\D<86>  & \C<86> )) | ((\[706]  & \[653] ) | ((~\[705]  & \[649] ) | ((\[705]  & \[650] ) | ((\[654]  & \key<224> ) | (\[651]  & \key<232> ))))),
  \[745]  = \D<66>  | \C<66> ,
  \KSi<118>  = \D<0> ,
  \[556]  = \new_D<88> ,
  \new_C<87>  = (\[647]  & (\D<87>  & \C<87> )) | ((\[704]  & \[653] ) | ((~\[703]  & \[649] ) | ((\[703]  & \[650] ) | ((\[654]  & \key<216> ) | (\[651]  & \key<224> ))))),
  \[746]  = (~\D<66>  & \C<66> ) | (\D<66>  & ~\C<66> ),
  \KSi<119>  = \D<3> ,
  \[557]  = \new_D<87> ,
  \new_C<88>  = (\[647]  & (\D<88>  & \C<88> )) | ((\[702]  & \[653] ) | ((~\[701]  & \[649] ) | ((\[701]  & \[650] ) | ((\[654]  & \key<208> ) | (\[651]  & \key<216> ))))),
  \[747]  = \D<65>  | \C<65> ,
  \[558]  = \new_D<86> ,
  \new_C<81>  = (\[647]  & (\D<81>  & \C<81> )) | ((\[716]  & \[653] ) | ((~\[715]  & \[649] ) | ((\[715]  & \[650] ) | ((\[654]  & \key<171> ) | (\[651]  & \key<179> ))))),
  \[748]  = (~\D<65>  & \C<65> ) | (\D<65>  & ~\C<65> ),
  \[559]  = \new_D<85> ,
  \new_C<82>  = (\[647]  & (\D<82>  & \C<82> )) | ((\[714]  & \[653] ) | ((~\[713]  & \[649] ) | ((\[713]  & \[650] ) | ((\[654]  & \key<163> ) | (\[651]  & \key<171> ))))),
  \[749]  = \D<64>  | \C<64> ,
  \new_C<83>  = (\[647]  & (\D<83>  & \C<83> )) | ((\[712]  & \[653] ) | ((~\[711]  & \[649] ) | ((\[711]  & \[650] ) | ((\[654]  & \key<248> ) | (\[651]  & \key<163> ))))),
  \new_C<84>  = (\[647]  & (\D<84>  & \C<84> )) | ((\[710]  & \[653] ) | ((~\[709]  & \[649] ) | ((\[709]  & \[650] ) | ((\[654]  & \key<240> ) | (\[651]  & \key<248> ))))),
  \KSi<140>  = \D<49> ,
  \KSi<141>  = \D<35> ,
  \new_C<80>  = (\[647]  & (\D<80>  & \C<80> )) | ((\[718]  & \[653] ) | ((~\[717]  & \[649] ) | ((\[717]  & \[650] ) | ((\[654]  & \key<179> ) | (\[651]  & \key<187> ))))),
  \KSi<142>  = \D<28> ,
  \[560]  = \new_D<84> ,
  \[750]  = (~\D<64>  & \C<64> ) | (\D<64>  & ~\C<64> ),
  \KSi<143>  = \D<31> ,
  \[561]  = \new_D<83> ,
  \[751]  = \D<63>  | \C<63> ,
  \KSi<144>  = \D<68> ,
  \new_D<99>  = (\[648]  & (\D<99>  & \C<99> )) | ((\[680]  & \[652] ) | ((~\[679]  & \[650] ) | ((\[679]  & \[649] ) | ((\[654]  & \key<252> ) | (\[651]  & \key<197> ))))),
  \[562]  = \new_D<82> ,
  \[752]  = (~\D<63>  & \C<63> ) | (\D<63>  & ~\C<63> ),
  \KSi<145>  = \D<79> ,
  \[563]  = \new_D<81> ,
  \[753]  = \D<62>  | \C<62> ,
  \KSi<146>  = \D<58> ,
  \[564]  = \new_D<80> ,
  \[754]  = (~\D<62>  & \C<62> ) | (\D<62>  & ~\C<62> ),
  \KSi<147>  = \D<64> ,
  \[565]  = \new_D<79> ,
  \[755]  = \D<61>  | \C<61> ,
  \$$COND1<0>8.1  = (\[879]  & (~\count<1>  & ~\count<2> )) | (\[880]  & ~\[879] ),
  \KSi<148>  = \D<74> ,
  \new_D<95>  = (\[648]  & (\D<95>  & \C<95> )) | ((\[688]  & \[652] ) | ((~\[687]  & \[650] ) | ((\[687]  & \[649] ) | ((\[654]  & \key<221> ) | (\[651]  & \key<229> ))))),
  \[566]  = \new_D<78> ,
  \[756]  = (~\D<61>  & \C<61> ) | (\D<61>  & ~\C<61> ),
  \KSi<149>  = \D<82> ,
  \new_D<96>  = (\[648]  & (\D<96>  & \C<96> )) | ((\[686]  & \[652] ) | ((~\[685]  & \[650] ) | ((\[685]  & \[649] ) | ((\[654]  & \key<213> ) | (\[651]  & \key<221> ))))),
  \[567]  = \new_D<77> ,
  \[757]  = \D<60>  | \C<60> ,
  \new_D<97>  = (\[648]  & (\D<97>  & \C<97> )) | ((\[684]  & \[652] ) | ((~\[683]  & \[650] ) | ((\[683]  & \[649] ) | ((\[654]  & \key<205> ) | (\[651]  & \key<213> )))));
always begin
  \D<0>  = \[644] ;
  \D<1>  = \[643] ;
  \D<2>  = \[642] ;
  \D<3>  = \[641] ;
  \D<4>  = \[640] ;
  \D<5>  = \[639] ;
  \D<6>  = \[638] ;
  \C<10>  = \[522] ;
  \D<7>  = \[637] ;
  \C<11>  = \[521] ;
  \D<8>  = \[636] ;
  \C<12>  = \[520] ;
  \D<9>  = \[635] ;
  \C<13>  = \[519] ;
  \C<14>  = \[518] ;
  \C<15>  = \[517] ;
  \C<16>  = \[516] ;
  \C<17>  = \[515] ;
  \C<18>  = \[514] ;
  \C<19>  = \[513] ;
  \C<20>  = \[512] ;
  \C<21>  = \[511] ;
  \C<22>  = \[510] ;
  \C<23>  = \[509] ;
  \C<24>  = \[508] ;
  \C<25>  = \[507] ;
  \C<26>  = \[506] ;
  \C<27>  = \[505] ;
  \C<28>  = \[504] ;
  \C<29>  = \[503] ;
  \C<30>  = \[502] ;
  \C<31>  = \[501] ;
  \C<32>  = \[500] ;
  \C<33>  = \[499] ;
  \C<34>  = \[498] ;
  \C<35>  = \[497] ;
  \C<36>  = \[496] ;
  \C<37>  = \[495] ;
  \C<38>  = \[494] ;
  \C<39>  = \[493] ;
  \C<40>  = \[492] ;
  \C<41>  = \[491] ;
  \C<42>  = \[490] ;
  \C<43>  = \[489] ;
  \C<44>  = \[488] ;
  \C<45>  = \[487] ;
  \C<46>  = \[486] ;
  \C<47>  = \[485] ;
  \C<48>  = \[484] ;
  \C<49>  = \[483] ;
  \C<50>  = \[482] ;
  \C<51>  = \[481] ;
  \C<52>  = \[480] ;
  \C<53>  = \[479] ;
  \C<54>  = \[478] ;
  \C<55>  = \[477] ;
  \C<56>  = \[476] ;
  \C<57>  = \[475] ;
  \C<58>  = \[474] ;
  \C<59>  = \[473] ;
  \C<60>  = \[472] ;
  \C<61>  = \[471] ;
  \C<62>  = \[470] ;
  \C<63>  = \[469] ;
  \C<64>  = \[468] ;
  \C<65>  = \[467] ;
  \C<66>  = \[466] ;
  \C<67>  = \[465] ;
  \C<68>  = \[464] ;
  \C<69>  = \[463] ;
  \C<70>  = \[462] ;
  \C<71>  = \[461] ;
  \C<72>  = \[460] ;
  \C<73>  = \[459] ;
  \C<74>  = \[458] ;
  \C<75>  = \[457] ;
  \C<76>  = \[456] ;
  \C<77>  = \[455] ;
  \C<78>  = \[454] ;
  \C<79>  = \[453] ;
  \C<80>  = \[452] ;
  \C<81>  = \[451] ;
  \C<82>  = \[450] ;
  \C<83>  = \[449] ;
  \C<84>  = \[448] ;
  \C<85>  = \[447] ;
  \C<86>  = \[446] ;
  \C<87>  = \[445] ;
  \C<88>  = \[444] ;
  \C<89>  = \[443] ;
  \C<90>  = \[442] ;
  \C<91>  = \[441] ;
  \D<10>  = \[634] ;
  \C<92>  = \[440] ;
  \D<11>  = \[633] ;
  \C<93>  = \[439] ;
  \D<12>  = \[632] ;
  \C<94>  = \[438] ;
  \D<13>  = \[631] ;
  \C<95>  = \[437] ;
  \D<14>  = \[630] ;
  \C<96>  = \[436] ;
  \D<15>  = \[629] ;
  \C<97>  = \[435] ;
  \D<16>  = \[628] ;
  \C<98>  = \[434] ;
  \D<17>  = \[627] ;
  \C<99>  = \[433] ;
  \D<18>  = \[626] ;
  \D<19>  = \[625] ;
  \D<20>  = \[624] ;
  \D<21>  = \[623] ;
  \D<22>  = \[622] ;
  \D<23>  = \[621] ;
  \D<24>  = \[620] ;
  \D<25>  = \[619] ;
  \D<26>  = \[618] ;
  \D<27>  = \[617] ;
  \D<28>  = \[616] ;
  \D<29>  = \[615] ;
  \D<30>  = \[614] ;
  \D<31>  = \[613] ;
  \D<32>  = \[612] ;
  \D<33>  = \[611] ;
  \D<34>  = \[610] ;
  \D<35>  = \[609] ;
  \D<36>  = \[608] ;
  \D<37>  = \[607] ;
  \D<38>  = \[606] ;
  \D<39>  = \[605] ;
  \D<40>  = \[604] ;
  \D<41>  = \[603] ;
  \D<42>  = \[602] ;
  \D<43>  = \[601] ;
  \D<44>  = \[600] ;
  \D<45>  = \[599] ;
  \D<46>  = \[598] ;
  \D<47>  = \[597] ;
  \D<48>  = \[596] ;
  \D<49>  = \[595] ;
  \D<50>  = \[594] ;
  \D<51>  = \[593] ;
  \D<52>  = \[592] ;
  \D<53>  = \[591] ;
  \D<54>  = \[590] ;
  \D<55>  = \[589] ;
  \D<56>  = \[588] ;
  \D<57>  = \[587] ;
  \D<58>  = \[586] ;
  \D<59>  = \[585] ;
  \D<60>  = \[584] ;
  \D<61>  = \[583] ;
  \D<62>  = \[582] ;
  \D<63>  = \[581] ;
  \D<64>  = \[580] ;
  \D<65>  = \[579] ;
  \D<66>  = \[578] ;
  \D<67>  = \[577] ;
  \D<68>  = \[576] ;
  \D<69>  = \[575] ;
  \C<100>  = \[432] ;
  \D<70>  = \[574] ;
  \C<101>  = \[431] ;
  \D<71>  = \[573] ;
  \C<102>  = \[430] ;
  \D<72>  = \[572] ;
  \C<103>  = \[429] ;
  \D<73>  = \[571] ;
  \C<104>  = \[428] ;
  \D<74>  = \[570] ;
  \C<105>  = \[427] ;
  \D<75>  = \[569] ;
  \C<106>  = \[426] ;
  \D<76>  = \[568] ;
  \C<107>  = \[425] ;
  \D<77>  = \[567] ;
  \C<108>  = \[424] ;
  \C<0>  = \[532] ;
  \D<78>  = \[566] ;
  \C<109>  = \[423] ;
  \C<1>  = \[531] ;
  \D<79>  = \[565] ;
  \C<2>  = \[530] ;
  \C<3>  = \[529] ;
  \C<4>  = \[528] ;
  \C<5>  = \[527] ;
  \C<6>  = \[526] ;
  \C<7>  = \[525] ;
  \C<110>  = \[422] ;
  \C<8>  = \[524] ;
  \D<80>  = \[564] ;
  \C<111>  = \[421] ;
  \C<9>  = \[523] ;
  \D<81>  = \[563] ;
  \D<82>  = \[562] ;
  \D<83>  = \[561] ;
  \D<84>  = \[560] ;
  \D<85>  = \[559] ;
  \D<86>  = \[558] ;
  \D<87>  = \[557] ;
  \D<88>  = \[556] ;
  \D<89>  = \[555] ;
  \D<90>  = \[554] ;
  \D<91>  = \[553] ;
  \D<92>  = \[552] ;
  \D<93>  = \[551] ;
  \D<94>  = \[550] ;
  \D<95>  = \[549] ;
  \D<96>  = \[548] ;
  \D<97>  = \[547] ;
  \D<98>  = \[546] ;
  \D<99>  = \[545] ;
  \D<100>  = \[544] ;
  \D<101>  = \[543] ;
  \D<102>  = \[542] ;
  \D<103>  = \[541] ;
  \D<104>  = \[540] ;
  \D<105>  = \[539] ;
  \D<106>  = \[538] ;
  \D<107>  = \[537] ;
  \D<108>  = \[536] ;
  \D<109>  = \[535] ;
  \D<110>  = \[534] ;
  \D<111>  = \[533] ;
end
initial begin
  \D<0>  = 0;
  \D<1>  = 0;
  \D<2>  = 0;
  \D<3>  = 0;
  \D<4>  = 0;
  \D<5>  = 0;
  \D<6>  = 0;
  \C<10>  = 0;
  \D<7>  = 0;
  \C<11>  = 0;
  \D<8>  = 0;
  \C<12>  = 0;
  \D<9>  = 0;
  \C<13>  = 0;
  \C<14>  = 0;
  \C<15>  = 0;
  \C<16>  = 0;
  \C<17>  = 0;
  \C<18>  = 0;
  \C<19>  = 0;
  \C<20>  = 0;
  \C<21>  = 0;
  \C<22>  = 0;
  \C<23>  = 0;
  \C<24>  = 0;
  \C<25>  = 0;
  \C<26>  = 0;
  \C<27>  = 0;
  \C<28>  = 0;
  \C<29>  = 0;
  \C<30>  = 0;
  \C<31>  = 0;
  \C<32>  = 0;
  \C<33>  = 0;
  \C<34>  = 0;
  \C<35>  = 0;
  \C<36>  = 0;
  \C<37>  = 0;
  \C<38>  = 0;
  \C<39>  = 0;
  \C<40>  = 0;
  \C<41>  = 0;
  \C<42>  = 0;
  \C<43>  = 0;
  \C<44>  = 0;
  \C<45>  = 0;
  \C<46>  = 0;
  \C<47>  = 0;
  \C<48>  = 0;
  \C<49>  = 0;
  \C<50>  = 0;
  \C<51>  = 0;
  \C<52>  = 0;
  \C<53>  = 0;
  \C<54>  = 0;
  \C<55>  = 0;
  \C<56>  = 0;
  \C<57>  = 0;
  \C<58>  = 0;
  \C<59>  = 0;
  \C<60>  = 0;
  \C<61>  = 0;
  \C<62>  = 0;
  \C<63>  = 0;
  \C<64>  = 0;
  \C<65>  = 0;
  \C<66>  = 0;
  \C<67>  = 0;
  \C<68>  = 0;
  \C<69>  = 0;
  \C<70>  = 0;
  \C<71>  = 0;
  \C<72>  = 0;
  \C<73>  = 0;
  \C<74>  = 0;
  \C<75>  = 0;
  \C<76>  = 0;
  \C<77>  = 0;
  \C<78>  = 0;
  \C<79>  = 0;
  \C<80>  = 0;
  \C<81>  = 0;
  \C<82>  = 0;
  \C<83>  = 0;
  \C<84>  = 0;
  \C<85>  = 0;
  \C<86>  = 0;
  \C<87>  = 0;
  \C<88>  = 0;
  \C<89>  = 0;
  \C<90>  = 0;
  \C<91>  = 0;
  \D<10>  = 0;
  \C<92>  = 0;
  \D<11>  = 0;
  \C<93>  = 0;
  \D<12>  = 0;
  \C<94>  = 0;
  \D<13>  = 0;
  \C<95>  = 0;
  \D<14>  = 0;
  \C<96>  = 0;
  \D<15>  = 0;
  \C<97>  = 0;
  \D<16>  = 0;
  \C<98>  = 0;
  \D<17>  = 0;
  \C<99>  = 0;
  \D<18>  = 0;
  \D<19>  = 0;
  \D<20>  = 0;
  \D<21>  = 0;
  \D<22>  = 0;
  \D<23>  = 0;
  \D<24>  = 0;
  \D<25>  = 0;
  \D<26>  = 0;
  \D<27>  = 0;
  \D<28>  = 0;
  \D<29>  = 0;
  \D<30>  = 0;
  \D<31>  = 0;
  \D<32>  = 0;
  \D<33>  = 0;
  \D<34>  = 0;
  \D<35>  = 0;
  \D<36>  = 0;
  \D<37>  = 0;
  \D<38>  = 0;
  \D<39>  = 0;
  \D<40>  = 0;
  \D<41>  = 0;
  \D<42>  = 0;
  \D<43>  = 0;
  \D<44>  = 0;
  \D<45>  = 0;
  \D<46>  = 0;
  \D<47>  = 0;
  \D<48>  = 0;
  \D<49>  = 0;
  \D<50>  = 0;
  \D<51>  = 0;
  \D<52>  = 0;
  \D<53>  = 0;
  \D<54>  = 0;
  \D<55>  = 0;
  \D<56>  = 0;
  \D<57>  = 0;
  \D<58>  = 0;
  \D<59>  = 0;
  \D<60>  = 0;
  \D<61>  = 0;
  \D<62>  = 0;
  \D<63>  = 0;
  \D<64>  = 0;
  \D<65>  = 0;
  \D<66>  = 0;
  \D<67>  = 0;
  \D<68>  = 0;
  \D<69>  = 0;
  \C<100>  = 0;
  \D<70>  = 0;
  \C<101>  = 0;
  \D<71>  = 0;
  \C<102>  = 0;
  \D<72>  = 0;
  \C<103>  = 0;
  \D<73>  = 0;
  \C<104>  = 0;
  \D<74>  = 0;
  \C<105>  = 0;
  \D<75>  = 0;
  \C<106>  = 0;
  \D<76>  = 0;
  \C<107>  = 0;
  \D<77>  = 0;
  \C<108>  = 0;
  \C<0>  = 0;
  \D<78>  = 0;
  \C<109>  = 0;
  \C<1>  = 0;
  \D<79>  = 0;
  \C<2>  = 0;
  \C<3>  = 0;
  \C<4>  = 0;
  \C<5>  = 0;
  \C<6>  = 0;
  \C<7>  = 0;
  \C<110>  = 0;
  \C<8>  = 0;
  \D<80>  = 0;
  \C<111>  = 0;
  \C<9>  = 0;
  \D<81>  = 0;
  \D<82>  = 0;
  \D<83>  = 0;
  \D<84>  = 0;
  \D<85>  = 0;
  \D<86>  = 0;
  \D<87>  = 0;
  \D<88>  = 0;
  \D<89>  = 0;
  \D<90>  = 0;
  \D<91>  = 0;
  \D<92>  = 0;
  \D<93>  = 0;
  \D<94>  = 0;
  \D<95>  = 0;
  \D<96>  = 0;
  \D<97>  = 0;
  \D<98>  = 0;
  \D<99>  = 0;
  \D<100>  = 0;
  \D<101>  = 0;
  \D<102>  = 0;
  \D<103>  = 0;
  \D<104>  = 0;
  \D<105>  = 0;
  \D<106>  = 0;
  \D<107>  = 0;
  \D<108>  = 0;
  \D<109>  = 0;
  \D<110>  = 0;
  \D<111>  = 0;
end
endmodule

