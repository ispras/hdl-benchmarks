//NOTE: no-implementation module stub

module GtCLK_MUX2 (
    output Z,
    input S,
    input A,
    input B
);

endmodule
