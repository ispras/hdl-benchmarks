module bitwise_nor_4_6_9(a, b, c);
  input [3:0] a;
  input [5:0] b;
  output [8:0] c;
  assign c = a ~| b;
endmodule
