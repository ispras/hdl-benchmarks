// IWLS benchmark module "i3" printed on Wed May 29 16:38:48 2002
module i3(\V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) , \V56(3) , \V28(3) , \V56(4) , \V28(4) , \V56(5) , \V28(5) , \V56(6) , \V28(6) , \V56(7) , \V28(7) , \V56(8) , \V28(8) , \V56(9) , \V28(9) , \V56(10) , \V28(10) , \V56(11) , \V28(11) , \V56(12) , \V28(12) , \V56(13) , \V28(13) , \V56(14) , \V28(14) , \V56(15) , \V28(15) , \V56(16) , \V28(16) , \V56(17) , \V28(17) , \V56(18) , \V28(18) , \V56(19) , \V28(19) , \V56(20) , \V28(20) , \V56(21) , \V28(21) , \V56(22) , \V28(22) , \V56(23) , \V28(23) , \V56(24) , \V28(24) , \V56(25) , \V28(25) , \V56(26) , \V28(26) , \V56(27) , \V28(27) , \V120(0) , \V88(0) , \V120(1) , \V88(1) , \V120(2) , \V88(2) , \V120(3) , \V88(3) , \V120(4) , \V88(4) , \V120(5) , \V88(5) , \V120(6) , \V88(6) , \V120(7) , \V88(7) , \V120(8) , \V88(8) , \V120(9) , \V88(9) , \V120(10) , \V88(10) , \V120(11) , \V88(11) , \V120(12) , \V88(12) , \V120(13) , \V88(13) , \V120(14) , \V88(14) , \V120(15) , \V88(15) , \V120(16) , \V88(16) , \V120(17) , \V88(17) , \V120(18) , \V88(18) , \V120(19) , \V88(19) , \V120(20) , \V88(20) , \V120(21) , \V88(21) , \V120(22) , \V88(22) , \V120(23) , \V88(23) , \V120(24) , \V88(24) , \V120(25) , \V88(25) , \V120(26) , \V88(26) , \V120(27) , \V88(27) , \V120(28) , \V88(28) , \V120(29) , \V88(29) , \V120(30) , \V88(30) , \V120(31) , \V88(31) , \V132(0) , \V126(0) , \V132(1) , \V126(1) , \V132(2) , \V126(2) , \V132(3) , \V126(3) , \V132(4) , \V126(4) , \V132(5) , \V126(5) , \V134(0) , \V134(1) , \V138(0) , \V138(1) , \V138(2) , \V138(3) );
input
  \V132(5) ,
  \V28(13) ,
  \V126(1) ,
  \V88(21) ,
  \V132(4) ,
  \V28(12) ,
  \V126(0) ,
  \V88(20) ,
  \V28(15) ,
  \V28(14) ,
  \V132(1) ,
  \V132(0) ,
  \V28(11) ,
  \V88(27) ,
  \V28(10) ,
  \V88(0) ,
  \V88(26) ,
  \V88(1) ,
  \V88(29) ,
  \V88(2) ,
  \V88(28) ,
  \V88(3) ,
  \V88(4) ,
  \V28(17) ,
  \V88(5) ,
  \V120(31) ,
  \V28(16) ,
  \V88(6) ,
  \V120(30) ,
  \V56(13) ,
  \V28(19) ,
  \V88(7) ,
  \V56(12) ,
  \V28(18) ,
  \V88(8) ,
  \V56(15) ,
  \V28(23) ,
  \V88(9) ,
  \V88(31) ,
  \V56(14) ,
  \V28(22) ,
  \V88(30) ,
  \V28(25) ,
  \V28(24) ,
  \V56(11) ,
  \V56(10) ,
  \V28(21) ,
  \V28(20) ,
  \V120(27) ,
  \V120(26) ,
  \V120(29) ,
  \V56(17) ,
  \V120(28) ,
  \V120(3) ,
  \V56(0) ,
  \V56(16) ,
  \V120(2) ,
  \V56(1) ,
  \V56(19) ,
  \V28(27) ,
  \V120(5) ,
  \V56(2) ,
  \V56(18) ,
  \V28(26) ,
  \V120(4) ,
  \V56(3) ,
  \V56(23) ,
  \V56(4) ,
  \V56(22) ,
  \V56(5) ,
  \V56(25) ,
  \V120(1) ,
  \V56(6) ,
  \V56(24) ,
  \V120(21) ,
  \V120(0) ,
  \V56(7) ,
  \V120(20) ,
  \V56(8) ,
  \V120(23) ,
  \V56(9) ,
  \V56(21) ,
  \V120(22) ,
  \V56(20) ,
  \V120(25) ,
  \V120(24) ,
  \V120(7) ,
  \V120(17) ,
  \V120(6) ,
  \V120(16) ,
  \V120(9) ,
  \V120(19) ,
  \V120(8) ,
  \V56(27) ,
  \V120(18) ,
  \V56(26) ,
  \V88(13) ,
  \V28(0) ,
  \V88(12) ,
  \V28(1) ,
  \V88(15) ,
  \V120(11) ,
  \V28(2) ,
  \V88(14) ,
  \V120(10) ,
  \V28(3) ,
  \V120(13) ,
  \V28(4) ,
  \V120(12) ,
  \V28(5) ,
  \V88(11) ,
  \V120(15) ,
  \V28(6) ,
  \V88(10) ,
  \V120(14) ,
  \V28(7) ,
  \V28(8) ,
  \V28(9) ,
  \V88(17) ,
  \V88(16) ,
  \V88(19) ,
  \V88(18) ,
  \V126(3) ,
  \V88(23) ,
  \V126(2) ,
  \V88(22) ,
  \V126(5) ,
  \V88(25) ,
  \V126(4) ,
  \V88(24) ,
  \V132(3) ,
  \V132(2) ;
output
  \V138(3) ,
  \V138(2) ,
  \V134(1) ,
  \V134(0) ,
  \V138(1) ,
  \V138(0) ;
wire
  \V202(7) ,
  \V202(6) ,
  \V202(9) ,
  \V202(8) ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \V170(11) ,
  \V170(10) ,
  \V170(13) ,
  \V186(3) ,
  \V170(12) ,
  \V154(11) ,
  \V186(2) ,
  \V170(15) ,
  \V154(10) ,
  \V186(5) ,
  \V170(14) ,
  \V154(13) ,
  \V186(4) ,
  \V154(12) ,
  \V154(15) ,
  \V154(14) ,
  \V186(1) ,
  \V186(0) ,
  \V202(11) ,
  \V202(10) ,
  \V202(13) ,
  \V202(12) ,
  \V186(7) ,
  \V202(15) ,
  \V186(6) ,
  \V202(14) ,
  \V186(9) ,
  \V186(8) ,
  \V154(3) ,
  \V154(2) ,
  \V154(5) ,
  \V154(4) ,
  \V154(1) ,
  \V154(0) ,
  \V170(3) ,
  \V170(2) ,
  \V170(5) ,
  \V170(4) ,
  \V154(7) ,
  \V154(6) ,
  \V154(9) ,
  \V186(11) ,
  \V170(1) ,
  \V154(8) ,
  \V186(10) ,
  \V170(0) ,
  \V186(13) ,
  \V186(12) ,
  \V202(3) ,
  \V186(15) ,
  \V202(2) ,
  \V186(14) ,
  \V202(5) ,
  \V170(7) ,
  \V202(4) ,
  \V170(6) ,
  \V170(9) ,
  \V170(8) ,
  \V202(1) ,
  \V202(0) ;
assign
  \V202(7)  = \V88(29)  | \V120(29) ,
  \V202(6)  = \V88(28)  | \V120(28) ,
  \V202(9)  = \V88(31)  | \V120(31) ,
  \V202(8)  = \V88(30)  | \V120(30) ,
  \[0]  = \V28(0)  | \V56(0) ,
  \[1]  = \V28(1)  | \V56(1) ,
  \[2]  = \V154(11)  & (\V154(10)  & (\V154(8)  & (\V154(9)  & (\V154(7)  & (\V154(5)  & (\V154(4)  & (\V154(6)  & (\V154(1)  & (\V154(0)  & (\V154(2)  & (\V154(3)  & (\V154(13)  & (\V154(12)  & (\V154(14)  & \V154(15) )))))))))))))),
  \[3]  = \V170(11)  & (\V170(10)  & (\V170(8)  & (\V170(9)  & (\V170(7)  & (\V170(5)  & (\V170(4)  & (\V170(6)  & (\V170(1)  & (\V170(0)  & (\V170(2)  & (\V170(3)  & (\V170(13)  & (\V170(12)  & (\V170(14)  & \V170(15) )))))))))))))),
  \[4]  = \V186(11)  & (\V186(10)  & (\V186(8)  & (\V186(9)  & (\V186(7)  & (\V186(5)  & (\V186(4)  & (\V186(6)  & (\V186(1)  & (\V186(0)  & (\V186(2)  & (\V186(3)  & (\V186(13)  & (\V186(12)  & (\V186(14)  & \V186(15) )))))))))))))),
  \[5]  = \V202(11)  & (\V202(10)  & (\V202(8)  & (\V202(9)  & (\V202(7)  & (\V202(5)  & (\V202(4)  & (\V202(6)  & (\V202(1)  & (\V202(0)  & (\V202(2)  & (\V202(3)  & (\V202(13)  & (\V202(12)  & (\V202(14)  & \V202(15) )))))))))))))),
  \V170(11)  = \V88(1)  | \V120(1) ,
  \V170(10)  = \V88(0)  | \V120(0) ,
  \V170(13)  = \V88(3)  | \V120(3) ,
  \V186(3)  = \V88(9)  | \V120(9) ,
  \V170(12)  = \V88(2)  | \V120(2) ,
  \V154(11)  = \V28(13)  | \V56(13) ,
  \V186(2)  = \V88(8)  | \V120(8) ,
  \V170(15)  = \V88(5)  | \V120(5) ,
  \V154(10)  = \V28(12)  | \V56(12) ,
  \V186(5)  = \V88(11)  | \V120(11) ,
  \V170(14)  = \V88(4)  | \V120(4) ,
  \V154(13)  = \V28(15)  | \V56(15) ,
  \V186(4)  = \V88(10)  | \V120(10) ,
  \V154(12)  = \V28(14)  | \V56(14) ,
  \V154(15)  = \V28(17)  | \V56(17) ,
  \V154(14)  = \V28(16)  | \V56(16) ,
  \V186(1)  = \V88(7)  | \V120(7) ,
  \V186(0)  = \V88(6)  | \V120(6) ,
  \V202(11)  = \V126(1)  | \V132(1) ,
  \V202(10)  = \V126(0)  | \V132(0) ,
  \V202(13)  = \V126(3)  | \V132(3) ,
  \V138(3)  = \[5] ,
  \V202(12)  = \V126(2)  | \V132(2) ,
  \V138(2)  = \[4] ,
  \V186(7)  = \V88(13)  | \V120(13) ,
  \V202(15)  = \V126(5)  | \V132(5) ,
  \V186(6)  = \V88(12)  | \V120(12) ,
  \V202(14)  = \V126(4)  | \V132(4) ,
  \V186(9)  = \V88(15)  | \V120(15) ,
  \V186(8)  = \V88(14)  | \V120(14) ,
  \V134(1)  = \[1] ,
  \V134(0)  = \[0] ,
  \V138(1)  = \[3] ,
  \V138(0)  = \[2] ,
  \V154(3)  = \V28(5)  | \V56(5) ,
  \V154(2)  = \V28(4)  | \V56(4) ,
  \V154(5)  = \V28(7)  | \V56(7) ,
  \V154(4)  = \V28(6)  | \V56(6) ,
  \V154(1)  = \V28(3)  | \V56(3) ,
  \V154(0)  = \V28(2)  | \V56(2) ,
  \V170(3)  = \V28(21)  | \V56(21) ,
  \V170(2)  = \V28(20)  | \V56(20) ,
  \V170(5)  = \V28(23)  | \V56(23) ,
  \V170(4)  = \V28(22)  | \V56(22) ,
  \V154(7)  = \V28(9)  | \V56(9) ,
  \V154(6)  = \V28(8)  | \V56(8) ,
  \V154(9)  = \V28(11)  | \V56(11) ,
  \V186(11)  = \V88(17)  | \V120(17) ,
  \V170(1)  = \V28(19)  | \V56(19) ,
  \V154(8)  = \V28(10)  | \V56(10) ,
  \V186(10)  = \V88(16)  | \V120(16) ,
  \V170(0)  = \V28(18)  | \V56(18) ,
  \V186(13)  = \V88(19)  | \V120(19) ,
  \V186(12)  = \V88(18)  | \V120(18) ,
  \V202(3)  = \V88(25)  | \V120(25) ,
  \V186(15)  = \V88(21)  | \V120(21) ,
  \V202(2)  = \V88(24)  | \V120(24) ,
  \V186(14)  = \V88(20)  | \V120(20) ,
  \V202(5)  = \V88(27)  | \V120(27) ,
  \V170(7)  = \V28(25)  | \V56(25) ,
  \V202(4)  = \V88(26)  | \V120(26) ,
  \V170(6)  = \V28(24)  | \V56(24) ,
  \V170(9)  = \V28(27)  | \V56(27) ,
  \V170(8)  = \V28(26)  | \V56(26) ,
  \V202(1)  = \V88(23)  | \V120(23) ,
  \V202(0)  = \V88(22)  | \V120(22) ;
endmodule

