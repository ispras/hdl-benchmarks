module cascade (midas_macys, kappa_rufus_outwire);
  input midas_macys;
  output kappa_rufus_outwire;
endmodule
