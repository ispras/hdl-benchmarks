module bitwise_and_4_1_1(a, b, c);
  input [3:0] a;
  input b;
  output c;
  assign c = a & b;
endmodule
