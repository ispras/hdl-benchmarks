//
// Conformal-LEC Version 15.10-d184 ( 07-Aug-2015) ( 64 bit executable)
//
module test ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 );
input 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 ;
output 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 ;

wire 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 , 
    n545 , 
    n546 , 
    n547 , 
    n548 , 
    n549 , 
    n550 , 
    n551 , 
    n552 , 
    n553 , 
    n554 ;
wire n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , 
     n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , 
     n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , 
     n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , 
     n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , 
     n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , 
     n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , 
     n49828 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , 
     n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , 
     n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , 
     n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , 
     n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , 
     n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , 
     n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , 
     n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , 
     n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , 
     n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , 
     n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , 
     n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , 
     n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n49956 , n683 , 
     n684 , n685 , n686 , n687 , n49962 , n689 , n49964 , n691 , n692 , n693 , 
     n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , 
     n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , 
     n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , 
     n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , 
     n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , 
     n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , 
     n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n50037 , 
     n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n50047 , 
     n774 , n50049 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , 
     n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , 
     n794 , n795 , n796 , n50071 , n798 , n50073 , n800 , n50075 , n50076 , n803 , 
     n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n50086 , n50087 , 
     n50088 , n50089 , n50090 , n50091 , n818 , n50093 , n820 , n50095 , n50096 , n823 , 
     n824 , n50099 , n826 , n50101 , n50102 , n829 , n50104 , n50105 , n832 , n833 , 
     n50108 , n50109 , n836 , n50111 , n50112 , n839 , n840 , n50115 , n50116 , n843 , 
     n50118 , n845 , n50120 , n50121 , n848 , n50123 , n850 , n50125 , n852 , n50127 , 
     n50128 , n50129 , n50130 , n50131 , n858 , n50133 , n50134 , n861 , n862 , n863 , 
     n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n50147 , 
     n874 , n50149 , n50150 , n877 , n50152 , n50153 , n50154 , n881 , n50156 , n50157 , 
     n884 , n50159 , n50160 , n50161 , n50162 , n889 , n50164 , n50165 , n892 , n50167 , 
     n50168 , n50169 , n896 , n50171 , n50172 , n899 , n50174 , n50175 , n902 , n50177 , 
     n904 , n50179 , n906 , n50181 , n908 , n909 , n50184 , n911 , n912 , n913 , 
     n914 , n50189 , n916 , n50191 , n918 , n919 , n50194 , n921 , n922 , n923 , 
     n50198 , n925 , n926 , n50201 , n928 , n50203 , n50204 , n50205 , n50206 , n50207 , 
     n50208 , n50209 , n50210 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , 
     n944 , n50219 , n946 , n50221 , n50222 , n949 , n50224 , n50225 , n50226 , n50227 , 
     n50228 , n955 , n50230 , n957 , n50232 , n50233 , n960 , n50235 , n50236 , n50237 , 
     n964 , n50239 , n50240 , n967 , n50242 , n50243 , n970 , n50245 , n50246 , n50247 , 
     n50248 , n50249 , n976 , n50251 , n50252 , n979 , n980 , n981 , n982 , n983 , 
     n984 , n50259 , n986 , n50261 , n50262 , n50263 , n50264 , n50265 , n992 , n50267 , 
     n50268 , n995 , n50270 , n997 , n50272 , n50273 , n1000 , n50275 , n50276 , n1003 , 
     n50278 , n50279 , n1006 , n50281 , n50282 , n50283 , n1010 , n1011 , n50286 , n1013 , 
     n1014 , n1015 , n1016 , n1017 , n50292 , n50293 , n50294 , n1021 , n50296 , n50297 , 
     n50298 , n50299 , n50300 , n1027 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , 
     n1034 , n1035 , n1036 , n50311 , n1038 , n1039 , n1040 , n1041 , n1042 , n50317 , 
     n1044 , n1045 , n1046 , n50321 , n50322 , n1049 , n50324 , n50325 , n50326 , n50327 , 
     n1054 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , 
     n1062 , n50339 , n50340 , n1065 , n1066 , n1067 , n1068 , n1069 , n50346 , n50347 , 
     n50348 , n50349 , n50350 , n1075 , n1076 , n50353 , n50354 , n50355 , n50356 , n50357 , 
     n1082 , n50359 , n50360 , n1085 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , 
     n50368 , n50369 , n50370 , n1095 , n50372 , n50373 , n50374 , n1099 , n1100 , n50377 , 
     n1102 , n50379 , n50380 , n50381 , n1106 , n1107 , n50384 , n50385 , n50386 , n50387 , 
     n50388 , n1113 , n50390 , n1115 , n1116 , n50393 , n50394 , n50395 , n50396 , n50397 , 
     n50398 , n1123 , n1124 , n50401 , n1126 , n50403 , n50404 , n50405 , n50406 , n50407 , 
     n50408 , n50409 , n50410 , n50411 , n1136 , n50413 , n50414 , n50415 , n50416 , n50417 , 
     n1142 , n50419 , n50420 , n1145 , n50422 , n50423 , n1148 , n50425 , n50426 , n50427 , 
     n50428 , n50429 , n1154 , n50431 , n50432 , n1157 , n50434 , n50435 , n1160 , n50437 , 
     n50438 , n50439 , n50440 , n50441 , n1166 , n50443 , n50444 , n1169 , n1170 , n50447 , 
     n1172 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , 
     n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , 
     n1177 , n1178 , n1179 , n1180 , n50472 , n1182 , n50474 , n50475 , n50476 , n1186 , 
     n50478 , n1188 , n1189 , n50481 , n1191 , n50483 , n1193 , n50485 , n50486 , n1196 , 
     n1197 , n1198 , n50490 , n50491 , n1201 , n50493 , n50494 , n50495 , n1205 , n50497 , 
     n1207 , n50499 , n50500 , n1210 , n1211 , n50503 , n1213 , n50505 , n50506 , n50507 , 
     n50508 , n1218 , n50510 , n1220 , n50512 , n50513 , n50514 , n1224 , n1225 , n50517 , 
     n50518 , n50519 , n50520 , n50521 , n1231 , n50523 , n50524 , n50525 , n1235 , n50527 , 
     n50528 , n50529 , n1239 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n1246 , 
     n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n1255 , n1256 , 
     n1257 , n1258 , n50550 , n50551 , n50552 , n50553 , n1263 , n50555 , n50556 , n50557 , 
     n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n1273 , n50565 , n1275 , n1276 , 
     n50568 , n1278 , n50570 , n1280 , n1281 , n50573 , n1283 , n50575 , n50576 , n1286 , 
     n50578 , n50579 , n1289 , n1290 , n1291 , n1292 , n50584 , n1294 , n1295 , n50587 , 
     n50588 , n50589 , n1299 , n50591 , n1301 , n1302 , n50594 , n50595 , n1305 , n50597 , 
     n50598 , n50599 , n1309 , n50601 , n1311 , n50603 , n50604 , n1314 , n50606 , n50607 , 
     n50608 , n1318 , n50610 , n50611 , n1321 , n50613 , n50614 , n50615 , n1325 , n50617 , 
     n50618 , n50619 , n1329 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , 
     n50628 , n1338 , n1339 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , 
     n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n1356 , 
     n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n50657 , 
     n1367 , n1368 , n1369 , n1370 , n1371 , n50663 , n1373 , n50665 , n50666 , n1376 , 
     n50668 , n50669 , n1379 , n50671 , n1381 , n50673 , n50674 , n1384 , n50676 , n50677 , 
     n1387 , n50679 , n1389 , n50681 , n50682 , n50683 , n50684 , n1394 , n50686 , n50687 , 
     n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n1403 , n1404 , n50696 , n50697 , 
     n50698 , n1408 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n1416 , 
     n1417 , n1418 , n50710 , n1420 , n50712 , n50713 , n50714 , n1424 , n50716 , n50717 , 
     n50718 , n50719 , n50720 , n50721 , n1431 , n50723 , n50724 , n50725 , n50726 , n50727 , 
     n1437 , n50729 , n50730 , n1440 , n50732 , n1442 , n50734 , n50735 , n50736 , n50737 , 
     n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n1453 , n50745 , n50746 , n50747 , 
     n50748 , n50749 , n1459 , n50751 , n50752 , n50753 , n50754 , n1464 , n50756 , n50757 , 
     n1467 , n50759 , n50760 , n1470 , n50762 , n1472 , n1473 , n50765 , n50766 , n50767 , 
     n50768 , n50769 , n50770 , n1480 , n50772 , n50773 , n1483 , n1484 , n50776 , n1486 , 
     n50778 , n1488 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , 
     n1497 , n50789 , n50790 , n50791 , n1501 , n1502 , n1503 , n1504 , n50796 , n1506 , 
     n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n1515 , n1516 , 
     n50808 , n1518 , n50810 , n50811 , n1521 , n50813 , n50814 , n50815 , n50816 , n50817 , 
     n50818 , n1528 , n1529 , n1530 , n1531 , n50823 , n1533 , n50825 , n50826 , n1536 , 
     n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , 
     n50838 , n50839 , n50840 , n50841 , n50842 , n1552 , n50844 , n1554 , n1555 , n50847 , 
     n50848 , n50849 , n1559 , n50851 , n50852 , n50853 , n50854 , n1564 , n1565 , n50857 , 
     n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , 
     n50868 , n50869 , n50870 , n1580 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , 
     n1587 , n50879 , n50880 , n1590 , n50882 , n50883 , n50884 , n1594 , n50886 , n1596 , 
     n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n1604 , n50896 , n1606 , 
     n50898 , n50899 , n1609 , n50901 , n50902 , n1612 , n1613 , n50905 , n1615 , n50907 , 
     n1617 , n50909 , n50910 , n50911 , n1621 , n50913 , n50914 , n1624 , n50916 , n50917 , 
     n1627 , n50919 , n50920 , n1630 , n50922 , n1632 , n1633 , n50925 , n50926 , n1636 , 
     n50928 , n1638 , n50930 , n1640 , n1641 , n50933 , n50934 , n1644 , n50936 , n50937 , 
     n50938 , n50939 , n1649 , n50941 , n50942 , n50943 , n1653 , n50945 , n50946 , n50947 , 
     n1657 , n1658 , n1659 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , 
     n50958 , n1668 , n1669 , n50961 , n50962 , n50963 , n50964 , n50965 , n1675 , n50967 , 
     n50968 , n1678 , n50970 , n1680 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , 
     n50978 , n50979 , n50980 , n50981 , n50982 , n1692 , n1693 , n50985 , n1695 , n1696 , 
     n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n50995 , n50996 , n50997 , 
     n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , 
     n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n1720 , 
     n51018 , n51019 , n51020 , n1724 , n51022 , n51023 , n1727 , n51025 , n51026 , n51027 , 
     n51028 , n51029 , n51030 , n51031 , n1735 , n51033 , n51034 , n1738 , n51036 , n51037 , 
     n51038 , n51039 , n51040 , n51041 , n1745 , n51043 , n51044 , n51045 , n51046 , n51047 , 
     n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n1754 , n51055 , n51056 , n51057 , 
     n1758 , n51059 , n51060 , n1761 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , 
     n1768 , n1769 , n51070 , n51071 , n51072 , n51073 , n1774 , n51075 , n51076 , n1777 , 
     n51078 , n51079 , n1780 , n1781 , n1782 , n51083 , n51084 , n1785 , n51086 , n51087 , 
     n1788 , n51089 , n51090 , n51091 , n51092 , n1793 , n51094 , n1795 , n51096 , n51097 , 
     n1798 , n1799 , n51100 , n1801 , n51102 , n51103 , n1804 , n51105 , n51106 , n1807 , 
     n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , 
     n1818 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , 
     n51128 , n51129 , n51130 , n51131 , n51132 , n1833 , n51134 , n51135 , n51136 , n51137 , 
     n51138 , n1839 , n51140 , n1840 , n51142 , n51143 , n51144 , n1844 , n51146 , n51147 , 
     n51148 , n51149 , n51150 , n51151 , n51152 , n1852 , n51154 , n51155 , n1855 , n51157 , 
     n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n1866 , 
     n1867 , n1868 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , 
     n51178 , n51179 , n51180 , n51181 , n1881 , n51183 , n51184 , n51185 , n51186 , n51187 , 
     n51188 , n51189 , n51190 , n51191 , n51192 , n1892 , n51194 , n51195 , n51196 , n51197 , 
     n51198 , n1898 , n51200 , n51201 , n1901 , n51203 , n51204 , n1904 , n51206 , n51207 , 
     n1907 , n51209 , n1909 , n51211 , n51212 , n51213 , n1913 , n51215 , n51216 , n51217 , 
     n51218 , n51219 , n51220 , n51221 , n1921 , n1922 , n51224 , n51225 , n51226 , n51227 , 
     n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n1933 , n51235 , n51236 , n51237 , 
     n1937 , n51239 , n51240 , n51241 , n1941 , n51243 , n51244 , n51245 , n51246 , n51247 , 
     n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n1955 , n1956 , 
     n51258 , n51259 , n1959 , n51261 , n1961 , n1962 , n51264 , n51265 , n51266 , n1966 , 
     n51268 , n51269 , n51270 , n51271 , n1971 , n51273 , n51274 , n51275 , n51276 , n51277 , 
     n51278 , n51279 , n51280 , n51281 , n1981 , n1982 , n51284 , n1983 , n51286 , n1985 , 
     n51288 , n1987 , n1988 , n51291 , n51292 , n1991 , n1992 , n51295 , n51296 , n1995 , 
     n51298 , n1997 , n51300 , n51301 , n51302 , n51303 , n51304 , n2003 , n51306 , n51307 , 
     n2006 , n51309 , n2008 , n51311 , n2010 , n2011 , n51314 , n51315 , n2014 , n2015 , 
     n51318 , n51319 , n2018 , n51321 , n51322 , n2021 , n51324 , n2023 , n51326 , n2025 , 
     n51328 , n51329 , n51330 , n51331 , n2030 , n51333 , n51334 , n2033 , n2034 , n51337 , 
     n51338 , n2037 , n2038 , n51341 , n51342 , n51343 , n51344 , n2043 , n51346 , n51347 , 
     n51348 , n51349 , n2048 , n51351 , n51352 , n2051 , n51354 , n51355 , n51356 , n51357 , 
     n2056 , n51359 , n51360 , n2059 , n2060 , n51363 , n51364 , n2063 , n2064 , n51367 , 
     n51368 , n2067 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , 
     n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n2082 , n51385 , n51386 , n51387 , 
     n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , 
     n51398 , n2097 , n51400 , n2099 , n2100 , n51403 , n2101 , n51405 , n51406 , n51407 , 
     n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n2111 , n51415 , n51416 , n51417 , 
     n51418 , n51419 , n51420 , n2118 , n51422 , n51423 , n2121 , n2122 , n51426 , n51427 , 
     n2125 , n51429 , n51430 , n51431 , n51432 , n51433 , n2130 , n2131 , n51436 , n51437 , 
     n51438 , n51439 , n51440 , n51441 , n2138 , n51443 , n51444 , n2141 , n51446 , n51447 , 
     n2144 , n2145 , n51450 , n2147 , n2148 , n2149 , n2150 , n51455 , n2152 , n2153 , 
     n51458 , n51459 , n51460 , n2157 , n51462 , n51463 , n51464 , n51465 , n2162 , n51467 , 
     n51468 , n2165 , n51470 , n51471 , n2168 , n51473 , n51474 , n2171 , n51476 , n51477 , 
     n2174 , n51479 , n51480 , n51481 , n51482 , n51483 , n2180 , n51485 , n51486 , n2183 , 
     n51488 , n51489 , n2186 , n51491 , n51492 , n51493 , n51494 , n2191 , n51496 , n51497 , 
     n51498 , n51499 , n2196 , n2197 , n2198 , n2199 , n2200 , n51505 , n51506 , n51507 , 
     n51508 , n2205 , n2206 , n51511 , n51512 , n2209 , n51514 , n51515 , n51516 , n51517 , 
     n2214 , n51519 , n51520 , n2217 , n2218 , n51523 , n2220 , n2221 , n2222 , n2223 , 
     n51528 , n51529 , n51530 , n2227 , n51532 , n51533 , n2230 , n51535 , n2232 , n2233 , 
     n2234 , n51539 , n51540 , n51541 , n51542 , n2239 , n51544 , n2241 , n2242 , n2243 , 
     n51548 , n51549 , n51550 , n51551 , n51552 , n2249 , n51554 , n51555 , n2252 , n2253 , 
     n2254 , n2255 , n51560 , n2257 , n51562 , n51563 , n51564 , n51565 , n2262 , n51567 , 
     n51568 , n2265 , n51570 , n2267 , n51572 , n51573 , n51574 , n2271 , n51576 , n2273 , 
     n51578 , n51579 , n51580 , n2277 , n51582 , n2279 , n51584 , n51585 , n2282 , n51587 , 
     n51588 , n2285 , n51590 , n2287 , n51592 , n2289 , n51594 , n51595 , n51596 , n51597 , 
     n51598 , n51599 , n2293 , n51601 , n51602 , n51603 , n2297 , n51605 , n51606 , n51607 , 
     n2301 , n51609 , n51610 , n51611 , n2305 , n51613 , n51614 , n51615 , n2309 , n51617 , 
     n51618 , n51619 , n51620 , n2314 , n2315 , n51623 , n51624 , n51625 , n2319 , n2320 , 
     n51628 , n2322 , n2323 , n2324 , n51632 , n2326 , n51634 , n2328 , n2329 , n2330 , 
     n2331 , n2332 , n2333 , n2334 , n2335 , n51643 , n2337 , n2338 , n2339 , n2340 , 
     n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , 
     n2351 , n2352 , n2353 , n51661 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , 
     n2361 , n2362 , n2363 , n2364 , n51672 , n2366 , n51674 , n51675 , n2369 , n2370 , 
     n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , 
     n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , 
     n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , 
     n51708 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , 
     n2411 , n2412 , n2413 , n2414 , n2415 , n51723 , n2417 , n2418 , n51726 , n2420 , 
     n2421 , n2422 , n2423 , n51731 , n2425 , n51733 , n51734 , n2428 , n51736 , n51737 , 
     n2431 , n51739 , n51740 , n51741 , n2435 , n51743 , n51744 , n51745 , n2439 , n51747 , 
     n51748 , n2442 , n51750 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n51757 , 
     n2451 , n2452 , n51760 , n51761 , n2455 , n51763 , n51764 , n2458 , n51766 , n51767 , 
     n2461 , n51769 , n51770 , n2464 , n51772 , n2466 , n2467 , n2468 , n2469 , n2470 , 
     n2471 , n2472 , n2473 , n2474 , n51782 , n2476 , n2477 , n2478 , n51786 , n2480 , 
     n51788 , n51789 , n2483 , n51791 , n51792 , n51793 , n51794 , n2488 , n51796 , n51797 , 
     n2491 , n51799 , n51800 , n2494 , n51802 , n51803 , n2497 , n51805 , n51806 , n51807 , 
     n51808 , n51809 , n2503 , n51811 , n51812 , n51813 , n51814 , n51815 , n2509 , n2510 , 
     n51818 , n2512 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n2520 , 
     n2521 , n51829 , n51830 , n2524 , n51832 , n51833 , n51834 , n2528 , n2529 , n2530 , 
     n2531 , n51839 , n2533 , n51841 , n51842 , n2536 , n51844 , n51845 , n2539 , n51847 , 
     n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n2547 , n51855 , n51856 , n2550 , 
     n51858 , n2552 , n2553 , n2554 , n51862 , n2556 , n51864 , n2558 , n51866 , n2560 , 
     n51868 , n2562 , n2563 , n2564 , n2565 , n2566 , n51874 , n51875 , n2569 , n51877 , 
     n51878 , n51879 , n51880 , n51881 , n2575 , n51883 , n51884 , n2578 , n51886 , n2580 , 
     n2581 , n2582 , n51890 , n2584 , n51892 , n51893 , n2587 , n51895 , n51896 , n2590 , 
     n2591 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , 
     n51908 , n2602 , n2603 , n51911 , n51912 , n2606 , n51914 , n51915 , n2609 , n2610 , 
     n2611 , n2612 , n2613 , n51921 , n51922 , n51923 , n51924 , n2618 , n51926 , n51927 , 
     n2621 , n51929 , n51930 , n2624 , n2625 , n51933 , n2627 , n51935 , n2629 , n51937 , 
     n51938 , n51939 , n51940 , n51941 , n2635 , n2636 , n51944 , n51945 , n51946 , n2640 , 
     n51948 , n2642 , n2643 , n51951 , n2645 , n51953 , n51954 , n51955 , n51956 , n2650 , 
     n51958 , n51959 , n51960 , n51961 , n51962 , n2656 , n2657 , n51965 , n2659 , n51967 , 
     n51968 , n51969 , n51970 , n51971 , n2665 , n51973 , n51974 , n51975 , n51976 , n51977 , 
     n2671 , n2672 , n2673 , n51981 , n2675 , n51983 , n2677 , n51985 , n51986 , n51987 , 
     n51988 , n2682 , n51990 , n51991 , n51992 , n51993 , n2687 , n51995 , n51996 , n2690 , 
     n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n2698 , n52006 , n52007 , 
     n2701 , n52009 , n2703 , n52011 , n52012 , n2706 , n52014 , n52015 , n2709 , n52017 , 
     n52018 , n52019 , n52020 , n52021 , n52022 , n2716 , n2717 , n52025 , n52026 , n52027 , 
     n2721 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n2728 , n52036 , n52037 , 
     n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , 
     n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n2748 , n2749 , n52057 , 
     n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , 
     n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , 
     n52078 , n52079 , n52080 , n52081 , n2775 , n52083 , n52084 , n52085 , n52086 , n52087 , 
     n52088 , n52089 , n52090 , n52091 , n2785 , n52093 , n52094 , n52095 , n52096 , n52097 , 
     n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n2797 , n52105 , n52106 , n52107 , 
     n52108 , n52109 , n52110 , n52111 , n52112 , n2806 , n52114 , n52115 , n52116 , n52117 , 
     n52118 , n52119 , n52120 , n52121 , n52122 , n2816 , n52124 , n52125 , n52126 , n2820 , 
     n52128 , n52129 , n2823 , n52131 , n52132 , n52133 , n2827 , n52135 , n52136 , n2830 , 
     n2831 , n52139 , n52140 , n2834 , n52142 , n2836 , n52144 , n52145 , n52146 , n2840 , 
     n2841 , n52149 , n52150 , n52151 , n52152 , n2846 , n52154 , n52155 , n2849 , n2850 , 
     n52158 , n2852 , n2853 , n52161 , n52162 , n52163 , n2857 , n52165 , n52166 , n2860 , 
     n52168 , n2862 , n52170 , n52171 , n2865 , n52173 , n52174 , n52175 , n52176 , n52177 , 
     n52178 , n52179 , n2873 , n52181 , n52182 , n52183 , n52184 , n52185 , n2879 , n52187 , 
     n52188 , n52189 , n2883 , n2884 , n52192 , n52193 , n52194 , n2888 , n2889 , n52197 , 
     n52198 , n52199 , n52200 , n52201 , n52202 , n2896 , n2897 , n52205 , n52206 , n2900 , 
     n52208 , n52209 , n52210 , n52211 , n52212 , n2906 , n52214 , n52215 , n52216 , n52217 , 
     n2911 , n52219 , n52220 , n52221 , n52222 , n2916 , n52224 , n52225 , n2919 , n52227 , 
     n52228 , n52229 , n52230 , n2924 , n52232 , n52233 , n52234 , n2928 , n52236 , n52237 , 
     n2931 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , 
     n2941 , n52249 , n52250 , n52251 , n52252 , n2946 , n2947 , n52255 , n2949 , n2950 , 
     n52258 , n2952 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , 
     n52268 , n2956 , n52270 , n52271 , n52272 , n2960 , n52274 , n2962 , n52276 , n52277 , 
     n2965 , n52279 , n52280 , n52281 , n52282 , n52283 , n2969 , n52285 , n2971 , n52287 , 
     n52288 , n52289 , n2975 , n52291 , n52292 , n2978 , n52294 , n52295 , n52296 , n52297 , 
     n52298 , n52299 , n52300 , n52301 , n52302 , n2988 , n52304 , n2990 , n2991 , n2992 , 
     n2993 , n52309 , n52310 , n52311 , n2997 , n52313 , n52314 , n52315 , n52316 , n52317 , 
     n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n3010 , n52326 , n52327 , 
     n52328 , n3014 , n52330 , n3016 , n52332 , n52333 , n52334 , n3020 , n3021 , n52337 , 
     n52338 , n52339 , n52340 , n52341 , n3027 , n52343 , n52344 , n52345 , n52346 , n52347 , 
     n52348 , n3032 , n52350 , n52351 , n3034 , n3035 , n52354 , n52355 , n52356 , n52357 , 
     n52358 , n52359 , n52360 , n3043 , n3044 , n3045 , n3046 , n52365 , n52366 , n52367 , 
     n52368 , n3051 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n3059 , 
     n52378 , n52379 , n3062 , n3063 , n52382 , n3065 , n52384 , n52385 , n52386 , n52387 , 
     n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , 
     n52398 , n52399 , n3082 , n52401 , n52402 , n3085 , n52404 , n52405 , n52406 , n52407 , 
     n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n3097 , n52417 , 
     n52418 , n52419 , n52420 , n3102 , n52422 , n52423 , n52424 , n52425 , n3107 , n52427 , 
     n52428 , n3110 , n52430 , n52431 , n52432 , n52433 , n52434 , n3116 , n52436 , n52437 , 
     n52438 , n3120 , n3121 , n52441 , n52442 , n52443 , n52444 , n3126 , n52446 , n3128 , 
     n3129 , n52449 , n52450 , n3132 , n52452 , n3134 , n3135 , n52455 , n3137 , n52457 , 
     n52458 , n52459 , n3141 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , 
     n52468 , n52469 , n3151 , n52471 , n52472 , n3154 , n52474 , n52475 , n52476 , n3158 , 
     n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n3166 , n52486 , n52487 , 
     n52488 , n52489 , n52490 , n52491 , n52492 , n3174 , n52494 , n52495 , n3177 , n52497 , 
     n52498 , n52499 , n3181 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , 
     n3189 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n3196 , n52516 , n52517 , 
     n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n3205 , n52525 , n52526 , n3208 , 
     n52528 , n52529 , n52530 , n3212 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , 
     n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , 
     n3229 , n3230 , n52550 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , 
     n3239 , n52559 , n3241 , n52561 , n3243 , n52563 , n52564 , n52565 , n52566 , n52567 , 
     n3249 , n52569 , n52570 , n3252 , n3253 , n52573 , n3255 , n3256 , n3257 , n3258 , 
     n52578 , n52579 , n3261 , n52581 , n52582 , n52583 , n52584 , n3266 , n3267 , n52587 , 
     n3269 , n3270 , n3271 , n3272 , n52592 , n52593 , n52594 , n3276 , n52596 , n52597 , 
     n52598 , n52599 , n3281 , n52601 , n52602 , n52603 , n52604 , n3286 , n52606 , n52607 , 
     n3289 , n3290 , n52610 , n3292 , n3293 , n3294 , n52614 , n52615 , n52616 , n52617 , 
     n52618 , n52619 , n52620 , n52621 , n52622 , n3304 , n52624 , n52625 , n52626 , n52627 , 
     n52628 , n52629 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , 
     n3319 , n3320 , n3321 , n52641 , n52642 , n52643 , n52644 , n52645 , n3327 , n52647 , 
     n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n3337 , n3338 , 
     n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n3346 , n3347 , n52667 , 
     n52668 , n52669 , n52670 , n3352 , n52672 , n52673 , n52674 , n3356 , n52676 , n52677 , 
     n52678 , n52679 , n52680 , n52681 , n3363 , n52683 , n52684 , n3366 , n3367 , n52687 , 
     n3369 , n52689 , n52690 , n52691 , n52692 , n52693 , n3375 , n3376 , n3377 , n3378 , 
     n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , 
     n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n52717 , 
     n52718 , n3400 , n52720 , n52721 , n52722 , n3404 , n3405 , n52725 , n3407 , n3408 , 
     n3409 , n3410 , n52730 , n52731 , n52732 , n52733 , n3415 , n3416 , n52736 , n52737 , 
     n52738 , n3420 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , 
     n3429 , n3430 , n52750 , n3432 , n52752 , n52753 , n52754 , n52755 , n52756 , n3438 , 
     n52758 , n52759 , n3441 , n52761 , n3443 , n52763 , n52764 , n52765 , n52766 , n52767 , 
     n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n3458 , 
     n52778 , n52779 , n52780 , n3462 , n52782 , n52783 , n52784 , n3466 , n52786 , n52787 , 
     n3469 , n3470 , n3471 , n3472 , n52792 , n52793 , n52794 , n3476 , n52796 , n52797 , 
     n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n3487 , n3488 , 
     n3489 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n3497 , n52817 , 
     n52818 , n3500 , n52820 , n52821 , n52822 , n52823 , n3505 , n3506 , n52826 , n3508 , 
     n3509 , n3510 , n3511 , n3512 , n52832 , n52833 , n52834 , n3516 , n52836 , n52837 , 
     n3519 , n3520 , n3521 , n52841 , n52842 , n52843 , n52844 , n3526 , n52846 , n52847 , 
     n52848 , n3530 , n52850 , n52851 , n52852 , n3534 , n52854 , n3536 , n52856 , n52857 , 
     n3539 , n3540 , n3541 , n52861 , n52862 , n52863 , n3545 , n3546 , n52866 , n52867 , 
     n52868 , n3550 , n52870 , n52871 , n52872 , n52873 , n3555 , n52875 , n52876 , n52877 , 
     n52878 , n3560 , n52880 , n52881 , n3563 , n3564 , n52884 , n52885 , n52886 , n3568 , 
     n52888 , n52889 , n52890 , n52891 , n3573 , n52893 , n52894 , n52895 , n52896 , n3578 , 
     n52898 , n52899 , n52900 , n52901 , n3583 , n52903 , n52904 , n3586 , n3587 , n52907 , 
     n3589 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n3598 , 
     n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , 
     n52928 , n52929 , n3611 , n3612 , n3613 , n3614 , n3615 , n52935 , n52936 , n3618 , 
     n52938 , n52939 , n3621 , n52941 , n52942 , n52943 , n52944 , n52945 , n3627 , n52947 , 
     n52948 , n3630 , n52950 , n3632 , n3633 , n3634 , n52954 , n52955 , n3637 , n52957 , 
     n52958 , n3640 , n52960 , n52961 , n3643 , n52963 , n52964 , n52965 , n3647 , n52967 , 
     n3649 , n3650 , n3651 , n3652 , n52972 , n3654 , n3655 , n3656 , n3657 , n3658 , 
     n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , 
     n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , 
     n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , 
     n3689 , n53009 , n53010 , n3692 , n53012 , n53013 , n3695 , n53015 , n53016 , n53017 , 
     n3699 , n53019 , n53020 , n3702 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , 
     n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , 
     n53038 , n53039 , n53040 , n3722 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , 
     n53048 , n3730 , n3731 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , 
     n3739 , n53059 , n53060 , n53061 , n3743 , n53063 , n53064 , n53065 , n53066 , n3748 , 
     n53068 , n53069 , n3751 , n53071 , n3753 , n53073 , n53074 , n3756 , n53076 , n53077 , 
     n53078 , n53079 , n53080 , n53081 , n3763 , n53083 , n53084 , n3766 , n53086 , n3768 , 
     n53088 , n53089 , n3771 , n53091 , n53092 , n3774 , n53094 , n53095 , n3777 , n3778 , 
     n53098 , n53099 , n3781 , n3782 , n3783 , n53103 , n53104 , n53105 , n53106 , n3788 , 
     n53108 , n53109 , n53110 , n53111 , n3792 , n53113 , n53114 , n53115 , n53116 , n3797 , 
     n53118 , n53119 , n3800 , n3801 , n53122 , n53123 , n3804 , n3805 , n3806 , n53127 , 
     n53128 , n53129 , n3810 , n53131 , n53132 , n53133 , n3814 , n53135 , n53136 , n53137 , 
     n53138 , n53139 , n53140 , n3821 , n3822 , n53143 , n53144 , n53145 , n3826 , n53147 , 
     n53148 , n3829 , n53150 , n53151 , n53152 , n53153 , n53154 , n3835 , n3836 , n53157 , 
     n53158 , n53159 , n3840 , n53161 , n53162 , n53163 , n53164 , n3845 , n53166 , n53167 , 
     n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n3854 , n53175 , n53176 , n53177 , 
     n53178 , n3859 , n53180 , n53181 , n53182 , n3863 , n53184 , n53185 , n53186 , n3867 , 
     n53188 , n53189 , n3870 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , 
     n53198 , n53199 , n53200 , n53201 , n3882 , n53203 , n3884 , n53205 , n53206 , n53207 , 
     n53208 , n53209 , n3890 , n53211 , n53212 , n53213 , n3894 , n53215 , n53216 , n3897 , 
     n53218 , n53219 , n53220 , n53221 , n3902 , n53223 , n53224 , n3905 , n53226 , n3907 , 
     n53228 , n3909 , n53230 , n53231 , n3912 , n53233 , n53234 , n3915 , n53236 , n53237 , 
     n53238 , n3919 , n3920 , n53241 , n53242 , n3923 , n53244 , n53245 , n3926 , n53247 , 
     n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n3937 , 
     n53258 , n53259 , n3940 , n3941 , n53262 , n3943 , n3944 , n3945 , n3946 , n53267 , 
     n53268 , n53269 , n53270 , n3951 , n53272 , n3953 , n53274 , n53275 , n53276 , n53277 , 
     n3958 , n53279 , n53280 , n3961 , n53282 , n3963 , n53284 , n3965 , n3966 , n53287 , 
     n53288 , n53289 , n3970 , n3971 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , 
     n3978 , n53299 , n53300 , n53301 , n3982 , n53303 , n3984 , n53305 , n53306 , n3987 , 
     n53308 , n53309 , n53310 , n53311 , n3992 , n53313 , n53314 , n53315 , n53316 , n3997 , 
     n3998 , n53319 , n53320 , n4001 , n4002 , n4003 , n53324 , n53325 , n4006 , n4007 , 
     n4008 , n53329 , n53330 , n4011 , n4012 , n4013 , n53334 , n53335 , n4016 , n4017 , 
     n4018 , n53339 , n53340 , n53341 , n53342 , n4023 , n53344 , n53345 , n53346 , n53347 , 
     n4028 , n4029 , n53350 , n53351 , n53352 , n4033 , n53354 , n53355 , n4036 , n4037 , 
     n53358 , n53359 , n4040 , n4041 , n4042 , n53363 , n53364 , n53365 , n53366 , n53367 , 
     n53368 , n4049 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , 
     n53378 , n53379 , n53380 , n4061 , n53382 , n53383 , n4064 , n4065 , n53386 , n53387 , 
     n53388 , n53389 , n4070 , n53391 , n4072 , n4073 , n53394 , n4075 , n53396 , n53397 , 
     n53398 , n4079 , n4080 , n4081 , n53402 , n53403 , n4084 , n53405 , n4086 , n53407 , 
     n53408 , n4089 , n53410 , n4091 , n4092 , n53413 , n53414 , n53415 , n53416 , n53417 , 
     n53418 , n53419 , n53420 , n4101 , n4102 , n53423 , n53424 , n53425 , n53426 , n53427 , 
     n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n4114 , n4115 , n53436 , n53437 , 
     n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n4126 , n53447 , 
     n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n4134 , n4135 , n53456 , n4137 , 
     n4138 , n4139 , n4140 , n4141 , n53462 , n4143 , n53464 , n53465 , n4146 , n4147 , 
     n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , 
     n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , 
     n4168 , n4169 , n4170 , n4171 , n4172 , n53493 , n53494 , n4175 , n53496 , n53497 , 
     n4178 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n4187 , 
     n4188 , n53509 , n4190 , n4191 , n53512 , n53513 , n4194 , n4195 , n4196 , n53517 , 
     n53518 , n53519 , n53520 , n4201 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , 
     n53528 , n53529 , n53530 , n4211 , n53532 , n53533 , n53534 , n53535 , n4216 , n53537 , 
     n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n4224 , n53545 , n4226 , n4227 , 
     n53548 , n4229 , n53550 , n4231 , n4232 , n53553 , n53554 , n53555 , n4235 , n53557 , 
     n53558 , n53559 , n53560 , n4240 , n53562 , n53563 , n53564 , n53565 , n4245 , n53567 , 
     n53568 , n4248 , n53570 , n53571 , n4251 , n4252 , n4253 , n53575 , n53576 , n53577 , 
     n53578 , n4258 , n53580 , n53581 , n4261 , n53583 , n53584 , n53585 , n4265 , n4266 , 
     n53588 , n4268 , n53590 , n53591 , n53592 , n53593 , n53594 , n4274 , n4275 , n4276 , 
     n4277 , n4278 , n53600 , n4280 , n4281 , n4282 , n4283 , n53605 , n4285 , n4286 , 
     n53608 , n4288 , n53610 , n4290 , n53612 , n53613 , n53614 , n53615 , n4295 , n53617 , 
     n53618 , n53619 , n53620 , n4300 , n53622 , n53623 , n53624 , n53625 , n4305 , n53627 , 
     n53628 , n53629 , n53630 , n53631 , n53632 , n4312 , n53634 , n53635 , n4315 , n53637 , 
     n4317 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n4324 , n4325 , n53647 , 
     n53648 , n4328 , n53650 , n53651 , n53652 , n4332 , n53654 , n4334 , n53656 , n53657 , 
     n4337 , n4338 , n53660 , n4340 , n53662 , n4342 , n53664 , n4344 , n53666 , n53667 , 
     n4347 , n53669 , n4349 , n53671 , n53672 , n53673 , n53674 , n53675 , n4355 , n53677 , 
     n53678 , n53679 , n4359 , n53681 , n4361 , n53683 , n53684 , n53685 , n53686 , n4366 , 
     n53688 , n53689 , n53690 , n53691 , n4371 , n53693 , n53694 , n4374 , n53696 , n53697 , 
     n53698 , n53699 , n4379 , n53701 , n4381 , n4382 , n53704 , n53705 , n53706 , n53707 , 
     n53708 , n53709 , n53710 , n53711 , n4391 , n53713 , n53714 , n4394 , n53716 , n53717 , 
     n4397 , n53719 , n4399 , n53721 , n53722 , n4402 , n4403 , n53725 , n4405 , n4406 , 
     n4407 , n4408 , n53730 , n4410 , n4411 , n4412 , n4413 , n53735 , n4415 , n4416 , 
     n4417 , n53739 , n53740 , n4420 , n53742 , n53743 , n4423 , n53745 , n53746 , n4426 , 
     n53748 , n4428 , n53750 , n53751 , n4431 , n4432 , n53754 , n53755 , n4435 , n4436 , 
     n4437 , n53759 , n53760 , n4440 , n4441 , n4442 , n53764 , n53765 , n4445 , n4446 , 
     n4447 , n53769 , n53770 , n53771 , n53772 , n4452 , n53774 , n53775 , n53776 , n53777 , 
     n4457 , n53779 , n53780 , n53781 , n53782 , n4462 , n53784 , n53785 , n4465 , n4466 , 
     n53788 , n53789 , n4469 , n4470 , n4471 , n53793 , n53794 , n53795 , n53796 , n4476 , 
     n4477 , n53799 , n53800 , n53801 , n4481 , n53803 , n53804 , n4484 , n4485 , n4486 , 
     n4487 , n53809 , n4489 , n4490 , n4491 , n4492 , n53814 , n53815 , n4495 , n53817 , 
     n53818 , n4498 , n4499 , n4500 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , 
     n53828 , n53829 , n53830 , n53831 , n4511 , n53833 , n53834 , n4514 , n4515 , n4516 , 
     n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n4525 , n53847 , 
     n53848 , n53849 , n53850 , n53851 , n4531 , n53853 , n53854 , n4534 , n53856 , n53857 , 
     n53858 , n53859 , n53860 , n53861 , n4541 , n53863 , n53864 , n53865 , n53866 , n4546 , 
     n53868 , n4548 , n53870 , n53871 , n53872 , n53873 , n4553 , n53875 , n4555 , n53877 , 
     n53878 , n4558 , n53880 , n53881 , n4561 , n53883 , n53884 , n4564 , n53886 , n53887 , 
     n53888 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , 
     n4577 , n53899 , n53900 , n4580 , n53902 , n53903 , n4583 , n53905 , n53906 , n4586 , 
     n53908 , n53909 , n4589 , n4590 , n53912 , n4592 , n4593 , n4594 , n4595 , n53917 , 
     n53918 , n53919 , n53920 , n4600 , n4601 , n53923 , n4603 , n4604 , n4605 , n4606 , 
     n53928 , n4608 , n4609 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , 
     n4617 , n53939 , n53940 , n53941 , n53942 , n4622 , n53944 , n53945 , n4625 , n53947 , 
     n53948 , n4628 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , 
     n53958 , n53959 , n53960 , n53961 , n53962 , n4642 , n53964 , n4644 , n4645 , n53967 , 
     n4647 , n53969 , n53970 , n53971 , n53972 , n4652 , n53974 , n53975 , n53976 , n53977 , 
     n4657 , n53979 , n4659 , n4660 , n53982 , n4662 , n53984 , n53985 , n53986 , n53987 , 
     n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n4675 , n53997 , 
     n53998 , n4678 , n4679 , n4680 , n54002 , n54003 , n54004 , n54005 , n4685 , n54007 , 
     n4687 , n4688 , n54010 , n54011 , n54012 , n54013 , n54014 , n4694 , n54016 , n54017 , 
     n54018 , n54019 , n4699 , n54021 , n54022 , n4702 , n54024 , n54025 , n4705 , n54027 , 
     n54028 , n4708 , n54030 , n54031 , n54032 , n54033 , n4713 , n54035 , n54036 , n4716 , 
     n4717 , n4718 , n54040 , n54041 , n54042 , n54043 , n4723 , n54045 , n54046 , n54047 , 
     n54048 , n4728 , n54050 , n54051 , n54052 , n4732 , n4733 , n54055 , n4735 , n4736 , 
     n54058 , n4738 , n54060 , n54061 , n54062 , n54063 , n4743 , n54065 , n54066 , n54067 , 
     n4747 , n4748 , n54070 , n54071 , n54072 , n54073 , n4753 , n54075 , n54076 , n54077 , 
     n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n4764 , n54086 , n54087 , 
     n4767 , n4768 , n4769 , n54091 , n54092 , n54093 , n4773 , n4774 , n4775 , n4776 , 
     n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n54105 , n4785 , n54107 , 
     n54108 , n54109 , n54110 , n4790 , n54112 , n4792 , n54114 , n54115 , n4795 , n4796 , 
     n54118 , n4798 , n4799 , n4800 , n4801 , n54123 , n4803 , n4804 , n54126 , n4806 , 
     n54128 , n54129 , n4809 , n4810 , n54132 , n4812 , n54134 , n54135 , n54136 , n54137 , 
     n54138 , n4818 , n54140 , n54141 , n54142 , n54143 , n54144 , n4824 , n4825 , n4826 , 
     n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n54157 , 
     n54158 , n54159 , n4839 , n4840 , n54162 , n4842 , n4843 , n4844 , n4845 , n54167 , 
     n54168 , n54169 , n54170 , n4850 , n4851 , n54173 , n4853 , n54175 , n54176 , n54177 , 
     n54178 , n54179 , n54180 , n54181 , n4861 , n4862 , n54184 , n54185 , n54186 , n4866 , 
     n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , 
     n54198 , n4878 , n54200 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , 
     n4887 , n4888 , n54210 , n54211 , n4891 , n54213 , n54214 , n54215 , n4895 , n4896 , 
     n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n4905 , n54227 , 
     n54228 , n4908 , n54230 , n54231 , n54232 , n4912 , n54234 , n54235 , n54236 , n54237 , 
     n4917 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n4925 , n4926 , 
     n54248 , n4928 , n54250 , n54251 , n4931 , n54253 , n54254 , n54255 , n54256 , n54257 , 
     n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n4944 , n54266 , n54267 , 
     n54268 , n54269 , n4949 , n54271 , n54272 , n54273 , n4953 , n4954 , n54276 , n4956 , 
     n4957 , n4958 , n4959 , n54281 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , 
     n4967 , n4968 , n4969 , n54291 , n4971 , n4972 , n54294 , n4974 , n4975 , n4976 , 
     n4977 , n54299 , n54300 , n54301 , n54302 , n4982 , n54304 , n54305 , n54306 , n54307 , 
     n54308 , n54309 , n54310 , n54311 , n4991 , n4992 , n54314 , n54315 , n54316 , n54317 , 
     n4997 , n54319 , n54320 , n54321 , n54322 , n5002 , n5003 , n54325 , n54326 , n54327 , 
     n54328 , n5008 , n54330 , n54331 , n54332 , n54333 , n5013 , n5014 , n54336 , n54337 , 
     n54338 , n54339 , n5019 , n54341 , n54342 , n54343 , n54344 , n5024 , n5025 , n54347 , 
     n54348 , n54349 , n5029 , n54351 , n54352 , n5032 , n5033 , n5034 , n5035 , n54357 , 
     n54358 , n54359 , n5039 , n54361 , n54362 , n54363 , n54364 , n54365 , n5045 , n54367 , 
     n5047 , n5048 , n54370 , n5050 , n54372 , n54373 , n5053 , n54375 , n54376 , n54377 , 
     n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n5063 , n5064 , n5065 , n5066 , 
     n5067 , n5068 , n5069 , n5070 , n5071 , n54393 , n5073 , n5074 , n54396 , n54397 , 
     n54398 , n54399 , n5079 , n5080 , n5081 , n54403 , n54404 , n54405 , n54406 , n5086 , 
     n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , 
     n54418 , n54419 , n54420 , n54421 , n5101 , n5102 , n5103 , n5104 , n54426 , n54427 , 
     n54428 , n54429 , n5109 , n5110 , n54432 , n5112 , n5113 , n5114 , n5115 , n54437 , 
     n54438 , n54439 , n5119 , n54441 , n54442 , n54443 , n5123 , n54445 , n54446 , n54447 , 
     n54448 , n54449 , n5129 , n5130 , n54452 , n54453 , n54454 , n5134 , n54456 , n54457 , 
     n54458 , n5138 , n54460 , n54461 , n54462 , n5142 , n54464 , n54465 , n54466 , n5146 , 
     n54468 , n54469 , n5149 , n54471 , n54472 , n5152 , n5153 , n5154 , n54476 , n54477 , 
     n54478 , n54479 , n54480 , n5160 , n54482 , n54483 , n5163 , n5164 , n5165 , n54487 , 
     n54488 , n54489 , n54490 , n54491 , n5171 , n54493 , n54494 , n5174 , n5175 , n5176 , 
     n54498 , n54499 , n5179 , n54501 , n54502 , n5182 , n54504 , n54505 , n54506 , n54507 , 
     n5187 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n5196 , 
     n54518 , n54519 , n54520 , n5200 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , 
     n54528 , n54529 , n5209 , n54531 , n54532 , n5212 , n54534 , n54535 , n5215 , n54537 , 
     n5217 , n54539 , n54540 , n5220 , n5221 , n54543 , n5223 , n5224 , n5225 , n5226 , 
     n54548 , n54549 , n54550 , n54551 , n5231 , n54553 , n54554 , n54555 , n5235 , n5236 , 
     n54558 , n54559 , n54560 , n54561 , n54562 , n5242 , n5243 , n54565 , n54566 , n54567 , 
     n54568 , n54569 , n54570 , n54571 , n5251 , n54573 , n54574 , n54575 , n54576 , n54577 , 
     n5257 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n5265 , n54587 , 
     n54588 , n5268 , n5269 , n5270 , n54592 , n54593 , n54594 , n54595 , n5275 , n54597 , 
     n54598 , n54599 , n54600 , n5280 , n5281 , n54603 , n54604 , n54605 , n54606 , n5286 , 
     n54608 , n54609 , n54610 , n54611 , n5291 , n5292 , n54614 , n54615 , n54616 , n5296 , 
     n54618 , n54619 , n5299 , n5300 , n5301 , n5302 , n54624 , n5304 , n5305 , n5306 , 
     n5307 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n5314 , n5315 , n54637 , 
     n54638 , n54639 , n5319 , n54641 , n54642 , n5322 , n5323 , n54645 , n54646 , n54647 , 
     n54648 , n5328 , n5329 , n5330 , n5331 , n54653 , n54654 , n54655 , n54656 , n54657 , 
     n54658 , n54659 , n54660 , n54661 , n5341 , n54663 , n54664 , n54665 , n54666 , n5346 , 
     n54668 , n54669 , n54670 , n5350 , n5351 , n54673 , n54674 , n54675 , n5355 , n54677 , 
     n54678 , n54679 , n5359 , n54681 , n54682 , n54683 , n54684 , n5364 , n54686 , n54687 , 
     n5367 , n54689 , n5369 , n54691 , n54692 , n5372 , n54694 , n54695 , n5375 , n54697 , 
     n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , 
     n54708 , n5388 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , 
     n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n5404 , n5405 , n54727 , 
     n54728 , n5408 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , 
     n54738 , n5418 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , 
     n54748 , n54749 , n5429 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , 
     n5437 , n54759 , n5439 , n54761 , n54762 , n5442 , n54764 , n54765 , n54766 , n54767 , 
     n5447 , n54769 , n54770 , n5450 , n54772 , n5452 , n54774 , n54775 , n54776 , n54777 , 
     n54778 , n5458 , n54780 , n54781 , n5461 , n54783 , n5463 , n54785 , n54786 , n54787 , 
     n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n5474 , n54796 , n54797 , 
     n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , 
     n54808 , n54809 , n54810 , n54811 , n54812 , n5492 , n5493 , n54815 , n5495 , n5496 , 
     n5497 , n5498 , n54820 , n54821 , n54822 , n5502 , n54824 , n54825 , n5505 , n54827 , 
     n54828 , n5508 , n54830 , n54831 , n54832 , n54833 , n5513 , n54835 , n54836 , n54837 , 
     n54838 , n54839 , n54840 , n54841 , n54842 , n5522 , n54844 , n5524 , n5525 , n54847 , 
     n5527 , n5528 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n5535 , n54857 , 
     n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n5545 , n5546 , 
     n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n5554 , n54876 , n54877 , 
     n5557 , n54879 , n54880 , n54881 , n54882 , n54883 , n5563 , n54885 , n5565 , n5566 , 
     n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n5574 , n54896 , n54897 , 
     n54898 , n54899 , n5579 , n54901 , n54902 , n5582 , n54904 , n5584 , n5585 , n54907 , 
     n54908 , n54909 , n5589 , n54911 , n54912 , n54913 , n54914 , n5594 , n54916 , n54917 , 
     n54918 , n54919 , n5599 , n54921 , n54922 , n5602 , n5603 , n54925 , n54926 , n54927 , 
     n5605 , n5606 , n54930 , n54931 , n54932 , n54933 , n54934 , n5612 , n54936 , n5614 , 
     n54938 , n54939 , n5617 , n54941 , n54942 , n54943 , n5621 , n54945 , n54946 , n54947 , 
     n54948 , n54949 , n54950 , n54951 , n54952 , n5630 , n5631 , n54955 , n54956 , n54957 , 
     n54958 , n5634 , n54960 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , 
     n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , 
     n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , 
     n5663 , n5664 , n5665 , n54991 , n54992 , n54993 , n54994 , n54995 , n5671 , n5672 , 
     n54998 , n5674 , n55000 , n55001 , n55002 , n55003 , n5679 , n55005 , n55006 , n55007 , 
     n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n5689 , n55015 , n55016 , n55017 , 
     n55018 , n55019 , n5695 , n5696 , n5697 , n55023 , n5699 , n55025 , n55026 , n5702 , 
     n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n5711 , n55037 , 
     n5713 , n55039 , n5715 , n55041 , n55042 , n55043 , n5719 , n55045 , n55046 , n5722 , 
     n55048 , n5724 , n55050 , n5726 , n5727 , n55053 , n5729 , n55055 , n5731 , n5732 , 
     n5733 , n5734 , n5735 , n55061 , n55062 , n5738 , n55064 , n55065 , n55066 , n55067 , 
     n5743 , n55069 , n55070 , n5746 , n55072 , n5748 , n55074 , n55075 , n5751 , n55077 , 
     n55078 , n55079 , n5755 , n55081 , n5757 , n55083 , n55084 , n55085 , n5761 , n55087 , 
     n55088 , n5764 , n55090 , n5766 , n5767 , n55093 , n5769 , n55095 , n55096 , n5772 , 
     n55098 , n55099 , n55100 , n5776 , n55102 , n55103 , n5779 , n55105 , n55106 , n55107 , 
     n5783 , n55109 , n5785 , n55111 , n55112 , n5788 , n55114 , n5790 , n55116 , n5792 , 
     n55118 , n5794 , n5795 , n5796 , n5797 , n55123 , n55124 , n55125 , n5801 , n55127 , 
     n55128 , n55129 , n5805 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , 
     n5813 , n55139 , n55140 , n5816 , n55142 , n55143 , n55144 , n5820 , n55146 , n5822 , 
     n55148 , n55149 , n5825 , n5826 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , 
     n55158 , n5834 , n5835 , n5836 , n5837 , n55163 , n5839 , n55165 , n5841 , n5842 , 
     n5843 , n55169 , n55170 , n5846 , n55172 , n5848 , n55174 , n55175 , n5851 , n55177 , 
     n5853 , n5854 , n5855 , n55181 , n5857 , n55183 , n5859 , n5860 , n55186 , n55187 , 
     n5863 , n5864 , n55190 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , 
     n55198 , n55199 , n5875 , n55201 , n55202 , n55203 , n5879 , n55205 , n55206 , n55207 , 
     n55208 , n5884 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , 
     n55218 , n5894 , n5895 , n55221 , n5897 , n5898 , n55224 , n5900 , n55226 , n5902 , 
     n55228 , n55229 , n55230 , n5906 , n55232 , n55233 , n55234 , n55235 , n5911 , n55237 , 
     n55238 , n55239 , n55240 , n55241 , n5917 , n5918 , n5919 , n55245 , n5921 , n5922 , 
     n55248 , n5924 , n55250 , n55251 , n5927 , n5928 , n55254 , n5930 , n5931 , n5932 , 
     n55258 , n5934 , n5935 , n5936 , n5937 , n5938 , n55264 , n5940 , n55266 , n55267 , 
     n5943 , n55269 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , 
     n5953 , n5954 , n5955 , n5956 , n5957 , n55283 , n55284 , n55285 , n55286 , n5962 , 
     n55288 , n55289 , n5965 , n55291 , n5967 , n5968 , n55294 , n55295 , n5971 , n5972 , 
     n55298 , n5974 , n55300 , n5976 , n55302 , n55303 , n5979 , n55305 , n5981 , n5982 , 
     n55308 , n5984 , n5985 , n5986 , n5987 , n55313 , n55314 , n5990 , n55316 , n55317 , 
     n5993 , n55319 , n55320 , n55321 , n55322 , n55323 , n5999 , n55325 , n55326 , n55327 , 
     n55328 , n55329 , n55330 , n55331 , n6007 , n55333 , n55334 , n6010 , n6011 , n55337 , 
     n55338 , n6014 , n55340 , n55341 , n6017 , n55343 , n55344 , n6020 , n55346 , n55347 , 
     n6023 , n55349 , n55350 , n6026 , n55352 , n55353 , n55354 , n55355 , n6031 , n6032 , 
     n55358 , n6034 , n55360 , n55361 , n55362 , n6038 , n6039 , n55365 , n6041 , n55367 , 
     n55368 , n6044 , n6045 , n6046 , n55372 , n55373 , n55374 , n6050 , n6051 , n55377 , 
     n6053 , n6054 , n55380 , n6056 , n55382 , n55383 , n6059 , n55385 , n55386 , n55387 , 
     n55388 , n55389 , n6065 , n55391 , n55392 , n55393 , n55394 , n55395 , n6071 , n55397 , 
     n6073 , n55399 , n55400 , n55401 , n6077 , n55403 , n55404 , n55405 , n6081 , n6082 , 
     n55408 , n55409 , n6085 , n55411 , n6087 , n55413 , n6089 , n55415 , n55416 , n6092 , 
     n55418 , n55419 , n6095 , n55421 , n6097 , n55423 , n55424 , n55425 , n55426 , n6102 , 
     n55428 , n55429 , n6105 , n6106 , n55432 , n6108 , n6109 , n55435 , n55436 , n55437 , 
     n55438 , n55439 , n6115 , n6116 , n55442 , n6118 , n55444 , n55445 , n6121 , n6122 , 
     n55448 , n6124 , n55450 , n6126 , n6127 , n55453 , n6129 , n55455 , n6131 , n6132 , 
     n55458 , n55459 , n6135 , n55461 , n55462 , n55463 , n6139 , n55465 , n6141 , n55467 , 
     n6143 , n55469 , n6145 , n55471 , n6147 , n55473 , n55474 , n6150 , n55476 , n55477 , 
     n6153 , n6154 , n55480 , n55481 , n6157 , n55483 , n55484 , n6160 , n55486 , n55487 , 
     n55488 , n6164 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , 
     n55498 , n6174 , n55500 , n6176 , n55502 , n55503 , n55504 , n6180 , n55506 , n6182 , 
     n6183 , n6184 , n6185 , n55511 , n55512 , n55513 , n55514 , n55515 , n6191 , n55517 , 
     n55518 , n6194 , n6195 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , 
     n55528 , n55529 , n55530 , n6206 , n6207 , n55533 , n55534 , n55535 , n55536 , n6212 , 
     n6213 , n55539 , n6215 , n55541 , n6217 , n6218 , n55544 , n6220 , n55546 , n55547 , 
     n6223 , n55549 , n55550 , n6226 , n6227 , n6228 , n6229 , n6230 , n55556 , n6232 , 
     n55558 , n55559 , n6235 , n55561 , n55562 , n6238 , n55564 , n6240 , n6241 , n6242 , 
     n6243 , n6244 , n55570 , n55571 , n6247 , n55573 , n55574 , n6250 , n55576 , n55577 , 
     n6253 , n55579 , n55580 , n55581 , n55582 , n6258 , n55584 , n55585 , n55586 , n6262 , 
     n6263 , n6264 , n6265 , n55591 , n55592 , n55593 , n55594 , n6270 , n55596 , n55597 , 
     n6273 , n55599 , n55600 , n6276 , n55602 , n55603 , n6279 , n55605 , n55606 , n6282 , 
     n55608 , n6284 , n55610 , n55611 , n55612 , n6288 , n55614 , n55615 , n6291 , n55617 , 
     n55618 , n55619 , n6295 , n55621 , n55622 , n6298 , n6299 , n55625 , n6301 , n6302 , 
     n55628 , n55629 , n55630 , n6306 , n55632 , n55633 , n55634 , n6310 , n6311 , n6312 , 
     n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n6319 , n6320 , n55646 , n6322 , 
     n55648 , n55649 , n55650 , n6326 , n6327 , n55653 , n6329 , n55655 , n6331 , n55657 , 
     n55658 , n55659 , n55660 , n55661 , n6337 , n55663 , n55664 , n55665 , n6341 , n55667 , 
     n55668 , n6344 , n6345 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n6352 , 
     n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , 
     n6363 , n55689 , n6365 , n55691 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , 
     n6373 , n55699 , n55700 , n6376 , n55702 , n6378 , n55704 , n6380 , n55706 , n55707 , 
     n55708 , n6384 , n55710 , n6386 , n55712 , n55713 , n6389 , n55715 , n6391 , n6392 , 
     n55718 , n6394 , n55720 , n6396 , n6397 , n6398 , n55724 , n55725 , n55726 , n6402 , 
     n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n6409 , n55735 , n55736 , n6412 , 
     n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , 
     n6423 , n6424 , n55750 , n6426 , n55752 , n55753 , n6429 , n6430 , n55756 , n6432 , 
     n55758 , n6434 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n6442 , 
     n6443 , n55769 , n6445 , n55771 , n55772 , n6448 , n55774 , n6450 , n55776 , n55777 , 
     n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n6459 , n6460 , n55786 , n55787 , 
     n6463 , n55789 , n55790 , n6466 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , 
     n55798 , n55799 , n6475 , n6476 , n6477 , n55803 , n6479 , n55805 , n55806 , n55807 , 
     n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n6491 , n6492 , 
     n6493 , n6494 , n55820 , n6496 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , 
     n6503 , n55829 , n55830 , n55831 , n55832 , n55833 , n6509 , n55835 , n55836 , n55837 , 
     n6513 , n6514 , n55840 , n55841 , n6517 , n6518 , n55844 , n55845 , n55846 , n55847 , 
     n55848 , n6524 , n6525 , n6526 , n55852 , n6528 , n55854 , n6530 , n55856 , n6532 , 
     n55858 , n6534 , n55860 , n6536 , n55862 , n55863 , n55864 , n6540 , n55866 , n6542 , 
     n6543 , n55869 , n6545 , n55871 , n6547 , n55873 , n55874 , n55875 , n6551 , n55877 , 
     n6553 , n6554 , n6555 , n6556 , n6557 , n55883 , n6559 , n55885 , n6561 , n55887 , 
     n55888 , n55889 , n55890 , n6566 , n6567 , n55893 , n55894 , n55895 , n6571 , n55897 , 
     n6573 , n55899 , n6575 , n6576 , n55902 , n55903 , n55904 , n6580 , n55906 , n55907 , 
     n6583 , n55909 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n55917 , 
     n55918 , n55919 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n55927 , 
     n55928 , n6603 , n55930 , n55931 , n55932 , n55933 , n55934 , n6609 , n6610 , n6611 , 
     n6612 , n6613 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , 
     n55948 , n55949 , n6616 , n55951 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , 
     n6624 , n6625 , n6626 , n6627 , n55962 , n6629 , n55964 , n55965 , n55966 , n55967 , 
     n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n6640 , n55975 , n55976 , n6643 , 
     n55978 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n55985 , n55986 , n55987 , 
     n55988 , n55989 , n55990 , n55991 , n55992 , n6659 , n55994 , n55995 , n55996 , n55997 , 
     n55998 , n6665 , n56000 , n6667 , n56002 , n6669 , n56004 , n56005 , n56006 , n6673 , 
     n56008 , n6675 , n56010 , n56011 , n56012 , n56013 , n6680 , n56015 , n6682 , n56017 , 
     n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , 
     n6694 , n6695 , n56030 , n56031 , n6698 , n56033 , n6700 , n56035 , n56036 , n56037 , 
     n56038 , n56039 , n6706 , n6707 , n56042 , n56043 , n56044 , n6711 , n56046 , n56047 , 
     n56048 , n56049 , n56050 , n56051 , n6718 , n56053 , n56054 , n6721 , n56056 , n6723 , 
     n6724 , n56059 , n6726 , n56061 , n56062 , n56063 , n56064 , n6731 , n56066 , n56067 , 
     n6734 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n6741 , n6742 , n56077 , 
     n6744 , n56079 , n56080 , n6747 , n56082 , n56083 , n56084 , n56085 , n6752 , n56087 , 
     n56088 , n56089 , n6756 , n56091 , n6758 , n56093 , n56094 , n6761 , n56096 , n56097 , 
     n56098 , n56099 , n6766 , n56101 , n56102 , n6769 , n56104 , n56105 , n6772 , n56107 , 
     n56108 , n6775 , n6776 , n56111 , n56112 , n6779 , n56114 , n56115 , n56116 , n56117 , 
     n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n6792 , n56127 , 
     n56128 , n6795 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n6803 , 
     n56138 , n56139 , n6806 , n56141 , n56142 , n6809 , n56144 , n6811 , n56146 , n56147 , 
     n56148 , n56149 , n56150 , n6817 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , 
     n6824 , n56159 , n56160 , n6827 , n56162 , n56163 , n6830 , n56165 , n56166 , n6833 , 
     n6834 , n6835 , n56170 , n6837 , n56172 , n56173 , n56174 , n6841 , n56176 , n56177 , 
     n6844 , n56179 , n6846 , n56181 , n6848 , n56183 , n6850 , n56185 , n6852 , n56187 , 
     n6854 , n56189 , n6856 , n56191 , n56192 , n56193 , n6860 , n56195 , n6862 , n56197 , 
     n56198 , n6865 , n56200 , n56201 , n6868 , n56203 , n56204 , n56205 , n56206 , n6873 , 
     n56208 , n56209 , n56210 , n56211 , n6878 , n6879 , n56214 , n6881 , n6882 , n6883 , 
     n6884 , n6885 , n56220 , n56221 , n6888 , n56223 , n56224 , n56225 , n56226 , n6893 , 
     n56228 , n56229 , n56230 , n56231 , n6898 , n56233 , n56234 , n6901 , n56236 , n6903 , 
     n56238 , n6905 , n56240 , n56241 , n6908 , n56243 , n6910 , n6911 , n56246 , n56247 , 
     n6914 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n6922 , n56257 , 
     n56258 , n6925 , n56260 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n56267 , 
     n56268 , n6935 , n56270 , n6937 , n6938 , n56273 , n6940 , n56275 , n56276 , n6943 , 
     n56278 , n56279 , n56280 , n56281 , n6948 , n56283 , n6950 , n6951 , n56286 , n56287 , 
     n6954 , n56289 , n56290 , n56291 , n6958 , n6959 , n56294 , n6961 , n56296 , n6963 , 
     n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n56305 , n6972 , n56307 , 
     n56308 , n56309 , n56310 , n56311 , n6978 , n6979 , n6980 , n56315 , n6982 , n6983 , 
     n56318 , n6985 , n56320 , n56321 , n6988 , n56323 , n6990 , n6991 , n6992 , n6993 , 
     n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n7001 , n7002 , n56337 , 
     n7004 , n56339 , n7006 , n56341 , n56342 , n7009 , n56344 , n56345 , n7012 , n7013 , 
     n56348 , n7015 , n7016 , n7017 , n7018 , n56353 , n7020 , n7021 , n56356 , n56357 , 
     n7024 , n56359 , n7026 , n7027 , n7028 , n7029 , n56364 , n7031 , n56366 , n7033 , 
     n56368 , n7035 , n7036 , n7037 , n7038 , n56373 , n7040 , n7041 , n56376 , n7043 , 
     n7044 , n56379 , n7046 , n7047 , n56382 , n7049 , n56384 , n56385 , n56386 , n7053 , 
     n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n7060 , n56395 , n56396 , n7063 , 
     n56398 , n56399 , n7066 , n7067 , n7068 , n7069 , n7070 , n56405 , n56406 , n7073 , 
     n7074 , n7075 , n7076 , n56411 , n56412 , n56413 , n7080 , n56415 , n7082 , n7083 , 
     n56418 , n56419 , n7086 , n56421 , n56422 , n7089 , n56424 , n56425 , n7092 , n7093 , 
     n56428 , n7095 , n7096 , n56431 , n56432 , n7099 , n7100 , n7101 , n56436 , n7103 , 
     n56438 , n56439 , n56440 , n7107 , n56442 , n7109 , n7110 , n7111 , n7112 , n56447 , 
     n7114 , n56449 , n7116 , n56451 , n56452 , n56453 , n7120 , n56455 , n56456 , n56457 , 
     n56458 , n56459 , n56460 , n7127 , n56462 , n7129 , n7130 , n56465 , n56466 , n56467 , 
     n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n7141 , n56476 , n7143 , 
     n56478 , n56479 , n7146 , n56481 , n56482 , n7149 , n56484 , n56485 , n56486 , n7153 , 
     n56488 , n7155 , n56490 , n56491 , n7158 , n56493 , n56494 , n7161 , n56496 , n7163 , 
     n7164 , n56499 , n7166 , n56501 , n7168 , n56503 , n7170 , n56505 , n56506 , n7173 , 
     n56508 , n56509 , n7176 , n7177 , n56512 , n7179 , n56514 , n7181 , n56516 , n7183 , 
     n56518 , n56519 , n7186 , n56521 , n7188 , n7189 , n56524 , n56525 , n7192 , n56527 , 
     n7194 , n56529 , n56530 , n56531 , n56532 , n56533 , n7200 , n56535 , n56536 , n7203 , 
     n7204 , n7205 , n7206 , n56541 , n56542 , n7209 , n56544 , n56545 , n56546 , n56547 , 
     n7214 , n7215 , n56550 , n7217 , n7218 , n56553 , n7220 , n56555 , n56556 , n7223 , 
     n56558 , n7225 , n56560 , n56561 , n7228 , n7229 , n7230 , n56565 , n56566 , n56567 , 
     n7234 , n7235 , n56570 , n7237 , n7238 , n56573 , n7240 , n7241 , n7242 , n7243 , 
     n7244 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , 
     n56588 , n56589 , n7256 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , 
     n56598 , n56599 , n56600 , n56601 , n7268 , n56603 , n7270 , n7271 , n7272 , n56607 , 
     n56608 , n7275 , n56610 , n7277 , n7278 , n7279 , n7280 , n7281 , n56616 , n56617 , 
     n7284 , n56619 , n56620 , n7287 , n56622 , n7289 , n56624 , n56625 , n56626 , n56627 , 
     n56628 , n7295 , n56630 , n56631 , n56632 , n56633 , n7300 , n56635 , n56636 , n7303 , 
     n56638 , n56639 , n7306 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , 
     n56648 , n56649 , n56650 , n7317 , n56652 , n56653 , n7320 , n56655 , n56656 , n7323 , 
     n56658 , n56659 , n56660 , n56661 , n7328 , n56663 , n56664 , n7331 , n7332 , n56667 , 
     n56668 , n56669 , n56670 , n7337 , n7338 , n56673 , n7340 , n56675 , n56676 , n7343 , 
     n56678 , n7345 , n56680 , n7347 , n7348 , n56683 , n56684 , n56685 , n7352 , n56687 , 
     n56688 , n56689 , n56690 , n7357 , n7358 , n7359 , n56694 , n56695 , n56696 , n56697 , 
     n56698 , n56699 , n7366 , n56701 , n56702 , n7369 , n56704 , n56705 , n7372 , n56707 , 
     n56708 , n7375 , n56710 , n7377 , n56712 , n56713 , n7380 , n56715 , n7382 , n56717 , 
     n7384 , n7385 , n56720 , n7387 , n56722 , n56723 , n56724 , n56725 , n56726 , n7393 , 
     n56728 , n56729 , n7396 , n56731 , n7398 , n7399 , n56734 , n7401 , n56736 , n56737 , 
     n56738 , n56739 , n56740 , n56741 , n7408 , n56743 , n7410 , n7411 , n56746 , n7413 , 
     n56748 , n7415 , n7416 , n7417 , n7418 , n56753 , n7420 , n56755 , n7422 , n7423 , 
     n56758 , n7425 , n56760 , n56761 , n7428 , n56763 , n56764 , n56765 , n56766 , n56767 , 
     n56768 , n56769 , n56770 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , 
     n7444 , n56779 , n7446 , n56781 , n7448 , n56783 , n56784 , n56785 , n56786 , n56787 , 
     n56788 , n7455 , n7456 , n56791 , n7458 , n56793 , n56794 , n7461 , n7462 , n56797 , 
     n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n7471 , n56806 , n56807 , 
     n56808 , n7475 , n7476 , n56811 , n7478 , n56813 , n56814 , n56815 , n56816 , n56817 , 
     n56818 , n7485 , n56820 , n56821 , n7488 , n56823 , n56824 , n56825 , n56826 , n7493 , 
     n7494 , n56829 , n7496 , n7497 , n7498 , n56833 , n7500 , n56835 , n56836 , n56837 , 
     n7504 , n56839 , n56840 , n56841 , n56842 , n56843 , n7510 , n56845 , n56846 , n56847 , 
     n56848 , n56849 , n7516 , n56851 , n56852 , n7519 , n56854 , n7521 , n56856 , n56857 , 
     n56858 , n56859 , n56860 , n7527 , n56862 , n56863 , n7530 , n7531 , n7532 , n56867 , 
     n56868 , n56869 , n56870 , n7537 , n56872 , n56873 , n7540 , n7541 , n7542 , n56877 , 
     n56878 , n7545 , n56880 , n7547 , n56882 , n56883 , n7550 , n56885 , n56886 , n7553 , 
     n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n7563 , 
     n56898 , n7565 , n56900 , n56901 , n7568 , n56903 , n7570 , n7571 , n56906 , n56907 , 
     n7574 , n56909 , n56910 , n7577 , n56912 , n56913 , n56914 , n56915 , n7582 , n56917 , 
     n7584 , n56919 , n7586 , n56921 , n7588 , n56923 , n56924 , n56925 , n56926 , n56927 , 
     n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n7601 , n7602 , n56937 , 
     n56938 , n56939 , n56940 , n56941 , n56942 , n7609 , n56944 , n56945 , n56946 , n56947 , 
     n56948 , n56949 , n7616 , n56951 , n56952 , n7619 , n56954 , n56955 , n56956 , n56957 , 
     n56958 , n56959 , n56960 , n7627 , n7628 , n56963 , n7630 , n56965 , n56966 , n56967 , 
     n56968 , n56969 , n56970 , n7637 , n56972 , n56973 , n56974 , n56975 , n7642 , n56977 , 
     n7644 , n56979 , n56980 , n56981 , n56982 , n7649 , n56984 , n7651 , n7652 , n56987 , 
     n56988 , n56989 , n56990 , n7657 , n7658 , n7659 , n7660 , n56995 , n56996 , n56997 , 
     n7664 , n56999 , n7666 , n57001 , n7668 , n57003 , n57004 , n57005 , n57006 , n57007 , 
     n57008 , n7675 , n57010 , n57011 , n7678 , n7679 , n57014 , n57015 , n57016 , n7683 , 
     n57018 , n57019 , n7686 , n57021 , n57022 , n57023 , n7690 , n57025 , n57026 , n7693 , 
     n7694 , n57029 , n7696 , n57031 , n57032 , n7699 , n7700 , n57035 , n57036 , n57037 , 
     n57038 , n57039 , n7706 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n7713 , 
     n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n7721 , n7722 , n57057 , 
     n7724 , n57059 , n57060 , n57061 , n57062 , n57063 , n7730 , n7731 , n57066 , n57067 , 
     n57068 , n57069 , n57070 , n7737 , n57072 , n57073 , n7740 , n57075 , n57076 , n57077 , 
     n57078 , n7745 , n57080 , n57081 , n7748 , n57083 , n57084 , n7751 , n7752 , n57087 , 
     n57088 , n7755 , n57090 , n7757 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , 
     n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , 
     n57108 , n57109 , n7776 , n57111 , n57112 , n7779 , n57114 , n57115 , n7782 , n57117 , 
     n57118 , n7785 , n57120 , n7787 , n57122 , n57123 , n7790 , n7791 , n57126 , n7793 , 
     n57128 , n57129 , n7796 , n57131 , n57132 , n7799 , n57134 , n7801 , n57136 , n7803 , 
     n57138 , n57139 , n7806 , n57141 , n57142 , n57143 , n57144 , n7811 , n57146 , n7813 , 
     n57148 , n7815 , n57150 , n57151 , n7818 , n57153 , n7820 , n7821 , n57156 , n57157 , 
     n57158 , n57159 , n57160 , n57161 , n7828 , n7829 , n57164 , n57165 , n7832 , n57167 , 
     n7834 , n7835 , n7836 , n57171 , n57172 , n57173 , n57174 , n7841 , n57176 , n57177 , 
     n7844 , n7845 , n7846 , n57181 , n57182 , n7849 , n57184 , n57185 , n7852 , n57187 , 
     n7854 , n57189 , n7856 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , 
     n57198 , n57199 , n57200 , n7867 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , 
     n57208 , n57209 , n7876 , n57211 , n57212 , n7879 , n57214 , n57215 , n57216 , n57217 , 
     n57218 , n7885 , n57220 , n57221 , n57222 , n57223 , n7890 , n57225 , n57226 , n7893 , 
     n57228 , n57229 , n7896 , n57231 , n57232 , n57233 , n57234 , n7901 , n57236 , n57237 , 
     n57238 , n57239 , n7906 , n57241 , n57242 , n7909 , n57244 , n7911 , n57246 , n57247 , 
     n57248 , n57249 , n57250 , n7917 , n57252 , n7919 , n57254 , n57255 , n57256 , n57257 , 
     n57258 , n7925 , n57260 , n7927 , n7928 , n57263 , n7930 , n7931 , n7932 , n57267 , 
     n7934 , n57269 , n57270 , n57271 , n57272 , n7939 , n57274 , n57275 , n57276 , n57277 , 
     n57278 , n7945 , n57280 , n7947 , n57282 , n57283 , n7950 , n57285 , n57286 , n57287 , 
     n57288 , n57289 , n57290 , n57291 , n7958 , n57293 , n7960 , n57295 , n57296 , n57297 , 
     n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , 
     n57308 , n7975 , n57310 , n57311 , n7978 , n7979 , n7980 , n57315 , n57316 , n7983 , 
     n57318 , n7985 , n57320 , n7987 , n57322 , n7989 , n7990 , n57325 , n57326 , n57327 , 
     n7994 , n57329 , n7996 , n7997 , n57332 , n57333 , n8000 , n57335 , n8002 , n57337 , 
     n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n8013 , 
     n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n8021 , n57356 , n57357 , 
     n8024 , n8025 , n8026 , n8027 , n8028 , n57363 , n8030 , n57365 , n57366 , n57367 , 
     n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n8043 , 
     n57378 , n8045 , n57380 , n8047 , n57382 , n8049 , n8050 , n57385 , n57386 , n8053 , 
     n57388 , n57389 , n8056 , n57391 , n57392 , n57393 , n8060 , n57395 , n8062 , n57397 , 
     n57398 , n57399 , n8066 , n8067 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , 
     n57408 , n57409 , n8076 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , 
     n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , 
     n57428 , n57429 , n57430 , n57431 , n8098 , n57433 , n57434 , n8101 , n57436 , n8103 , 
     n8104 , n57439 , n57440 , n57441 , n57442 , n8109 , n8110 , n57445 , n57446 , n57447 , 
     n57448 , n57449 , n8116 , n57451 , n57452 , n57453 , n57454 , n57455 , n8122 , n57457 , 
     n8124 , n8125 , n57460 , n57461 , n57462 , n8129 , n57464 , n57465 , n57466 , n57467 , 
     n8134 , n57469 , n57470 , n57471 , n8138 , n8139 , n57474 , n8141 , n57476 , n8143 , 
     n57478 , n8145 , n8146 , n57481 , n8148 , n57483 , n8150 , n8151 , n8152 , n8153 , 
     n8154 , n8155 , n8156 , n8157 , n57492 , n8159 , n8160 , n8161 , n8162 , n8163 , 
     n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n57504 , n8171 , n57506 , n57507 , 
     n8174 , n57509 , n57510 , n57511 , n8178 , n57513 , n57514 , n57515 , n57516 , n57517 , 
     n57518 , n57519 , n8186 , n8187 , n8188 , n57523 , n57524 , n8191 , n8192 , n8193 , 
     n8194 , n8195 , n57530 , n8197 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , 
     n8204 , n57539 , n8206 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n8213 , 
     n57548 , n8215 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n8222 , n8223 , 
     n8224 , n8225 , n8226 , n8227 , n8228 , n57563 , n8230 , n57565 , n8232 , n57567 , 
     n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n57574 , n57575 , n8242 , n57577 , 
     n8244 , n57579 , n57580 , n8247 , n8248 , n57583 , n8250 , n57585 , n57586 , n57587 , 
     n8254 , n57589 , n8256 , n57591 , n57592 , n8259 , n57594 , n57595 , n8262 , n8263 , 
     n8264 , n57599 , n57600 , n8267 , n57602 , n8269 , n8270 , n8271 , n8272 , n8273 , 
     n8274 , n8275 , n8276 , n8277 , n8278 , n57613 , n57614 , n57615 , n57616 , n57617 , 
     n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n8290 , n57625 , n57626 , n57627 , 
     n57628 , n57629 , n57630 , n57631 , n8298 , n57633 , n57634 , n57635 , n57636 , n57637 , 
     n57638 , n8305 , n57640 , n8307 , n57642 , n57643 , n8310 , n8311 , n57646 , n8313 , 
     n57648 , n8315 , n8316 , n57651 , n57652 , n8319 , n57654 , n8321 , n8322 , n57657 , 
     n8324 , n57659 , n57660 , n8327 , n57662 , n8329 , n8330 , n57665 , n57666 , n8333 , 
     n8334 , n57669 , n8336 , n8337 , n57672 , n57673 , n8340 , n8341 , n57676 , n8343 , 
     n57678 , n57679 , n57680 , n8347 , n8348 , n8349 , n57684 , n8351 , n57686 , n57687 , 
     n8354 , n57689 , n8356 , n8357 , n8358 , n8359 , n57694 , n57695 , n8362 , n57697 , 
     n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n57705 , n57706 , n8373 , 
     n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , 
     n8384 , n57719 , n57720 , n57721 , n57722 , n8389 , n57724 , n57725 , n8392 , n8393 , 
     n8394 , n8395 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n8402 , n57737 , 
     n57738 , n8405 , n57740 , n57741 , n8408 , n57743 , n8410 , n57745 , n8412 , n57747 , 
     n57748 , n57749 , n8416 , n57751 , n8418 , n57753 , n57754 , n8421 , n57756 , n57757 , 
     n57758 , n8425 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n8432 , n57767 , 
     n57768 , n8435 , n57770 , n57771 , n8438 , n8439 , n57774 , n57775 , n8442 , n57777 , 
     n57778 , n8445 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n8452 , n57787 , 
     n57788 , n8455 , n57790 , n8457 , n8458 , n57793 , n8460 , n57795 , n8462 , n57797 , 
     n57798 , n8465 , n57800 , n57801 , n8468 , n57803 , n8470 , n57805 , n57806 , n8473 , 
     n57808 , n57809 , n57810 , n8477 , n57812 , n57813 , n57814 , n57815 , n57816 , n8483 , 
     n57818 , n57819 , n8486 , n57821 , n57822 , n8489 , n57824 , n57825 , n8492 , n57827 , 
     n57828 , n8495 , n57830 , n57831 , n8498 , n57833 , n57834 , n57835 , n57836 , n8503 , 
     n8504 , n57839 , n57840 , n8507 , n57842 , n57843 , n57844 , n8511 , n57846 , n8513 , 
     n8514 , n8515 , n8516 , n8517 , n8518 , n57853 , n8520 , n57855 , n8522 , n8523 , 
     n57858 , n8525 , n57860 , n57861 , n8528 , n57863 , n57864 , n8531 , n57866 , n57867 , 
     n8534 , n57869 , n57870 , n8537 , n57872 , n57873 , n8540 , n57875 , n57876 , n57877 , 
     n57878 , n57879 , n57880 , n57881 , n8548 , n57883 , n57884 , n8551 , n57886 , n57887 , 
     n8554 , n57889 , n57890 , n8557 , n57892 , n8559 , n8560 , n57895 , n8562 , n57897 , 
     n8564 , n57899 , n8566 , n8567 , n57902 , n57903 , n8570 , n57905 , n57906 , n8573 , 
     n57908 , n8575 , n8576 , n57911 , n8578 , n8579 , n57914 , n8581 , n8582 , n8583 , 
     n8584 , n8585 , n8586 , n57921 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , 
     n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n57934 , n8601 , n57936 , n57937 , 
     n57938 , n8605 , n57940 , n57941 , n8608 , n57943 , n57944 , n8611 , n8612 , n57947 , 
     n8614 , n57949 , n57950 , n8617 , n57952 , n8619 , n8620 , n57955 , n8622 , n8623 , 
     n8624 , n8625 , n57960 , n8627 , n57962 , n8629 , n57964 , n57965 , n57966 , n57967 , 
     n57968 , n57969 , n57970 , n8637 , n8638 , n8639 , n8640 , n8641 , n57976 , n57977 , 
     n8644 , n57979 , n57980 , n8647 , n8648 , n8649 , n8650 , n57985 , n8652 , n57987 , 
     n57988 , n57989 , n8656 , n57991 , n8658 , n8659 , n57994 , n57995 , n57996 , n57997 , 
     n57998 , n57999 , n58000 , n58001 , n58002 , n8669 , n58004 , n58005 , n58006 , n8673 , 
     n58008 , n58009 , n8676 , n58011 , n58012 , n8679 , n58014 , n8681 , n8682 , n8683 , 
     n8684 , n58019 , n8686 , n8687 , n8688 , n58023 , n8690 , n58025 , n58026 , n58027 , 
     n58028 , n58029 , n8696 , n58031 , n58032 , n8699 , n8700 , n8701 , n8702 , n58037 , 
     n8704 , n58039 , n8706 , n58041 , n8708 , n8709 , n58044 , n8711 , n58046 , n58047 , 
     n58048 , n8715 , n58050 , n58051 , n8718 , n58053 , n58054 , n8721 , n58056 , n58057 , 
     n8724 , n58059 , n8726 , n58061 , n58062 , n8729 , n58064 , n8731 , n58066 , n58067 , 
     n8734 , n58069 , n8736 , n58071 , n8738 , n58073 , n8740 , n58075 , n8742 , n8743 , 
     n8744 , n8745 , n58080 , n58081 , n58082 , n8749 , n58084 , n58085 , n58086 , n8753 , 
     n58088 , n8755 , n58090 , n58091 , n8758 , n8759 , n8760 , n8761 , n58096 , n8763 , 
     n8764 , n8765 , n8766 , n8767 , n8768 , n58103 , n8770 , n58105 , n58106 , n58107 , 
     n8774 , n58109 , n8776 , n58111 , n58112 , n8779 , n58114 , n58115 , n8782 , n58117 , 
     n58118 , n8785 , n8786 , n8787 , n58122 , n8789 , n58124 , n8791 , n58126 , n8793 , 
     n58128 , n58129 , n58130 , n58131 , n58132 , n8799 , n58134 , n8801 , n8802 , n8803 , 
     n58138 , n8805 , n58140 , n58141 , n58142 , n8809 , n58144 , n58145 , n8812 , n58147 , 
     n8814 , n58149 , n58150 , n8817 , n8818 , n58153 , n8820 , n58155 , n58156 , n8823 , 
     n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n8832 , n58167 , 
     n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n8840 , n8841 , n58176 , n8843 , 
     n8844 , n8845 , n8846 , n8847 , n58182 , n8849 , n58184 , n58185 , n58186 , n58187 , 
     n58188 , n8855 , n8856 , n58191 , n8858 , n58193 , n8860 , n8861 , n58196 , n58197 , 
     n8864 , n58199 , n58200 , n8867 , n58202 , n58203 , n58204 , n8871 , n58206 , n58207 , 
     n8874 , n58209 , n58210 , n8877 , n58212 , n8879 , n58214 , n58215 , n58216 , n8883 , 
     n58218 , n58219 , n58220 , n58221 , n8888 , n8889 , n58224 , n58225 , n8892 , n58227 , 
     n58228 , n8895 , n8896 , n58231 , n58232 , n58233 , n8900 , n58235 , n58236 , n58237 , 
     n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n8910 , n58245 , n58246 , n58247 , 
     n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n8923 , 
     n58258 , n58259 , n8926 , n58261 , n58262 , n8929 , n58264 , n58265 , n8932 , n58267 , 
     n58268 , n58269 , n58270 , n58271 , n8938 , n58273 , n58274 , n58275 , n58276 , n58277 , 
     n8944 , n58279 , n58280 , n58281 , n58282 , n58283 , n8950 , n8951 , n8952 , n8953 , 
     n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n58294 , n58295 , n8962 , n58297 , 
     n58298 , n58299 , n58300 , n8967 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , 
     n58308 , n58309 , n8976 , n58311 , n58312 , n8979 , n58314 , n58315 , n8982 , n58317 , 
     n58318 , n8985 , n8986 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n8993 , 
     n58328 , n58329 , n8996 , n58331 , n8998 , n58333 , n9000 , n58335 , n58336 , n58337 , 
     n9004 , n9005 , n58340 , n9007 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , 
     n9014 , n58349 , n58350 , n58351 , n58352 , n9019 , n58354 , n58355 , n9022 , n9023 , 
     n58358 , n9025 , n58360 , n9027 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , 
     n9034 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n9042 , n58377 , 
     n58378 , n9045 , n9046 , n9047 , n58382 , n58383 , n9050 , n58385 , n58386 , n58387 , 
     n9054 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n9062 , n58397 , 
     n9064 , n9065 , n58400 , n58401 , n9068 , n58403 , n9070 , n58405 , n9072 , n58407 , 
     n58408 , n9075 , n58410 , n9077 , n58412 , n9079 , n9080 , n9081 , n58416 , n58417 , 
     n9084 , n58419 , n9086 , n58421 , n9088 , n58423 , n58424 , n9091 , n58426 , n58427 , 
     n58428 , n58429 , n58430 , n58431 , n9098 , n58433 , n9100 , n58435 , n58436 , n9103 , 
     n58438 , n9105 , n9106 , n58441 , n58442 , n58443 , n9110 , n58445 , n9112 , n58447 , 
     n9114 , n9115 , n58450 , n9117 , n58452 , n9119 , n58454 , n58455 , n9122 , n58457 , 
     n58458 , n9125 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , 
     n58468 , n58469 , n9136 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , 
     n9144 , n9145 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , 
     n58488 , n58489 , n58490 , n9157 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , 
     n58498 , n58499 , n58500 , n9167 , n58502 , n9169 , n9170 , n9171 , n9172 , n9173 , 
     n58508 , n9175 , n58510 , n9177 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , 
     n58518 , n9185 , n9186 , n58521 , n58522 , n9189 , n58524 , n9191 , n58526 , n58527 , 
     n58528 , n58529 , n58530 , n9197 , n58532 , n58533 , n58534 , n9201 , n58536 , n58537 , 
     n9204 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n9212 , n9213 , 
     n9214 , n58549 , n58550 , n58551 , n9218 , n58553 , n58554 , n9221 , n58556 , n58557 , 
     n58558 , n9225 , n58560 , n58561 , n9228 , n58563 , n9230 , n58565 , n58566 , n58567 , 
     n58568 , n9235 , n58570 , n58571 , n9238 , n9239 , n58574 , n9241 , n9242 , n9243 , 
     n58578 , n9245 , n58580 , n58581 , n9248 , n58583 , n9250 , n9251 , n58586 , n9253 , 
     n58588 , n58589 , n9256 , n9257 , n58592 , n58593 , n58594 , n58595 , n9262 , n58597 , 
     n58598 , n9265 , n58600 , n58601 , n9268 , n58603 , n58604 , n9271 , n58606 , n9273 , 
     n9274 , n58609 , n9276 , n58611 , n58612 , n58613 , n58614 , n58615 , n9282 , n58617 , 
     n58618 , n9285 , n58620 , n9287 , n9288 , n58623 , n9290 , n58625 , n9292 , n58627 , 
     n9294 , n9295 , n9296 , n9297 , n58632 , n58633 , n9300 , n58635 , n58636 , n9303 , 
     n9304 , n9305 , n58640 , n9307 , n58642 , n9309 , n9310 , n9311 , n58646 , n9313 , 
     n58648 , n58649 , n58650 , n58651 , n9318 , n58653 , n58654 , n9321 , n58656 , n58657 , 
     n9324 , n58659 , n58660 , n58661 , n58662 , n58663 , n9330 , n58665 , n58666 , n9333 , 
     n9334 , n58669 , n58670 , n58671 , n9338 , n58673 , n58674 , n9341 , n58676 , n9343 , 
     n9344 , n58679 , n58680 , n58681 , n58682 , n9349 , n58684 , n58685 , n58686 , n58687 , 
     n58688 , n9355 , n58690 , n58691 , n9358 , n58693 , n58694 , n58695 , n58696 , n58697 , 
     n9364 , n58699 , n58700 , n9367 , n58702 , n58703 , n9370 , n9371 , n9372 , n9373 , 
     n9374 , n58709 , n58710 , n9377 , n58712 , n9379 , n58714 , n9381 , n9382 , n58717 , 
     n9384 , n9385 , n58720 , n58721 , n9388 , n58723 , n58724 , n58725 , n58726 , n58727 , 
     n58728 , n58729 , n58730 , n9397 , n58732 , n58733 , n58734 , n58735 , n9402 , n58737 , 
     n9404 , n58739 , n9406 , n9407 , n58742 , n9409 , n58744 , n9411 , n9412 , n9413 , 
     n9414 , n9415 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n9422 , n58757 , 
     n9424 , n58759 , n58760 , n9427 , n58762 , n9429 , n9430 , n58765 , n9432 , n58767 , 
     n58768 , n9435 , n58770 , n9437 , n58772 , n58773 , n58774 , n58775 , n58776 , n9443 , 
     n58778 , n9445 , n58780 , n9447 , n58782 , n58783 , n9450 , n58785 , n9452 , n58787 , 
     n9454 , n58789 , n9456 , n9457 , n58792 , n58793 , n9460 , n9461 , n58796 , n58797 , 
     n9464 , n58799 , n9466 , n9467 , n58802 , n58803 , n58804 , n9471 , n9472 , n58807 , 
     n9474 , n58809 , n9476 , n58811 , n9478 , n58813 , n9480 , n58815 , n58816 , n58817 , 
     n58818 , n9485 , n58820 , n58821 , n58822 , n58823 , n9490 , n58825 , n58826 , n58827 , 
     n9494 , n9495 , n58830 , n58831 , n58832 , n58833 , n9500 , n58835 , n58836 , n58837 , 
     n58838 , n58839 , n58840 , n58841 , n58842 , n9509 , n58844 , n58845 , n58846 , n58847 , 
     n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , 
     n58858 , n58859 , n58860 , n9527 , n9528 , n58863 , n58864 , n9531 , n58866 , n58867 , 
     n58868 , n58869 , n9536 , n58871 , n9538 , n58873 , n9540 , n9541 , n9542 , n9543 , 
     n9544 , n58879 , n9546 , n9547 , n58882 , n58883 , n58884 , n9550 , n58886 , n58887 , 
     n9553 , n58889 , n58890 , n58891 , n58892 , n58893 , n9559 , n58895 , n9561 , n58897 , 
     n9563 , n9564 , n9565 , n58901 , n58902 , n9566 , n58904 , n58905 , n9569 , n58907 , 
     n9571 , n9572 , n58910 , n58911 , n9575 , n9576 , n9577 , n9578 , n9579 , n58917 , 
     n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , 
     n9587 , n58929 , n58930 , n9590 , n58932 , n9592 , n58934 , n58935 , n58936 , n9596 , 
     n58938 , n9598 , n58940 , n58941 , n9601 , n58943 , n58944 , n58945 , n58946 , n9605 , 
     n58948 , n9607 , n9608 , n9609 , n58952 , n9611 , n9612 , n58955 , n58956 , n58957 , 
     n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n9619 , n58967 , 
     n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , 
     n9624 , n58979 , n9626 , n58981 , n58982 , n58983 , n58984 , n9631 , n58986 , n58987 , 
     n58988 , n58989 , n9634 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , 
     n58998 , n58999 , n59000 , n9637 , n59002 , n59003 , n59004 , n9641 , n59006 , n59007 , 
     n59008 , n59009 , n9646 , n59011 , n9648 , n59013 , n59014 , n59015 , n59016 , n9653 , 
     n59018 , n9655 , n59020 , n59021 , n9658 , n59023 , n59024 , n59025 , n9661 , n59027 , 
     n59028 , n9664 , n59030 , n59031 , n59032 , n9668 , n9669 , n59035 , n59036 , n59037 , 
     n59038 , n59039 , n9675 , n59041 , n9677 , n59043 , n59044 , n59045 , n9681 , n9682 , 
     n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n9690 , n9691 , n9692 , 
     n59058 , n9694 , n59060 , n59061 , n59062 , n9698 , n59064 , n59065 , n59066 , n59067 , 
     n59068 , n59069 , n59070 , n9706 , n59072 , n9708 , n59074 , n9710 , n59076 , n9712 , 
     n59078 , n59079 , n9715 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , 
     n9721 , n59089 , n59090 , n59091 , n59092 , n59093 , n9727 , n59095 , n59096 , n9730 , 
     n9731 , n9732 , n59100 , n59101 , n9735 , n59103 , n9737 , n9738 , n59106 , n9740 , 
     n59108 , n59109 , n9743 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , 
     n59118 , n59119 , n59120 , n9754 , n59122 , n59123 , n9757 , n9758 , n59126 , n9760 , 
     n59128 , n59129 , n9763 , n59131 , n59132 , n59133 , n9766 , n9767 , n9768 , n59137 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n59143 , n59144 , n59145 , n59146 , n9779 , 
     n9780 , n59149 , n59150 , n59151 , n59152 , n9785 , n9786 , n59155 , n59156 , n9789 , 
     n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n9796 , n59165 , n59166 , n59167 , 
     n9800 , n59169 , n59170 , n9803 , n59172 , n59173 , n59174 , n59175 , n9808 , n9809 , 
     n59178 , n9811 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n9816 , n9817 , 
     n59188 , n59189 , n59190 , n59191 , n9822 , n59193 , n59194 , n59195 , n59196 , n9827 , 
     n59198 , n59199 , n9830 , n9831 , n59202 , n9833 , n9834 , n59205 , n9836 , n59207 , 
     n9838 , n59209 , n59210 , n9841 , n59212 , n59213 , n59214 , n59215 , n59216 , n9847 , 
     n59218 , n59219 , n9850 , n59221 , n59222 , n59223 , n9854 , n59225 , n9856 , n9857 , 
     n59228 , n9859 , n59230 , n59231 , n59232 , n59233 , n9864 , n59235 , n9866 , n9867 , 
     n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n9877 , 
     n59248 , n59249 , n59250 , n59251 , n9882 , n59253 , n59254 , n59255 , n59256 , n59257 , 
     n9888 , n59259 , n9890 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n9897 , 
     n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n9906 , n59277 , 
     n9908 , n9909 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , 
     n59288 , n9919 , n59290 , n9921 , n9922 , n9923 , n59294 , n59295 , n9926 , n59297 , 
     n9928 , n59299 , n59300 , n59301 , n9932 , n59303 , n59304 , n9935 , n59306 , n59307 , 
     n59308 , n59309 , n59310 , n59311 , n9942 , n59313 , n59314 , n9945 , n59316 , n59317 , 
     n9948 , n59319 , n59320 , n59321 , n9952 , n59323 , n59324 , n9955 , n59326 , n9957 , 
     n9958 , n59329 , n59330 , n9961 , n9962 , n59333 , n59334 , n9965 , n59336 , n59337 , 
     n9968 , n59339 , n59340 , n59341 , n59342 , n9973 , n59344 , n9975 , n59346 , n59347 , 
     n59348 , n59349 , n59350 , n9981 , n59352 , n59353 , n59354 , n59355 , n59356 , n9987 , 
     n9988 , n59359 , n59360 , n59361 , n59362 , n59363 , n9994 , n59365 , n59366 , n59367 , 
     n59368 , n59369 , n59370 , n59371 , n10002 , n10003 , n59374 , n59375 , n10005 , n59377 , 
     n59378 , n59379 , n59380 , n10010 , n59382 , n59383 , n59384 , n59385 , n10015 , n10016 , 
     n59388 , n10018 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n10025 , n59397 , 
     n59398 , n59399 , n10029 , n59401 , n59402 , n10032 , n59404 , n59405 , n59406 , n10036 , 
     n59408 , n59409 , n59410 , n10040 , n59412 , n59413 , n10043 , n59415 , n59416 , n10046 , 
     n10047 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n10054 , n10055 , n59427 , 
     n59428 , n59429 , n59430 , n59431 , n59432 , n10062 , n59434 , n10064 , n59436 , n10066 , 
     n10067 , n59439 , n59440 , n59441 , n59442 , n59443 , n10073 , n59445 , n59446 , n59447 , 
     n59448 , n59449 , n59450 , n10080 , n59452 , n59453 , n59454 , n10084 , n59456 , n10086 , 
     n59458 , n59459 , n59460 , n59461 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , 
     n10097 , n10098 , n10099 , n59471 , n10101 , n59473 , n10103 , n10104 , n10105 , n10106 , 
     n59478 , n10108 , n59480 , n59481 , n59482 , n10112 , n59484 , n10114 , n10115 , n10116 , 
     n59488 , n59489 , n10119 , n59491 , n10121 , n59493 , n10123 , n59495 , n10125 , n59497 , 
     n10127 , n10128 , n10129 , n59501 , n10131 , n10132 , n59504 , n59505 , n10135 , n59507 , 
     n59508 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , 
     n10147 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n10155 , n10156 , 
     n10157 , n10158 , n10159 , n10160 , n59532 , n59533 , n10163 , n59535 , n10165 , n59537 , 
     n10167 , n10168 , n10169 , n59541 , n10171 , n59543 , n10173 , n59545 , n59546 , n10176 , 
     n59548 , n59549 , n10179 , n59551 , n10181 , n59553 , n59554 , n10184 , n59556 , n59557 , 
     n10187 , n59559 , n59560 , n10190 , n59562 , n10192 , n59564 , n59565 , n10195 , n59567 , 
     n59568 , n10198 , n59570 , n59571 , n10201 , n10202 , n59574 , n59575 , n59576 , n59577 , 
     n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , 
     n59588 , n59589 , n10219 , n59591 , n59592 , n10222 , n59594 , n10224 , n59596 , n10226 , 
     n59598 , n10228 , n10229 , n10230 , n59602 , n59603 , n59604 , n10234 , n59606 , n59607 , 
     n10237 , n59609 , n59610 , n10240 , n59612 , n59613 , n10243 , n59615 , n59616 , n10246 , 
     n59618 , n10248 , n10249 , n59621 , n10251 , n59623 , n59624 , n59625 , n59626 , n59627 , 
     n59628 , n59629 , n59630 , n59631 , n59632 , n10262 , n59634 , n59635 , n10264 , n10265 , 
     n59638 , n59639 , n59640 , n59641 , n10270 , n59643 , n59644 , n59645 , n59646 , n59647 , 
     n59648 , n59649 , n10278 , n59651 , n59652 , n59653 , n59654 , n59655 , n10284 , n59657 , 
     n59658 , n10287 , n59660 , n59661 , n59662 , n59663 , n10292 , n10293 , n59666 , n59667 , 
     n10296 , n10297 , n10298 , n59671 , n59672 , n59673 , n59674 , n10301 , n59676 , n10303 , 
     n10304 , n10305 , n59680 , n10307 , n59682 , n59683 , n59684 , n59685 , n10312 , n59687 , 
     n10314 , n10315 , n59690 , n10317 , n59692 , n10319 , n59694 , n59695 , n59696 , n59697 , 
     n59698 , n59699 , n59700 , n59701 , n59702 , n10329 , n59704 , n59705 , n59706 , n59707 , 
     n10334 , n10335 , n59710 , n10337 , n10338 , n59713 , n59714 , n10341 , n59716 , n10343 , 
     n59718 , n59719 , n59720 , n10347 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , 
     n59728 , n59729 , n59730 , n10357 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , 
     n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n10371 , n59746 , n59747 , 
     n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n10381 , n59756 , n10383 , 
     n59758 , n10385 , n10386 , n59761 , n10388 , n59763 , n10390 , n59765 , n59766 , n59767 , 
     n10394 , n59769 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , 
     n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , 
     n10414 , n59789 , n59790 , n59791 , n59792 , n59793 , n10420 , n59795 , n10422 , n59797 , 
     n59798 , n10425 , n59800 , n59801 , n59802 , n10429 , n59804 , n59805 , n10432 , n10433 , 
     n59808 , n10435 , n59810 , n10437 , n59812 , n59813 , n59814 , n10441 , n59816 , n10443 , 
     n59818 , n10445 , n59820 , n10447 , n59822 , n10449 , n59824 , n10451 , n59826 , n10453 , 
     n10454 , n59829 , n10456 , n59831 , n59832 , n59833 , n10460 , n59835 , n59836 , n10463 , 
     n10464 , n59839 , n59840 , n10467 , n10468 , n59843 , n59844 , n59845 , n59846 , n59847 , 
     n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , 
     n59858 , n10485 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , 
     n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n10500 , n59875 , n10502 , n59877 , 
     n59878 , n59879 , n10506 , n59881 , n59882 , n10509 , n59884 , n59885 , n10512 , n59887 , 
     n10514 , n59889 , n59890 , n59891 , n10518 , n10519 , n10520 , n10521 , n59896 , n10523 , 
     n59898 , n10525 , n59900 , n10527 , n59902 , n10529 , n59904 , n10531 , n10532 , n59907 , 
     n59908 , n10535 , n10536 , n59911 , n59912 , n59913 , n59914 , n59915 , n10542 , n59917 , 
     n59918 , n10545 , n10546 , n59921 , n59922 , n59923 , n59924 , n59925 , n10552 , n59927 , 
     n59928 , n10555 , n10556 , n59931 , n59932 , n10559 , n59934 , n10561 , n59936 , n10563 , 
     n59938 , n59939 , n10566 , n59941 , n59942 , n10569 , n59944 , n59945 , n59946 , n10573 , 
     n59948 , n59949 , n10576 , n10577 , n59952 , n59953 , n59954 , n59955 , n59956 , n10583 , 
     n10584 , n59959 , n59960 , n10587 , n10588 , n59963 , n59964 , n10591 , n59966 , n10593 , 
     n10594 , n10595 , n10596 , n59971 , n59972 , n10599 , n10600 , n59975 , n59976 , n10603 , 
     n59978 , n59979 , n59980 , n59981 , n59982 , n10609 , n59984 , n10611 , n59986 , n10613 , 
     n59988 , n10615 , n10616 , n10617 , n10618 , n10619 , n59994 , n59995 , n59996 , n10623 , 
     n10624 , n59999 , n60000 , n10627 , n60002 , n60003 , n10630 , n60005 , n60006 , n10633 , 
     n10634 , n10635 , n60010 , n60011 , n10638 , n10639 , n10640 , n60015 , n60016 , n10643 , 
     n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , 
     n60028 , n60029 , n60030 , n10657 , n10658 , n10659 , n10660 , n10661 , n60036 , n10663 , 
     n60038 , n60039 , n10666 , n10667 , n60042 , n10669 , n60044 , n60045 , n60046 , n60047 , 
     n10674 , n60049 , n10676 , n60051 , n60052 , n10679 , n60054 , n60055 , n10682 , n60057 , 
     n60058 , n10685 , n60060 , n60061 , n60062 , n10689 , n60064 , n60065 , n10692 , n10693 , 
     n60068 , n10695 , n60070 , n10697 , n10698 , n10699 , n10700 , n10701 , n60076 , n60077 , 
     n10704 , n60079 , n60080 , n60081 , n10708 , n60083 , n10710 , n10711 , n60086 , n60087 , 
     n60088 , n60089 , n10716 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , 
     n60098 , n60099 , n60100 , n60101 , n10728 , n60103 , n60104 , n60105 , n60106 , n10733 , 
     n10734 , n60109 , n60110 , n10737 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , 
     n60118 , n60119 , n60120 , n60121 , n60122 , n10749 , n60124 , n60125 , n10752 , n60127 , 
     n60128 , n10755 , n60130 , n60131 , n10758 , n60133 , n60134 , n10761 , n60136 , n60137 , 
     n10764 , n60139 , n60140 , n60141 , n60142 , n60143 , n10770 , n60145 , n60146 , n10773 , 
     n60148 , n10775 , n60150 , n10777 , n60152 , n60153 , n10780 , n10781 , n60156 , n60157 , 
     n10784 , n60159 , n60160 , n10787 , n10788 , n10789 , n10790 , n60165 , n10792 , n10793 , 
     n60168 , n10795 , n60170 , n60171 , n10798 , n60173 , n60174 , n60175 , n10802 , n60177 , 
     n60178 , n60179 , n10806 , n60181 , n10808 , n60183 , n60184 , n60185 , n60186 , n60187 , 
     n60188 , n10815 , n60190 , n60191 , n60192 , n60193 , n10820 , n60195 , n60196 , n10823 , 
     n60198 , n60199 , n60200 , n10827 , n60202 , n60203 , n10830 , n10831 , n60206 , n10833 , 
     n60208 , n10835 , n60210 , n60211 , n60212 , n10839 , n60214 , n60215 , n10842 , n60217 , 
     n60218 , n10845 , n60220 , n60221 , n10848 , n60223 , n60224 , n10851 , n60226 , n10853 , 
     n60228 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n60236 , n10863 , 
     n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n10873 , 
     n60248 , n60249 , n60250 , n60251 , n60252 , n10879 , n60254 , n60255 , n10882 , n60257 , 
     n60258 , n60259 , n60260 , n60261 , n60262 , n10889 , n60264 , n60265 , n60266 , n60267 , 
     n60268 , n60269 , n10896 , n60271 , n10898 , n60273 , n10900 , n60275 , n60276 , n60277 , 
     n60278 , n60279 , n60280 , n60281 , n10908 , n60283 , n60284 , n60285 , n60286 , n10913 , 
     n10914 , n60289 , n10916 , n60291 , n10918 , n60293 , n60294 , n10921 , n60296 , n60297 , 
     n60298 , n60299 , n10926 , n60301 , n60302 , n10929 , n10930 , n60305 , n60306 , n10933 , 
     n60308 , n60309 , n10936 , n60311 , n60312 , n10939 , n60314 , n10941 , n10942 , n10943 , 
     n60318 , n10945 , n60320 , n60321 , n10948 , n60323 , n60324 , n10951 , n10952 , n10953 , 
     n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n60334 , n60335 , n60336 , n10963 , 
     n60338 , n60339 , n10966 , n60341 , n60342 , n10969 , n10970 , n60345 , n10972 , n10973 , 
     n60348 , n60349 , n10976 , n60351 , n60352 , n10979 , n60354 , n60355 , n60356 , n10983 , 
     n60358 , n10985 , n10986 , n10987 , n10988 , n60363 , n10990 , n60365 , n10992 , n10993 , 
     n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , 
     n11004 , n60379 , n11006 , n60381 , n11008 , n11009 , n11010 , n11011 , n11012 , n60387 , 
     n11014 , n60389 , n60390 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , 
     n60398 , n11025 , n60400 , n60401 , n11028 , n60403 , n60404 , n11031 , n11032 , n11033 , 
     n11034 , n60409 , n60410 , n11037 , n60412 , n60413 , n11040 , n60415 , n60416 , n60417 , 
     n11044 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n11053 , 
     n60428 , n11055 , n60430 , n60431 , n60432 , n60433 , n60434 , n11061 , n60436 , n11063 , 
     n60438 , n60439 , n11066 , n60441 , n60442 , n11069 , n11070 , n60445 , n60446 , n60447 , 
     n60448 , n60449 , n60450 , n60451 , n11078 , n11079 , n11080 , n11081 , n11082 , n60457 , 
     n60458 , n11085 , n11086 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , 
     n11094 , n11095 , n60470 , n60471 , n60472 , n11099 , n60474 , n11101 , n60476 , n60477 , 
     n60478 , n11105 , n60480 , n11107 , n60482 , n11109 , n11110 , n60485 , n11112 , n60487 , 
     n60488 , n11115 , n11116 , n60491 , n60492 , n11119 , n60494 , n60495 , n11122 , n11123 , 
     n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n11130 , n60505 , n60506 , n11133 , 
     n11134 , n60509 , n11136 , n60511 , n60512 , n11139 , n60514 , n60515 , n60516 , n11143 , 
     n11144 , n60519 , n11146 , n60521 , n11148 , n60523 , n60524 , n60525 , n11152 , n60527 , 
     n60528 , n11155 , n11156 , n60531 , n60532 , n11159 , n60534 , n60535 , n60536 , n60537 , 
     n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n11173 , 
     n11174 , n11175 , n11176 , n60551 , n11178 , n11179 , n60554 , n11181 , n60556 , n60557 , 
     n11184 , n11185 , n60560 , n11187 , n11188 , n60563 , n11190 , n11191 , n60566 , n11193 , 
     n60568 , n11195 , n60570 , n11197 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , 
     n60578 , n60579 , n60580 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , 
     n11214 , n11215 , n11216 , n11217 , n60592 , n11219 , n60594 , n60595 , n60596 , n60597 , 
     n60598 , n11225 , n60600 , n60601 , n11228 , n60603 , n11230 , n11231 , n11232 , n11233 , 
     n60608 , n60609 , n11236 , n60611 , n60612 , n11239 , n60614 , n11241 , n11242 , n11243 , 
     n11244 , n60619 , n11246 , n60621 , n11248 , n11249 , n11250 , n11251 , n60626 , n11253 , 
     n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , 
     n11264 , n11265 , n11266 , n11267 , n60642 , n11269 , n60644 , n60645 , n11272 , n60647 , 
     n60648 , n11275 , n11276 , n60651 , n11278 , n11279 , n11280 , n11281 , n60656 , n11283 , 
     n60658 , n60659 , n11286 , n60661 , n11288 , n60663 , n60664 , n11291 , n60666 , n60667 , 
     n11294 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , 
     n60678 , n11305 , n60680 , n60681 , n11308 , n60683 , n60684 , n11311 , n60686 , n60687 , 
     n60688 , n60689 , n60690 , n60691 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , 
     n60698 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , 
     n11334 , n60709 , n11336 , n60711 , n60712 , n11339 , n60714 , n60715 , n11342 , n11343 , 
     n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , 
     n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , 
     n11364 , n60739 , n11366 , n60741 , n60742 , n11369 , n60744 , n60745 , n11372 , n60747 , 
     n60748 , n60749 , n60750 , n60751 , n60752 , n11379 , n11380 , n60755 , n11382 , n60757 , 
     n60758 , n60759 , n60760 , n60761 , n11388 , n60763 , n60764 , n60765 , n60766 , n60767 , 
     n60768 , n60769 , n60770 , n60771 , n11398 , n11399 , n11400 , n60775 , n11402 , n60777 , 
     n11404 , n11405 , n11406 , n60781 , n11408 , n60783 , n60784 , n11411 , n60786 , n60787 , 
     n11414 , n60789 , n60790 , n11417 , n60792 , n60793 , n11420 , n60795 , n11422 , n11423 , 
     n60798 , n11425 , n60800 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n60807 , 
     n60808 , n11435 , n60810 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , 
     n11444 , n60819 , n11446 , n60821 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , 
     n11454 , n11455 , n11456 , n60831 , n11458 , n11459 , n11460 , n11461 , n60836 , n60837 , 
     n60838 , n11465 , n60840 , n60841 , n11468 , n60843 , n60844 , n60845 , n11472 , n11473 , 
     n11474 , n60849 , n60850 , n60851 , n60852 , n11479 , n60854 , n11481 , n11482 , n11483 , 
     n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n60865 , n11492 , n60867 , 
     n11494 , n11495 , n60870 , n60871 , n11498 , n60873 , n11500 , n60875 , n60876 , n11503 , 
     n60878 , n11505 , n11506 , n60881 , n60882 , n11509 , n60884 , n11511 , n11512 , n11513 , 
     n11514 , n60889 , n60890 , n11517 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , 
     n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n60906 , n11533 , 
     n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n60916 , n60917 , 
     n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n11553 , 
     n60928 , n11555 , n60930 , n60931 , n11558 , n60933 , n11560 , n11561 , n11562 , n11563 , 
     n11564 , n11565 , n60940 , n60941 , n11568 , n60943 , n11570 , n60945 , n60946 , n60947 , 
     n60948 , n60949 , n60950 , n11577 , n11578 , n60953 , n60954 , n60955 , n11582 , n60957 , 
     n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n11590 , n60965 , n60966 , n60967 , 
     n11594 , n60969 , n11596 , n60971 , n60972 , n60973 , n11600 , n11601 , n11602 , n11603 , 
     n11604 , n60979 , n11606 , n60981 , n11608 , n11609 , n11610 , n11611 , n11612 , n60987 , 
     n11614 , n60989 , n11616 , n11617 , n60992 , n11619 , n60994 , n11621 , n11622 , n11623 , 
     n11624 , n11625 , n11626 , n61001 , n11628 , n61003 , n61004 , n61005 , n61006 , n61007 , 
     n11634 , n61009 , n11636 , n61011 , n11638 , n11639 , n61014 , n11641 , n61016 , n61017 , 
     n11644 , n61019 , n61020 , n61021 , n11648 , n61023 , n61024 , n11651 , n61026 , n61027 , 
     n11654 , n61029 , n61030 , n11657 , n61032 , n11659 , n11660 , n61035 , n11662 , n61037 , 
     n11664 , n61039 , n61040 , n11667 , n61042 , n11669 , n11670 , n11671 , n11672 , n11673 , 
     n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , 
     n11684 , n11685 , n11686 , n11687 , n61062 , n11689 , n61064 , n11691 , n11692 , n11693 , 
     n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n61077 , 
     n11704 , n61079 , n61080 , n11707 , n61082 , n11709 , n61084 , n11711 , n61086 , n11713 , 
     n61088 , n11715 , n11716 , n61091 , n61092 , n11719 , n61094 , n11721 , n61096 , n11723 , 
     n61098 , n11725 , n11726 , n11727 , n11728 , n61103 , n11730 , n11731 , n61106 , n61107 , 
     n11734 , n61109 , n61110 , n11737 , n61112 , n11739 , n61114 , n11741 , n61116 , n11743 , 
     n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n61125 , n61126 , n11753 , 
     n61128 , n61129 , n11756 , n61131 , n61132 , n11759 , n61134 , n61135 , n11762 , n11763 , 
     n11764 , n61139 , n11766 , n61141 , n11768 , n11769 , n11770 , n11771 , n61146 , n61147 , 
     n11774 , n61149 , n61150 , n11777 , n61152 , n61153 , n11780 , n61155 , n61156 , n61157 , 
     n61158 , n61159 , n11786 , n61161 , n11788 , n61163 , n11790 , n11791 , n11792 , n11793 , 
     n61168 , n11795 , n11796 , n11797 , n11798 , n61173 , n11800 , n61175 , n11802 , n61177 , 
     n61178 , n11805 , n61180 , n11807 , n61182 , n11809 , n61184 , n61185 , n61186 , n61187 , 
     n61188 , n11815 , n61190 , n11817 , n11818 , n11819 , n11820 , n11821 , n61196 , n61197 , 
     n11824 , n61199 , n61200 , n61201 , n61202 , n11829 , n11830 , n61205 , n61206 , n61207 , 
     n61208 , n11835 , n61210 , n11837 , n61212 , n61213 , n61214 , n11841 , n61216 , n11843 , 
     n11844 , n11845 , n11846 , n11847 , n11848 , n61223 , n11850 , n61225 , n61226 , n61227 , 
     n11854 , n61229 , n11856 , n11857 , n61232 , n61233 , n11860 , n11861 , n61236 , n61237 , 
     n61238 , n61239 , n61240 , n61241 , n11868 , n11869 , n61244 , n11871 , n61246 , n61247 , 
     n61248 , n61249 , n11876 , n61251 , n61252 , n61253 , n11880 , n61255 , n61256 , n11883 , 
     n61258 , n61259 , n61260 , n11887 , n61262 , n61263 , n11890 , n61265 , n61266 , n11893 , 
     n11894 , n11895 , n61270 , n61271 , n11898 , n61273 , n11900 , n11901 , n11902 , n61277 , 
     n11904 , n61279 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n61287 , 
     n11914 , n61289 , n11916 , n11917 , n61292 , n11919 , n61294 , n11921 , n11922 , n61297 , 
     n61298 , n11925 , n61300 , n11927 , n61302 , n61303 , n11930 , n61305 , n61306 , n61307 , 
     n61308 , n61309 , n11936 , n61311 , n61312 , n11939 , n11940 , n11941 , n11942 , n11943 , 
     n61318 , n11945 , n11946 , n61321 , n61322 , n11949 , n61324 , n61325 , n11952 , n61327 , 
     n61328 , n61329 , n61330 , n61331 , n11958 , n11959 , n61334 , n61335 , n11962 , n61337 , 
     n11964 , n11965 , n61340 , n11967 , n61342 , n61343 , n11970 , n61345 , n11972 , n61347 , 
     n11974 , n61349 , n61350 , n11977 , n61352 , n11979 , n11980 , n61355 , n11982 , n61357 , 
     n11984 , n61359 , n61360 , n11987 , n61362 , n61363 , n11990 , n61365 , n61366 , n61367 , 
     n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n12002 , n12003 , 
     n12004 , n12005 , n12006 , n12007 , n61382 , n12009 , n61384 , n12011 , n61386 , n12013 , 
     n61388 , n12015 , n61390 , n12017 , n61392 , n12019 , n12020 , n12021 , n12022 , n12023 , 
     n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n61404 , n61405 , n12032 , n61407 , 
     n12034 , n61409 , n12036 , n12037 , n61412 , n61413 , n12040 , n61415 , n61416 , n12043 , 
     n61418 , n61419 , n12046 , n12047 , n61422 , n61423 , n12050 , n61425 , n61426 , n61427 , 
     n61428 , n61429 , n12056 , n61431 , n61432 , n61433 , n12060 , n12061 , n12062 , n61437 , 
     n12064 , n12065 , n12066 , n61441 , n61442 , n12069 , n61444 , n61445 , n61446 , n61447 , 
     n61448 , n12075 , n61450 , n61451 , n12078 , n61453 , n61454 , n61455 , n61456 , n12083 , 
     n12084 , n12085 , n12086 , n61461 , n12088 , n12089 , n61464 , n61465 , n61466 , n61467 , 
     n12094 , n12095 , n12096 , n12097 , n61472 , n12099 , n12100 , n61475 , n61476 , n12103 , 
     n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n12110 , n61485 , n12112 , n12113 , 
     n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n61494 , n12121 , n61496 , n61497 , 
     n12124 , n12125 , n61500 , n12127 , n61502 , n12129 , n61504 , n61505 , n12132 , n61507 , 
     n61508 , n61509 , n61510 , n12137 , n61512 , n61513 , n12140 , n61515 , n61516 , n61517 , 
     n61518 , n12145 , n61520 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , 
     n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , 
     n61538 , n12165 , n61540 , n61541 , n61542 , n61543 , n61544 , n12171 , n61546 , n12173 , 
     n12174 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n12181 , n12182 , n61557 , 
     n12184 , n61559 , n61560 , n61561 , n12188 , n61563 , n61564 , n61565 , n61566 , n61567 , 
     n61568 , n12195 , n61570 , n61571 , n12198 , n61573 , n61574 , n61575 , n12202 , n61577 , 
     n61578 , n61579 , n61580 , n12207 , n61582 , n61583 , n61584 , n61585 , n12212 , n61587 , 
     n61588 , n12215 , n61590 , n61591 , n61592 , n12219 , n61594 , n61595 , n12222 , n61597 , 
     n12224 , n61599 , n61600 , n61601 , n12228 , n61603 , n12230 , n61605 , n61606 , n12233 , 
     n61608 , n12235 , n12236 , n61611 , n12238 , n61613 , n61614 , n61615 , n12242 , n61617 , 
     n12244 , n61619 , n12246 , n61621 , n12248 , n12249 , n12250 , n61625 , n61626 , n12253 , 
     n61628 , n61629 , n61630 , n61631 , n12258 , n61633 , n12260 , n12261 , n12262 , n61637 , 
     n61638 , n12265 , n61640 , n12267 , n61642 , n12269 , n12270 , n61645 , n12272 , n61647 , 
     n12274 , n12275 , n12276 , n12277 , n61652 , n12279 , n61654 , n61655 , n12282 , n61657 , 
     n61658 , n12285 , n61660 , n12287 , n12288 , n61663 , n61664 , n12291 , n61666 , n61667 , 
     n61668 , n61669 , n61670 , n61671 , n12298 , n61673 , n12300 , n12301 , n12302 , n12303 , 
     n12304 , n12305 , n12306 , n12307 , n12308 , n61683 , n12310 , n12311 , n61686 , n12313 , 
     n61688 , n61689 , n61690 , n12317 , n12318 , n12319 , n61694 , n61695 , n12322 , n61697 , 
     n61698 , n12325 , n61700 , n61701 , n12328 , n61703 , n61704 , n12331 , n61706 , n61707 , 
     n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n61715 , n61716 , n12343 , 
     n61718 , n12345 , n61720 , n12347 , n61722 , n12349 , n12350 , n12351 , n61726 , n61727 , 
     n12354 , n12355 , n12356 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n12363 , 
     n12364 , n61739 , n61740 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n61747 , 
     n61748 , n61749 , n61750 , n12377 , n12378 , n61753 , n12380 , n61755 , n61756 , n61757 , 
     n12384 , n61759 , n12386 , n61761 , n61762 , n61763 , n12390 , n61765 , n61766 , n12393 , 
     n61768 , n61769 , n12396 , n12397 , n12398 , n12399 , n61774 , n12401 , n12402 , n61777 , 
     n61778 , n61779 , n61780 , n12407 , n12408 , n12409 , n61784 , n12411 , n12412 , n61787 , 
     n61788 , n12415 , n61790 , n12417 , n61792 , n12419 , n12420 , n12421 , n12422 , n12423 , 
     n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n61807 , 
     n61808 , n61809 , n12433 , n12434 , n12435 , n61813 , n12437 , n61815 , n12439 , n12440 , 
     n12441 , n12442 , n12443 , n61821 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , 
     n12451 , n12452 , n61830 , n12454 , n61832 , n12456 , n12457 , n61835 , n61836 , n12460 , 
     n61838 , n61839 , n12463 , n61841 , n61842 , n61843 , n12467 , n61845 , n61846 , n12470 , 
     n12471 , n61849 , n12473 , n61851 , n61852 , n12476 , n12477 , n61855 , n61856 , n12480 , 
     n12481 , n61859 , n61860 , n12484 , n61862 , n61863 , n12487 , n12488 , n12489 , n12490 , 
     n12491 , n12492 , n12493 , n61871 , n12495 , n61873 , n12497 , n12498 , n12499 , n61877 , 
     n12501 , n61879 , n12503 , n61881 , n12505 , n12506 , n61884 , n61885 , n12509 , n12510 , 
     n61888 , n12512 , n61890 , n61891 , n61892 , n12516 , n12517 , n12518 , n61896 , n12520 , 
     n61898 , n61899 , n12523 , n61901 , n61902 , n12526 , n61904 , n61905 , n61906 , n61907 , 
     n61908 , n61909 , n12533 , n61911 , n12535 , n12536 , n12537 , n12538 , n61916 , n61917 , 
     n12541 , n61919 , n12543 , n61921 , n61922 , n12546 , n61924 , n61925 , n12549 , n61927 , 
     n61928 , n61929 , n61930 , n12554 , n61932 , n12556 , n12557 , n61935 , n61936 , n12560 , 
     n12561 , n12562 , n61940 , n12564 , n61942 , n12566 , n12567 , n61945 , n12569 , n12570 , 
     n12571 , n61949 , n61950 , n61951 , n12575 , n61953 , n61954 , n61955 , n61956 , n61957 , 
     n61958 , n61959 , n12583 , n61961 , n61962 , n61963 , n61964 , n12588 , n61966 , n61967 , 
     n12591 , n61969 , n61970 , n61971 , n12595 , n61973 , n12597 , n61975 , n61976 , n61977 , 
     n61978 , n61979 , n61980 , n12604 , n61982 , n12606 , n12607 , n12608 , n12609 , n12610 , 
     n12611 , n61989 , n61990 , n61991 , n12615 , n61993 , n12617 , n12618 , n12619 , n12620 , 
     n61998 , n12622 , n62000 , n62001 , n12625 , n62003 , n62004 , n62005 , n62006 , n12630 , 
     n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n12637 , n62015 , n62016 , n62017 , 
     n12641 , n62019 , n12643 , n62021 , n62022 , n62023 , n62024 , n62025 , n12645 , n62027 , 
     n62028 , n12648 , n12649 , n12650 , n62032 , n12652 , n12653 , n12654 , n12655 , n12656 , 
     n62038 , n62039 , n62040 , n12657 , n12658 , n12659 , n62044 , n12661 , n62046 , n12663 , 
     n62048 , n12665 , n12666 , n62051 , n62052 , n62053 , n62054 , n62055 , n12672 , n62057 , 
     n62058 , n12675 , n62060 , n12677 , n62062 , n12679 , n12680 , n12681 , n12682 , n12683 , 
     n62068 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n62075 , n12692 , n62077 , 
     n12694 , n12695 , n12696 , n12697 , n12698 , n62083 , n12700 , n62085 , n62086 , n62087 , 
     n62088 , n62089 , n12706 , n12707 , n62092 , n62093 , n12710 , n62095 , n62096 , n12713 , 
     n62098 , n62099 , n12716 , n12717 , n62102 , n62103 , n12720 , n62105 , n62106 , n12723 , 
     n12724 , n62109 , n62110 , n12727 , n62112 , n62113 , n12730 , n12731 , n62116 , n12733 , 
     n62118 , n62119 , n12736 , n62121 , n62122 , n12739 , n12740 , n12741 , n12742 , n12743 , 
     n12744 , n12745 , n62130 , n12747 , n62132 , n12749 , n12750 , n62135 , n62136 , n62137 , 
     n12754 , n62139 , n12756 , n12757 , n12758 , n12759 , n62144 , n12761 , n62146 , n12763 , 
     n12764 , n12765 , n12766 , n12767 , n62152 , n62153 , n62154 , n12771 , n62156 , n62157 , 
     n62158 , n12775 , n12776 , n62161 , n12778 , n62163 , n62164 , n12781 , n62166 , n12783 , 
     n62168 , n62169 , n62170 , n12787 , n62172 , n62173 , n62174 , n62175 , n12792 , n62177 , 
     n62178 , n12795 , n62180 , n12797 , n12798 , n12799 , n62184 , n62185 , n12802 , n62187 , 
     n12804 , n62189 , n62190 , n12807 , n62192 , n62193 , n12810 , n12811 , n62196 , n62197 , 
     n62198 , n12815 , n62200 , n62201 , n12818 , n62203 , n12820 , n12821 , n62206 , n62207 , 
     n12824 , n62209 , n12826 , n62211 , n62212 , n12829 , n62214 , n62215 , n12832 , n12833 , 
     n12834 , n62219 , n62220 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n62227 , 
     n12844 , n62229 , n12846 , n62231 , n12848 , n62233 , n62234 , n62235 , n12852 , n62237 , 
     n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , 
     n12864 , n12865 , n62250 , n12867 , n62252 , n12869 , n12870 , n12871 , n12872 , n12873 , 
     n12874 , n12875 , n12876 , n12877 , n12878 , n62263 , n12880 , n12881 , n12882 , n12883 , 
     n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n62274 , n12891 , n12892 , n62277 , 
     n12894 , n62279 , n12896 , n62281 , n12898 , n12899 , n12900 , n62285 , n62286 , n12903 , 
     n12904 , n62289 , n12906 , n62291 , n62292 , n62293 , n62294 , n12911 , n62296 , n12913 , 
     n12914 , n12915 , n12916 , n62301 , n62302 , n62303 , n12920 , n62305 , n12922 , n62307 , 
     n62308 , n12925 , n62310 , n12927 , n12928 , n62313 , n62314 , n12931 , n62316 , n12933 , 
     n62318 , n62319 , n12936 , n62321 , n62322 , n12939 , n62324 , n62325 , n12942 , n62327 , 
     n62328 , n62329 , n62330 , n12947 , n12948 , n12949 , n12950 , n62335 , n62336 , n12953 , 
     n62338 , n12955 , n12956 , n62341 , n62342 , n12959 , n12960 , n62345 , n12962 , n62347 , 
     n12964 , n62349 , n12966 , n12967 , n62352 , n62353 , n12970 , n12971 , n12972 , n62357 , 
     n62358 , n62359 , n12976 , n62361 , n62362 , n62363 , n62364 , n62365 , n12982 , n12983 , 
     n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n12992 , n62377 , 
     n62378 , n62379 , n62380 , n62381 , n62382 , n12999 , n13000 , n13001 , n13002 , n13003 , 
     n13004 , n13005 , n13006 , n62391 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , 
     n62398 , n62399 , n13016 , n62401 , n13018 , n13019 , n13020 , n62405 , n13022 , n62407 , 
     n13024 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n13031 , n62416 , n13033 , 
     n62418 , n13035 , n62420 , n62421 , n13038 , n62423 , n62424 , n62425 , n13042 , n62427 , 
     n62428 , n13045 , n13046 , n62431 , n13048 , n13049 , n62434 , n62435 , n62436 , n62437 , 
     n13054 , n62439 , n62440 , n13057 , n13058 , n13059 , n13060 , n62445 , n62446 , n62447 , 
     n62448 , n62449 , n62450 , n62451 , n62452 , n13069 , n62454 , n62455 , n62456 , n13073 , 
     n62458 , n13075 , n62460 , n13077 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , 
     n13084 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , 
     n13094 , n62479 , n13096 , n62481 , n62482 , n13099 , n62484 , n62485 , n13102 , n62487 , 
     n13104 , n62489 , n62490 , n62491 , n13108 , n62493 , n13110 , n62495 , n62496 , n62497 , 
     n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n13121 , n13122 , n62507 , 
     n13124 , n62509 , n62510 , n13127 , n13128 , n62513 , n62514 , n13131 , n13132 , n62517 , 
     n62518 , n62519 , n13136 , n13137 , n13138 , n62523 , n13140 , n62525 , n62526 , n62527 , 
     n13144 , n62529 , n13146 , n62531 , n62532 , n13149 , n62534 , n13151 , n13152 , n62537 , 
     n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n13160 , n62545 , n62546 , n13163 , 
     n62548 , n13165 , n62550 , n62551 , n13168 , n62553 , n13170 , n13171 , n13172 , n13173 , 
     n13174 , n13175 , n13176 , n62561 , n13178 , n62563 , n13180 , n62565 , n62566 , n13183 , 
     n62568 , n13185 , n62570 , n62571 , n13188 , n13189 , n13190 , n13191 , n62576 , n13193 , 
     n62578 , n62579 , n13196 , n62581 , n13198 , n13199 , n13200 , n13201 , n13202 , n62587 , 
     n62588 , n62589 , n13206 , n62591 , n13208 , n62593 , n13210 , n62595 , n62596 , n13213 , 
     n62598 , n62599 , n13216 , n13217 , n13218 , n62603 , n62604 , n13221 , n62606 , n62607 , 
     n62608 , n62609 , n62610 , n13227 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , 
     n62618 , n13235 , n62620 , n13237 , n62622 , n62623 , n62624 , n62625 , n13242 , n13243 , 
     n62628 , n62629 , n62630 , n13247 , n62632 , n62633 , n62634 , n62635 , n62636 , n13253 , 
     n62638 , n62639 , n62640 , n13257 , n62642 , n62643 , n13260 , n13261 , n62646 , n62647 , 
     n13264 , n13265 , n62650 , n13267 , n62652 , n62653 , n62654 , n13271 , n62656 , n13273 , 
     n62658 , n62659 , n13276 , n62661 , n62662 , n13279 , n13280 , n13281 , n13282 , n62667 , 
     n62668 , n13285 , n62670 , n62671 , n13288 , n62673 , n62674 , n62675 , n62676 , n13293 , 
     n62678 , n13295 , n62680 , n13297 , n62682 , n62683 , n13300 , n62685 , n13302 , n62687 , 
     n62688 , n13305 , n62690 , n13307 , n62692 , n13309 , n62694 , n62695 , n62696 , n62697 , 
     n62698 , n62699 , n62700 , n62701 , n13318 , n13319 , n62704 , n13321 , n62706 , n62707 , 
     n62708 , n62709 , n13326 , n13327 , n62712 , n13329 , n62714 , n62715 , n62716 , n13333 , 
     n13334 , n13335 , n62720 , n13337 , n62722 , n13339 , n13340 , n62725 , n13342 , n62727 , 
     n62728 , n62729 , n62730 , n62731 , n13348 , n13349 , n62734 , n62735 , n13352 , n13353 , 
     n13354 , n62739 , n62740 , n13357 , n62742 , n13359 , n62744 , n13361 , n62746 , n62747 , 
     n13364 , n13365 , n62750 , n13367 , n13368 , n62753 , n62754 , n13371 , n62756 , n62757 , 
     n13374 , n13375 , n62760 , n62761 , n13378 , n62763 , n62764 , n62765 , n62766 , n62767 , 
     n13384 , n62769 , n13386 , n62771 , n62772 , n13389 , n13390 , n62775 , n13392 , n62777 , 
     n62778 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , 
     n62788 , n13405 , n62790 , n13407 , n62792 , n13409 , n13410 , n62795 , n13412 , n62797 , 
     n62798 , n62799 , n13416 , n62801 , n62802 , n13419 , n62804 , n13421 , n62806 , n62807 , 
     n13424 , n62809 , n13426 , n62811 , n62812 , n62813 , n62814 , n13431 , n62816 , n62817 , 
     n13434 , n62819 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , 
     n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n62835 , n13452 , n13453 , 
     n62838 , n62839 , n62840 , n62841 , n13458 , n62843 , n13460 , n62845 , n13462 , n13463 , 
     n13464 , n13465 , n13466 , n13467 , n62852 , n13469 , n62854 , n13471 , n13472 , n62857 , 
     n13474 , n13475 , n13476 , n13477 , n62862 , n13479 , n62864 , n13481 , n62866 , n62867 , 
     n13484 , n13485 , n62870 , n62871 , n13488 , n62873 , n62874 , n13491 , n62876 , n62877 , 
     n13494 , n13495 , n62880 , n13497 , n62882 , n13499 , n13500 , n13501 , n62886 , n13503 , 
     n62888 , n62889 , n13506 , n62891 , n13508 , n13509 , n13510 , n13511 , n62896 , n13513 , 
     n13514 , n13515 , n13516 , n62901 , n13518 , n62903 , n62904 , n62905 , n13522 , n62907 , 
     n62908 , n13525 , n62910 , n62911 , n13528 , n62913 , n13530 , n62915 , n13532 , n62917 , 
     n13534 , n62919 , n13536 , n62921 , n62922 , n62923 , n13540 , n62925 , n13542 , n13543 , 
     n62928 , n13545 , n13546 , n13547 , n13548 , n62933 , n13550 , n62935 , n62936 , n13553 , 
     n13554 , n62939 , n62940 , n13557 , n62942 , n62943 , n13560 , n62945 , n13562 , n13563 , 
     n13564 , n13565 , n62950 , n13567 , n62952 , n13569 , n13570 , n13571 , n13572 , n13573 , 
     n13574 , n13575 , n62960 , n13576 , n62962 , n13578 , n62964 , n13580 , n62966 , n13582 , 
     n13583 , n13584 , n13585 , n62971 , n62972 , n13588 , n62974 , n13590 , n62976 , n62977 , 
     n62978 , n13594 , n62980 , n62981 , n13597 , n13598 , n62984 , n13600 , n62986 , n13602 , 
     n62988 , n13604 , n62990 , n62991 , n13607 , n62993 , n62994 , n13610 , n13611 , n13612 , 
     n13613 , n13614 , n13615 , n63001 , n13617 , n13618 , n63004 , n13620 , n63006 , n13622 , 
     n63008 , n13624 , n63010 , n13626 , n13627 , n13628 , n13629 , n63015 , n13631 , n13632 , 
     n13633 , n13634 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , 
     n63028 , n63029 , n63030 , n13646 , n13647 , n13648 , n13649 , n63035 , n63036 , n63037 , 
     n13653 , n63039 , n63040 , n13656 , n13657 , n63043 , n63044 , n63045 , n13661 , n13662 , 
     n63048 , n13664 , n13665 , n63051 , n63052 , n63053 , n63054 , n13670 , n63056 , n63057 , 
     n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , 
     n63068 , n13684 , n63070 , n63071 , n13687 , n63073 , n63074 , n63075 , n63076 , n63077 , 
     n63078 , n13694 , n13695 , n63081 , n63082 , n63083 , n63084 , n13699 , n63086 , n63087 , 
     n13702 , n63089 , n13704 , n13705 , n13706 , n63093 , n63094 , n13709 , n63096 , n63097 , 
     n13712 , n63099 , n63100 , n13715 , n63102 , n63103 , n63104 , n63105 , n63106 , n13721 , 
     n63108 , n13723 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n13726 , 
     n63118 , n13728 , n63120 , n13730 , n13731 , n13732 , n13733 , n13734 , n63126 , n63127 , 
     n63128 , n63129 , n13739 , n63131 , n63132 , n63133 , n63134 , n63135 , n13745 , n63137 , 
     n13747 , n63139 , n63140 , n13750 , n63142 , n63143 , n13753 , n63145 , n63146 , n13756 , 
     n13757 , n63149 , n13759 , n13760 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , 
     n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , 
     n13777 , n63169 , n13779 , n13780 , n63172 , n63173 , n13783 , n13784 , n63176 , n63177 , 
     n13787 , n13788 , n13789 , n63181 , n63182 , n13792 , n13793 , n63185 , n63186 , n13796 , 
     n63188 , n63189 , n13799 , n63191 , n63192 , n13802 , n13803 , n63195 , n63196 , n63197 , 
     n63198 , n63199 , n13809 , n63201 , n63202 , n63203 , n63204 , n63205 , n13815 , n13816 , 
     n63208 , n63209 , n63210 , n13820 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , 
     n63218 , n63219 , n63220 , n13830 , n63222 , n63223 , n63224 , n13834 , n63226 , n13836 , 
     n13837 , n63229 , n63230 , n13840 , n13841 , n63233 , n63234 , n13844 , n63236 , n13846 , 
     n63238 , n63239 , n63240 , n63241 , n13851 , n13852 , n63244 , n13854 , n13855 , n13856 , 
     n63248 , n63249 , n63250 , n63251 , n13861 , n63253 , n63254 , n13864 , n63256 , n63257 , 
     n63258 , n63259 , n63260 , n13870 , n63262 , n63263 , n63264 , n13874 , n63266 , n63267 , 
     n13877 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n13884 , n63276 , n63277 , 
     n13887 , n63279 , n63280 , n13890 , n63282 , n63283 , n63284 , n63285 , n13895 , n63287 , 
     n63288 , n63289 , n63290 , n63291 , n63292 , n13902 , n63294 , n13904 , n13905 , n63297 , 
     n13907 , n63299 , n63300 , n13910 , n63302 , n13912 , n13913 , n13914 , n63306 , n13916 , 
     n13917 , n13918 , n63310 , n13920 , n13921 , n13922 , n63314 , n63315 , n63316 , n63317 , 
     n63318 , n63319 , n63320 , n13930 , n13931 , n13932 , n13933 , n63325 , n13935 , n63327 , 
     n13937 , n63329 , n13939 , n63331 , n13941 , n13942 , n63334 , n13944 , n63336 , n13946 , 
     n63338 , n63339 , n13949 , n63341 , n63342 , n13952 , n63344 , n13954 , n63346 , n63347 , 
     n63348 , n63349 , n63350 , n63351 , n63352 , n13959 , n63354 , n63355 , n13962 , n63357 , 
     n63358 , n63359 , n13966 , n63361 , n63362 , n63363 , n63364 , n13971 , n63366 , n63367 , 
     n63368 , n13975 , n13976 , n13977 , n63372 , n13979 , n63374 , n63375 , n13982 , n13983 , 
     n63378 , n13985 , n63380 , n13987 , n63382 , n63383 , n63384 , n63385 , n13992 , n63387 , 
     n63388 , n13995 , n63390 , n63391 , n63392 , n63393 , n14000 , n14001 , n63396 , n63397 , 
     n14004 , n63399 , n14006 , n14007 , n63402 , n14009 , n63404 , n14011 , n14012 , n63407 , 
     n63408 , n14015 , n63410 , n63411 , n14018 , n63413 , n63414 , n14021 , n63416 , n14023 , 
     n63418 , n14025 , n14026 , n14027 , n14028 , n63423 , n63424 , n63425 , n14032 , n63427 , 
     n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n14040 , n63435 , n14042 , n14043 , 
     n63438 , n14045 , n63440 , n14047 , n14048 , n14049 , n63444 , n14051 , n63446 , n14053 , 
     n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , 
     n14060 , n63459 , n14062 , n14063 , n63462 , n14065 , n63464 , n63465 , n14068 , n14069 , 
     n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , 
     n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , 
     n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , 
     n14072 , n63499 , n14074 , n14075 , n14076 , n14077 , n63504 , n63505 , n14080 , n63507 , 
     n14082 , n63509 , n63510 , n63511 , n14086 , n63513 , n63514 , n63515 , n14090 , n63517 , 
     n14092 , n63519 , n63520 , n14095 , n63522 , n63523 , n14098 , n14099 , n63526 , n14101 , 
     n63528 , n14103 , n63530 , n63531 , n14106 , n63533 , n63534 , n63535 , n63536 , n63537 , 
     n14112 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n14119 , n14120 , n63547 , 
     n14122 , n63549 , n63550 , n63551 , n63552 , n63553 , n14128 , n63555 , n63556 , n63557 , 
     n63558 , n63559 , n14134 , n63561 , n63562 , n14137 , n63564 , n63565 , n63566 , n63567 , 
     n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , 
     n14152 , n63579 , n14154 , n63581 , n63582 , n63583 , n14158 , n63585 , n63586 , n14161 , 
     n14162 , n14163 , n63590 , n63591 , n14166 , n14167 , n14168 , n14169 , n14170 , n63597 , 
     n14172 , n63599 , n63600 , n63601 , n14176 , n63603 , n14178 , n63605 , n14180 , n63607 , 
     n14182 , n14183 , n14184 , n63611 , n14186 , n63613 , n63614 , n14189 , n14190 , n14191 , 
     n14192 , n63619 , n63620 , n63621 , n14196 , n63623 , n63624 , n63625 , n63626 , n63627 , 
     n14202 , n14203 , n63630 , n63631 , n14206 , n63633 , n63634 , n63635 , n63636 , n14211 , 
     n63638 , n14213 , n63640 , n63641 , n14216 , n14217 , n63644 , n14219 , n63646 , n63647 , 
     n63648 , n63649 , n63650 , n14225 , n14226 , n63653 , n63654 , n63655 , n63656 , n63657 , 
     n63658 , n63659 , n63660 , n63661 , n63662 , n14237 , n63664 , n63665 , n14240 , n63667 , 
     n63668 , n63669 , n63670 , n14245 , n14246 , n14247 , n14248 , n14249 , n63676 , n14251 , 
     n63678 , n63679 , n63680 , n63681 , n14256 , n63683 , n63684 , n14259 , n63686 , n63687 , 
     n14262 , n14263 , n14264 , n14265 , n63692 , n14267 , n63694 , n63695 , n14270 , n63697 , 
     n63698 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n63705 , n63706 , n14281 , 
     n63708 , n14283 , n14284 , n63711 , n14286 , n14287 , n14288 , n14289 , n63716 , n63717 , 
     n63718 , n14293 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , 
     n14302 , n63729 , n14304 , n14305 , n14306 , n63733 , n63734 , n63735 , n14310 , n63737 , 
     n63738 , n63739 , n14314 , n63741 , n63742 , n63743 , n14318 , n63745 , n14319 , n14320 , 
     n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , 
     n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n14321 , 
     n63768 , n63769 , n14324 , n14325 , n63772 , n63773 , n63774 , n14329 , n14330 , n14331 , 
     n14332 , n63779 , n63780 , n63781 , n14336 , n63783 , n63784 , n63785 , n14340 , n63787 , 
     n63788 , n63789 , n14344 , n14345 , n63792 , n63793 , n14347 , n63795 , n14349 , n14350 , 
     n14351 , n14352 , n63800 , n14354 , n63802 , n63803 , n63804 , n63805 , n63806 , n14360 , 
     n14361 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , 
     n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , 
     n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , 
     n63838 , n63839 , n63840 , n14369 , n63842 , n14371 , n63844 , n63845 , n14374 , n63847 , 
     n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , 
     n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , 
     n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , 
     n63878 , n63879 , n63880 , n14394 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , 
     n63888 , n63889 , n63890 , n14399 , n14400 , n14401 , n14402 , n14403 , n63896 , n14405 , 
     n14406 , n14407 , n14408 , n63901 , n63902 , n63903 , n63904 , n63905 , n14414 , n63907 , 
     n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n14421 , n63917 , 
     n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n14432 , 
     n63928 , n63929 , n63930 , n63931 , n63932 , n14438 , n63934 , n63935 , n14441 , n63937 , 
     n63938 , n63939 , n14445 , n63941 , n63942 , n14448 , n63944 , n63945 , n63946 , n63947 , 
     n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n14457 , 
     n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n14462 , n63965 , n14464 , n14465 , 
     n63968 , n14467 , n14468 , n63971 , n63972 , n63973 , n14472 , n63975 , n63976 , n63977 , 
     n14476 , n63979 , n63980 , n63981 , n14480 , n63983 , n63984 , n63985 , n14484 , n14485 , 
     n63988 , n14487 , n14488 , n63991 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , 
     n63998 , n63999 , n64000 , n14496 , n14497 , n14498 , n64004 , n64005 , n14501 , n64007 , 
     n14503 , n14504 , n14505 , n64011 , n64012 , n64013 , n64014 , n14507 , n14508 , n14509 , 
     n14510 , n14511 , n14512 , n64021 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
     n14519 , n14520 , n14521 , n14522 , n14523 , n64033 , n14524 , n14525 , n14526 , n14527 , 
     n14528 , n64039 , n64040 , n64041 , n64042 , n14529 , n14530 , n14531 , n14532 , n14533 , 
     n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , 
     n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , 
     n14554 , n64069 , n64070 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n64077 , 
     n64078 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , 
     n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , 
     n14580 , n14581 , n14582 , n14583 , n14584 , n64103 , n64104 , n64105 , n14588 , n14589 , 
     n14590 , n14591 , n64110 , n14593 ;
buf ( n370  , n0 );
buf ( n371  , n1 );
buf ( n372  , n2 );
buf ( n373  , n3 );
buf ( n374  , n4 );
buf ( n375  , n5 );
buf ( n376  , n6 );
buf ( n377  , n7 );
buf ( n378  , n8 );
buf ( n379  , n9 );
buf ( n380  , n10 );
buf ( n381  , n11 );
buf ( n382  , n12 );
buf ( n383  , n13 );
buf ( n384  , n14 );
buf ( n385  , n15 );
buf ( n386  , n16 );
buf ( n387  , n17 );
buf ( n388  , n18 );
buf ( n389  , n19 );
buf ( n390  , n20 );
buf ( n391  , n21 );
buf ( n392  , n22 );
buf ( n393  , n23 );
buf ( n394  , n24 );
buf ( n395  , n25 );
buf ( n396  , n26 );
buf ( n397  , n27 );
buf ( n398  , n28 );
buf ( n399  , n29 );
buf ( n400  , n30 );
buf ( n401  , n31 );
buf ( n402  , n32 );
buf ( n403  , n33 );
buf ( n404  , n34 );
buf ( n405  , n35 );
buf ( n406  , n36 );
buf ( n407  , n37 );
buf ( n408  , n38 );
buf ( n409  , n39 );
buf ( n410  , n40 );
buf ( n411  , n41 );
buf ( n412  , n42 );
buf ( n413  , n43 );
buf ( n414  , n44 );
buf ( n415  , n45 );
buf ( n416  , n46 );
buf ( n417  , n47 );
buf ( n418  , n48 );
buf ( n419  , n49 );
buf ( n420  , n50 );
buf ( n421  , n51 );
buf ( n422  , n52 );
buf ( n423  , n53 );
buf ( n424  , n54 );
buf ( n425  , n55 );
buf ( n56 , n426 );
buf ( n57 , n427 );
buf ( n58 , n428 );
buf ( n59 , n429 );
buf ( n60 , n430 );
buf ( n61 , n431 );
buf ( n62 , n432 );
buf ( n63 , n433 );
buf ( n64 , n434 );
buf ( n65 , n435 );
buf ( n66 , n436 );
buf ( n67 , n437 );
buf ( n68 , n438 );
buf ( n69 , n439 );
buf ( n70 , n440 );
buf ( n71 , n441 );
buf ( n72 , n442 );
buf ( n73 , n443 );
buf ( n74 , n444 );
buf ( n75 , n445 );
buf ( n76 , n446 );
buf ( n77 , n447 );
buf ( n78 , n448 );
buf ( n79 , n449 );
buf ( n80 , n450 );
buf ( n81 , n451 );
buf ( n82 , n452 );
buf ( n83 , n453 );
buf ( n84 , n454 );
buf ( n85 , n455 );
buf ( n86 , n456 );
buf ( n87 , n457 );
buf ( n88 , n458 );
buf ( n89 , n459 );
buf ( n90 , n460 );
buf ( n91 , n461 );
buf ( n92 , n462 );
buf ( n93 , n463 );
buf ( n94 , n464 );
buf ( n95 , n465 );
buf ( n96 , n466 );
buf ( n97 , n467 );
buf ( n98 , n468 );
buf ( n99 , n469 );
buf ( n100 , n470 );
buf ( n101 , n471 );
buf ( n102 , n472 );
buf ( n103 , n473 );
buf ( n104 , n474 );
buf ( n105 , n475 );
buf ( n106 , n476 );
buf ( n107 , n477 );
buf ( n108 , n478 );
buf ( n109 , n479 );
buf ( n110 , n480 );
buf ( n111 , n481 );
buf ( n112 , n482 );
buf ( n113 , n483 );
buf ( n114 , n484 );
buf ( n115 , n485 );
buf ( n116 , n486 );
buf ( n117 , n487 );
buf ( n118 , n488 );
buf ( n119 , n489 );
buf ( n120 , n490 );
buf ( n121 , n491 );
buf ( n122 , n492 );
buf ( n123 , n493 );
buf ( n124 , n494 );
buf ( n125 , n495 );
buf ( n126 , n496 );
buf ( n127 , n497 );
buf ( n128 , n498 );
buf ( n129 , n499 );
buf ( n130 , n500 );
buf ( n131 , n501 );
buf ( n132 , n502 );
buf ( n133 , n503 );
buf ( n134 , n504 );
buf ( n135 , n505 );
buf ( n136 , n506 );
buf ( n137 , n507 );
buf ( n138 , n508 );
buf ( n139 , n509 );
buf ( n140 , n510 );
buf ( n141 , n511 );
buf ( n142 , n512 );
buf ( n143 , n513 );
buf ( n144 , n514 );
buf ( n145 , n515 );
buf ( n146 , n516 );
buf ( n147 , n517 );
buf ( n148 , n518 );
buf ( n149 , n519 );
buf ( n150 , n520 );
buf ( n151 , n521 );
buf ( n152 , n522 );
buf ( n153 , n523 );
buf ( n154 , n524 );
buf ( n155 , n525 );
buf ( n156 , n526 );
buf ( n157 , n527 );
buf ( n158 , n528 );
buf ( n159 , n529 );
buf ( n160 , n530 );
buf ( n161 , n531 );
buf ( n162 , n532 );
buf ( n163 , n533 );
buf ( n164 , n534 );
buf ( n165 , n535 );
buf ( n166 , n536 );
buf ( n167 , n537 );
buf ( n168 , n538 );
buf ( n169 , n539 );
buf ( n170 , n540 );
buf ( n171 , n541 );
buf ( n172 , n542 );
buf ( n173 , n543 );
buf ( n174 , n544 );
buf ( n175 , n545 );
buf ( n176 , n546 );
buf ( n177 , n547 );
buf ( n178 , n548 );
buf ( n179 , n549 );
buf ( n180 , n550 );
buf ( n181 , n551 );
buf ( n182 , n552 );
buf ( n183 , n553 );
buf ( n184 , n554 );
buf ( n426 , 1'b0 );
buf ( n427 , 1'b0 );
buf ( n428 , 1'b0 );
buf ( n429 , 1'b0 );
buf ( n430 , 1'b0 );
buf ( n431 , 1'b0 );
buf ( n432 , 1'b0 );
buf ( n433 , 1'b0 );
buf ( n434 , 1'b0 );
buf ( n435 , 1'b0 );
buf ( n436 , 1'b0 );
buf ( n437 , 1'b0 );
buf ( n438 , 1'b0 );
buf ( n439 , 1'b0 );
buf ( n440 , 1'b0 );
buf ( n441 , 1'b0 );
buf ( n442 , 1'b0 );
buf ( n443 , 1'b0 );
buf ( n444 , 1'b0 );
buf ( n445 , 1'b0 );
buf ( n446 , 1'b0 );
buf ( n447 , 1'b0 );
buf ( n448 , 1'b0 );
buf ( n449 , 1'b0 );
buf ( n450 , 1'b0 );
buf ( n451 , 1'b0 );
buf ( n452 , 1'b0 );
buf ( n453 , 1'b0 );
buf ( n454 , 1'b0 );
buf ( n455 , 1'b0 );
buf ( n456 , 1'b0 );
buf ( n457 , 1'b0 );
buf ( n458 , 1'b0 );
buf ( n459 , 1'b0 );
buf ( n460 , 1'b0 );
buf ( n461 , 1'b0 );
buf ( n462 , 1'b0 );
buf ( n463 , 1'b0 );
buf ( n464 , 1'b0 );
buf ( n465 , 1'b0 );
buf ( n466 , 1'b0 );
buf ( n467 , 1'b0 );
buf ( n468 , 1'b0 );
buf ( n469 , 1'b0 );
buf ( n470 , 1'b0 );
buf ( n471 , 1'b0 );
buf ( n472 , 1'b0 );
buf ( n473 , 1'b0 );
buf ( n474 , 1'b0 );
buf ( n475 , 1'b0 );
buf ( n476 , 1'b0 );
buf ( n477 , 1'b0 );
buf ( n478 , 1'b0 );
buf ( n479 , 1'b0 );
buf ( n480 , 1'b0 );
buf ( n481 , 1'b0 );
buf ( n482 , 1'b0 );
buf ( n483 , 1'b0 );
buf ( n484 , 1'b0 );
buf ( n485 , 1'b0 );
buf ( n486 , 1'b0 );
buf ( n487 , 1'b0 );
buf ( n488 , 1'b0 );
buf ( n489 , 1'b0 );
buf ( n490 , n63535 );
buf ( n491 , n14484 );
buf ( n492 , n63423 );
buf ( n493 , n64005 );
buf ( n494 , n63470 );
buf ( n495 , n14546 );
buf ( n496 , n14526 );
buf ( n497 , n64040 );
buf ( n498 , n63557 );
buf ( n499 , n63581 );
buf ( n500 , n63733 );
buf ( n501 , n63733 );
buf ( n502 , n63733 );
buf ( n503 , n63733 );
buf ( n504 , n63733 );
buf ( n505 , n63733 );
buf ( n506 , n14448 );
buf ( n507 , n14448 );
buf ( n508 , n14448 );
buf ( n509 , n14448 );
buf ( n510 , n14448 );
buf ( n511 , n14448 );
buf ( n512 , n14448 );
buf ( n513 , n14448 );
buf ( n514 , n14448 );
buf ( n515 , n14448 );
buf ( n516 , n14448 );
buf ( n517 , n14448 );
buf ( n518 , n14448 );
buf ( n519 , n14448 );
buf ( n520 , n14448 );
buf ( n521 , n14448 );
buf ( n522 , n14448 );
buf ( n523 , n14448 );
buf ( n524 , n14448 );
buf ( n525 , n14448 );
buf ( n526 , n14448 );
buf ( n527 , n14448 );
buf ( n528 , n14448 );
buf ( n529 , n63619 );
buf ( n530 , n63973 );
buf ( n531 , n64021 );
buf ( n532 , n63640 );
buf ( n533 , n14561 );
buf ( n534 , n63999 );
buf ( n535 , n63716 );
buf ( n536 , n63692 );
buf ( n537 , n14584 );
buf ( n538 , n63764 );
buf ( n539 , n63779 );
buf ( n540 , n14361 );
buf ( n541 , n14593 );
buf ( n542 , n14556 );
buf ( n543 , n64110 );
buf ( n544 , n63836 );
buf ( n545 , n14578 );
buf ( n546 , n63870 );
buf ( n547 , n63884 );
buf ( n548 , n14538 );
buf ( n549 , n63909 );
buf ( n550 , n14574 );
buf ( n551 , n63932 );
buf ( n552 , n63917 );
buf ( n553 , n63920 );
buf ( n554 , n14567 );
and ( n49826 , n373 , n374 );
and ( n49827 , n373 , n49826 );
nand ( n49828 , n371 , n376 );
not ( n555 , n49828 );
and ( n556 , n370 , n377 );
xor ( n557 , n555 , n556 );
and ( n558 , n372 , n375 );
and ( n559 , n557 , n558 );
and ( n560 , n555 , n556 );
or ( n561 , n559 , n560 );
xor ( n562 , n49827 , n561 );
nand ( n563 , n372 , n374 );
not ( n564 , n563 );
and ( n565 , n371 , n375 );
xor ( n566 , n564 , n565 );
and ( n567 , n370 , n376 );
xor ( n568 , n566 , n567 );
xor ( n569 , n562 , n568 );
not ( n570 , n569 );
xor ( n571 , n373 , n49826 );
nand ( n572 , n373 , n375 );
not ( n573 , n572 );
nand ( n574 , n372 , n376 );
not ( n575 , n574 );
and ( n576 , n573 , n575 );
xor ( n577 , n571 , n576 );
xor ( n578 , n555 , n556 );
xor ( n579 , n578 , n558 );
and ( n580 , n577 , n579 );
and ( n581 , n571 , n576 );
or ( n582 , n580 , n581 );
not ( n583 , n582 );
nand ( n584 , n570 , n583 );
not ( n585 , n584 );
and ( n586 , n374 , n377 );
xor ( n587 , n375 , n586 );
and ( n588 , n375 , n376 );
nand ( n589 , n587 , n588 );
nand ( n590 , n376 , n377 );
not ( n591 , n590 );
nand ( n592 , n375 , n377 );
not ( n593 , n592 );
nand ( n594 , n591 , n593 );
and ( n595 , n589 , n594 );
and ( n596 , n375 , n586 );
nand ( n597 , n374 , n376 );
and ( n598 , n373 , n377 );
and ( n599 , n597 , n598 );
not ( n600 , n597 );
nand ( n601 , n373 , n377 );
and ( n602 , n600 , n601 );
or ( n603 , n599 , n602 );
nor ( n604 , n596 , n603 );
nor ( n605 , n595 , n604 );
nand ( n606 , n603 , n596 );
not ( n607 , n606 );
nor ( n608 , n605 , n607 );
nand ( n609 , n372 , n377 );
not ( n610 , n609 );
and ( n611 , n373 , n376 );
xor ( n612 , n610 , n611 );
and ( n613 , n374 , n375 );
not ( n614 , n374 );
nor ( n615 , n613 , n614 );
xor ( n616 , n612 , n615 );
and ( n617 , n373 , n376 , n374 , n377 );
nor ( n618 , n616 , n617 );
or ( n619 , n608 , n618 );
nand ( n620 , n617 , n616 );
nand ( n621 , n619 , n620 );
and ( n622 , n371 , n377 );
xor ( n623 , n573 , n575 );
xor ( n624 , n622 , n623 );
and ( n625 , n374 , n375 );
xor ( n626 , n624 , n625 );
not ( n627 , n626 );
xor ( n628 , n610 , n611 );
and ( n629 , n628 , n615 );
and ( n630 , n610 , n611 );
or ( n631 , n629 , n630 );
not ( n632 , n631 );
nand ( n633 , n627 , n632 );
and ( n634 , n621 , n633 );
nor ( n635 , n627 , n632 );
nor ( n636 , n634 , n635 );
xor ( n637 , n571 , n576 );
xor ( n638 , n637 , n579 );
xor ( n639 , n622 , n623 );
and ( n640 , n639 , n625 );
and ( n641 , n622 , n623 );
or ( n642 , n640 , n641 );
buf ( n643 , n642 );
nor ( n644 , n638 , n643 );
or ( n645 , n636 , n644 );
nand ( n646 , n638 , n642 );
nand ( n647 , n645 , n646 );
not ( n648 , n647 );
or ( n649 , n585 , n648 );
not ( n650 , n583 );
not ( n651 , n570 );
nand ( n652 , n650 , n651 );
nand ( n653 , n649 , n652 );
xor ( n654 , n49827 , n561 );
and ( n655 , n654 , n568 );
and ( n656 , n49827 , n561 );
or ( n657 , n655 , n656 );
buf ( n658 , n657 );
and ( n659 , n371 , n374 );
xor ( n660 , n564 , n565 );
and ( n661 , n660 , n567 );
and ( n662 , n564 , n565 );
or ( n663 , n661 , n662 );
xor ( n664 , n659 , n663 );
and ( n665 , n372 , n373 );
xor ( n666 , n372 , n665 );
and ( n667 , n370 , n375 );
xor ( n668 , n666 , n667 );
xor ( n669 , n664 , n668 );
buf ( n670 , n669 );
and ( n671 , n658 , n670 );
not ( n672 , n658 );
not ( n673 , n670 );
and ( n674 , n672 , n673 );
nor ( n675 , n671 , n674 );
and ( n676 , n653 , n675 );
not ( n677 , n653 );
not ( n678 , n675 );
and ( n679 , n677 , n678 );
nor ( n680 , n676 , n679 );
buf ( n681 , n680 );
buf ( n49956 , n681 );
not ( n683 , n618 );
nand ( n684 , n683 , n620 );
not ( n685 , n608 );
xor ( n686 , n684 , n685 );
not ( n687 , n686 );
buf ( n49962 , n687 );
nand ( n689 , n49956 , n49962 );
buf ( n49964 , n689 );
xor ( n691 , n659 , n663 );
and ( n692 , n691 , n668 );
and ( n693 , n659 , n663 );
or ( n694 , n692 , n693 );
not ( n695 , n694 );
and ( n696 , n371 , n373 );
and ( n697 , n370 , n374 );
xor ( n698 , n696 , n697 );
xor ( n699 , n372 , n665 );
and ( n700 , n699 , n667 );
and ( n701 , n372 , n665 );
or ( n702 , n700 , n701 );
xor ( n703 , n698 , n702 );
not ( n704 , n703 );
nand ( n705 , n695 , n704 );
not ( n706 , n705 );
not ( n707 , n647 );
not ( n708 , n669 );
not ( n709 , n657 );
and ( n710 , n708 , n709 );
nor ( n711 , n569 , n582 );
nor ( n712 , n710 , n711 );
not ( n713 , n712 );
or ( n714 , n707 , n713 );
and ( n715 , n708 , n709 );
nand ( n716 , n569 , n582 );
nor ( n717 , n715 , n716 );
nor ( n718 , n709 , n708 );
nor ( n719 , n717 , n718 );
nand ( n720 , n714 , n719 );
not ( n721 , n720 );
or ( n722 , n706 , n721 );
nand ( n723 , n694 , n703 );
buf ( n724 , n723 );
nand ( n725 , n722 , n724 );
xor ( n726 , n696 , n697 );
and ( n727 , n726 , n702 );
and ( n728 , n696 , n697 );
or ( n729 , n727 , n728 );
and ( n730 , n371 , n372 );
xor ( n731 , n371 , n730 );
and ( n732 , n370 , n373 );
xor ( n733 , n731 , n732 );
nand ( n734 , n729 , n733 );
or ( n735 , n729 , n733 );
nand ( n736 , n734 , n735 );
and ( n737 , n725 , n736 );
not ( n738 , n725 );
not ( n739 , n736 );
and ( n740 , n738 , n739 );
nor ( n741 , n737 , n740 );
not ( n742 , n741 );
or ( n743 , n587 , n588 );
nand ( n744 , n743 , n589 );
not ( n745 , n744 );
and ( n746 , n594 , n745 );
not ( n747 , n594 );
and ( n748 , n747 , n744 );
or ( n749 , n746 , n748 );
nand ( n750 , n742 , n749 );
xor ( n751 , n49964 , n750 );
nand ( n752 , n694 , n703 );
and ( n753 , n752 , n705 );
not ( n754 , n753 );
buf ( n755 , n720 );
not ( n756 , n755 );
not ( n757 , n756 );
or ( n758 , n754 , n757 );
not ( n759 , n753 );
nand ( n760 , n759 , n755 );
nand ( n761 , n758 , n760 );
buf ( n762 , n761 );
buf ( n50037 , n762 );
not ( n764 , n604 );
nand ( n765 , n764 , n606 );
not ( n766 , n765 );
nand ( n767 , n594 , n589 );
not ( n768 , n767 );
or ( n769 , n766 , n768 );
or ( n770 , n767 , n765 );
nand ( n771 , n769 , n770 );
buf ( n772 , n771 );
buf ( n50047 , n772 );
nand ( n774 , n50037 , n50047 );
buf ( n50049 , n774 );
and ( n776 , n751 , n50049 );
and ( n777 , n49964 , n750 );
or ( n778 , n776 , n777 );
nor ( n779 , n694 , n703 );
not ( n780 , n735 );
nor ( n781 , n779 , n780 );
not ( n782 , n781 );
xor ( n783 , n371 , n730 );
and ( n784 , n783 , n732 );
and ( n785 , n371 , n730 );
or ( n786 , n784 , n785 );
not ( n787 , n786 );
nand ( n788 , n370 , n372 );
nand ( n789 , n787 , n788 );
not ( n790 , n789 );
not ( n791 , n790 );
nand ( n792 , n791 , n370 );
nor ( n793 , n782 , n792 );
not ( n794 , n793 );
not ( n795 , n755 );
or ( n796 , n794 , n795 );
not ( n50071 , n792 );
or ( n798 , n752 , n780 );
not ( n50073 , n798 );
and ( n800 , n50071 , n50073 );
or ( n50075 , n734 , n790 );
not ( n50076 , n788 );
nand ( n803 , n50076 , n786 );
nand ( n804 , n50075 , n803 );
not ( n805 , n804 );
not ( n806 , n371 );
nand ( n807 , n805 , n806 );
and ( n808 , n807 , n370 );
nor ( n809 , n800 , n808 );
nand ( n810 , n796 , n809 );
buf ( n811 , n810 );
buf ( n50086 , n811 );
and ( n50087 , n590 , n376 );
buf ( n50088 , n50087 );
nand ( n50089 , n50086 , n50088 );
buf ( n50090 , n50089 );
buf ( n50091 , n50090 );
not ( n818 , n50091 );
not ( n50093 , n582 );
not ( n820 , n651 );
or ( n50095 , n50093 , n820 );
nand ( n50096 , n50095 , n584 );
buf ( n823 , n647 );
xnor ( n824 , n50096 , n823 );
buf ( n50099 , n824 );
not ( n826 , n50099 );
buf ( n50101 , n826 );
buf ( n50102 , n50101 );
not ( n829 , n50102 );
buf ( n50104 , n829 );
buf ( n50105 , n50104 );
not ( n832 , n50105 );
and ( n833 , n818 , n832 );
buf ( n50108 , n50090 );
buf ( n50109 , n50101 );
not ( n836 , n50109 );
buf ( n50111 , n836 );
buf ( n50112 , n50111 );
and ( n839 , n50108 , n50112 );
nor ( n840 , n833 , n839 );
buf ( n50115 , n840 );
buf ( n50116 , n824 );
not ( n843 , n635 );
nand ( n50118 , n843 , n633 );
not ( n845 , n50118 );
buf ( n50120 , n621 );
not ( n50121 , n50120 );
or ( n848 , n845 , n50121 );
or ( n50123 , n50118 , n50120 );
nand ( n850 , n848 , n50123 );
buf ( n50125 , n850 );
buf ( n852 , n50125 );
buf ( n50127 , n852 );
buf ( n50128 , n50127 );
nand ( n50129 , n50116 , n50128 );
buf ( n50130 , n50129 );
buf ( n50131 , n50130 );
not ( n858 , n50131 );
buf ( n50133 , n858 );
buf ( n50134 , n50133 );
not ( n861 , n50134 );
nand ( n862 , n735 , n789 );
nor ( n863 , n779 , n862 );
not ( n864 , n863 );
not ( n865 , n720 );
or ( n866 , n864 , n865 );
not ( n867 , n723 );
not ( n868 , n862 );
and ( n869 , n867 , n868 );
nor ( n870 , n869 , n804 );
nand ( n871 , n866 , n870 );
nand ( n872 , n806 , n370 );
and ( n50147 , n871 , n872 );
not ( n874 , n871 );
not ( n50149 , n872 );
and ( n50150 , n874 , n50149 );
nor ( n877 , n50147 , n50150 );
not ( n50152 , n877 );
buf ( n50153 , n50152 );
buf ( n50154 , n50087 );
nand ( n881 , n50153 , n50154 );
buf ( n50156 , n881 );
buf ( n50157 , n50156 );
not ( n884 , n50157 );
buf ( n50159 , n884 );
buf ( n50160 , n50159 );
not ( n50161 , n50160 );
or ( n50162 , n861 , n50161 );
not ( n889 , n50130 );
not ( n50164 , n50156 );
or ( n50165 , n889 , n50164 );
and ( n892 , n789 , n803 );
not ( n50167 , n781 );
not ( n50168 , n755 );
or ( n50169 , n50167 , n50168 );
and ( n896 , n798 , n734 );
nand ( n50171 , n50169 , n896 );
xor ( n50172 , n892 , n50171 );
and ( n899 , n590 , n593 );
not ( n50174 , n590 );
and ( n50175 , n50174 , n592 );
or ( n902 , n899 , n50175 );
and ( n50177 , n50172 , n902 );
nand ( n904 , n50165 , n50177 );
buf ( n50179 , n904 );
nand ( n906 , n50162 , n50179 );
buf ( n50181 , n906 );
xor ( n908 , n50115 , n50181 );
xor ( n909 , n778 , n908 );
buf ( n50184 , n909 );
nand ( n911 , n50156 , n50133 );
nand ( n912 , n50159 , n50130 );
nand ( n913 , n911 , n912 );
not ( n914 , n913 );
buf ( n50189 , n50172 );
buf ( n916 , n50189 );
buf ( n50191 , n916 );
nand ( n918 , n50191 , n902 );
not ( n919 , n918 );
not ( n50194 , n919 );
or ( n921 , n914 , n50194 );
nand ( n922 , n912 , n911 , n918 );
nand ( n923 , n921 , n922 );
buf ( n50198 , n923 );
xor ( n925 , n49964 , n750 );
xor ( n926 , n925 , n50049 );
buf ( n50201 , n926 );
nand ( n928 , n50198 , n50201 );
buf ( n50203 , n928 );
buf ( n50204 , n50203 );
not ( n50205 , n50204 );
buf ( n50206 , n811 );
buf ( n50207 , n377 );
nand ( n50208 , n50206 , n50207 );
buf ( n50209 , n50208 );
buf ( n50210 , n636 );
not ( n937 , n50210 );
xnor ( n938 , n638 , n642 );
nand ( n939 , n937 , n938 );
not ( n940 , n938 );
nand ( n941 , n940 , n50210 );
nand ( n942 , n939 , n941 );
buf ( n943 , n942 );
xor ( n944 , n50209 , n943 );
buf ( n50219 , n944 );
not ( n946 , n50219 );
buf ( n50221 , n946 );
buf ( n50222 , n50221 );
not ( n949 , n50222 );
buf ( n50224 , n50152 );
buf ( n50225 , n50224 );
buf ( n50226 , n50225 );
buf ( n50227 , n50226 );
buf ( n50228 , n942 );
not ( n955 , n50228 );
buf ( n50230 , n955 );
not ( n957 , n50230 );
buf ( n50232 , n957 );
buf ( n50233 , n687 );
and ( n960 , n50232 , n50233 );
buf ( n50235 , n960 );
buf ( n50236 , n50235 );
buf ( n50237 , n377 );
nand ( n964 , n50227 , n50236 , n50237 );
buf ( n50239 , n964 );
buf ( n50240 , n50239 );
not ( n967 , n50240 );
buf ( n50242 , n967 );
buf ( n50243 , n50242 );
not ( n970 , n50243 );
or ( n50245 , n949 , n970 );
buf ( n50246 , n944 );
not ( n50247 , n50246 );
buf ( n50248 , n50239 );
not ( n50249 , n50248 );
or ( n976 , n50247 , n50249 );
buf ( n50251 , n681 );
buf ( n50252 , n749 );
and ( n979 , n50251 , n50252 );
buf ( n980 , n979 );
buf ( n981 , n980 );
and ( n982 , n725 , n736 );
not ( n983 , n725 );
and ( n984 , n983 , n739 );
nor ( n50259 , n982 , n984 );
not ( n986 , n50259 );
and ( n50261 , n986 , n50087 );
buf ( n50262 , n50261 );
xor ( n50263 , n981 , n50262 );
buf ( n50264 , n762 );
buf ( n50265 , n902 );
and ( n992 , n50264 , n50265 );
buf ( n50267 , n992 );
buf ( n50268 , n50267 );
and ( n995 , n50263 , n50268 );
and ( n50270 , n981 , n50262 );
or ( n997 , n995 , n50270 );
buf ( n50272 , n997 );
buf ( n50273 , n50272 );
nand ( n1000 , n976 , n50273 );
buf ( n50275 , n1000 );
buf ( n50276 , n50275 );
nand ( n1003 , n50245 , n50276 );
buf ( n50278 , n1003 );
buf ( n50279 , n50278 );
not ( n1006 , n50279 );
or ( n50281 , n50205 , n1006 );
or ( n50282 , n923 , n926 );
buf ( n50283 , n50282 );
nand ( n1010 , n50281 , n50283 );
buf ( n1011 , n1010 );
buf ( n50286 , n1011 );
not ( n1013 , n941 );
not ( n1014 , n939 );
or ( n1015 , n1013 , n1014 );
nand ( n1016 , n1015 , n50127 );
not ( n1017 , n1016 );
buf ( n50292 , n1017 );
buf ( n50293 , n681 );
buf ( n50294 , n772 );
nand ( n1021 , n50293 , n50294 );
buf ( n50296 , n1021 );
buf ( n50297 , n50296 );
not ( n50298 , n50297 );
buf ( n50299 , n50298 );
buf ( n50300 , n50299 );
xor ( n1027 , n50292 , n50300 );
buf ( n50302 , n687 );
not ( n50303 , n50302 );
buf ( n50304 , n50101 );
nor ( n50305 , n50303 , n50304 );
buf ( n50306 , n50305 );
buf ( n50307 , n50306 );
and ( n1034 , n1027 , n50307 );
and ( n1035 , n50292 , n50300 );
or ( n1036 , n1034 , n1035 );
buf ( n50311 , n1036 );
not ( n1038 , n50311 );
and ( n1039 , n811 , n943 , n377 );
not ( n1040 , n1039 );
nand ( n1041 , n1038 , n1040 );
not ( n1042 , n1041 );
not ( n50317 , n902 );
nor ( n1044 , n50317 , n50259 );
buf ( n1045 , n1044 );
not ( n1046 , n753 );
not ( n50321 , n756 );
or ( n50322 , n1046 , n50321 );
nand ( n1049 , n50322 , n760 );
and ( n50324 , n749 , n1049 );
buf ( n50325 , n50324 );
xor ( n50326 , n1045 , n50325 );
buf ( n50327 , n50172 );
not ( n1054 , n50327 );
buf ( n50329 , n50087 );
not ( n50330 , n50329 );
buf ( n50331 , n50330 );
buf ( n50332 , n50331 );
nor ( n50333 , n1054 , n50332 );
buf ( n50334 , n50333 );
buf ( n50335 , n50334 );
and ( n50336 , n50326 , n50335 );
and ( n50337 , n1045 , n50325 );
or ( n1062 , n50336 , n50337 );
buf ( n50339 , n1062 );
not ( n50340 , n50339 );
or ( n1065 , n1042 , n50340 );
and ( n1066 , n50311 , n1039 );
not ( n1067 , n1066 );
nand ( n1068 , n1065 , n1067 );
not ( n1069 , n1068 );
buf ( n50346 , n772 );
not ( n50347 , n50346 );
buf ( n50348 , n50347 );
nor ( n50349 , n741 , n50348 );
not ( n50350 , n50349 );
not ( n1075 , n50350 );
not ( n1076 , n50230 );
buf ( n50353 , n1076 );
buf ( n50354 , n50101 );
not ( n50355 , n50354 );
buf ( n50356 , n50355 );
buf ( n50357 , n50356 );
nand ( n1082 , n50353 , n50357 );
buf ( n50359 , n1082 );
buf ( n50360 , n50359 );
not ( n1085 , n50360 );
buf ( n50362 , n681 );
buf ( n50363 , n50127 );
nand ( n50364 , n50362 , n50363 );
buf ( n50365 , n50364 );
buf ( n50366 , n50365 );
not ( n50367 , n50366 );
buf ( n50368 , n50367 );
buf ( n50369 , n50368 );
not ( n50370 , n50369 );
or ( n1095 , n1085 , n50370 );
buf ( n50372 , n50359 );
buf ( n50373 , n50368 );
or ( n50374 , n50372 , n50373 );
nand ( n1099 , n1095 , n50374 );
buf ( n1100 , n1099 );
not ( n50377 , n1100 );
or ( n1102 , n1075 , n50377 );
or ( n50379 , n1100 , n50350 );
nand ( n50380 , n1102 , n50379 );
buf ( n50381 , n50152 );
not ( n1106 , n50381 );
buf ( n1107 , n1106 );
buf ( n50384 , n1107 );
not ( n50385 , n50384 );
buf ( n50386 , n50385 );
buf ( n50387 , n50386 );
buf ( n50388 , n902 );
nand ( n1113 , n50387 , n50388 );
buf ( n50390 , n1113 );
not ( n1115 , n50390 );
buf ( n1116 , n1049 );
buf ( n50393 , n1116 );
buf ( n50394 , n687 );
and ( n50395 , n50393 , n50394 );
buf ( n50396 , n50395 );
not ( n50397 , n50396 );
or ( n50398 , n1115 , n50397 );
nand ( n1123 , n761 , n687 );
buf ( n1124 , n1123 );
buf ( n50401 , n50152 );
not ( n1126 , n50401 );
buf ( n50403 , n902 );
not ( n50404 , n50403 );
buf ( n50405 , n50404 );
buf ( n50406 , n50405 );
nor ( n50407 , n1126 , n50406 );
buf ( n50408 , n50407 );
buf ( n50409 , n50408 );
nand ( n50410 , n1124 , n50409 );
buf ( n50411 , n50410 );
nand ( n1136 , n50398 , n50411 );
buf ( n50413 , n50172 );
buf ( n50414 , n749 );
and ( n50415 , n50413 , n50414 );
buf ( n50416 , n50415 );
not ( n50417 , n50416 );
and ( n1142 , n1136 , n50417 );
not ( n50419 , n1136 );
and ( n50420 , n50419 , n50416 );
nor ( n1145 , n1142 , n50420 );
and ( n50422 , n50380 , n1145 );
not ( n50423 , n50380 );
not ( n1148 , n1145 );
and ( n50425 , n50423 , n1148 );
nor ( n50426 , n50422 , n50425 );
not ( n50427 , n50426 );
or ( n50428 , n1069 , n50427 );
or ( n50429 , n50426 , n1068 );
nand ( n1154 , n50428 , n50429 );
buf ( n50431 , n1154 );
xor ( n50432 , n50184 , n50286 );
xor ( n1157 , n50432 , n50431 );
buf ( n50434 , n1157 );
xor ( n50435 , n50184 , n50286 );
and ( n1160 , n50435 , n50431 );
and ( n50437 , n50184 , n50286 );
or ( n50438 , n1160 , n50437 );
buf ( n50439 , n50438 );
buf ( n50440 , n942 );
buf ( n50441 , n749 );
nand ( n1166 , n50440 , n50441 );
buf ( n50443 , n1166 );
buf ( n50444 , n50443 );
not ( n1169 , n50444 );
buf ( n1170 , n1169 );
buf ( n50447 , n1170 );
not ( n1172 , n50447 );
buf ( n50449 , n681 );
buf ( n50450 , n50087 );
nand ( n50451 , n50449 , n50450 );
buf ( n50452 , n50451 );
buf ( n50453 , n50452 );
not ( n50454 , n50453 );
buf ( n50455 , n50454 );
buf ( n50456 , n50455 );
not ( n50457 , n50456 );
or ( n50458 , n1172 , n50457 );
buf ( n50459 , n50443 );
not ( n50460 , n50459 );
buf ( n50461 , n50452 );
not ( n50462 , n50461 );
or ( n50463 , n50460 , n50462 );
not ( n50464 , n902 );
nor ( n50465 , n50464 , n50101 );
buf ( n50466 , n50465 );
nand ( n50467 , n50463 , n50466 );
buf ( n1177 , n50467 );
buf ( n1178 , n1177 );
nand ( n1179 , n50458 , n1178 );
buf ( n1180 , n1179 );
buf ( n50472 , n1180 );
not ( n1182 , n50472 );
buf ( n50474 , n1182 );
buf ( n50475 , n50474 );
not ( n50476 , n50127 );
not ( n1186 , n50476 );
nand ( n50478 , n50172 , n377 );
not ( n1188 , n50478 );
or ( n1189 , n1186 , n1188 );
or ( n50481 , n50478 , n50476 );
nand ( n1191 , n1189 , n50481 );
buf ( n50483 , n1191 );
or ( n1193 , n50475 , n50483 );
buf ( n50485 , n1193 );
buf ( n50486 , n50485 );
not ( n1196 , n50474 );
not ( n1197 , n1191 );
or ( n1198 , n1196 , n1197 );
buf ( n50490 , n50127 );
buf ( n50491 , n687 );
and ( n1201 , n50490 , n50491 );
buf ( n50493 , n1201 );
buf ( n50494 , n50493 );
buf ( n50495 , n681 );
not ( n1205 , n50495 );
buf ( n50497 , n50405 );
nor ( n1207 , n1205 , n50497 );
buf ( n50499 , n1207 );
buf ( n50500 , n50499 );
xor ( n1210 , n50494 , n50500 );
buf ( n1211 , n1116 );
buf ( n50503 , n50087 );
and ( n1213 , n1211 , n50503 );
buf ( n50505 , n1213 );
buf ( n50506 , n50505 );
xor ( n50507 , n1210 , n50506 );
buf ( n50508 , n50507 );
nand ( n1218 , n1198 , n50508 );
buf ( n50510 , n1218 );
nand ( n1220 , n50486 , n50510 );
buf ( n50512 , n1220 );
buf ( n50513 , n50512 );
buf ( n50514 , n50104 );
buf ( n1224 , n772 );
and ( n1225 , n50514 , n1224 );
buf ( n50517 , n1225 );
buf ( n50518 , n50517 );
buf ( n50519 , n50191 );
buf ( n50520 , n50127 );
buf ( n50521 , n377 );
and ( n1231 , n50519 , n50520 , n50521 );
buf ( n50523 , n1231 );
buf ( n50524 , n50523 );
xor ( n50525 , n50518 , n50524 );
and ( n1235 , n50386 , n377 );
and ( n50527 , n50235 , n1235 );
not ( n50528 , n50235 );
nand ( n50529 , n50226 , n377 );
and ( n1239 , n50528 , n50529 );
nor ( n50531 , n50527 , n1239 );
buf ( n50532 , n50531 );
xor ( n50533 , n50525 , n50532 );
buf ( n50534 , n50533 );
buf ( n50535 , n50534 );
xor ( n50536 , n50494 , n50500 );
and ( n1246 , n50536 , n50506 );
and ( n50538 , n50494 , n50500 );
or ( n50539 , n1246 , n50538 );
buf ( n50540 , n50539 );
buf ( n50541 , n50540 );
xor ( n50542 , n981 , n50262 );
xor ( n50543 , n50542 , n50268 );
buf ( n50544 , n50543 );
buf ( n50545 , n50544 );
xor ( n1255 , n50541 , n50545 );
not ( n1256 , n50259 );
nand ( n1257 , n1256 , n377 );
not ( n1258 , n1257 );
buf ( n50550 , n50127 );
buf ( n50551 , n772 );
nand ( n50552 , n50550 , n50551 );
buf ( n50553 , n50552 );
not ( n1263 , n50553 );
and ( n50555 , n1258 , n1263 );
not ( n50556 , n50555 );
buf ( n50557 , n50111 );
buf ( n50558 , n749 );
and ( n50559 , n50557 , n50558 );
buf ( n50560 , n50559 );
not ( n50561 , n50560 );
buf ( n50562 , n1076 );
buf ( n50563 , n772 );
and ( n1273 , n50562 , n50563 );
buf ( n50565 , n1273 );
not ( n1275 , n50565 );
nand ( n1276 , n50561 , n1275 );
not ( n50568 , n1276 );
or ( n1278 , n50556 , n50568 );
not ( n50570 , n1275 );
nand ( n1280 , n50570 , n50560 );
nand ( n1281 , n1278 , n1280 );
buf ( n50573 , n1281 );
xor ( n1283 , n1255 , n50573 );
buf ( n50575 , n1283 );
buf ( n50576 , n50575 );
xor ( n1286 , n50513 , n50535 );
xor ( n50578 , n1286 , n50576 );
buf ( n50579 , n50578 );
xor ( n1289 , n50513 , n50535 );
and ( n1290 , n1289 , n50576 );
and ( n1291 , n50513 , n50535 );
or ( n1292 , n1290 , n1291 );
buf ( n50584 , n1292 );
xor ( n1294 , n50565 , n50560 );
xor ( n1295 , n1294 , n50555 );
buf ( n50587 , n1295 );
nor ( n50588 , n50331 , n50101 );
not ( n50589 , n50588 );
not ( n1299 , n50405 );
nand ( n50591 , n1299 , n942 );
nand ( n1301 , n772 , n687 );
nand ( n1302 , n50591 , n1301 );
not ( n50594 , n1302 );
or ( n50595 , n50589 , n50594 );
nor ( n1305 , n50591 , n1301 );
not ( n50597 , n1305 );
nand ( n50598 , n50595 , n50597 );
not ( n50599 , n50553 );
not ( n1309 , n1258 );
or ( n50601 , n50599 , n1309 );
not ( n1311 , n50553 );
nand ( n50603 , n1311 , n1257 );
nand ( n50604 , n50601 , n50603 );
xor ( n1314 , n50598 , n50604 );
buf ( n50606 , n687 );
buf ( n50607 , n762 );
buf ( n50608 , n377 );
and ( n1318 , n50607 , n50608 );
buf ( n50610 , n1318 );
buf ( n50611 , n50610 );
and ( n1321 , n50606 , n50611 );
buf ( n50613 , n1321 );
and ( n50614 , n1314 , n50613 );
and ( n50615 , n50598 , n50604 );
or ( n1325 , n50614 , n50615 );
buf ( n50617 , n1325 );
buf ( n50618 , n50474 );
buf ( n50619 , n1191 );
xor ( n1329 , n50618 , n50619 );
buf ( n50621 , n50508 );
xor ( n50622 , n1329 , n50621 );
buf ( n50623 , n50622 );
buf ( n50624 , n50623 );
xor ( n50625 , n50587 , n50617 );
xor ( n50626 , n50625 , n50624 );
buf ( n50627 , n50626 );
xor ( n50628 , n50587 , n50617 );
and ( n1338 , n50628 , n50624 );
and ( n1339 , n50587 , n50617 );
or ( n50631 , n1338 , n1339 );
buf ( n50632 , n50631 );
xor ( n50633 , n50465 , n1170 );
xor ( n50634 , n50633 , n50455 );
buf ( n50635 , n50634 );
buf ( n50636 , n50127 );
buf ( n50637 , n749 );
and ( n50638 , n50636 , n50637 );
buf ( n50639 , n50638 );
buf ( n50640 , n50639 );
buf ( n50641 , n681 );
buf ( n50642 , n50641 );
buf ( n50643 , n377 );
nand ( n50644 , n50642 , n50643 );
buf ( n50645 , n50644 );
buf ( n50646 , n50645 );
buf ( n1356 , n687 );
buf ( n1357 , n749 );
nand ( n1358 , n1356 , n1357 );
buf ( n1359 , n1358 );
buf ( n1360 , n1359 );
nor ( n1361 , n50646 , n1360 );
buf ( n1362 , n1361 );
buf ( n1363 , n1362 );
xor ( n1364 , n50640 , n1363 );
xor ( n1365 , n50606 , n50611 );
buf ( n50657 , n1365 );
buf ( n1367 , n50657 );
and ( n1368 , n1364 , n1367 );
and ( n1369 , n50640 , n1363 );
or ( n1370 , n1368 , n1369 );
buf ( n1371 , n1370 );
buf ( n50663 , n1371 );
xor ( n1373 , n50598 , n50604 );
xor ( n50665 , n1373 , n50613 );
buf ( n50666 , n50665 );
xor ( n1376 , n50635 , n50663 );
xor ( n50668 , n1376 , n50666 );
buf ( n50669 , n50668 );
xor ( n1379 , n50635 , n50663 );
and ( n50671 , n1379 , n50666 );
and ( n1381 , n50635 , n50663 );
or ( n50673 , n50671 , n1381 );
buf ( n50674 , n50673 );
xor ( n1384 , n50292 , n50300 );
xor ( n50676 , n1384 , n50307 );
buf ( n50677 , n50676 );
buf ( n1387 , n50677 );
xor ( n50679 , n1045 , n50325 );
xor ( n1389 , n50679 , n50335 );
buf ( n50681 , n1389 );
buf ( n50682 , n50681 );
xor ( n50683 , n50518 , n50524 );
and ( n50684 , n50683 , n50532 );
and ( n1394 , n50518 , n50524 );
or ( n50686 , n50684 , n1394 );
buf ( n50687 , n50686 );
buf ( n50688 , n50687 );
xor ( n50689 , n1387 , n50682 );
xor ( n50690 , n50689 , n50688 );
buf ( n50691 , n50690 );
xor ( n50692 , n1387 , n50682 );
and ( n50693 , n50692 , n50688 );
and ( n1403 , n1387 , n50682 );
or ( n1404 , n50693 , n1403 );
buf ( n50696 , n1404 );
xor ( n50697 , n50541 , n50545 );
and ( n50698 , n50697 , n50573 );
and ( n1408 , n50541 , n50545 );
or ( n50700 , n50698 , n1408 );
buf ( n50701 , n50700 );
buf ( n50702 , n942 );
buf ( n50703 , n824 );
nand ( n50704 , n50702 , n50703 );
buf ( n50705 , n50704 );
buf ( n50706 , n50705 );
buf ( n1416 , n50365 );
nand ( n1417 , n50706 , n1416 );
buf ( n1418 , n1417 );
buf ( n50710 , n1418 );
not ( n1420 , n50710 );
buf ( n50712 , n50349 );
not ( n50713 , n50712 );
or ( n50714 , n1420 , n50713 );
not ( n1424 , n50705 );
nand ( n50716 , n1424 , n50368 );
buf ( n50717 , n50716 );
nand ( n50718 , n50714 , n50717 );
buf ( n50719 , n50718 );
buf ( n50720 , n50719 );
buf ( n50721 , n811 );
buf ( n1431 , n50356 );
buf ( n50723 , n50087 );
and ( n50724 , n50721 , n1431 , n50723 );
buf ( n50725 , n50724 );
buf ( n50726 , n50725 );
buf ( n50727 , n50408 );
not ( n1437 , n50727 );
buf ( n50729 , n50396 );
not ( n50730 , n50729 );
or ( n1440 , n1437 , n50730 );
buf ( n50732 , n50390 );
not ( n1442 , n50732 );
buf ( n50734 , n1123 );
not ( n50735 , n50734 );
or ( n50736 , n1442 , n50735 );
buf ( n50737 , n50416 );
nand ( n50738 , n50736 , n50737 );
buf ( n50739 , n50738 );
buf ( n50740 , n50739 );
nand ( n50741 , n1440 , n50740 );
buf ( n50742 , n50741 );
buf ( n50743 , n50742 );
xor ( n1453 , n50720 , n50726 );
xor ( n50745 , n1453 , n50743 );
buf ( n50746 , n50745 );
xor ( n50747 , n50720 , n50726 );
and ( n50748 , n50747 , n50743 );
and ( n50749 , n50720 , n50726 );
or ( n1459 , n50748 , n50749 );
buf ( n50751 , n1459 );
buf ( n50752 , n50191 );
not ( n50753 , n50752 );
buf ( n50754 , n50259 );
not ( n1464 , n50754 );
buf ( n50756 , n1464 );
buf ( n50757 , n50756 );
not ( n1467 , n50757 );
buf ( n50759 , n1467 );
buf ( n50760 , n50759 );
nor ( n1470 , n50753 , n50760 );
buf ( n50762 , n1470 );
buf ( n1472 , n50762 );
buf ( n1473 , n811 );
buf ( n50765 , n50356 );
and ( n50766 , n1473 , n50765 );
buf ( n50767 , n50766 );
buf ( n50768 , n50767 );
buf ( n50769 , n50191 );
buf ( n50770 , n762 );
nand ( n1480 , n50769 , n50770 );
buf ( n50772 , n1480 );
buf ( n50773 , n50772 );
not ( n1483 , n50773 );
buf ( n1484 , n1483 );
buf ( n50776 , n1484 );
xor ( n1486 , n50768 , n50776 );
buf ( n50778 , n50386 );
buf ( n1488 , n50778 );
buf ( n50780 , n1488 );
buf ( n50781 , n50780 );
buf ( n50782 , n50641 );
and ( n50783 , n50781 , n50782 );
buf ( n50784 , n50783 );
buf ( n50785 , n50784 );
and ( n50786 , n1486 , n50785 );
and ( n50787 , n50768 , n50776 );
or ( n1497 , n50786 , n50787 );
buf ( n50789 , n1497 );
buf ( n50790 , n50789 );
buf ( n50791 , n50191 );
buf ( n1501 , n811 );
buf ( n1502 , n50641 );
and ( n1503 , n1501 , n1502 );
buf ( n1504 , n1503 );
buf ( n50796 , n1504 );
xor ( n1506 , n50791 , n50796 );
buf ( n50798 , n50780 );
buf ( n50799 , n762 );
and ( n50800 , n50798 , n50799 );
buf ( n50801 , n50800 );
buf ( n50802 , n50801 );
xor ( n50803 , n1506 , n50802 );
buf ( n50804 , n50803 );
buf ( n50805 , n50804 );
xor ( n1515 , n1472 , n50790 );
xor ( n1516 , n1515 , n50805 );
buf ( n50808 , n1516 );
xor ( n1518 , n1472 , n50790 );
and ( n50810 , n1518 , n50805 );
and ( n50811 , n1472 , n50790 );
or ( n1521 , n50810 , n50811 );
buf ( n50813 , n1521 );
buf ( n50814 , n50127 );
buf ( n50815 , n50087 );
nand ( n50816 , n50814 , n50815 );
buf ( n50817 , n50816 );
buf ( n50818 , n50817 );
buf ( n1528 , n687 );
buf ( n1529 , n902 );
nand ( n1530 , n1528 , n1529 );
buf ( n1531 , n1530 );
buf ( n50823 , n1531 );
and ( n1533 , n50818 , n50823 );
buf ( n50825 , n772 );
buf ( n50826 , n749 );
and ( n1536 , n50825 , n50826 );
buf ( n50828 , n1536 );
buf ( n50829 , n50828 );
not ( n50830 , n50829 );
buf ( n50831 , n50830 );
buf ( n50832 , n50831 );
nor ( n50833 , n1533 , n50832 );
buf ( n50834 , n50833 );
buf ( n50835 , n50834 );
buf ( n50836 , n50817 );
buf ( n50837 , n1531 );
nor ( n50838 , n50836 , n50837 );
buf ( n50839 , n50838 );
buf ( n50840 , n50839 );
or ( n50841 , n50835 , n50840 );
buf ( n50842 , n50841 );
buf ( n1552 , n50842 );
buf ( n50844 , n1359 );
not ( n1554 , n50844 );
buf ( n1555 , n1554 );
buf ( n50847 , n1555 );
not ( n50848 , n50847 );
buf ( n50849 , n50645 );
not ( n1559 , n50849 );
or ( n50851 , n50848 , n1559 );
buf ( n50852 , n50645 );
buf ( n50853 , n1555 );
or ( n50854 , n50852 , n50853 );
nand ( n1564 , n50851 , n50854 );
buf ( n1565 , n1564 );
buf ( n50857 , n1565 );
buf ( n50858 , n50127 );
buf ( n50859 , n902 );
and ( n50860 , n50858 , n50859 );
buf ( n50861 , n50860 );
buf ( n50862 , n50861 );
buf ( n50863 , n943 );
buf ( n50864 , n50087 );
and ( n50865 , n50863 , n50864 );
buf ( n50866 , n50865 );
buf ( n50867 , n50866 );
xor ( n50868 , n50862 , n50867 );
buf ( n50869 , n50111 );
buf ( n50870 , n377 );
nand ( n1580 , n50869 , n50870 );
buf ( n50872 , n1580 );
buf ( n50873 , n50872 );
buf ( n50874 , n50348 );
nor ( n50875 , n50873 , n50874 );
buf ( n50876 , n50875 );
buf ( n50877 , n50876 );
xor ( n1587 , n50868 , n50877 );
buf ( n50879 , n1587 );
buf ( n50880 , n50879 );
xor ( n1590 , n1552 , n50857 );
xor ( n50882 , n1590 , n50880 );
buf ( n50883 , n50882 );
xor ( n50884 , n1552 , n50857 );
and ( n1594 , n50884 , n50880 );
and ( n50886 , n1552 , n50857 );
or ( n1596 , n1594 , n50886 );
buf ( n50888 , n1596 );
buf ( n50889 , n50191 );
buf ( n50890 , n50111 );
and ( n50891 , n50889 , n50890 );
buf ( n50892 , n50891 );
buf ( n50893 , n50892 );
nand ( n50894 , n50152 , n50127 );
not ( n1604 , n50894 );
not ( n50896 , n1604 );
nand ( n1606 , n681 , n1116 );
not ( n50898 , n1606 );
not ( n50899 , n50898 );
or ( n1609 , n50896 , n50899 );
not ( n50901 , n1606 );
not ( n50902 , n50894 );
or ( n1612 , n50901 , n50902 );
and ( n1613 , n50172 , n943 );
nand ( n50905 , n1612 , n1613 );
nand ( n1615 , n1609 , n50905 );
buf ( n50907 , n1615 );
and ( n1617 , n742 , n50104 );
xor ( n50909 , n762 , n1617 );
buf ( n50910 , n811 );
buf ( n50911 , n687 );
and ( n1621 , n50910 , n50911 );
buf ( n50913 , n1621 );
and ( n50914 , n50909 , n50913 );
and ( n1624 , n762 , n1617 );
or ( n50916 , n50914 , n1624 );
buf ( n50917 , n50916 );
xor ( n1627 , n50893 , n50907 );
xor ( n50919 , n1627 , n50917 );
buf ( n50920 , n50919 );
xor ( n1630 , n50893 , n50907 );
and ( n50922 , n1630 , n50917 );
and ( n1632 , n50893 , n50907 );
or ( n1633 , n50922 , n1632 );
buf ( n50925 , n1633 );
buf ( n50926 , n50817 );
not ( n1636 , n50926 );
buf ( n50928 , n50828 );
not ( n1638 , n50928 );
buf ( n50930 , n1531 );
not ( n1640 , n50930 );
or ( n1641 , n1638 , n1640 );
buf ( n50933 , n1531 );
buf ( n50934 , n50828 );
or ( n1644 , n50933 , n50934 );
nand ( n50936 , n1641 , n1644 );
buf ( n50937 , n50936 );
buf ( n50938 , n50937 );
not ( n50939 , n50938 );
or ( n1649 , n1636 , n50939 );
buf ( n50941 , n50937 );
buf ( n50942 , n50817 );
or ( n50943 , n50941 , n50942 );
nand ( n1653 , n1649 , n50943 );
buf ( n50945 , n1653 );
buf ( n50946 , n50945 );
buf ( n50947 , n957 );
buf ( n1657 , n377 );
and ( n1658 , n50947 , n1657 );
buf ( n1659 , n1658 );
buf ( n50951 , n772 );
buf ( n50952 , n902 );
and ( n50953 , n50951 , n50952 );
buf ( n50954 , n50953 );
and ( n50955 , n1659 , n50954 );
buf ( n50956 , n50955 );
buf ( n50957 , n50872 );
buf ( n50958 , n50348 );
and ( n1668 , n50957 , n50958 );
not ( n1669 , n50957 );
buf ( n50961 , n772 );
and ( n50962 , n1669 , n50961 );
nor ( n50963 , n1668 , n50962 );
buf ( n50964 , n50963 );
buf ( n50965 , n50964 );
xor ( n1675 , n50946 , n50956 );
xor ( n50967 , n1675 , n50965 );
buf ( n50968 , n50967 );
xor ( n1678 , n50946 , n50956 );
and ( n50970 , n1678 , n50965 );
and ( n1680 , n50946 , n50956 );
or ( n50972 , n50970 , n1680 );
buf ( n50973 , n50972 );
buf ( n50974 , n50386 );
buf ( n50975 , n50356 );
and ( n50976 , n50974 , n50975 );
buf ( n50977 , n50976 );
buf ( n50978 , n50977 );
buf ( n50979 , n50191 );
buf ( n50980 , n50641 );
and ( n50981 , n50979 , n50980 );
buf ( n50982 , n50981 );
buf ( n1692 , n50982 );
not ( n1693 , n741 );
nand ( n50985 , n50641 , n1693 );
buf ( n1695 , n50985 );
not ( n1696 , n1695 );
buf ( n1697 , n811 );
buf ( n1698 , n50127 );
nand ( n1699 , n1697 , n1698 );
buf ( n1700 , n1699 );
buf ( n1701 , n1700 );
not ( n1702 , n1701 );
or ( n1703 , n1696 , n1702 );
buf ( n50995 , n50386 );
not ( n50996 , n50995 );
buf ( n50997 , n50230 );
nor ( n50998 , n50996 , n50997 );
buf ( n50999 , n50998 );
buf ( n51000 , n50999 );
nand ( n51001 , n1703 , n51000 );
buf ( n51002 , n51001 );
buf ( n51003 , n51002 );
buf ( n51004 , n1700 );
not ( n51005 , n51004 );
buf ( n51006 , n50985 );
not ( n51007 , n51006 );
buf ( n51008 , n51007 );
buf ( n51009 , n51008 );
nand ( n51010 , n51005 , n51009 );
buf ( n51011 , n51010 );
buf ( n51012 , n51011 );
nand ( n51013 , n51003 , n51012 );
buf ( n51014 , n51013 );
buf ( n51015 , n51014 );
xor ( n51016 , n50978 , n1692 );
xor ( n1720 , n51016 , n51015 );
buf ( n51018 , n1720 );
xor ( n51019 , n50978 , n1692 );
and ( n51020 , n51019 , n51015 );
and ( n1724 , n50978 , n1692 );
or ( n51022 , n51020 , n1724 );
buf ( n51023 , n51022 );
xor ( n1727 , n50640 , n1363 );
xor ( n51025 , n1727 , n1367 );
buf ( n51026 , n51025 );
buf ( n51027 , n50386 );
buf ( n51028 , n687 );
and ( n51029 , n51027 , n51028 );
buf ( n51030 , n51029 );
buf ( n51031 , n51030 );
not ( n1735 , n51031 );
buf ( n51033 , n50191 );
buf ( n51034 , n50127 );
nand ( n1738 , n51033 , n51034 );
buf ( n51036 , n1738 );
buf ( n51037 , n51036 );
nand ( n51038 , n1735 , n51037 );
buf ( n51039 , n51038 );
buf ( n51040 , n51039 );
nand ( n51041 , n50386 , n772 );
not ( n1745 , n51041 );
buf ( n51043 , n762 );
buf ( n51044 , n957 );
and ( n51045 , n51043 , n51044 );
buf ( n51046 , n51045 );
not ( n51047 , n51046 );
not ( n51048 , n51047 );
or ( n51049 , n1745 , n51048 );
buf ( n51050 , n50172 );
buf ( n51051 , n687 );
and ( n51052 , n51050 , n51051 );
buf ( n51053 , n51052 );
nand ( n1754 , n51049 , n51053 );
not ( n51055 , n51047 );
not ( n51056 , n51041 );
nand ( n51057 , n51055 , n51056 );
nand ( n1758 , n1754 , n51057 );
buf ( n51059 , n1758 );
buf ( n51060 , n51036 );
not ( n1761 , n51060 );
buf ( n51062 , n51030 );
nand ( n51063 , n1761 , n51062 );
buf ( n51064 , n51063 );
buf ( n51065 , n51064 );
not ( n51066 , n51040 );
not ( n51067 , n51059 );
or ( n1768 , n51066 , n51067 );
nand ( n1769 , n1768 , n51065 );
buf ( n51070 , n1769 );
xor ( n51071 , n50768 , n50776 );
xor ( n51072 , n51071 , n50785 );
buf ( n51073 , n51072 );
xor ( n1774 , n50791 , n50796 );
and ( n51075 , n1774 , n50802 );
and ( n51076 , n50791 , n50796 );
or ( n1777 , n51075 , n51076 );
buf ( n51078 , n1777 );
xor ( n51079 , n50862 , n50867 );
and ( n1780 , n51079 , n50877 );
and ( n1781 , n50862 , n50867 );
or ( n1782 , n1780 , n1781 );
buf ( n51083 , n1782 );
not ( n51084 , n681 );
nor ( n1785 , n51084 , n50230 );
buf ( n51086 , n1785 );
nand ( n51087 , n742 , n687 );
buf ( n1788 , n51087 );
not ( n51089 , n1788 );
buf ( n51090 , n51089 );
buf ( n51091 , n51090 );
buf ( n51092 , n811 );
not ( n1793 , n51092 );
buf ( n51094 , n50405 );
nor ( n1795 , n1793 , n51094 );
buf ( n51096 , n1795 );
buf ( n51097 , n51096 );
xor ( n1798 , n51086 , n51091 );
xor ( n1799 , n1798 , n51097 );
buf ( n51100 , n1799 );
xor ( n1801 , n51086 , n51091 );
and ( n51102 , n1801 , n51097 );
and ( n51103 , n51086 , n51091 );
or ( n1804 , n51102 , n51103 );
buf ( n51105 , n1804 );
buf ( n51106 , n50641 );
and ( n1807 , n986 , n50127 );
buf ( n51108 , n1807 );
buf ( n51109 , n811 );
buf ( n51110 , n749 );
and ( n51111 , n51109 , n51110 );
buf ( n51112 , n51111 );
buf ( n51113 , n51112 );
xor ( n51114 , n51106 , n51108 );
xor ( n51115 , n51114 , n51113 );
buf ( n51116 , n51115 );
xor ( n51117 , n51106 , n51108 );
and ( n1818 , n51117 , n51113 );
and ( n51119 , n51106 , n51108 );
or ( n51120 , n1818 , n51119 );
buf ( n51121 , n51120 );
buf ( n51122 , n749 );
buf ( n51123 , n749 );
buf ( n51124 , n902 );
nand ( n51125 , n51123 , n51124 );
buf ( n51126 , n51125 );
buf ( n51127 , n51126 );
buf ( n51128 , n50127 );
buf ( n51129 , n377 );
nand ( n51130 , n51128 , n51129 );
buf ( n51131 , n51130 );
buf ( n51132 , n51131 );
xor ( n1833 , n51122 , n51127 );
xor ( n51134 , n1833 , n51132 );
buf ( n51135 , n51134 );
buf ( n51136 , n944 );
buf ( n51137 , n50221 );
buf ( n51138 , n50242 );
and ( n1839 , n51138 , n51137 );
not ( n51140 , n51138 );
and ( n1840 , n51140 , n51136 );
nor ( n51142 , n1839 , n1840 );
buf ( n51143 , n51142 );
buf ( n51144 , n50759 );
not ( n1844 , n51144 );
buf ( n51146 , n1844 );
buf ( n51147 , n51146 );
buf ( n51148 , n811 );
buf ( n51149 , n1076 );
nand ( n51150 , n51148 , n51149 );
buf ( n51151 , n51150 );
buf ( n51152 , n51151 );
not ( n1852 , n51152 );
buf ( n51154 , n1852 );
buf ( n51155 , n51154 );
buf ( n1855 , n762 );
buf ( n51157 , n50756 );
and ( n51158 , n1855 , n51157 );
buf ( n51159 , n51158 );
buf ( n51160 , n51159 );
not ( n51161 , n51160 );
buf ( n51162 , n51161 );
buf ( n51163 , n51162 );
not ( n51164 , n51147 );
not ( n51165 , n51155 );
or ( n51166 , n51164 , n51165 );
nand ( n1866 , n51166 , n51163 );
buf ( n1867 , n1866 );
buf ( n1868 , n404 );
buf ( n51170 , n749 );
buf ( n51171 , n377 );
and ( n51172 , n51170 , n51171 );
buf ( n51173 , n51172 );
buf ( n51174 , n51173 );
xor ( n51175 , n1868 , n51174 );
buf ( n51176 , n51175 );
and ( n51177 , n1868 , n51174 );
buf ( n51178 , n51177 );
buf ( n51179 , n402 );
buf ( n51180 , n687 );
buf ( n51181 , n377 );
and ( n1881 , n51180 , n51181 );
buf ( n51183 , n1881 );
buf ( n51184 , n51183 );
xor ( n51185 , n51179 , n51184 );
buf ( n51186 , n51185 );
and ( n51187 , n51179 , n51184 );
buf ( n51188 , n51187 );
buf ( n51189 , n403 );
buf ( n51190 , n902 );
xor ( n51191 , n51189 , n51190 );
buf ( n51192 , n51191 );
and ( n1892 , n51189 , n51190 );
buf ( n51194 , n1892 );
buf ( n51195 , n405 );
buf ( n51196 , n50087 );
xor ( n51197 , n51195 , n51196 );
buf ( n51198 , n51197 );
and ( n1898 , n51195 , n51196 );
buf ( n51200 , n1898 );
buf ( n51201 , n51131 );
not ( n1901 , n51201 );
buf ( n51203 , n1901 );
buf ( n51204 , n50780 );
buf ( n1904 , n51204 );
buf ( n51206 , n1904 );
buf ( n51207 , n51206 );
buf ( n1907 , n811 );
buf ( n51209 , n1907 );
and ( n1909 , n51207 , n51209 );
buf ( n51211 , n1909 );
buf ( n51212 , n50191 );
buf ( n51213 , n1907 );
and ( n1913 , n51212 , n51213 );
buf ( n51215 , n1913 );
buf ( n51216 , n51146 );
buf ( n51217 , n1907 );
nand ( n51218 , n51216 , n51217 );
buf ( n51219 , n51218 );
buf ( n51220 , n50152 );
buf ( n51221 , n749 );
and ( n1921 , n51220 , n51221 );
buf ( n1922 , n1921 );
buf ( n51224 , n772 );
buf ( n51225 , n377 );
and ( n51226 , n51224 , n51225 );
buf ( n51227 , n51226 );
buf ( n51228 , n772 );
buf ( n51229 , n50087 );
and ( n51230 , n51228 , n51229 );
buf ( n51231 , n51230 );
buf ( n51232 , n50191 );
buf ( n51233 , n51206 );
nand ( n1933 , n51232 , n51233 );
buf ( n51235 , n1933 );
buf ( n51236 , n1049 );
buf ( n51237 , n50127 );
and ( n1937 , n51236 , n51237 );
buf ( n51239 , n1937 );
buf ( n51240 , n50641 );
buf ( n51241 , n50111 );
and ( n1941 , n51240 , n51241 );
buf ( n51243 , n1941 );
buf ( n51244 , n749 );
buf ( n51245 , n50087 );
and ( n51246 , n51244 , n51245 );
buf ( n51247 , n51246 );
buf ( n51248 , n50172 );
buf ( n51249 , n772 );
and ( n51250 , n51248 , n51249 );
buf ( n51251 , n51250 );
buf ( n51252 , n762 );
buf ( n51253 , n1907 );
and ( n51254 , n51252 , n51253 );
buf ( n51255 , n51254 );
not ( n1955 , n51255 );
not ( n1956 , n1955 );
buf ( n51258 , n50780 );
buf ( n51259 , n50756 );
and ( n1959 , n51258 , n51259 );
buf ( n51261 , n1959 );
not ( n1961 , n51261 );
and ( n1962 , n1956 , n1961 );
and ( n51264 , n1955 , n51261 );
nor ( n51265 , n1962 , n51264 );
not ( n51266 , n51078 );
xor ( n1966 , n51265 , n51266 );
or ( n51268 , n50813 , n1966 );
not ( n51269 , n51268 );
buf ( n51270 , n51269 );
not ( n51271 , n51270 );
nand ( n1971 , n1966 , n50813 );
buf ( n51273 , n1971 );
nand ( n51274 , n51271 , n51273 );
buf ( n51275 , n51274 );
buf ( n51276 , n51275 );
buf ( n51277 , n51275 );
not ( n51278 , n51277 );
buf ( n51279 , n51278 );
buf ( n51280 , n51279 );
buf ( n51281 , n50669 );
and ( n1981 , n1305 , n50588 );
not ( n1982 , n1302 );
and ( n51284 , n1982 , n50588 );
nor ( n1983 , n1981 , n51284 );
not ( n51286 , n50588 );
not ( n1985 , n50591 );
and ( n51288 , n51286 , n1985 , n1301 );
nor ( n1987 , n50588 , n1985 , n1301 );
nor ( n1988 , n51288 , n1987 );
nand ( n51291 , n1983 , n1988 );
xor ( n51292 , n51291 , n51083 );
and ( n1991 , n51292 , n51026 );
and ( n1992 , n51291 , n51083 );
or ( n51295 , n1991 , n1992 );
buf ( n51296 , n51295 );
nor ( n1995 , n51281 , n51296 );
buf ( n51298 , n1995 );
xor ( n1997 , n51291 , n51083 );
xor ( n51300 , n1997 , n51026 );
buf ( n51301 , n51300 );
buf ( n51302 , n50888 );
nand ( n51303 , n51301 , n51302 );
buf ( n51304 , n51303 );
or ( n2003 , n51298 , n51304 );
buf ( n51306 , n50669 );
buf ( n51307 , n51295 );
nand ( n2006 , n51306 , n51307 );
buf ( n51309 , n2006 );
nand ( n2008 , n2003 , n51309 );
not ( n51311 , n2008 );
not ( n2010 , n50674 );
not ( n2011 , n2010 );
not ( n51314 , n50627 );
not ( n51315 , n51314 );
or ( n2014 , n2011 , n51315 );
not ( n2015 , n50579 );
not ( n51318 , n50632 );
nand ( n51319 , n2015 , n51318 );
nand ( n2018 , n2014 , n51319 );
not ( n51321 , n2018 );
not ( n51322 , n51321 );
or ( n2021 , n51311 , n51322 );
and ( n51324 , n50627 , n50674 );
not ( n2023 , n50579 );
nand ( n51326 , n2023 , n51318 );
and ( n2025 , n51324 , n51326 );
buf ( n51328 , n50579 );
buf ( n51329 , n50632 );
and ( n51330 , n51328 , n51329 );
buf ( n51331 , n51330 );
nor ( n2030 , n2025 , n51331 );
nand ( n51333 , n2021 , n2030 );
not ( n51334 , n51333 );
or ( n2033 , n51188 , n51231 );
not ( n2034 , n2033 );
not ( n51337 , n51135 );
or ( n51338 , n2034 , n51337 );
nand ( n2037 , n51188 , n51231 );
nand ( n2038 , n51338 , n2037 );
buf ( n51341 , n2038 );
not ( n51342 , n51341 );
and ( n51343 , n687 , n50087 );
xor ( n51344 , n51343 , n50954 );
xnor ( n2043 , n51344 , n1659 );
not ( n51346 , n749 );
not ( n51347 , n51203 );
or ( n51348 , n51346 , n51347 );
nand ( n51349 , n51348 , n51126 );
xnor ( n2048 , n2043 , n51349 );
buf ( n51351 , n2048 );
not ( n51352 , n51351 );
or ( n2051 , n51342 , n51352 );
buf ( n51354 , n2048 );
buf ( n51355 , n2038 );
or ( n51356 , n51354 , n51355 );
xor ( n51357 , n51188 , n51231 );
xor ( n2056 , n51357 , n51135 );
buf ( n51359 , n2056 );
not ( n51360 , n51194 );
not ( n2059 , n51247 );
nand ( n2060 , n51360 , n2059 );
not ( n51363 , n2060 );
not ( n51364 , n51186 );
or ( n2063 , n51363 , n51364 );
nand ( n2064 , n51247 , n51194 );
nand ( n51367 , n2063 , n2064 );
buf ( n51368 , n51367 );
nand ( n2067 , n51356 , n51359 , n51368 );
buf ( n51370 , n2067 );
buf ( n51371 , n51370 );
nand ( n51372 , n2051 , n51371 );
buf ( n51373 , n51372 );
not ( n51374 , n51373 );
buf ( n51375 , n50883 );
buf ( n51376 , n50973 );
nor ( n51377 , n51375 , n51376 );
buf ( n51378 , n51377 );
buf ( n51379 , n51378 );
buf ( n51380 , n50968 );
not ( n51381 , n51343 );
xnor ( n51382 , n50954 , n1659 );
not ( n51383 , n51382 );
not ( n2082 , n51383 );
or ( n51385 , n51381 , n2082 );
not ( n51386 , n51343 );
nand ( n51387 , n51386 , n51382 );
nand ( n51388 , n51387 , n51349 );
nand ( n51389 , n51385 , n51388 );
buf ( n51390 , n51389 );
nor ( n51391 , n51380 , n51390 );
buf ( n51392 , n51391 );
buf ( n51393 , n51392 );
nor ( n51394 , n51379 , n51393 );
buf ( n51395 , n51394 );
not ( n51396 , n51395 );
or ( n51397 , n51374 , n51396 );
buf ( n51398 , n51378 );
not ( n2097 , n51398 );
buf ( n51400 , n2097 );
and ( n2099 , n51400 , n50968 , n51389 );
and ( n2100 , n50883 , n50973 );
nor ( n51403 , n2099 , n2100 );
nand ( n2101 , n51397 , n51403 );
buf ( n51405 , n51300 );
buf ( n51406 , n50888 );
nor ( n51407 , n51405 , n51406 );
buf ( n51408 , n51407 );
nor ( n51409 , n51408 , n51298 );
nand ( n51410 , n2101 , n51321 , n51409 );
and ( n51411 , n51192 , n51227 );
buf ( n51412 , n51411 );
and ( n51413 , n51194 , n2059 );
not ( n2111 , n51194 );
and ( n51415 , n2111 , n51247 );
nor ( n51416 , n51413 , n51415 );
xnor ( n51417 , n51416 , n51186 );
buf ( n51418 , n51417 );
or ( n51419 , n51412 , n51418 );
buf ( n51420 , n51419 );
xor ( n2118 , n51192 , n51227 );
and ( n51422 , n51420 , n2118 , n51178 );
and ( n51423 , n51417 , n51411 );
nor ( n2121 , n51422 , n51423 );
not ( n2122 , n2121 );
buf ( n51426 , n902 );
buf ( n51427 , n51198 );
or ( n2125 , n51426 , n51427 );
buf ( n51429 , n51176 );
buf ( n51430 , n51200 );
or ( n51431 , n51429 , n51430 );
buf ( n51432 , n51431 );
buf ( n51433 , n51432 );
nand ( n2130 , n2125 , n51433 );
buf ( n2131 , n2130 );
and ( n51436 , n406 , n407 , n408 );
nand ( n51437 , n51436 , n377 , n409 );
or ( n51438 , n2131 , n51437 );
buf ( n51439 , n51432 );
buf ( n51440 , n902 );
buf ( n51441 , n51198 );
and ( n2138 , n51439 , n51440 , n51441 );
buf ( n51443 , n51176 );
buf ( n51444 , n51200 );
and ( n2141 , n51443 , n51444 );
nor ( n51446 , n2138 , n2141 );
buf ( n51447 , n51446 );
nand ( n2144 , n51438 , n51447 );
not ( n2145 , n2144 );
or ( n51450 , n2118 , n51178 );
nand ( n2147 , n51450 , n51420 );
nor ( n2148 , n2145 , n2147 );
or ( n2149 , n2122 , n2148 );
or ( n2150 , n2038 , n2048 );
or ( n51455 , n2056 , n51367 );
nand ( n2152 , n2149 , n2150 , n51455 );
nor ( n2153 , n51392 , n51378 , n2152 );
nand ( n51458 , n51321 , n51409 , n2153 );
nand ( n51459 , n51334 , n51410 , n51458 );
buf ( n51460 , n51459 );
not ( n2157 , n51460 );
not ( n51462 , n50439 );
not ( n51463 , n51462 );
not ( n51464 , n1068 );
not ( n51465 , n50380 );
nand ( n2162 , n51465 , n1145 );
not ( n51467 , n2162 );
or ( n51468 , n51464 , n51467 );
buf ( n2165 , n50380 );
nand ( n51470 , n2165 , n1148 );
nand ( n51471 , n51468 , n51470 );
xor ( n2168 , n50746 , n51471 );
buf ( n51473 , n51239 );
xor ( n51474 , n1922 , n51473 );
xor ( n2171 , n51474 , n51251 );
and ( n51476 , n2171 , n51100 );
not ( n51477 , n2171 );
not ( n2174 , n51100 );
and ( n51479 , n51477 , n2174 );
nor ( n51480 , n51476 , n51479 );
buf ( n51481 , n50133 );
not ( n51482 , n51481 );
buf ( n51483 , n50159 );
not ( n2180 , n51483 );
or ( n51485 , n51482 , n2180 );
buf ( n51486 , n904 );
nand ( n2183 , n51485 , n51486 );
buf ( n51488 , n2183 );
not ( n51489 , n51488 );
not ( n2186 , n50115 );
not ( n51491 , n2186 );
or ( n51492 , n51489 , n51491 );
buf ( n51493 , n2186 );
buf ( n51494 , n50181 );
nor ( n2191 , n51493 , n51494 );
buf ( n51496 , n2191 );
or ( n51497 , n778 , n51496 );
nand ( n51498 , n51492 , n51497 );
and ( n51499 , n51480 , n51498 );
not ( n2196 , n51480 );
not ( n2197 , n51498 );
and ( n2198 , n2196 , n2197 );
nor ( n2199 , n51499 , n2198 );
xor ( n2200 , n2168 , n2199 );
buf ( n51505 , n2200 );
not ( n51506 , n51505 );
buf ( n51507 , n51506 );
not ( n51508 , n51507 );
or ( n2205 , n51463 , n51508 );
buf ( n2206 , n50434 );
not ( n51511 , n2206 );
buf ( n51512 , n51511 );
not ( n2209 , n1039 );
nand ( n51514 , n2209 , n50311 );
not ( n51515 , n51514 );
nand ( n51516 , n1038 , n1039 );
not ( n51517 , n51516 );
or ( n2214 , n51515 , n51517 );
not ( n51519 , n50339 );
nand ( n51520 , n2214 , n51519 );
nand ( n2217 , n50339 , n1066 );
not ( n2218 , n1041 );
nand ( n51523 , n50339 , n2218 );
nand ( n2220 , n51520 , n2217 , n51523 );
xor ( n2221 , n2220 , n50696 );
not ( n2222 , n50278 );
not ( n2223 , n926 );
and ( n51528 , n923 , n2223 );
not ( n51529 , n923 );
and ( n51530 , n51529 , n926 );
nor ( n2227 , n51528 , n51530 );
not ( n51532 , n2227 );
or ( n51533 , n2222 , n51532 );
or ( n2230 , n50278 , n2227 );
nand ( n51535 , n51533 , n2230 );
and ( n2232 , n2221 , n51535 );
and ( n2233 , n2220 , n50696 );
or ( n2234 , n2232 , n2233 );
buf ( n51539 , n2234 );
not ( n51540 , n51539 );
buf ( n51541 , n51540 );
nand ( n51542 , n51512 , n51541 );
nand ( n2239 , n2205 , n51542 );
buf ( n51544 , n2239 );
not ( n2241 , n51544 );
buf ( n2242 , n2241 );
buf ( n2243 , n2242 );
buf ( n51548 , n51143 );
buf ( n51549 , n50272 );
xor ( n51550 , n51548 , n51549 );
buf ( n51551 , n51550 );
not ( n51552 , n50701 );
and ( n2249 , n51551 , n51552 );
not ( n51554 , n51551 );
and ( n51555 , n51554 , n50701 );
or ( n2252 , n2249 , n51555 );
and ( n2253 , n2252 , n50691 );
not ( n2254 , n2252 );
not ( n2255 , n50691 );
and ( n51560 , n2254 , n2255 );
nor ( n2257 , n2253 , n51560 );
not ( n51562 , n2257 );
not ( n51563 , n50584 );
and ( n51564 , n51562 , n51563 );
xor ( n51565 , n2220 , n50696 );
xor ( n2262 , n51565 , n51535 );
not ( n51567 , n2262 );
not ( n51568 , n51551 );
nand ( n2265 , n51568 , n51552 );
not ( n51570 , n2265 );
not ( n2267 , n50691 );
or ( n51572 , n51570 , n2267 );
nand ( n51573 , n51551 , n50701 );
nand ( n51574 , n51572 , n51573 );
not ( n2271 , n51574 );
and ( n51576 , n51567 , n2271 );
nor ( n2273 , n51564 , n51576 );
buf ( n51578 , n2273 );
nand ( n51579 , n2243 , n51578 );
buf ( n51580 , n51579 );
not ( n2277 , n51580 );
buf ( n51582 , n51498 );
not ( n2279 , n51582 );
not ( n51584 , n2171 );
nand ( n51585 , n2174 , n51584 );
buf ( n2282 , n51585 );
not ( n51587 , n2282 );
or ( n51588 , n2279 , n51587 );
nand ( n2285 , n51100 , n2171 );
buf ( n51590 , n2285 );
nand ( n2287 , n51588 , n51590 );
buf ( n51592 , n2287 );
buf ( n2289 , n51105 );
buf ( n51594 , n1922 );
not ( n51595 , n51594 );
not ( n51596 , n51595 );
not ( n51597 , n51473 );
not ( n51598 , n51597 );
or ( n51599 , n51596 , n51598 );
nand ( n2293 , n51599 , n51251 );
nand ( n51601 , n51473 , n51594 );
nand ( n51602 , n2293 , n51601 );
nand ( n51603 , n51243 , n2289 , n51602 );
not ( n2297 , n51243 );
and ( n51605 , n51602 , n2297 );
not ( n51606 , n2289 );
nand ( n51607 , n51605 , n51606 );
not ( n2301 , n51602 );
nand ( n51609 , n51606 , n2301 , n51243 );
nand ( n51610 , n2301 , n2289 , n2297 );
nand ( n51611 , n51603 , n51607 , n51609 , n51610 );
xor ( n2305 , n51592 , n51611 );
not ( n51613 , n51046 );
not ( n51614 , n51041 );
or ( n51615 , n51613 , n51614 );
nand ( n2309 , n51047 , n51056 );
nand ( n51617 , n51615 , n2309 );
and ( n51618 , n51617 , n51053 );
not ( n51619 , n51617 );
not ( n51620 , n51053 );
and ( n2314 , n51619 , n51620 );
nor ( n2315 , n51618 , n2314 );
not ( n51623 , n2315 );
xor ( n51624 , n51116 , n51623 );
xnor ( n51625 , n51624 , n50751 );
xor ( n2319 , n2305 , n51625 );
not ( n2320 , n2319 );
xor ( n51628 , n50746 , n51471 );
and ( n2322 , n51628 , n2199 );
and ( n2323 , n50746 , n51471 );
or ( n2324 , n2322 , n2323 );
buf ( n51632 , n2324 );
not ( n2326 , n51632 );
buf ( n51634 , n2326 );
nand ( n2328 , n2320 , n51634 );
nand ( n2329 , n1116 , n50104 );
not ( n2330 , n2329 );
not ( n2331 , n2330 );
nand ( n2332 , n1693 , n942 );
not ( n2333 , n2332 );
not ( n2334 , n2333 );
or ( n2335 , n2331 , n2334 );
not ( n51643 , n2329 );
not ( n2337 , n2332 );
or ( n2338 , n51643 , n2337 );
nand ( n2339 , n811 , n772 );
not ( n2340 , n2339 );
nand ( n2341 , n2338 , n2340 );
nand ( n2342 , n2335 , n2341 );
xor ( n2343 , n762 , n1617 );
xor ( n2344 , n2343 , n50913 );
xor ( n2345 , n2342 , n2344 );
and ( n2346 , n50898 , n1604 );
not ( n2347 , n50898 );
and ( n2348 , n2347 , n50894 );
nor ( n2349 , n2346 , n2348 );
nand ( n2350 , n50191 , n943 );
not ( n2351 , n2350 );
and ( n2352 , n2349 , n2351 );
not ( n2353 , n2349 );
and ( n51661 , n2353 , n2350 );
nor ( n2355 , n2352 , n51661 );
xor ( n2356 , n2345 , n2355 );
xor ( n2357 , n51070 , n2356 );
not ( n2358 , n2333 );
not ( n2359 , n2330 );
not ( n2360 , n2340 );
or ( n2361 , n2359 , n2360 );
nand ( n2362 , n2339 , n2329 );
nand ( n2363 , n2361 , n2362 );
not ( n2364 , n2363 );
or ( n51672 , n2358 , n2364 );
or ( n2366 , n2333 , n2363 );
nand ( n51674 , n51672 , n2366 );
not ( n51675 , n51674 );
not ( n2369 , n51121 );
nand ( n2370 , n51675 , n2369 );
not ( n2371 , n2370 );
not ( n2372 , n51602 );
not ( n2373 , n51105 );
nand ( n2374 , n2373 , n2297 );
not ( n2375 , n2374 );
or ( n2376 , n2372 , n2375 );
nand ( n2377 , n2289 , n51243 );
nand ( n2378 , n2376 , n2377 );
not ( n2379 , n2378 );
or ( n2380 , n2371 , n2379 );
nand ( n2381 , n51121 , n51674 );
nand ( n2382 , n2380 , n2381 );
and ( n2383 , n2357 , n2382 );
and ( n2384 , n51070 , n2356 );
or ( n2385 , n2383 , n2384 );
xor ( n2386 , n51008 , n1700 );
xnor ( n2387 , n2386 , n50999 );
xor ( n2388 , n2387 , n50920 );
xor ( n2389 , n2342 , n2344 );
and ( n2390 , n2389 , n2355 );
and ( n2391 , n2342 , n2344 );
or ( n2392 , n2390 , n2391 );
xor ( n2393 , n2388 , n2392 );
or ( n2394 , n2385 , n2393 );
xor ( n2395 , n51030 , n51036 );
not ( n2396 , n1758 );
and ( n2397 , n2395 , n2396 );
not ( n2398 , n2395 );
and ( n2399 , n2398 , n1758 );
nor ( n2400 , n2397 , n2399 );
not ( n51708 , n51116 );
not ( n2402 , n2315 );
or ( n2403 , n51708 , n2402 );
not ( n2404 , n51116 );
not ( n2405 , n2404 );
not ( n2406 , n51623 );
or ( n2407 , n2405 , n2406 );
nand ( n2408 , n2407 , n50751 );
nand ( n2409 , n2403 , n2408 );
xor ( n2410 , n2400 , n2409 );
not ( n2411 , n51121 );
not ( n2412 , n51674 );
or ( n2413 , n2411 , n2412 );
nand ( n2414 , n51675 , n2369 );
nand ( n2415 , n2413 , n2414 );
not ( n51723 , n2378 );
and ( n2417 , n2415 , n51723 );
not ( n2418 , n2415 );
and ( n51726 , n2418 , n2378 );
nor ( n2420 , n2417 , n51726 );
and ( n2421 , n2410 , n2420 );
and ( n2422 , n2400 , n2409 );
or ( n2423 , n2421 , n2422 );
buf ( n51731 , n2423 );
not ( n2425 , n51731 );
buf ( n51733 , n2425 );
xor ( n51734 , n51070 , n2356 );
xor ( n2428 , n51734 , n2382 );
not ( n51736 , n2428 );
nand ( n51737 , n51733 , n51736 );
xor ( n2431 , n2400 , n2409 );
xor ( n51739 , n2431 , n2420 );
not ( n51740 , n51739 );
xor ( n51741 , n51592 , n51611 );
and ( n2435 , n51741 , n51625 );
and ( n51743 , n51592 , n51611 );
or ( n51744 , n2435 , n51743 );
not ( n51745 , n51744 );
nand ( n2439 , n51740 , n51745 );
nand ( n51747 , n2328 , n2394 , n51737 , n2439 );
not ( n51748 , n51747 );
nand ( n2442 , n2277 , n51748 );
not ( n51750 , n1867 );
not ( n2444 , n51073 );
or ( n2445 , n51750 , n2444 );
or ( n2446 , n51073 , n1867 );
nand ( n2447 , n2446 , n51023 );
nand ( n2448 , n2445 , n2447 );
nor ( n2449 , n50808 , n2448 );
buf ( n51757 , n2449 );
not ( n2451 , n51757 );
not ( n2452 , n2387 );
not ( n51760 , n2452 );
not ( n51761 , n50920 );
not ( n2455 , n51761 );
or ( n51763 , n51760 , n2455 );
nand ( n51764 , n51763 , n2392 );
not ( n2458 , n2452 );
nand ( n51766 , n2458 , n50920 );
nand ( n51767 , n51764 , n51766 );
buf ( n2461 , n51767 );
xor ( n51769 , n50756 , n51151 );
xor ( n51770 , n51769 , n51159 );
xor ( n2464 , n51770 , n51018 );
xnor ( n51772 , n2464 , n50925 );
buf ( n2466 , n51772 );
nor ( n2467 , n2461 , n2466 );
not ( n2468 , n51018 );
buf ( n2469 , n51770 );
nor ( n2470 , n2468 , n2469 );
not ( n2471 , n2470 );
xor ( n2472 , n1867 , n51023 );
xnor ( n2473 , n2472 , n51073 );
nand ( n2474 , n2468 , n2469 );
nand ( n51782 , n2474 , n50925 );
nand ( n2476 , n2471 , n2473 , n51782 );
not ( n2477 , n2476 );
nor ( n2478 , n2467 , n2477 );
buf ( n51786 , n2478 );
buf ( n2480 , n51786 );
buf ( n51788 , n2480 );
buf ( n51789 , n51788 );
nand ( n2483 , n2451 , n51789 );
buf ( n51791 , n2483 );
nor ( n51792 , n2442 , n51791 );
buf ( n51793 , n51792 );
not ( n51794 , n51793 );
or ( n2488 , n2157 , n51794 );
not ( n51796 , n2473 );
and ( n51797 , n2474 , n50925 );
nor ( n2491 , n51797 , n2470 );
not ( n51799 , n2491 );
nand ( n51800 , n51796 , n51799 );
nand ( n2494 , n51772 , n51767 );
not ( n51802 , n2494 );
nand ( n51803 , n51802 , n2476 );
nand ( n2497 , n51800 , n51803 );
buf ( n51805 , n2497 );
not ( n51806 , n51805 );
buf ( n51807 , n51806 );
buf ( n51808 , n51807 );
buf ( n51809 , n2449 );
or ( n2503 , n51808 , n51809 );
nand ( n51811 , n2448 , n50808 );
buf ( n51812 , n51811 );
nand ( n51813 , n2503 , n51812 );
buf ( n51814 , n51813 );
not ( n51815 , n51814 );
not ( n2509 , n51815 );
not ( n2510 , n51791 );
nor ( n51818 , n2385 , n2393 );
not ( n2512 , n51818 );
buf ( n51820 , n2428 );
buf ( n51821 , n2423 );
nand ( n51822 , n51820 , n51821 );
buf ( n51823 , n51822 );
not ( n51824 , n51823 );
and ( n51825 , n2512 , n51824 );
buf ( n51826 , n2385 );
buf ( n2520 , n51826 );
buf ( n2521 , n2520 );
buf ( n51829 , n2393 );
and ( n51830 , n2521 , n51829 );
nor ( n2524 , n51825 , n51830 );
not ( n51832 , n2524 );
not ( n51833 , n51832 );
not ( n51834 , n51818 );
nand ( n2528 , n51733 , n51736 );
nand ( n2529 , n51834 , n2528 );
nand ( n2530 , n51833 , n2529 );
nand ( n2531 , n2510 , n2530 );
not ( n51839 , n2531 );
or ( n2533 , n2509 , n51839 );
not ( n51841 , n51574 );
not ( n51842 , n2262 );
and ( n2536 , n51841 , n51842 );
buf ( n51844 , n2262 );
buf ( n51845 , n51574 );
nand ( n2539 , n51844 , n51845 );
buf ( n51847 , n2539 );
buf ( n51848 , n50584 );
buf ( n51849 , n2257 );
nand ( n51850 , n51848 , n51849 );
buf ( n51851 , n51850 );
and ( n51852 , n51847 , n51851 );
nor ( n51853 , n2536 , n51852 );
not ( n2547 , n51853 );
not ( n51855 , n2239 );
not ( n51856 , n51855 );
or ( n2550 , n2547 , n51856 );
buf ( n51858 , n50434 );
buf ( n2552 , n2234 );
and ( n2553 , n51858 , n2552 );
buf ( n2554 , n2553 );
not ( n51862 , n2200 );
nand ( n2556 , n51862 , n51462 );
and ( n51864 , n2554 , n2556 );
buf ( n2558 , n2200 );
buf ( n51866 , n50439 );
and ( n2560 , n2558 , n51866 );
buf ( n51868 , n2560 );
nor ( n2562 , n51864 , n51868 );
nand ( n2563 , n2550 , n2562 );
buf ( n2564 , n2563 );
not ( n2565 , n51739 );
nand ( n2566 , n2565 , n51745 );
and ( n51874 , n2566 , n2328 );
buf ( n51875 , n51874 );
nand ( n2569 , n2564 , n51875 );
buf ( n51877 , n51739 );
buf ( n51878 , n51744 );
nand ( n51879 , n51877 , n51878 );
buf ( n51880 , n51879 );
not ( n51881 , n51880 );
nand ( n2575 , n2324 , n2319 );
not ( n51883 , n2575 );
or ( n51884 , n51881 , n51883 );
nand ( n2578 , n51884 , n2566 );
not ( n51886 , n2578 );
nor ( n2580 , n51832 , n51886 );
nand ( n2581 , n2569 , n51815 , n2580 );
nand ( n2582 , n2533 , n2581 );
buf ( n51890 , n2582 );
nand ( n2584 , n2488 , n51890 );
buf ( n51892 , n2584 );
buf ( n51893 , n51892 );
and ( n2587 , n51893 , n51280 );
not ( n51895 , n51893 );
and ( n51896 , n51895 , n51276 );
nor ( n2590 , n2587 , n51896 );
buf ( n2591 , n2590 );
buf ( n51899 , n2528 );
buf ( n51900 , n51823 );
nand ( n51901 , n51899 , n51900 );
buf ( n51902 , n51901 );
buf ( n51903 , n51902 );
buf ( n51904 , n51902 );
not ( n51905 , n51904 );
buf ( n51906 , n51905 );
buf ( n51907 , n51906 );
not ( n51908 , n51886 );
not ( n2602 , n2008 );
not ( n2603 , n51321 );
or ( n51911 , n2602 , n2603 );
nand ( n51912 , n51911 , n2030 );
not ( n2606 , n51912 );
nand ( n51914 , n2606 , n51410 , n51458 );
buf ( n51915 , n51874 );
not ( n2609 , n51915 );
buf ( n2610 , n2242 );
buf ( n2611 , n2273 );
nand ( n2612 , n2610 , n2611 );
buf ( n2613 , n2612 );
buf ( n51921 , n2613 );
nor ( n51922 , n2609 , n51921 );
buf ( n51923 , n51922 );
nand ( n51924 , n51914 , n51923 );
nand ( n2618 , n2564 , n51875 );
nand ( n51926 , n51908 , n51924 , n2618 );
buf ( n51927 , n51926 );
and ( n2621 , n51927 , n51907 );
not ( n51929 , n51927 );
and ( n51930 , n51929 , n51903 );
nor ( n2624 , n2621 , n51930 );
buf ( n2625 , n2624 );
nand ( n51933 , n51803 , n51800 );
not ( n2627 , n51268 );
nor ( n51935 , n2627 , n2449 );
nand ( n2629 , n51933 , n51935 );
buf ( n51937 , n2629 );
not ( n51938 , n51937 );
buf ( n51939 , n51912 );
nor ( n51940 , n51938 , n51939 );
buf ( n51941 , n51940 );
buf ( n2635 , n51941 );
buf ( n2636 , n51410 );
buf ( n51944 , n51458 );
not ( n51945 , n51261 );
nand ( n51946 , n51945 , n1955 );
not ( n2640 , n51946 );
not ( n51948 , n51266 );
not ( n2642 , n51948 );
or ( n2643 , n2640 , n2642 );
nand ( n51951 , n51255 , n51261 );
nand ( n2645 , n2643 , n51951 );
buf ( n51953 , n2645 );
buf ( n51954 , n51235 );
not ( n51955 , n51219 );
xor ( n51956 , n51206 , n51955 );
xnor ( n2650 , n51954 , n51956 );
buf ( n51958 , n2650 );
nand ( n51959 , n51953 , n51958 );
buf ( n51960 , n51959 );
buf ( n51961 , n51960 );
not ( n51962 , n51961 );
or ( n2656 , n51269 , n51811 );
nand ( n2657 , n2656 , n1971 );
buf ( n51965 , n2657 );
nor ( n2659 , n51962 , n51965 );
buf ( n51967 , n2659 );
buf ( n51968 , n51967 );
nand ( n51969 , n2635 , n2636 , n51944 , n51968 );
buf ( n51970 , n51969 );
buf ( n51971 , n51459 );
not ( n2665 , n2442 );
buf ( n51973 , n2665 );
buf ( n51974 , n51788 );
nand ( n51975 , n51971 , n51973 , n51974 );
buf ( n51976 , n51975 );
not ( n51977 , n51748 );
not ( n2671 , n2563 );
or ( n2672 , n51977 , n2671 );
not ( n2673 , n2578 );
not ( n51981 , n2529 );
and ( n2675 , n2673 , n51981 );
nor ( n51983 , n2675 , n51832 );
nand ( n2677 , n2672 , n51983 );
buf ( n51985 , n2677 );
not ( n51986 , n51985 );
buf ( n51987 , n51986 );
buf ( n51988 , n2564 );
buf ( n2682 , n51874 );
buf ( n51990 , n2528 );
and ( n51991 , n2682 , n51990 );
buf ( n51992 , n51991 );
buf ( n51993 , n51992 );
buf ( n2687 , n2528 );
not ( n51995 , n2687 );
buf ( n51996 , n51995 );
or ( n2690 , n51996 , n2578 );
nand ( n51998 , n2690 , n51823 );
buf ( n51999 , n51998 );
and ( n52000 , n51988 , n51993 );
nor ( n52001 , n52000 , n51999 );
buf ( n52002 , n52001 );
not ( n52003 , n51219 );
nand ( n52004 , n52003 , n51206 );
not ( n2698 , n51215 );
and ( n52006 , n52004 , n51954 , n2698 );
nor ( n52007 , n51960 , n52006 );
nand ( n2701 , n52004 , n51954 );
buf ( n52009 , n2701 );
buf ( n2703 , n51215 );
nand ( n52011 , n52009 , n2703 );
buf ( n52012 , n52011 );
not ( n2706 , n52012 );
nor ( n52014 , n52007 , n2706 );
buf ( n52015 , n52014 );
not ( n2709 , n51811 );
nand ( n52017 , n2709 , n51268 );
nand ( n52018 , n52015 , n52017 , n1971 );
buf ( n52019 , n52018 );
buf ( n52020 , n51580 );
buf ( n52021 , n2629 );
not ( n52022 , n52019 );
nand ( n2716 , n52022 , n52020 , n52021 );
buf ( n2717 , n2716 );
buf ( n52025 , n2657 );
buf ( n52026 , n2629 );
not ( n52027 , n52025 );
nand ( n2721 , n52027 , n52026 );
buf ( n52029 , n2721 );
not ( n52030 , n52015 );
buf ( n52031 , n52030 );
buf ( n52032 , n1907 );
buf ( n52033 , n51211 );
and ( n52034 , n52031 , n52032 );
nor ( n2728 , n52034 , n52033 );
buf ( n52036 , n2728 );
buf ( n52037 , n2449 );
buf ( n52038 , n51811 );
not ( n52039 , n52037 );
nand ( n52040 , n52039 , n52038 );
buf ( n52041 , n52040 );
buf ( n52042 , n2645 );
buf ( n52043 , n2650 );
or ( n52044 , n52042 , n52043 );
buf ( n52045 , n52044 );
buf ( n52046 , n52045 );
not ( n52047 , n52046 );
buf ( n52048 , n52047 );
buf ( n52049 , n1971 );
buf ( n52050 , n51960 );
and ( n52051 , n52049 , n52050 );
buf ( n52052 , n52051 );
buf ( n52053 , n51992 );
buf ( n52054 , n2613 );
not ( n2748 , n52053 );
nor ( n2749 , n2748 , n52054 );
buf ( n52057 , n2749 );
buf ( n52058 , n51269 );
buf ( n52059 , n2449 );
or ( n52060 , n52058 , n52059 );
buf ( n52061 , n52060 );
buf ( n52062 , n409 );
buf ( n52063 , n415 );
and ( n52064 , n52062 , n52063 );
buf ( n52065 , n52064 );
buf ( n52066 , n52065 );
buf ( n52067 , n407 );
buf ( n52068 , n417 );
and ( n52069 , n52067 , n52068 );
buf ( n52070 , n52069 );
buf ( n52071 , n52070 );
buf ( n52072 , n408 );
buf ( n52073 , n416 );
and ( n52074 , n52072 , n52073 );
buf ( n52075 , n52074 );
buf ( n52076 , n52075 );
xor ( n52077 , n52066 , n52071 );
xor ( n52078 , n52077 , n52076 );
buf ( n52079 , n52078 );
xor ( n52080 , n52066 , n52071 );
and ( n52081 , n52080 , n52076 );
and ( n2775 , n52066 , n52071 );
or ( n52083 , n52081 , n2775 );
buf ( n52084 , n52083 );
buf ( n52085 , n391 );
buf ( n52086 , n393 );
and ( n52087 , n52085 , n52086 );
buf ( n52088 , n52087 );
buf ( n52089 , n52088 );
buf ( n52090 , n392 );
buf ( n52091 , n393 );
nand ( n2785 , n52090 , n52091 );
buf ( n52093 , n2785 );
buf ( n52094 , n52093 );
buf ( n52095 , n409 );
buf ( n52096 , n416 );
nand ( n52097 , n52095 , n52096 );
buf ( n52098 , n52097 );
buf ( n52099 , n52098 );
nor ( n52100 , n52094 , n52099 );
buf ( n52101 , n52100 );
buf ( n52102 , n52101 );
buf ( n52103 , 1'b0 );
xor ( n2797 , n52089 , n52102 );
xor ( n52105 , n2797 , n52103 );
buf ( n52106 , n52105 );
and ( n52107 , n52089 , n52102 );
or ( n52108 , 1'b0 , n52107 );
buf ( n52109 , n52108 );
xor ( n52110 , n52089 , n52102 );
buf ( n52111 , n408 );
buf ( n52112 , n415 );
and ( n2806 , n52111 , n52112 );
buf ( n52114 , n2806 );
buf ( n52115 , n52114 );
buf ( n52116 , n407 );
buf ( n52117 , n416 );
and ( n52118 , n52116 , n52117 );
buf ( n52119 , n52118 );
buf ( n52120 , n52119 );
buf ( n52121 , n406 );
buf ( n52122 , n417 );
and ( n2816 , n52121 , n52122 );
buf ( n52124 , n2816 );
buf ( n52125 , n52124 );
xor ( n52126 , n52115 , n52120 );
xor ( n2820 , n52126 , n52125 );
buf ( n52128 , n2820 );
xor ( n52129 , n52115 , n52120 );
and ( n2823 , n52129 , n52125 );
and ( n52131 , n52115 , n52120 );
or ( n52132 , n2823 , n52131 );
buf ( n52133 , n52132 );
nand ( n2827 , n393 , n391 );
not ( n52135 , n2827 );
nand ( n52136 , n393 , n392 );
not ( n2830 , n52136 );
or ( n2831 , n52135 , n2830 );
nand ( n52139 , n393 , n391 );
nand ( n52140 , n393 , n392 );
or ( n2834 , n52139 , n52140 );
nand ( n52142 , n2831 , n2834 );
not ( n2836 , n52142 );
buf ( n52144 , n2836 );
buf ( n52145 , n409 );
buf ( n52146 , n414 );
nand ( n2840 , n52145 , n52146 );
buf ( n2841 , n2840 );
buf ( n52149 , n2841 );
not ( n52150 , n52149 );
buf ( n52151 , n390 );
buf ( n52152 , n393 );
nand ( n2846 , n52151 , n52152 );
buf ( n52154 , n2846 );
buf ( n52155 , n52154 );
not ( n2849 , n52155 );
buf ( n2850 , n2849 );
buf ( n52158 , n2850 );
not ( n2852 , n52158 );
or ( n2853 , n52150 , n2852 );
buf ( n52161 , n2850 );
buf ( n52162 , n2841 );
or ( n52163 , n52161 , n52162 );
nand ( n2857 , n2853 , n52163 );
buf ( n52165 , n2857 );
buf ( n52166 , n52165 );
and ( n2860 , n52140 , n392 );
buf ( n52168 , n2860 );
xor ( n2862 , n52144 , n52166 );
xor ( n52170 , n2862 , n52168 );
buf ( n52171 , n52170 );
xor ( n2865 , n52144 , n52166 );
and ( n52173 , n2865 , n52168 );
and ( n52174 , n52144 , n52166 );
or ( n52175 , n52173 , n52174 );
buf ( n52176 , n52175 );
buf ( n52177 , n52084 );
buf ( n52178 , n52128 );
buf ( n52179 , n52109 );
xor ( n2873 , n52177 , n52178 );
xor ( n52181 , n2873 , n52179 );
buf ( n52182 , n52181 );
xor ( n52183 , n52177 , n52178 );
and ( n52184 , n52183 , n52179 );
and ( n52185 , n52177 , n52178 );
or ( n2879 , n52184 , n52185 );
buf ( n52187 , n2879 );
buf ( n52188 , n407 );
buf ( n52189 , n415 );
and ( n2883 , n52188 , n52189 );
buf ( n2884 , n2883 );
buf ( n52192 , n2884 );
buf ( n52193 , n409 );
buf ( n52194 , n413 );
and ( n2888 , n52193 , n52194 );
buf ( n2889 , n2888 );
buf ( n52197 , n2889 );
buf ( n52198 , n406 );
buf ( n52199 , n416 );
and ( n52200 , n52198 , n52199 );
buf ( n52201 , n52200 );
buf ( n52202 , n52201 );
xor ( n2896 , n52192 , n52197 );
xor ( n2897 , n2896 , n52202 );
buf ( n52205 , n2897 );
xor ( n52206 , n52192 , n52197 );
and ( n2900 , n52206 , n52202 );
and ( n52208 , n52192 , n52197 );
or ( n52209 , n2900 , n52208 );
buf ( n52210 , n52209 );
buf ( n52211 , n405 );
buf ( n52212 , n417 );
and ( n2906 , n52211 , n52212 );
buf ( n52214 , n2906 );
buf ( n52215 , n52214 );
buf ( n52216 , n408 );
buf ( n52217 , n414 );
and ( n2911 , n52216 , n52217 );
buf ( n52219 , n2911 );
buf ( n52220 , n52219 );
buf ( n52221 , n389 );
buf ( n52222 , n393 );
and ( n2916 , n52221 , n52222 );
buf ( n52224 , n2916 );
buf ( n52225 , n52224 );
xor ( n2919 , n52220 , n52225 );
buf ( n52227 , n2919 );
buf ( n52228 , n52227 );
buf ( n52229 , n2860 );
buf ( n52230 , n391 );
and ( n2924 , n52229 , n52230 );
buf ( n52232 , n2924 );
buf ( n52233 , n52232 );
xor ( n52234 , n52215 , n52228 );
xor ( n2928 , n52234 , n52233 );
buf ( n52236 , n2928 );
xor ( n52237 , n52215 , n52228 );
and ( n2931 , n52237 , n52233 );
and ( n52239 , n52215 , n52228 );
or ( n52240 , n2931 , n52239 );
buf ( n52241 , n52240 );
buf ( n52242 , n52154 );
buf ( n52243 , n2841 );
nor ( n52244 , n52242 , n52243 );
buf ( n52245 , n52244 );
buf ( n52246 , n52245 );
buf ( n52247 , n2836 );
buf ( n2941 , n392 );
and ( n52249 , n52247 , n2941 );
buf ( n52250 , n52249 );
buf ( n52251 , n52250 );
buf ( n52252 , n52133 );
xor ( n2946 , n52246 , n52251 );
xor ( n2947 , n2946 , n52252 );
buf ( n52255 , n2947 );
xor ( n2949 , n52246 , n52251 );
and ( n2950 , n2949 , n52252 );
and ( n52258 , n52246 , n52251 );
or ( n2952 , n2950 , n52258 );
buf ( n52260 , n2952 );
buf ( n52261 , n52205 );
buf ( n52262 , n52176 );
buf ( n52263 , n52236 );
xor ( n52264 , n52261 , n52262 );
xor ( n52265 , n52264 , n52263 );
buf ( n52266 , n52265 );
xor ( n52267 , n52261 , n52262 );
and ( n52268 , n52267 , n52263 );
and ( n2956 , n52261 , n52262 );
or ( n52270 , n52268 , n2956 );
buf ( n52271 , n52270 );
not ( n52272 , n390 );
not ( n2960 , n393 );
or ( n52274 , n52272 , n2960 );
not ( n2962 , n391 );
nand ( n52276 , n52274 , n2962 );
nand ( n52277 , n390 , n393 , n391 );
nand ( n2965 , n52276 , n52277 );
nand ( n52279 , n391 , n392 );
nor ( n52280 , n2965 , n52279 );
not ( n52281 , n52280 );
nand ( n52282 , n2965 , n52279 );
and ( n52283 , n52281 , n52282 );
not ( n2969 , n52139 );
and ( n52285 , n392 , n393 );
nand ( n2971 , n2969 , n52285 );
not ( n52287 , n2971 );
and ( n52288 , n52283 , n52287 );
not ( n52289 , n52283 );
and ( n2975 , n52289 , n2971 );
nor ( n52291 , n52288 , n2975 );
buf ( n52292 , n52291 );
buf ( n2978 , n52292 );
buf ( n52294 , n2978 );
buf ( n52295 , n52294 );
buf ( n52296 , n393 );
and ( n52297 , n52295 , n52296 );
buf ( n52298 , n52297 );
buf ( n52299 , n52298 );
buf ( n52300 , n52255 );
buf ( n52301 , n52187 );
xor ( n52302 , n52299 , n52300 );
xor ( n2988 , n52302 , n52301 );
buf ( n52304 , n2988 );
xor ( n2990 , n52299 , n52300 );
and ( n2991 , n2990 , n52301 );
and ( n2992 , n52299 , n52300 );
or ( n2993 , n2991 , n2992 );
buf ( n52309 , n2993 );
buf ( n52310 , n407 );
buf ( n52311 , n414 );
and ( n2997 , n52310 , n52311 );
buf ( n52313 , n2997 );
buf ( n52314 , n52313 );
buf ( n52315 , n408 );
buf ( n52316 , n413 );
and ( n52317 , n52315 , n52316 );
buf ( n52318 , n52317 );
buf ( n52319 , n52318 );
buf ( n52320 , n409 );
buf ( n52321 , n412 );
and ( n52322 , n52320 , n52321 );
buf ( n52323 , n52322 );
buf ( n52324 , n52323 );
xor ( n3010 , n52314 , n52319 );
xor ( n52326 , n3010 , n52324 );
buf ( n52327 , n52326 );
xor ( n52328 , n52314 , n52319 );
and ( n3014 , n52328 , n52324 );
and ( n52330 , n52314 , n52319 );
or ( n3016 , n3014 , n52330 );
buf ( n52332 , n3016 );
buf ( n52333 , n388 );
buf ( n52334 , n393 );
and ( n3020 , n52333 , n52334 );
buf ( n3021 , n3020 );
buf ( n52337 , n3021 );
buf ( n52338 , n404 );
buf ( n52339 , n417 );
and ( n52340 , n52338 , n52339 );
buf ( n52341 , n52340 );
buf ( n3027 , n52341 );
buf ( n52343 , n2860 );
buf ( n52344 , n390 );
and ( n52345 , n52343 , n52344 );
buf ( n52346 , n52345 );
buf ( n52347 , n52346 );
xor ( n52348 , n52337 , n3027 );
xor ( n3032 , n52348 , n52347 );
buf ( n52350 , n3032 );
xor ( n52351 , n52337 , n3027 );
and ( n3034 , n52351 , n52347 );
and ( n3035 , n52337 , n3027 );
or ( n52354 , n3034 , n3035 );
buf ( n52355 , n52354 );
buf ( n52356 , n405 );
buf ( n52357 , n416 );
and ( n52358 , n52356 , n52357 );
buf ( n52359 , n52358 );
buf ( n52360 , n52359 );
buf ( n3043 , n406 );
buf ( n3044 , n415 );
and ( n3045 , n3043 , n3044 );
buf ( n3046 , n3045 );
buf ( n52365 , n3046 );
xor ( n52366 , n52360 , n52365 );
buf ( n52367 , n52366 );
buf ( n52368 , n52367 );
buf ( n3051 , n2836 );
buf ( n52370 , n391 );
and ( n52371 , n3051 , n52370 );
buf ( n52372 , n52371 );
buf ( n52373 , n52372 );
and ( n52374 , n52220 , n52225 );
buf ( n52375 , n52374 );
buf ( n52376 , n52375 );
xor ( n3059 , n52368 , n52373 );
xor ( n52378 , n3059 , n52376 );
buf ( n52379 , n52378 );
xor ( n3062 , n52368 , n52373 );
and ( n3063 , n3062 , n52376 );
and ( n52382 , n52368 , n52373 );
or ( n3065 , n3063 , n52382 );
buf ( n52384 , n3065 );
buf ( n52385 , n52210 );
buf ( n52386 , n52327 );
buf ( n52387 , n52350 );
xor ( n52388 , n52385 , n52386 );
xor ( n52389 , n52388 , n52387 );
buf ( n52390 , n52389 );
xor ( n52391 , n52385 , n52386 );
and ( n52392 , n52391 , n52387 );
and ( n52393 , n52385 , n52386 );
or ( n52394 , n52392 , n52393 );
buf ( n52395 , n52394 );
buf ( n52396 , n52241 );
buf ( n52397 , n52260 );
buf ( n52398 , n52379 );
xor ( n52399 , n52396 , n52397 );
xor ( n3082 , n52399 , n52398 );
buf ( n52401 , n3082 );
xor ( n52402 , n52396 , n52397 );
and ( n3085 , n52402 , n52398 );
and ( n52404 , n52396 , n52397 );
or ( n52405 , n3085 , n52404 );
buf ( n52406 , n52405 );
buf ( n52407 , n52294 );
buf ( n52408 , n392 );
and ( n52409 , n52407 , n52408 );
buf ( n52410 , n52409 );
buf ( n52411 , n52410 );
and ( n52412 , n52285 , n391 , n393 );
not ( n52413 , n52412 );
nand ( n52414 , n52413 , n52281 );
nand ( n52415 , n390 , n392 );
not ( n3097 , n52415 );
nand ( n52417 , n389 , n393 );
not ( n52418 , n52417 );
or ( n52419 , n3097 , n52418 );
nand ( n52420 , n390 , n392 , n393 , n389 );
nand ( n3102 , n52419 , n52420 );
nand ( n52422 , n393 , n390 , n391 );
nand ( n52423 , n3102 , n52422 );
buf ( n52424 , n52423 );
not ( n52425 , n3102 );
not ( n3107 , n52422 );
nand ( n52427 , n52425 , n3107 );
nand ( n52428 , n52424 , n52427 );
xnor ( n3110 , n52414 , n52428 );
buf ( n52430 , n3110 );
buf ( n52431 , n52430 );
buf ( n52432 , n52431 );
buf ( n52433 , n52432 );
buf ( n52434 , n393 );
and ( n3116 , n52433 , n52434 );
buf ( n52436 , n3116 );
buf ( n52437 , n52436 );
buf ( n52438 , n52390 );
xor ( n3120 , n52411 , n52437 );
xor ( n3121 , n3120 , n52438 );
buf ( n52441 , n3121 );
xor ( n52442 , n52411 , n52437 );
and ( n52443 , n52442 , n52438 );
and ( n52444 , n52411 , n52437 );
or ( n3126 , n52443 , n52444 );
buf ( n52446 , n3126 );
buf ( n3128 , n52271 );
buf ( n3129 , n52401 );
buf ( n52449 , n52441 );
xor ( n52450 , n3128 , n3129 );
xor ( n3132 , n52450 , n52449 );
buf ( n52452 , n3132 );
xor ( n3134 , n3128 , n3129 );
and ( n3135 , n3134 , n52449 );
and ( n52455 , n3128 , n3129 );
or ( n3137 , n3135 , n52455 );
buf ( n52457 , n3137 );
buf ( n52458 , n409 );
buf ( n52459 , n411 );
and ( n3141 , n52458 , n52459 );
buf ( n52461 , n3141 );
buf ( n52462 , n52461 );
buf ( n52463 , n387 );
buf ( n52464 , n393 );
and ( n52465 , n52463 , n52464 );
buf ( n52466 , n52465 );
buf ( n52467 , n52466 );
buf ( n52468 , n405 );
buf ( n52469 , n415 );
and ( n3151 , n52468 , n52469 );
buf ( n52471 , n3151 );
buf ( n52472 , n52471 );
xor ( n3154 , n52462 , n52467 );
xor ( n52474 , n3154 , n52472 );
buf ( n52475 , n52474 );
xor ( n52476 , n52462 , n52467 );
and ( n3158 , n52476 , n52472 );
and ( n52478 , n52462 , n52467 );
or ( n52479 , n3158 , n52478 );
buf ( n52480 , n52479 );
buf ( n52481 , n407 );
buf ( n52482 , n413 );
and ( n52483 , n52481 , n52482 );
buf ( n52484 , n52483 );
buf ( n3166 , n52484 );
buf ( n52486 , n408 );
buf ( n52487 , n412 );
and ( n52488 , n52486 , n52487 );
buf ( n52489 , n52488 );
buf ( n52490 , n52489 );
buf ( n52491 , n406 );
buf ( n52492 , n414 );
and ( n3174 , n52491 , n52492 );
buf ( n52494 , n3174 );
buf ( n52495 , n52494 );
xor ( n3177 , n3166 , n52490 );
xor ( n52497 , n3177 , n52495 );
buf ( n52498 , n52497 );
xor ( n52499 , n3166 , n52490 );
and ( n3181 , n52499 , n52495 );
and ( n52501 , n3166 , n52490 );
or ( n52502 , n3181 , n52501 );
buf ( n52503 , n52502 );
buf ( n52504 , n2836 );
buf ( n52505 , n390 );
and ( n52506 , n52504 , n52505 );
buf ( n52507 , n52506 );
buf ( n3189 , n52507 );
buf ( n52509 , n403 );
buf ( n52510 , n417 );
and ( n52511 , n52509 , n52510 );
buf ( n52512 , n52511 );
buf ( n52513 , n52512 );
buf ( n52514 , n404 );
buf ( n3196 , n416 );
and ( n52516 , n52514 , n3196 );
buf ( n52517 , n52516 );
buf ( n52518 , n52517 );
xor ( n52519 , n52513 , n52518 );
buf ( n52520 , n52519 );
buf ( n52521 , n52520 );
buf ( n52522 , n2860 );
buf ( n52523 , n389 );
and ( n3205 , n52522 , n52523 );
buf ( n52525 , n3205 );
buf ( n52526 , n52525 );
xor ( n3208 , n3189 , n52521 );
xor ( n52528 , n3208 , n52526 );
buf ( n52529 , n52528 );
xor ( n52530 , n3189 , n52521 );
and ( n3212 , n52530 , n52526 );
and ( n52532 , n3189 , n52521 );
or ( n52533 , n3212 , n52532 );
buf ( n52534 , n52533 );
and ( n52535 , n52360 , n52365 );
buf ( n52536 , n52535 );
buf ( n52537 , n52536 );
buf ( n3219 , n52332 );
buf ( n3220 , n52475 );
xor ( n3221 , n52537 , n3219 );
xor ( n3222 , n3221 , n3220 );
buf ( n3223 , n3222 );
xor ( n3224 , n52537 , n3219 );
and ( n3225 , n3224 , n3220 );
and ( n3226 , n52537 , n3219 );
or ( n3227 , n3225 , n3226 );
buf ( n3228 , n3227 );
buf ( n3229 , n52498 );
buf ( n3230 , n52355 );
buf ( n52550 , n52384 );
xor ( n3232 , n3229 , n3230 );
xor ( n3233 , n3232 , n52550 );
buf ( n3234 , n3233 );
xor ( n3235 , n3229 , n3230 );
and ( n3236 , n3235 , n52550 );
and ( n3237 , n3229 , n3230 );
or ( n3238 , n3236 , n3237 );
buf ( n3239 , n3238 );
buf ( n52559 , n52291 );
not ( n3241 , n52559 );
buf ( n52561 , n2962 );
nor ( n3243 , n3241 , n52561 );
buf ( n52563 , n3243 );
buf ( n52564 , n52563 );
buf ( n52565 , n52529 );
buf ( n52566 , n3110 );
buf ( n52567 , n392 );
and ( n3249 , n52566 , n52567 );
buf ( n52569 , n3249 );
buf ( n52570 , n52569 );
xor ( n3252 , n52564 , n52565 );
xor ( n3253 , n3252 , n52570 );
buf ( n52573 , n3253 );
xor ( n3255 , n52564 , n52565 );
and ( n3256 , n3255 , n52570 );
and ( n3257 , n52564 , n52565 );
or ( n3258 , n3256 , n3257 );
buf ( n52578 , n3258 );
buf ( n52579 , n3223 );
nand ( n3261 , n2962 , n390 );
not ( n52581 , n3261 );
nand ( n52582 , n392 , n393 , n389 , n390 );
not ( n52583 , n52582 );
xor ( n52584 , n52581 , n52583 );
nand ( n3266 , n388 , n393 );
not ( n3267 , n3266 );
nand ( n52587 , n389 , n392 );
not ( n3269 , n52587 );
or ( n3270 , n3267 , n3269 );
nand ( n3271 , n389 , n392 , n388 , n393 );
nand ( n3272 , n3270 , n3271 );
not ( n52592 , n3272 );
xnor ( n52593 , n52584 , n52592 );
nand ( n52594 , n52280 , n52423 );
nand ( n3276 , n52423 , n52412 );
nand ( n52596 , n52594 , n3276 , n52427 );
buf ( n52597 , n52596 );
and ( n52598 , n52593 , n52597 );
not ( n52599 , n52598 );
not ( n3281 , n52581 );
not ( n52601 , n3272 );
not ( n52602 , n52601 );
or ( n52603 , n3281 , n52602 );
nand ( n52604 , n3272 , n3261 );
nand ( n3286 , n52603 , n52604 );
not ( n52606 , n3286 );
buf ( n52607 , n52606 );
nor ( n3289 , n52607 , n52582 );
nor ( n3290 , n52583 , n3286 );
or ( n52610 , n3289 , n3290 );
not ( n3292 , n52597 );
nand ( n3293 , n52610 , n3292 );
nand ( n3294 , n52599 , n3293 );
buf ( n52614 , n3294 );
buf ( n52615 , n393 );
and ( n52616 , n52614 , n52615 );
buf ( n52617 , n52616 );
buf ( n52618 , n52617 );
buf ( n52619 , n52395 );
xor ( n52620 , n52579 , n52618 );
xor ( n52621 , n52620 , n52619 );
buf ( n52622 , n52621 );
xor ( n3304 , n52579 , n52618 );
and ( n52624 , n3304 , n52619 );
and ( n52625 , n52579 , n52618 );
or ( n52626 , n52624 , n52625 );
buf ( n52627 , n52626 );
buf ( n52628 , n52406 );
buf ( n52629 , n3234 );
buf ( n3311 , n52573 );
xor ( n3312 , n52628 , n52629 );
xor ( n3313 , n3312 , n3311 );
buf ( n3314 , n3313 );
xor ( n3315 , n52628 , n52629 );
and ( n3316 , n3315 , n3311 );
and ( n3317 , n52628 , n52629 );
or ( n3318 , n3316 , n3317 );
buf ( n3319 , n3318 );
buf ( n3320 , n52446 );
buf ( n3321 , n52622 );
buf ( n52641 , n3314 );
xor ( n52642 , n3320 , n3321 );
xor ( n52643 , n52642 , n52641 );
buf ( n52644 , n52643 );
xor ( n52645 , n3320 , n3321 );
and ( n3327 , n52645 , n52641 );
and ( n52647 , n3320 , n3321 );
or ( n52648 , n3327 , n52647 );
buf ( n52649 , n52648 );
buf ( n52650 , n406 );
buf ( n52651 , n413 );
and ( n52652 , n52650 , n52651 );
buf ( n52653 , n52652 );
buf ( n52654 , n52653 );
buf ( n52655 , n403 );
buf ( n3337 , n416 );
and ( n3338 , n52655 , n3337 );
buf ( n52658 , n3338 );
buf ( n52659 , n52658 );
buf ( n52660 , n404 );
buf ( n52661 , n415 );
and ( n52662 , n52660 , n52661 );
buf ( n52663 , n52662 );
buf ( n52664 , n52663 );
xor ( n3346 , n52654 , n52659 );
xor ( n3347 , n3346 , n52664 );
buf ( n52667 , n3347 );
xor ( n52668 , n52654 , n52659 );
and ( n52669 , n52668 , n52664 );
and ( n52670 , n52654 , n52659 );
or ( n3352 , n52669 , n52670 );
buf ( n52672 , n3352 );
buf ( n52673 , n409 );
buf ( n52674 , n410 );
and ( n3356 , n52673 , n52674 );
buf ( n52676 , n3356 );
buf ( n52677 , n52676 );
and ( n52678 , n405 , n414 );
buf ( n52679 , n52678 );
buf ( n52680 , n407 );
buf ( n52681 , n412 );
and ( n3363 , n52680 , n52681 );
buf ( n52683 , n3363 );
buf ( n52684 , n52683 );
xor ( n3366 , n52677 , n52679 );
xor ( n3367 , n3366 , n52684 );
buf ( n52687 , n3367 );
xor ( n3369 , n52677 , n52679 );
and ( n52689 , n3369 , n52684 );
and ( n52690 , n52677 , n52679 );
or ( n52691 , n52689 , n52690 );
buf ( n52692 , n52691 );
buf ( n52693 , n3319 );
buf ( n3375 , n52578 );
not ( n3376 , n52596 );
nand ( n3377 , n3286 , n52582 );
not ( n3378 , n3377 );
or ( n3379 , n3376 , n3378 );
nand ( n3380 , n52606 , n52583 );
nand ( n3381 , n3379 , n3380 );
buf ( n3382 , n3381 );
not ( n3383 , n3382 );
not ( n3384 , n3383 );
nand ( n3385 , n389 , n392 );
nand ( n3386 , n388 , n393 );
nand ( n3387 , n3385 , n3386 );
not ( n3388 , n3387 );
not ( n3389 , n52581 );
or ( n3390 , n3388 , n3389 );
or ( n3391 , n3386 , n3385 );
nand ( n3392 , n3390 , n3391 );
not ( n3393 , n3392 );
nand ( n3394 , n390 , n391 );
nand ( n3395 , n387 , n393 );
not ( n3396 , n3395 );
xor ( n3397 , n3394 , n3396 );
nand ( n52717 , n389 , n391 );
not ( n52718 , n52717 );
nand ( n3400 , n388 , n392 );
not ( n52720 , n3400 );
or ( n52721 , n52718 , n52720 );
nand ( n52722 , n392 , n389 , n391 , n388 );
nand ( n3404 , n52721 , n52722 );
xnor ( n3405 , n3397 , n3404 );
and ( n52725 , n3393 , n3405 );
not ( n3407 , n3393 );
not ( n3408 , n3405 );
and ( n3409 , n3407 , n3408 );
nor ( n3410 , n52725 , n3409 );
not ( n52730 , n3410 );
or ( n52731 , n3384 , n52730 );
not ( n52732 , n3410 );
nand ( n52733 , n52732 , n3382 );
nand ( n3415 , n52731 , n52733 );
not ( n3416 , n3415 );
not ( n52736 , n3416 );
buf ( n52737 , n52736 );
buf ( n52738 , n393 );
and ( n3420 , n52737 , n52738 );
buf ( n52740 , n3420 );
buf ( n52741 , n52740 );
xor ( n52742 , n3375 , n52741 );
buf ( n52743 , n52534 );
buf ( n52744 , n52294 );
buf ( n52745 , n390 );
and ( n52746 , n52744 , n52745 );
buf ( n52747 , n52746 );
buf ( n3429 , n52747 );
xor ( n3430 , n52743 , n3429 );
buf ( n52750 , n2860 );
buf ( n3432 , n388 );
and ( n52752 , n52750 , n3432 );
buf ( n52753 , n52752 );
buf ( n52754 , n52753 );
buf ( n52755 , n2836 );
buf ( n52756 , n389 );
and ( n3438 , n52755 , n52756 );
buf ( n52758 , n3438 );
buf ( n52759 , n52758 );
xor ( n3441 , n52754 , n52759 );
buf ( n52761 , n52480 );
xor ( n3443 , n3441 , n52761 );
buf ( n52763 , n3443 );
buf ( n52764 , n52763 );
xor ( n52765 , n3430 , n52764 );
buf ( n52766 , n52765 );
buf ( n52767 , n52766 );
xor ( n52768 , n52742 , n52767 );
buf ( n52769 , n52768 );
buf ( n52770 , n52769 );
buf ( n52771 , n52627 );
buf ( n52772 , n408 );
buf ( n52773 , n411 );
and ( n52774 , n52772 , n52773 );
buf ( n52775 , n52774 );
buf ( n52776 , n52775 );
and ( n3458 , n386 , n393 );
and ( n52778 , n402 , n417 );
xor ( n52779 , n3458 , n52778 );
buf ( n52780 , n52779 );
xor ( n3462 , n52776 , n52780 );
and ( n52782 , n52513 , n52518 );
buf ( n52783 , n52782 );
buf ( n52784 , n52783 );
xor ( n3466 , n3462 , n52784 );
buf ( n52786 , n3466 );
buf ( n52787 , n52786 );
buf ( n3469 , n3110 );
buf ( n3470 , n391 );
and ( n3471 , n3469 , n3470 );
buf ( n3472 , n3471 );
buf ( n52792 , n3472 );
xor ( n52793 , n52787 , n52792 );
buf ( n52794 , n3228 );
xor ( n3476 , n52793 , n52794 );
buf ( n52796 , n3476 );
buf ( n52797 , n52796 );
xor ( n52798 , n52771 , n52797 );
buf ( n52799 , n3239 );
buf ( n52800 , n3294 );
buf ( n52801 , n392 );
and ( n52802 , n52800 , n52801 );
buf ( n52803 , n52802 );
buf ( n52804 , n52803 );
xor ( n52805 , n52799 , n52804 );
buf ( n3487 , n52503 );
buf ( n3488 , n52687 );
xor ( n3489 , n3487 , n3488 );
buf ( n52809 , n52667 );
xor ( n52810 , n3489 , n52809 );
buf ( n52811 , n52810 );
buf ( n52812 , n52811 );
xor ( n52813 , n52805 , n52812 );
buf ( n52814 , n52813 );
buf ( n52815 , n52814 );
xor ( n3497 , n52798 , n52815 );
buf ( n52817 , n3497 );
buf ( n52818 , n52817 );
xor ( n3500 , n52693 , n52770 );
xor ( n52820 , n3500 , n52818 );
buf ( n52821 , n52820 );
xor ( n52822 , n52693 , n52770 );
and ( n52823 , n52822 , n52818 );
and ( n3505 , n52693 , n52770 );
or ( n3506 , n52823 , n3505 );
buf ( n52826 , n3506 );
xor ( n3508 , n52776 , n52780 );
and ( n3509 , n3508 , n52784 );
and ( n3510 , n52776 , n52780 );
or ( n3511 , n3509 , n3510 );
buf ( n3512 , n3511 );
xor ( n52832 , n52754 , n52759 );
and ( n52833 , n52832 , n52761 );
and ( n52834 , n52754 , n52759 );
or ( n3516 , n52833 , n52834 );
buf ( n52836 , n3516 );
xor ( n52837 , n3487 , n3488 );
and ( n3519 , n52837 , n52809 );
and ( n3520 , n3487 , n3488 );
or ( n3521 , n3519 , n3520 );
buf ( n52841 , n3521 );
xor ( n52842 , n52743 , n3429 );
and ( n52843 , n52842 , n52764 );
and ( n52844 , n52743 , n3429 );
or ( n3526 , n52843 , n52844 );
buf ( n52846 , n3526 );
xor ( n52847 , n52787 , n52792 );
and ( n52848 , n52847 , n52794 );
and ( n3530 , n52787 , n52792 );
or ( n52850 , n52848 , n3530 );
buf ( n52851 , n52850 );
xor ( n52852 , n52799 , n52804 );
and ( n3534 , n52852 , n52812 );
and ( n52854 , n52799 , n52804 );
or ( n3536 , n3534 , n52854 );
buf ( n52856 , n3536 );
xor ( n52857 , n3375 , n52741 );
and ( n3539 , n52857 , n52767 );
and ( n3540 , n3375 , n52741 );
or ( n3541 , n3539 , n3540 );
buf ( n52861 , n3541 );
xor ( n52862 , n52771 , n52797 );
and ( n52863 , n52862 , n52815 );
and ( n3545 , n52771 , n52797 );
or ( n3546 , n52863 , n3545 );
buf ( n52866 , n3546 );
buf ( n52867 , n408 );
buf ( n52868 , n410 );
and ( n3550 , n52867 , n52868 );
buf ( n52870 , n3550 );
buf ( n52871 , n52870 );
buf ( n52872 , n403 );
buf ( n52873 , n415 );
and ( n3555 , n52872 , n52873 );
buf ( n52875 , n3555 );
buf ( n52876 , n52875 );
buf ( n52877 , n404 );
buf ( n52878 , n414 );
and ( n3560 , n52877 , n52878 );
buf ( n52880 , n3560 );
buf ( n52881 , n52880 );
xor ( n3563 , n52871 , n52876 );
xor ( n3564 , n3563 , n52881 );
buf ( n52884 , n3564 );
xor ( n52885 , n52871 , n52876 );
and ( n52886 , n52885 , n52881 );
and ( n3568 , n52871 , n52876 );
or ( n52888 , n52886 , n3568 );
buf ( n52889 , n52888 );
buf ( n52890 , n402 );
buf ( n52891 , n416 );
and ( n3573 , n52890 , n52891 );
buf ( n52893 , n3573 );
buf ( n52894 , n52893 );
buf ( n52895 , n407 );
buf ( n52896 , n411 );
and ( n3578 , n52895 , n52896 );
buf ( n52898 , n3578 );
buf ( n52899 , n52898 );
buf ( n52900 , n405 );
buf ( n52901 , n413 );
and ( n3583 , n52900 , n52901 );
buf ( n52903 , n3583 );
buf ( n52904 , n52903 );
xor ( n3586 , n52894 , n52899 );
xor ( n3587 , n3586 , n52904 );
buf ( n52907 , n3587 );
xor ( n3589 , n52894 , n52899 );
and ( n52909 , n3589 , n52904 );
and ( n52910 , n52894 , n52899 );
or ( n52911 , n52909 , n52910 );
buf ( n52912 , n52911 );
buf ( n52913 , n52907 );
buf ( n52914 , n52884 );
xor ( n52915 , n52913 , n52914 );
buf ( n52916 , n3512 );
xor ( n3598 , n52915 , n52916 );
buf ( n52918 , n3598 );
buf ( n52919 , n52918 );
buf ( n52920 , n3294 );
buf ( n52921 , n391 );
and ( n52922 , n52920 , n52921 );
buf ( n52923 , n52922 );
buf ( n52924 , n52923 );
xor ( n52925 , n52919 , n52924 );
buf ( n52926 , n52846 );
xor ( n52927 , n52925 , n52926 );
buf ( n52928 , n52927 );
buf ( n52929 , n52928 );
buf ( n3611 , n52861 );
buf ( n3612 , n3415 );
buf ( n3613 , n392 );
and ( n3614 , n3612 , n3613 );
buf ( n3615 , n3614 );
buf ( n52935 , n3615 );
buf ( n52936 , n52851 );
xor ( n3618 , n52935 , n52936 );
buf ( n52938 , n406 );
buf ( n52939 , n412 );
and ( n3621 , n52938 , n52939 );
buf ( n52941 , n3621 );
buf ( n52942 , n52941 );
and ( n52943 , n3458 , n52778 );
buf ( n52944 , n52943 );
xor ( n52945 , n52942 , n52944 );
not ( n3627 , n388 );
nor ( n52947 , n52142 , n3627 );
buf ( n52948 , n52947 );
xor ( n3630 , n52945 , n52948 );
buf ( n52950 , n3630 );
buf ( n3632 , n52950 );
buf ( n3633 , n52836 );
xor ( n3634 , n3632 , n3633 );
buf ( n52954 , n52294 );
buf ( n52955 , n389 );
and ( n3637 , n52954 , n52955 );
buf ( n52957 , n3637 );
buf ( n52958 , n52957 );
xor ( n3640 , n3634 , n52958 );
buf ( n52960 , n3640 );
buf ( n52961 , n52960 );
xor ( n3643 , n3618 , n52961 );
buf ( n52963 , n3643 );
buf ( n52964 , n52963 );
xor ( n52965 , n52929 , n3611 );
xor ( n3647 , n52965 , n52964 );
buf ( n52967 , n3647 );
xor ( n3649 , n52929 , n3611 );
and ( n3650 , n3649 , n52964 );
and ( n3651 , n52929 , n3611 );
or ( n3652 , n3650 , n3651 );
buf ( n52972 , n3652 );
not ( n3654 , n3394 );
not ( n3655 , n3654 );
not ( n3656 , n3396 );
or ( n3657 , n3655 , n3656 );
nand ( n3658 , n3657 , n3404 );
nand ( n3659 , n3395 , n3394 );
nand ( n3660 , n3658 , n3659 );
not ( n3661 , n3660 );
not ( n3662 , n3661 );
nand ( n3663 , n386 , n393 );
nand ( n3664 , n388 , n391 );
and ( n3665 , n3663 , n3664 );
not ( n3666 , n3663 );
and ( n3667 , n388 , n391 );
and ( n3668 , n3666 , n3667 );
nor ( n3669 , n3665 , n3668 );
nand ( n3670 , n387 , n392 );
not ( n3671 , n3670 );
and ( n3672 , n3669 , n3671 );
not ( n3673 , n3669 );
and ( n3674 , n3673 , n3670 );
nor ( n3675 , n3672 , n3674 );
nand ( n3676 , n389 , n391 , n388 , n392 );
not ( n3677 , n3676 );
not ( n3678 , n390 );
nand ( n3679 , n3678 , n389 );
not ( n3680 , n3679 );
xnor ( n3681 , n3677 , n3680 );
and ( n3682 , n3675 , n3681 );
not ( n3683 , n3675 );
not ( n3684 , n3681 );
and ( n3685 , n3683 , n3684 );
nor ( n3686 , n3682 , n3685 );
not ( n3687 , n3686 );
not ( n3688 , n3687 );
or ( n3689 , n3662 , n3688 );
nand ( n53009 , n3686 , n3660 );
buf ( n53010 , n53009 );
nand ( n3692 , n3689 , n53010 );
nand ( n53012 , n3405 , n3393 );
not ( n53013 , n53012 );
not ( n3695 , n3381 );
or ( n53015 , n53013 , n3695 );
nand ( n53016 , n3408 , n3392 );
nand ( n53017 , n53015 , n53016 );
buf ( n3699 , n53017 );
not ( n53019 , n3699 );
and ( n53020 , n3692 , n53019 );
not ( n3702 , n3692 );
and ( n53022 , n3702 , n3699 );
nor ( n53023 , n53020 , n53022 );
buf ( n53024 , n53023 );
buf ( n53025 , n393 );
and ( n53026 , n53024 , n53025 );
buf ( n53027 , n53026 );
buf ( n53028 , n53027 );
buf ( n53029 , n52841 );
buf ( n53030 , n3110 );
buf ( n53031 , n390 );
and ( n53032 , n53030 , n53031 );
buf ( n53033 , n53032 );
buf ( n53034 , n53033 );
xor ( n53035 , n53029 , n53034 );
buf ( n53036 , n2860 );
buf ( n53037 , n387 );
and ( n53038 , n53036 , n53037 );
buf ( n53039 , n53038 );
buf ( n53040 , n53039 );
buf ( n3722 , n52672 );
xor ( n53042 , n53040 , n3722 );
buf ( n53043 , n52692 );
xor ( n53044 , n53042 , n53043 );
buf ( n53045 , n53044 );
buf ( n53046 , n53045 );
xor ( n53047 , n53035 , n53046 );
buf ( n53048 , n53047 );
buf ( n3730 , n53048 );
xor ( n3731 , n53028 , n3730 );
buf ( n53051 , n52856 );
xor ( n53052 , n3731 , n53051 );
buf ( n53053 , n53052 );
buf ( n53054 , n53053 );
buf ( n53055 , n52866 );
buf ( n53056 , n52967 );
xor ( n53057 , n53054 , n53055 );
xor ( n3739 , n53057 , n53056 );
buf ( n53059 , n3739 );
xor ( n53060 , n53054 , n53055 );
and ( n53061 , n53060 , n53056 );
and ( n3743 , n53054 , n53055 );
or ( n53063 , n53061 , n3743 );
buf ( n53064 , n53063 );
xor ( n53065 , n52942 , n52944 );
and ( n53066 , n53065 , n52948 );
and ( n3748 , n52942 , n52944 );
or ( n53068 , n53066 , n3748 );
buf ( n53069 , n53068 );
xor ( n3751 , n53040 , n3722 );
and ( n53071 , n3751 , n53043 );
and ( n3753 , n53040 , n3722 );
or ( n53073 , n53071 , n3753 );
buf ( n53074 , n53073 );
xor ( n3756 , n52913 , n52914 );
and ( n53076 , n3756 , n52916 );
and ( n53077 , n52913 , n52914 );
or ( n53078 , n53076 , n53077 );
buf ( n53079 , n53078 );
xor ( n53080 , n3632 , n3633 );
and ( n53081 , n53080 , n52958 );
and ( n3763 , n3632 , n3633 );
or ( n53083 , n53081 , n3763 );
buf ( n53084 , n53083 );
xor ( n3766 , n53029 , n53034 );
and ( n53086 , n3766 , n53046 );
and ( n3768 , n53029 , n53034 );
or ( n53088 , n53086 , n3768 );
buf ( n53089 , n53088 );
xor ( n3771 , n52919 , n52924 );
and ( n53091 , n3771 , n52926 );
and ( n53092 , n52919 , n52924 );
or ( n3774 , n53091 , n53092 );
buf ( n53094 , n3774 );
xor ( n53095 , n52935 , n52936 );
and ( n3777 , n53095 , n52961 );
and ( n3778 , n52935 , n52936 );
or ( n53098 , n3777 , n3778 );
buf ( n53099 , n53098 );
xor ( n3781 , n53028 , n3730 );
and ( n3782 , n3781 , n53051 );
and ( n3783 , n53028 , n3730 );
or ( n53103 , n3782 , n3783 );
buf ( n53104 , n53103 );
buf ( n53105 , n402 );
buf ( n53106 , n415 );
and ( n3788 , n53105 , n53106 );
buf ( n53108 , n3788 );
buf ( n53109 , n53108 );
buf ( n53110 , n403 );
buf ( n53111 , n414 );
and ( n3792 , n53110 , n53111 );
buf ( n53113 , n3792 );
buf ( n53114 , n53113 );
buf ( n53115 , n406 );
buf ( n53116 , n411 );
and ( n3797 , n53115 , n53116 );
buf ( n53118 , n3797 );
buf ( n53119 , n53118 );
xor ( n3800 , n53109 , n53114 );
xor ( n3801 , n3800 , n53119 );
buf ( n53122 , n3801 );
xor ( n53123 , n53109 , n53114 );
and ( n3804 , n53123 , n53119 );
and ( n3805 , n53109 , n53114 );
or ( n3806 , n3804 , n3805 );
buf ( n53127 , n3806 );
buf ( n53128 , n404 );
buf ( n53129 , n413 );
and ( n3810 , n53128 , n53129 );
buf ( n53131 , n3810 );
buf ( n53132 , n53131 );
nand ( n53133 , n405 , n412 );
not ( n3814 , n53133 );
buf ( n53135 , n3814 );
buf ( n53136 , n407 );
buf ( n53137 , n410 );
and ( n53138 , n53136 , n53137 );
buf ( n53139 , n53138 );
buf ( n53140 , n53139 );
xor ( n3821 , n53132 , n53135 );
xor ( n3822 , n3821 , n53140 );
buf ( n53143 , n3822 );
xor ( n53144 , n53132 , n53135 );
and ( n53145 , n53144 , n53140 );
and ( n3826 , n53132 , n53135 );
or ( n53147 , n53145 , n3826 );
buf ( n53148 , n53147 );
buf ( n3829 , n53104 );
buf ( n53150 , n53089 );
buf ( n53151 , n3415 );
buf ( n53152 , n391 );
and ( n53153 , n53151 , n53152 );
buf ( n53154 , n53153 );
buf ( n3835 , n53154 );
xor ( n3836 , n53150 , n3835 );
buf ( n53157 , n53069 );
buf ( n53158 , n2860 );
buf ( n53159 , n386 );
and ( n3840 , n53158 , n53159 );
buf ( n53161 , n3840 );
buf ( n53162 , n53161 );
buf ( n53163 , n2836 );
buf ( n53164 , n387 );
and ( n3845 , n53163 , n53164 );
buf ( n53166 , n3845 );
buf ( n53167 , n53166 );
xor ( n53168 , n53162 , n53167 );
buf ( n53169 , n52912 );
xor ( n53170 , n53168 , n53169 );
buf ( n53171 , n53170 );
buf ( n53172 , n53171 );
xor ( n53173 , n53157 , n53172 );
and ( n3854 , n52294 , n388 );
buf ( n53175 , n3854 );
xor ( n53176 , n53173 , n53175 );
buf ( n53177 , n53176 );
buf ( n53178 , n53177 );
xor ( n3859 , n3836 , n53178 );
buf ( n53180 , n3859 );
buf ( n53181 , n53180 );
buf ( n53182 , n53023 );
buf ( n3863 , n53182 );
buf ( n53184 , n3863 );
buf ( n53185 , n53184 );
buf ( n53186 , n392 );
and ( n3867 , n53185 , n53186 );
buf ( n53188 , n3867 );
buf ( n53189 , n53188 );
buf ( n3870 , n53074 );
buf ( n53191 , n52432 );
buf ( n53192 , n389 );
and ( n53193 , n53191 , n53192 );
buf ( n53194 , n53193 );
buf ( n53195 , n53194 );
xor ( n53196 , n3870 , n53195 );
buf ( n53197 , n53079 );
xor ( n53198 , n53196 , n53197 );
buf ( n53199 , n53198 );
buf ( n53200 , n53199 );
xor ( n53201 , n53189 , n53200 );
not ( n3882 , n53009 );
not ( n53203 , n53017 );
or ( n3884 , n3882 , n53203 );
nand ( n53205 , n3687 , n3661 );
nand ( n53206 , n3884 , n53205 );
buf ( n53207 , n53206 );
nand ( n53208 , n3676 , n3679 );
not ( n53209 , n53208 );
not ( n3890 , n3675 );
or ( n53211 , n53209 , n3890 );
nand ( n53212 , n3677 , n3680 );
nand ( n53213 , n53211 , n53212 );
not ( n3894 , n53213 );
nand ( n53215 , n389 , n390 );
nand ( n53216 , n388 , n391 );
not ( n3897 , n53216 );
not ( n53218 , n3670 );
or ( n53219 , n3897 , n53218 );
and ( n53220 , n386 , n393 );
nand ( n53221 , n53219 , n53220 );
not ( n3902 , n3664 );
nand ( n53223 , n3902 , n3671 );
and ( n53224 , n53221 , n53223 );
xor ( n3905 , n53215 , n53224 );
and ( n53226 , n386 , n392 );
not ( n3907 , n53226 );
and ( n53228 , n388 , n390 );
nand ( n3909 , n387 , n391 );
nand ( n53230 , n53228 , n3909 );
and ( n53231 , n387 , n391 );
nand ( n3912 , n388 , n390 );
nand ( n53233 , n53231 , n3912 );
nand ( n53234 , n53230 , n53233 );
not ( n3915 , n53234 );
or ( n53236 , n3907 , n3915 );
not ( n53237 , n392 );
not ( n53238 , n386 );
nor ( n3919 , n53237 , n53238 );
not ( n3920 , n3919 );
nand ( n53241 , n53233 , n53230 , n3920 );
nand ( n53242 , n53236 , n53241 );
xor ( n3923 , n3905 , n53242 );
nor ( n53244 , n3894 , n3923 );
not ( n53245 , n53244 );
nand ( n3926 , n3923 , n3894 );
nand ( n53247 , n53245 , n3926 );
xnor ( n53248 , n53207 , n53247 );
buf ( n53249 , n53248 );
buf ( n53250 , n53249 );
buf ( n53251 , n53250 );
buf ( n53252 , n53251 );
buf ( n53253 , n393 );
and ( n53254 , n53252 , n53253 );
buf ( n53255 , n53254 );
buf ( n53256 , n53255 );
xor ( n3937 , n53201 , n53256 );
buf ( n53258 , n3937 );
buf ( n53259 , n53258 );
xor ( n3940 , n3829 , n53181 );
xor ( n3941 , n3940 , n53259 );
buf ( n53262 , n3941 );
xor ( n3943 , n3829 , n53181 );
and ( n3944 , n3943 , n53259 );
and ( n3945 , n3829 , n53181 );
or ( n3946 , n3944 , n3945 );
buf ( n53267 , n3946 );
buf ( n53268 , n53094 );
buf ( n53269 , n52889 );
buf ( n53270 , n53143 );
xor ( n3951 , n53269 , n53270 );
buf ( n53272 , n53122 );
xor ( n3953 , n3951 , n53272 );
buf ( n53274 , n3953 );
buf ( n53275 , n53274 );
buf ( n53276 , n3294 );
buf ( n53277 , n390 );
and ( n3958 , n53276 , n53277 );
buf ( n53279 , n3958 );
buf ( n53280 , n53279 );
xor ( n3961 , n53275 , n53280 );
buf ( n53282 , n53084 );
xor ( n3963 , n3961 , n53282 );
buf ( n53284 , n3963 );
buf ( n3965 , n53284 );
xor ( n3966 , n53268 , n3965 );
buf ( n53287 , n53099 );
xor ( n53288 , n3966 , n53287 );
buf ( n53289 , n53288 );
buf ( n3970 , n53289 );
buf ( n3971 , n52972 );
buf ( n53292 , n53262 );
xor ( n53293 , n3970 , n3971 );
xor ( n53294 , n53293 , n53292 );
buf ( n53295 , n53294 );
xor ( n53296 , n3970 , n3971 );
and ( n53297 , n53296 , n53292 );
and ( n3978 , n3970 , n3971 );
or ( n53299 , n53297 , n3978 );
buf ( n53300 , n53299 );
xor ( n53301 , n53162 , n53167 );
and ( n3982 , n53301 , n53169 );
and ( n53303 , n53162 , n53167 );
or ( n3984 , n3982 , n53303 );
buf ( n53305 , n3984 );
xor ( n53306 , n53269 , n53270 );
and ( n3987 , n53306 , n53272 );
and ( n53308 , n53269 , n53270 );
or ( n53309 , n3987 , n53308 );
buf ( n53310 , n53309 );
xor ( n53311 , n53157 , n53172 );
and ( n3992 , n53311 , n53175 );
and ( n53313 , n53157 , n53172 );
or ( n53314 , n3992 , n53313 );
buf ( n53315 , n53314 );
xor ( n53316 , n3870 , n53195 );
and ( n3997 , n53316 , n53197 );
and ( n3998 , n3870 , n53195 );
or ( n53319 , n3997 , n3998 );
buf ( n53320 , n53319 );
xor ( n4001 , n53275 , n53280 );
and ( n4002 , n4001 , n53282 );
and ( n4003 , n53275 , n53280 );
or ( n53324 , n4002 , n4003 );
buf ( n53325 , n53324 );
xor ( n4006 , n53150 , n3835 );
and ( n4007 , n4006 , n53178 );
and ( n4008 , n53150 , n3835 );
or ( n53329 , n4007 , n4008 );
buf ( n53330 , n53329 );
xor ( n4011 , n53189 , n53200 );
and ( n4012 , n4011 , n53256 );
and ( n4013 , n53189 , n53200 );
or ( n53334 , n4012 , n4013 );
buf ( n53335 , n53334 );
xor ( n4016 , n53268 , n3965 );
and ( n4017 , n4016 , n53287 );
and ( n4018 , n53268 , n3965 );
or ( n53339 , n4017 , n4018 );
buf ( n53340 , n53339 );
buf ( n53341 , n406 );
buf ( n53342 , n410 );
and ( n4023 , n53341 , n53342 );
buf ( n53344 , n4023 );
buf ( n53345 , n53344 );
buf ( n53346 , n404 );
buf ( n53347 , n412 );
and ( n4028 , n53346 , n53347 );
buf ( n4029 , n4028 );
buf ( n53350 , n4029 );
buf ( n53351 , n405 );
buf ( n53352 , n411 );
and ( n4033 , n53351 , n53352 );
buf ( n53354 , n4033 );
buf ( n53355 , n53354 );
xor ( n4036 , n53345 , n53350 );
xor ( n4037 , n4036 , n53355 );
buf ( n53358 , n4037 );
xor ( n53359 , n53345 , n53350 );
and ( n4040 , n53359 , n53355 );
and ( n4041 , n53345 , n53350 );
or ( n4042 , n4040 , n4041 );
buf ( n53363 , n4042 );
buf ( n53364 , n2836 );
buf ( n53365 , n386 );
and ( n53366 , n53364 , n53365 );
buf ( n53367 , n53366 );
buf ( n53368 , n53367 );
buf ( n4049 , n402 );
buf ( n53370 , n414 );
and ( n53371 , n4049 , n53370 );
buf ( n53372 , n53371 );
buf ( n53373 , n53372 );
buf ( n53374 , n403 );
buf ( n53375 , n413 );
and ( n53376 , n53374 , n53375 );
buf ( n53377 , n53376 );
buf ( n53378 , n53377 );
xor ( n53379 , n53373 , n53378 );
buf ( n53380 , n53379 );
buf ( n4061 , n53380 );
buf ( n53382 , n4061 );
buf ( n53383 , n53148 );
xor ( n4064 , n53368 , n53382 );
xor ( n4065 , n4064 , n53383 );
buf ( n53386 , n4065 );
xor ( n53387 , n53368 , n53382 );
and ( n53388 , n53387 , n53383 );
and ( n53389 , n53368 , n53382 );
or ( n4070 , n53388 , n53389 );
buf ( n53391 , n4070 );
buf ( n4072 , n53330 );
buf ( n4073 , n53315 );
buf ( n53394 , n52291 );
not ( n4075 , n53394 );
buf ( n53396 , n387 );
not ( n53397 , n53396 );
buf ( n53398 , n53397 );
buf ( n4079 , n53398 );
nor ( n4080 , n4075 , n4079 );
buf ( n4081 , n4080 );
buf ( n53402 , n4081 );
buf ( n53403 , n53386 );
xor ( n4084 , n53402 , n53403 );
buf ( n53405 , n53310 );
xor ( n4086 , n4084 , n53405 );
buf ( n53407 , n4086 );
buf ( n53408 , n53407 );
xor ( n4089 , n4073 , n53408 );
not ( n53410 , n52736 );
buf ( n4091 , n53410 );
buf ( n4092 , n390 );
not ( n53413 , n4092 );
buf ( n53414 , n53413 );
buf ( n53415 , n53414 );
nor ( n53416 , n4091 , n53415 );
buf ( n53417 , n53416 );
buf ( n53418 , n53417 );
xor ( n53419 , n4089 , n53418 );
buf ( n53420 , n53419 );
buf ( n4101 , n53420 );
xor ( n4102 , n4072 , n4101 );
buf ( n53423 , n53335 );
xor ( n53424 , n4102 , n53423 );
buf ( n53425 , n53424 );
buf ( n53426 , n53425 );
buf ( n53427 , n53267 );
buf ( n53428 , n53023 );
not ( n53429 , n53428 );
buf ( n53430 , n2962 );
nor ( n53431 , n53429 , n53430 );
buf ( n53432 , n53431 );
buf ( n53433 , n53432 );
buf ( n4114 , n53320 );
xor ( n4115 , n53433 , n4114 );
buf ( n53436 , n53325 );
xor ( n53437 , n4115 , n53436 );
buf ( n53438 , n53437 );
buf ( n53439 , n53438 );
buf ( n53440 , n53251 );
buf ( n53441 , n392 );
and ( n53442 , n53440 , n53441 );
buf ( n53443 , n53442 );
buf ( n53444 , n53443 );
buf ( n53445 , n52432 );
buf ( n4126 , n388 );
and ( n53447 , n53445 , n4126 );
buf ( n53448 , n53447 );
buf ( n53449 , n53448 );
buf ( n53450 , n3294 );
buf ( n53451 , n389 );
and ( n53452 , n53450 , n53451 );
buf ( n53453 , n53452 );
buf ( n4134 , n53453 );
xor ( n4135 , n53449 , n4134 );
buf ( n53456 , n53127 );
buf ( n4137 , n53358 );
xor ( n4138 , n53456 , n4137 );
buf ( n4139 , n53305 );
xor ( n4140 , n4138 , n4139 );
buf ( n4141 , n4140 );
buf ( n53462 , n4141 );
xor ( n4143 , n4135 , n53462 );
buf ( n53464 , n4143 );
buf ( n53465 , n53464 );
xor ( n4146 , n53444 , n53465 );
and ( n4147 , n53207 , n3926 );
buf ( n4148 , n53244 );
nor ( n4149 , n4147 , n4148 );
xor ( n4150 , n53215 , n53224 );
and ( n4151 , n4150 , n53242 );
and ( n4152 , n53215 , n53224 );
or ( n4153 , n4151 , n4152 );
nand ( n4154 , n387 , n390 );
not ( n4155 , n3919 );
nand ( n4156 , n3912 , n3909 );
not ( n4157 , n4156 );
or ( n4158 , n4155 , n4157 );
nand ( n4159 , n53228 , n53231 );
nand ( n4160 , n4158 , n4159 );
xor ( n4161 , n4154 , n4160 );
nand ( n4162 , n386 , n391 );
not ( n4163 , n388 );
nor ( n4164 , n4163 , n389 );
xor ( n4165 , n4162 , n4164 );
xnor ( n4166 , n4161 , n4165 );
xnor ( n4167 , n4153 , n4166 );
and ( n4168 , n4149 , n4167 );
not ( n4169 , n4149 );
not ( n4170 , n4167 );
and ( n4171 , n4169 , n4170 );
nor ( n4172 , n4168 , n4171 );
buf ( n53493 , n4172 );
buf ( n53494 , n393 );
and ( n4175 , n53493 , n53494 );
buf ( n53496 , n4175 );
buf ( n53497 , n53496 );
xor ( n4178 , n4146 , n53497 );
buf ( n53499 , n4178 );
buf ( n53500 , n53499 );
xor ( n53501 , n53439 , n53500 );
buf ( n53502 , n53340 );
xor ( n53503 , n53501 , n53502 );
buf ( n53504 , n53503 );
buf ( n53505 , n53504 );
xor ( n53506 , n53426 , n53427 );
xor ( n4187 , n53506 , n53505 );
buf ( n4188 , n4187 );
xor ( n53509 , n53426 , n53427 );
and ( n4190 , n53509 , n53505 );
and ( n4191 , n53426 , n53427 );
or ( n53512 , n4190 , n4191 );
buf ( n53513 , n53512 );
xor ( n4194 , n53456 , n4137 );
and ( n4195 , n4194 , n4139 );
and ( n4196 , n53456 , n4137 );
or ( n53517 , n4195 , n4196 );
buf ( n53518 , n53517 );
xor ( n53519 , n53402 , n53403 );
and ( n53520 , n53519 , n53405 );
and ( n4201 , n53402 , n53403 );
or ( n53522 , n53520 , n4201 );
buf ( n53523 , n53522 );
xor ( n53524 , n53449 , n4134 );
and ( n53525 , n53524 , n53462 );
and ( n53526 , n53449 , n4134 );
or ( n53527 , n53525 , n53526 );
buf ( n53528 , n53527 );
xor ( n53529 , n4073 , n53408 );
and ( n53530 , n53529 , n53418 );
and ( n4211 , n4073 , n53408 );
or ( n53532 , n53530 , n4211 );
buf ( n53533 , n53532 );
xor ( n53534 , n53433 , n4114 );
and ( n53535 , n53534 , n53436 );
and ( n4216 , n53433 , n4114 );
or ( n53537 , n53535 , n4216 );
buf ( n53538 , n53537 );
xor ( n53539 , n53444 , n53465 );
and ( n53540 , n53539 , n53497 );
and ( n53541 , n53444 , n53465 );
or ( n53542 , n53540 , n53541 );
buf ( n53543 , n53542 );
xor ( n4224 , n4072 , n4101 );
and ( n53545 , n4224 , n53423 );
and ( n4226 , n4072 , n4101 );
or ( n4227 , n53545 , n4226 );
buf ( n53548 , n4227 );
xor ( n4229 , n53439 , n53500 );
and ( n53550 , n4229 , n53502 );
and ( n4231 , n53439 , n53500 );
or ( n4232 , n53550 , n4231 );
buf ( n53553 , n4232 );
buf ( n53554 , n402 );
buf ( n53555 , n413 );
and ( n4235 , n53554 , n53555 );
buf ( n53557 , n4235 );
buf ( n53558 , n53557 );
buf ( n53559 , n403 );
buf ( n53560 , n412 );
and ( n4240 , n53559 , n53560 );
buf ( n53562 , n4240 );
buf ( n53563 , n53562 );
buf ( n53564 , n404 );
buf ( n53565 , n411 );
and ( n4245 , n53564 , n53565 );
buf ( n53567 , n4245 );
buf ( n53568 , n53567 );
xor ( n4248 , n53558 , n53563 );
xor ( n53570 , n4248 , n53568 );
buf ( n53571 , n53570 );
xor ( n4251 , n53558 , n53563 );
and ( n4252 , n4251 , n53568 );
and ( n4253 , n53558 , n53563 );
or ( n53575 , n4252 , n4253 );
buf ( n53576 , n53575 );
buf ( n53577 , n405 );
buf ( n53578 , n410 );
and ( n4258 , n53577 , n53578 );
buf ( n53580 , n4258 );
buf ( n53581 , n53580 );
and ( n4261 , n53373 , n53378 );
buf ( n53583 , n4261 );
buf ( n53584 , n53583 );
buf ( n53585 , n53363 );
xor ( n4265 , n53581 , n53584 );
xor ( n4266 , n4265 , n53585 );
buf ( n53588 , n4266 );
xor ( n4268 , n53581 , n53584 );
and ( n53590 , n4268 , n53585 );
and ( n53591 , n53581 , n53584 );
or ( n53592 , n53590 , n53591 );
buf ( n53593 , n53592 );
buf ( n53594 , n53538 );
buf ( n4274 , n53523 );
buf ( n4275 , n52291 );
buf ( n4276 , n386 );
and ( n4277 , n4275 , n4276 );
buf ( n4278 , n4277 );
buf ( n53600 , n4278 );
buf ( n4280 , n3110 );
buf ( n4281 , n387 );
and ( n4282 , n4280 , n4281 );
buf ( n4283 , n4282 );
buf ( n53605 , n4283 );
xor ( n4285 , n53600 , n53605 );
not ( n4286 , n52598 );
and ( n53608 , n3293 , n4286 );
nor ( n4288 , n53608 , n3627 );
buf ( n53610 , n4288 );
xor ( n4290 , n4285 , n53610 );
buf ( n53612 , n4290 );
buf ( n53613 , n53612 );
xor ( n53614 , n4274 , n53613 );
buf ( n53615 , n53023 );
not ( n4295 , n53615 );
buf ( n53617 , n53414 );
nor ( n53618 , n4295 , n53617 );
buf ( n53619 , n53618 );
buf ( n53620 , n53619 );
xor ( n4300 , n53614 , n53620 );
buf ( n53622 , n4300 );
buf ( n53623 , n53622 );
xor ( n53624 , n53594 , n53623 );
buf ( n53625 , n53543 );
xor ( n4305 , n53624 , n53625 );
buf ( n53627 , n4305 );
buf ( n53628 , n53627 );
buf ( n53629 , n53553 );
buf ( n53630 , n53528 );
buf ( n53631 , n53251 );
buf ( n53632 , n391 );
and ( n4312 , n53631 , n53632 );
buf ( n53634 , n4312 );
buf ( n53635 , n53634 );
xor ( n4315 , n53630 , n53635 );
buf ( n53637 , n4172 );
buf ( n4317 , n53637 );
buf ( n53639 , n4317 );
and ( n53640 , n53639 , n392 );
buf ( n53641 , n53640 );
xor ( n53642 , n4315 , n53641 );
buf ( n53643 , n53642 );
buf ( n53644 , n53643 );
buf ( n4324 , n53533 );
and ( n4325 , n4153 , n4166 );
and ( n53647 , n3923 , n3894 );
nor ( n53648 , n4325 , n53647 );
not ( n4328 , n53648 );
not ( n53650 , n53206 );
or ( n53651 , n4328 , n53650 );
not ( n53652 , n4153 );
not ( n4332 , n4166 );
and ( n53654 , n53652 , n4332 );
nand ( n4334 , n4153 , n4166 );
and ( n53656 , n4334 , n53244 );
nor ( n53657 , n53654 , n53656 );
nand ( n4337 , n53651 , n53657 );
buf ( n4338 , n4337 );
not ( n53660 , n388 );
not ( n4340 , n4162 );
nor ( n53662 , n4340 , n389 );
nor ( n4342 , n53660 , n53662 );
not ( n53664 , n4342 );
not ( n4344 , n53664 );
nand ( n53666 , n386 , n390 );
not ( n53667 , n53666 );
nand ( n4347 , n387 , n389 );
not ( n53669 , n4347 );
not ( n4349 , n53669 );
or ( n53671 , n53667 , n4349 );
or ( n53672 , n53666 , n53669 );
nand ( n53673 , n53671 , n53672 );
not ( n53674 , n53673 );
and ( n53675 , n4344 , n53674 );
and ( n4355 , n53664 , n53673 );
nor ( n53677 , n53675 , n4355 );
not ( n53678 , n4154 );
not ( n53679 , n4165 );
or ( n4359 , n53678 , n53679 );
nand ( n53681 , n4359 , n4160 );
or ( n4361 , n4165 , n4154 );
and ( n53683 , n53681 , n4361 );
nor ( n53684 , n53677 , n53683 );
not ( n53685 , n53684 );
nand ( n53686 , n53677 , n53683 );
nand ( n4366 , n53685 , n53686 );
nor ( n53688 , n4338 , n4366 );
not ( n53689 , n53688 );
nand ( n53690 , n4338 , n4366 );
nand ( n53691 , n53689 , n53690 );
and ( n4371 , n53691 , n393 );
buf ( n53693 , n4371 );
xor ( n53694 , n4324 , n53693 );
buf ( n4374 , n53518 );
buf ( n53696 , n53571 );
buf ( n53697 , n53391 );
xor ( n53698 , n53696 , n53697 );
buf ( n53699 , n53588 );
xor ( n4379 , n53698 , n53699 );
buf ( n53701 , n4379 );
buf ( n4381 , n53701 );
xor ( n4382 , n4374 , n4381 );
buf ( n53704 , n53410 );
buf ( n53705 , n389 );
not ( n53706 , n53705 );
buf ( n53707 , n53706 );
buf ( n53708 , n53707 );
nor ( n53709 , n53704 , n53708 );
buf ( n53710 , n53709 );
buf ( n53711 , n53710 );
xor ( n4391 , n4382 , n53711 );
buf ( n53713 , n4391 );
buf ( n53714 , n53713 );
xor ( n4394 , n53694 , n53714 );
buf ( n53716 , n4394 );
buf ( n53717 , n53716 );
xor ( n4397 , n53644 , n53717 );
buf ( n53719 , n53548 );
xor ( n4399 , n4397 , n53719 );
buf ( n53721 , n4399 );
buf ( n53722 , n53721 );
xor ( n4402 , n53628 , n53629 );
xor ( n4403 , n4402 , n53722 );
buf ( n53725 , n4403 );
xor ( n4405 , n53628 , n53629 );
and ( n4406 , n4405 , n53722 );
and ( n4407 , n53628 , n53629 );
or ( n4408 , n4406 , n4407 );
buf ( n53730 , n4408 );
xor ( n4410 , n53696 , n53697 );
and ( n4411 , n4410 , n53699 );
and ( n4412 , n53696 , n53697 );
or ( n4413 , n4411 , n4412 );
buf ( n53735 , n4413 );
xor ( n4415 , n53600 , n53605 );
and ( n4416 , n4415 , n53610 );
and ( n4417 , n53600 , n53605 );
or ( n53739 , n4416 , n4417 );
buf ( n53740 , n53739 );
xor ( n4420 , n4374 , n4381 );
and ( n53742 , n4420 , n53711 );
and ( n53743 , n4374 , n4381 );
or ( n4423 , n53742 , n53743 );
buf ( n53745 , n4423 );
xor ( n53746 , n4274 , n53613 );
and ( n4426 , n53746 , n53620 );
and ( n53748 , n4274 , n53613 );
or ( n4428 , n4426 , n53748 );
buf ( n53750 , n4428 );
xor ( n53751 , n53630 , n53635 );
and ( n4431 , n53751 , n53641 );
and ( n4432 , n53630 , n53635 );
or ( n53754 , n4431 , n4432 );
buf ( n53755 , n53754 );
xor ( n4435 , n4324 , n53693 );
and ( n4436 , n4435 , n53714 );
and ( n4437 , n4324 , n53693 );
or ( n53759 , n4436 , n4437 );
buf ( n53760 , n53759 );
xor ( n4440 , n53594 , n53623 );
and ( n4441 , n4440 , n53625 );
and ( n4442 , n53594 , n53623 );
or ( n53764 , n4441 , n4442 );
buf ( n53765 , n53764 );
xor ( n4445 , n53644 , n53717 );
and ( n4446 , n4445 , n53719 );
and ( n4447 , n53644 , n53717 );
or ( n53769 , n4446 , n4447 );
buf ( n53770 , n53769 );
buf ( n53771 , n402 );
buf ( n53772 , n412 );
and ( n4452 , n53771 , n53772 );
buf ( n53774 , n4452 );
buf ( n53775 , n53774 );
buf ( n53776 , n403 );
buf ( n53777 , n411 );
and ( n4457 , n53776 , n53777 );
buf ( n53779 , n4457 );
buf ( n53780 , n53779 );
buf ( n53781 , n404 );
buf ( n53782 , n410 );
and ( n4462 , n53781 , n53782 );
buf ( n53784 , n4462 );
buf ( n53785 , n53784 );
xor ( n4465 , n53775 , n53780 );
xor ( n4466 , n4465 , n53785 );
buf ( n53788 , n4466 );
xor ( n53789 , n53775 , n53780 );
and ( n4469 , n53789 , n53785 );
and ( n4470 , n53775 , n53780 );
or ( n4471 , n4469 , n4470 );
buf ( n53793 , n4471 );
buf ( n53794 , n53576 );
buf ( n53795 , n53788 );
buf ( n53796 , n53593 );
xor ( n4476 , n53794 , n53795 );
xor ( n4477 , n4476 , n53796 );
buf ( n53799 , n4477 );
xor ( n53800 , n53794 , n53795 );
and ( n53801 , n53800 , n53796 );
and ( n4481 , n53794 , n53795 );
or ( n53803 , n53801 , n4481 );
buf ( n53804 , n53803 );
buf ( n4484 , n52432 );
buf ( n4485 , n386 );
and ( n4486 , n4484 , n4485 );
buf ( n4487 , n4486 );
buf ( n53809 , n4487 );
buf ( n4489 , n3294 );
buf ( n4490 , n387 );
and ( n4491 , n4489 , n4490 );
buf ( n4492 , n4491 );
buf ( n53814 , n4492 );
buf ( n53815 , n53735 );
xor ( n4495 , n53809 , n53814 );
xor ( n53817 , n4495 , n53815 );
buf ( n53818 , n53817 );
xor ( n4498 , n53809 , n53814 );
and ( n4499 , n4498 , n53815 );
and ( n4500 , n53809 , n53814 );
or ( n53822 , n4499 , n4500 );
buf ( n53823 , n53822 );
buf ( n53824 , n53799 );
buf ( n53825 , n3415 );
buf ( n53826 , n388 );
and ( n53827 , n53825 , n53826 );
buf ( n53828 , n53827 );
buf ( n53829 , n53828 );
buf ( n53830 , n53740 );
xor ( n53831 , n53824 , n53829 );
xor ( n4511 , n53831 , n53830 );
buf ( n53833 , n4511 );
xor ( n53834 , n53824 , n53829 );
and ( n4514 , n53834 , n53830 );
and ( n4515 , n53824 , n53829 );
or ( n4516 , n4514 , n4515 );
buf ( n53838 , n4516 );
buf ( n53839 , n53184 );
not ( n53840 , n53839 );
buf ( n53841 , n53707 );
nor ( n53842 , n53840 , n53841 );
buf ( n53843 , n53842 );
buf ( n53844 , n53843 );
buf ( n53845 , n53818 );
buf ( n4525 , n53251 );
buf ( n53847 , n390 );
and ( n53848 , n4525 , n53847 );
buf ( n53849 , n53848 );
buf ( n53850 , n53849 );
xor ( n53851 , n53844 , n53845 );
xor ( n4531 , n53851 , n53850 );
buf ( n53853 , n4531 );
xor ( n53854 , n53844 , n53845 );
and ( n4534 , n53854 , n53850 );
and ( n53856 , n53844 , n53845 );
or ( n53857 , n4534 , n53856 );
buf ( n53858 , n53857 );
buf ( n53859 , n53745 );
buf ( n53860 , n53639 );
buf ( n53861 , n391 );
and ( n4541 , n53860 , n53861 );
buf ( n53863 , n4541 );
buf ( n53864 , n53863 );
buf ( n53865 , n53833 );
xor ( n53866 , n53859 , n53864 );
xor ( n4546 , n53866 , n53865 );
buf ( n53868 , n4546 );
xor ( n4548 , n53859 , n53864 );
and ( n53870 , n4548 , n53865 );
and ( n53871 , n53859 , n53864 );
or ( n53872 , n53870 , n53871 );
buf ( n53873 , n53872 );
buf ( n4553 , n53750 );
nand ( n53875 , n4347 , n53666 );
not ( n4555 , n53875 );
not ( n53877 , n4342 );
or ( n53878 , n4555 , n53877 );
not ( n4558 , n53666 );
nand ( n53880 , n4558 , n53669 );
nand ( n53881 , n53878 , n53880 );
and ( n4561 , n386 , n389 );
xor ( n53883 , n387 , n4561 );
and ( n53884 , n387 , n388 );
xor ( n4564 , n53883 , n53884 );
nor ( n53886 , n53881 , n4564 );
not ( n53887 , n53886 );
nand ( n53888 , n4564 , n53881 );
nand ( n4568 , n53887 , n53888 );
not ( n4569 , n4568 );
and ( n4570 , n4337 , n53686 );
nor ( n4571 , n4570 , n53684 );
not ( n4572 , n4571 );
not ( n4573 , n4572 );
or ( n4574 , n4569 , n4573 );
not ( n4575 , n4568 );
nand ( n4576 , n4575 , n4571 );
nand ( n4577 , n4574 , n4576 );
buf ( n53899 , n4577 );
buf ( n53900 , n393 );
and ( n4580 , n53899 , n53900 );
buf ( n53902 , n4580 );
buf ( n53903 , n53902 );
not ( n4583 , n53691 );
buf ( n53905 , n4583 );
buf ( n53906 , n53237 );
nor ( n4586 , n53905 , n53906 );
buf ( n53908 , n4586 );
buf ( n53909 , n53908 );
xor ( n4589 , n4553 , n53903 );
xor ( n4590 , n4589 , n53909 );
buf ( n53912 , n4590 );
xor ( n4592 , n4553 , n53903 );
and ( n4593 , n4592 , n53909 );
and ( n4594 , n4553 , n53903 );
or ( n4595 , n4593 , n4594 );
buf ( n53917 , n4595 );
buf ( n53918 , n53853 );
buf ( n53919 , n53755 );
buf ( n53920 , n53760 );
xor ( n4600 , n53918 , n53919 );
xor ( n4601 , n4600 , n53920 );
buf ( n53923 , n4601 );
xor ( n4603 , n53918 , n53919 );
and ( n4604 , n4603 , n53920 );
and ( n4605 , n53918 , n53919 );
or ( n4606 , n4604 , n4605 );
buf ( n53928 , n4606 );
buf ( n4608 , n53868 );
buf ( n4609 , n53912 );
buf ( n53931 , n53765 );
xor ( n53932 , n4608 , n4609 );
xor ( n53933 , n53932 , n53931 );
buf ( n53934 , n53933 );
xor ( n53935 , n4608 , n4609 );
and ( n53936 , n53935 , n53931 );
and ( n53937 , n4608 , n4609 );
or ( n4617 , n53936 , n53937 );
buf ( n53939 , n4617 );
buf ( n53940 , n53923 );
buf ( n53941 , n53770 );
buf ( n53942 , n53934 );
xor ( n4622 , n53940 , n53941 );
xor ( n53944 , n4622 , n53942 );
buf ( n53945 , n53944 );
xor ( n4625 , n53940 , n53941 );
and ( n53947 , n4625 , n53942 );
and ( n53948 , n53940 , n53941 );
or ( n4628 , n53947 , n53948 );
buf ( n53950 , n4628 );
buf ( n53951 , n402 );
buf ( n53952 , n411 );
and ( n53953 , n53951 , n53952 );
buf ( n53954 , n53953 );
buf ( n53955 , n53954 );
buf ( n53956 , n403 );
buf ( n53957 , n410 );
and ( n53958 , n53956 , n53957 );
buf ( n53959 , n53958 );
buf ( n53960 , n53959 );
buf ( n53961 , n53793 );
xor ( n53962 , n53955 , n53960 );
xor ( n4642 , n53962 , n53961 );
buf ( n53964 , n4642 );
xor ( n4644 , n53955 , n53960 );
and ( n4645 , n4644 , n53961 );
and ( n53967 , n53955 , n53960 );
or ( n4647 , n4645 , n53967 );
buf ( n53969 , n4647 );
buf ( n53970 , n53964 );
buf ( n53971 , n3294 );
buf ( n53972 , n386 );
and ( n4652 , n53971 , n53972 );
buf ( n53974 , n4652 );
buf ( n53975 , n53974 );
buf ( n53976 , n53804 );
xor ( n53977 , n53970 , n53975 );
xor ( n4657 , n53977 , n53976 );
buf ( n53979 , n4657 );
xor ( n4659 , n53970 , n53975 );
and ( n4660 , n4659 , n53976 );
and ( n53982 , n53970 , n53975 );
or ( n4662 , n4660 , n53982 );
buf ( n53984 , n4662 );
buf ( n53985 , n3415 );
buf ( n53986 , n387 );
and ( n53987 , n53985 , n53986 );
buf ( n53988 , n53987 );
buf ( n53989 , n53988 );
buf ( n53990 , n53184 );
buf ( n53991 , n388 );
and ( n53992 , n53990 , n53991 );
buf ( n53993 , n53992 );
buf ( n53994 , n53993 );
buf ( n53995 , n53823 );
xor ( n4675 , n53989 , n53994 );
xor ( n53997 , n4675 , n53995 );
buf ( n53998 , n53997 );
xor ( n4678 , n53989 , n53994 );
and ( n4679 , n4678 , n53995 );
and ( n4680 , n53989 , n53994 );
or ( n54002 , n4679 , n4680 );
buf ( n54003 , n54002 );
buf ( n54004 , n53248 );
buf ( n54005 , n389 );
and ( n4685 , n54004 , n54005 );
buf ( n54007 , n4685 );
buf ( n4687 , n54007 );
buf ( n4688 , n53979 );
buf ( n54010 , n4172 );
buf ( n54011 , n390 );
and ( n54012 , n54010 , n54011 );
buf ( n54013 , n54012 );
buf ( n54014 , n54013 );
xor ( n4694 , n4687 , n4688 );
xor ( n54016 , n4694 , n54014 );
buf ( n54017 , n54016 );
xor ( n54018 , n4687 , n4688 );
and ( n54019 , n54018 , n54014 );
and ( n4699 , n4687 , n4688 );
or ( n54021 , n54019 , n4699 );
buf ( n54022 , n54021 );
and ( n4702 , n4577 , n392 );
buf ( n54024 , n4702 );
not ( n54025 , n53688 );
nand ( n4705 , n54025 , n53690 );
buf ( n54027 , n4705 );
buf ( n54028 , n391 );
and ( n4708 , n54027 , n54028 );
buf ( n54030 , n4708 );
buf ( n54031 , n54030 );
buf ( n54032 , n53838 );
xor ( n54033 , n54024 , n54031 );
xor ( n4713 , n54033 , n54032 );
buf ( n54035 , n4713 );
xor ( n54036 , n54024 , n54031 );
and ( n4716 , n54036 , n54032 );
and ( n4717 , n54024 , n54031 );
or ( n4718 , n4716 , n4717 );
buf ( n54040 , n4718 );
buf ( n54041 , n53998 );
buf ( n54042 , n53858 );
not ( n54043 , n53886 );
not ( n4723 , n54043 );
not ( n54045 , n4572 );
or ( n54046 , n4723 , n54045 );
nand ( n54047 , n54046 , n53888 );
xor ( n54048 , n387 , n4561 );
and ( n4728 , n54048 , n53884 );
and ( n54050 , n387 , n4561 );
or ( n54051 , n4728 , n54050 );
and ( n54052 , n386 , n388 );
nor ( n4732 , n54051 , n54052 );
not ( n4733 , n4732 );
nand ( n54055 , n54051 , n54052 );
nand ( n4735 , n4733 , n54055 );
xnor ( n4736 , n54047 , n4735 );
buf ( n54058 , n4736 );
buf ( n4738 , n54058 );
buf ( n54060 , n4738 );
and ( n54061 , n54060 , n393 );
buf ( n54062 , n54061 );
xor ( n54063 , n54041 , n54042 );
xor ( n4743 , n54063 , n54062 );
buf ( n54065 , n4743 );
xor ( n54066 , n54041 , n54042 );
and ( n54067 , n54066 , n54062 );
and ( n4747 , n54041 , n54042 );
or ( n4748 , n54067 , n4747 );
buf ( n54070 , n4748 );
buf ( n54071 , n54017 );
buf ( n54072 , n53917 );
buf ( n54073 , n53873 );
xor ( n4753 , n54071 , n54072 );
xor ( n54075 , n4753 , n54073 );
buf ( n54076 , n54075 );
xor ( n54077 , n54071 , n54072 );
and ( n54078 , n54077 , n54073 );
and ( n54079 , n54071 , n54072 );
or ( n54080 , n54078 , n54079 );
buf ( n54081 , n54080 );
buf ( n54082 , n54035 );
buf ( n54083 , n54065 );
buf ( n54084 , n53928 );
xor ( n4764 , n54082 , n54083 );
xor ( n54086 , n4764 , n54084 );
buf ( n54087 , n54086 );
xor ( n4767 , n54082 , n54083 );
and ( n4768 , n4767 , n54084 );
and ( n4769 , n54082 , n54083 );
or ( n54091 , n4768 , n4769 );
buf ( n54092 , n54091 );
buf ( n54093 , n54076 );
buf ( n4773 , n53939 );
buf ( n4774 , n54087 );
xor ( n4775 , n54093 , n4773 );
xor ( n4776 , n4775 , n4774 );
buf ( n4777 , n4776 );
xor ( n4778 , n54093 , n4773 );
and ( n4779 , n4778 , n4774 );
and ( n4780 , n54093 , n4773 );
or ( n4781 , n4779 , n4780 );
buf ( n4782 , n4781 );
buf ( n4783 , n402 );
buf ( n54105 , n410 );
and ( n4785 , n4783 , n54105 );
buf ( n54107 , n4785 );
buf ( n54108 , n54107 );
buf ( n54109 , n53969 );
buf ( n54110 , n386 );
not ( n4790 , n54110 );
buf ( n54112 , n3416 );
nor ( n4792 , n4790 , n54112 );
buf ( n54114 , n4792 );
buf ( n54115 , n54114 );
xor ( n4795 , n54108 , n54109 );
xor ( n4796 , n4795 , n54115 );
buf ( n54118 , n4796 );
xor ( n4798 , n54108 , n54109 );
and ( n4799 , n4798 , n54115 );
and ( n4800 , n54108 , n54109 );
or ( n4801 , n4799 , n4800 );
buf ( n54123 , n4801 );
not ( n4803 , n53023 );
nor ( n4804 , n4803 , n53398 );
buf ( n54126 , n4804 );
and ( n4806 , n53248 , n388 );
buf ( n54128 , n4806 );
buf ( n54129 , n53984 );
xor ( n4809 , n54126 , n54128 );
xor ( n4810 , n4809 , n54129 );
buf ( n54132 , n4810 );
xor ( n4812 , n54126 , n54128 );
and ( n54134 , n4812 , n54129 );
and ( n54135 , n54126 , n54128 );
or ( n54136 , n54134 , n54135 );
buf ( n54137 , n54136 );
buf ( n54138 , n54118 );
buf ( n4818 , n53639 );
buf ( n54140 , n389 );
and ( n54141 , n4818 , n54140 );
buf ( n54142 , n54141 );
buf ( n54143 , n54142 );
buf ( n54144 , n53691 );
buf ( n4824 , n390 );
and ( n4825 , n54144 , n4824 );
buf ( n4826 , n4825 );
buf ( n4827 , n4826 );
xor ( n4828 , n54138 , n54143 );
xor ( n4829 , n4828 , n4827 );
buf ( n4830 , n4829 );
xor ( n4831 , n54138 , n54143 );
and ( n4832 , n4831 , n4827 );
and ( n4833 , n54138 , n54143 );
or ( n4834 , n4832 , n4833 );
buf ( n4835 , n4834 );
and ( n54157 , n4577 , n391 );
buf ( n54158 , n54157 );
nor ( n54159 , n53886 , n4732 );
not ( n4839 , n54159 );
not ( n4840 , n4572 );
or ( n54162 , n4839 , n4840 );
or ( n4842 , n53888 , n4732 );
nand ( n4843 , n4842 , n54055 );
not ( n4844 , n4843 );
nand ( n4845 , n54162 , n4844 );
not ( n54167 , n4845 );
nor ( n54168 , n53238 , n387 );
not ( n54169 , n54168 );
nand ( n54170 , n54167 , n54169 );
nand ( n4850 , n4845 , n54168 );
nand ( n4851 , n54170 , n4850 , n393 );
buf ( n54173 , n4851 );
not ( n4853 , n54173 );
buf ( n54175 , n4853 );
buf ( n54176 , n54175 );
buf ( n54177 , n54003 );
xor ( n54178 , n54158 , n54176 );
xor ( n54179 , n54178 , n54177 );
buf ( n54180 , n54179 );
xor ( n54181 , n54158 , n54176 );
and ( n4861 , n54181 , n54177 );
and ( n4862 , n54158 , n54176 );
or ( n54184 , n4861 , n4862 );
buf ( n54185 , n54184 );
buf ( n54186 , n54022 );
and ( n4866 , n54060 , n392 );
buf ( n54188 , n4866 );
buf ( n54189 , n54132 );
xor ( n54190 , n54186 , n54188 );
xor ( n54191 , n54190 , n54189 );
buf ( n54192 , n54191 );
xor ( n54193 , n54186 , n54188 );
and ( n54194 , n54193 , n54189 );
and ( n54195 , n54186 , n54188 );
or ( n54196 , n54194 , n54195 );
buf ( n54197 , n54196 );
buf ( n54198 , n54040 );
buf ( n4878 , n4830 );
buf ( n54200 , n54070 );
xor ( n4880 , n54198 , n4878 );
xor ( n4881 , n4880 , n54200 );
buf ( n4882 , n4881 );
xor ( n4883 , n54198 , n4878 );
and ( n4884 , n4883 , n54200 );
and ( n4885 , n54198 , n4878 );
or ( n4886 , n4884 , n4885 );
buf ( n4887 , n4886 );
buf ( n4888 , n54180 );
buf ( n54210 , n54192 );
buf ( n54211 , n54081 );
xor ( n4891 , n4888 , n54210 );
xor ( n54213 , n4891 , n54211 );
buf ( n54214 , n54213 );
xor ( n54215 , n4888 , n54210 );
and ( n4895 , n54215 , n54211 );
and ( n4896 , n4888 , n54210 );
or ( n54218 , n4895 , n4896 );
buf ( n54219 , n54218 );
buf ( n54220 , n4882 );
buf ( n54221 , n54092 );
buf ( n54222 , n54214 );
xor ( n54223 , n54220 , n54221 );
xor ( n54224 , n54223 , n54222 );
buf ( n54225 , n54224 );
xor ( n4905 , n54220 , n54221 );
and ( n54227 , n4905 , n54222 );
and ( n54228 , n54220 , n54221 );
or ( n4908 , n54227 , n54228 );
buf ( n54230 , n4908 );
buf ( n54231 , n53184 );
buf ( n54232 , n386 );
and ( n4912 , n54231 , n54232 );
buf ( n54234 , n4912 );
buf ( n54235 , n54234 );
buf ( n54236 , n53251 );
buf ( n54237 , n387 );
and ( n4917 , n54236 , n54237 );
buf ( n54239 , n4917 );
buf ( n54240 , n54239 );
buf ( n54241 , n4172 );
buf ( n54242 , n388 );
and ( n54243 , n54241 , n54242 );
buf ( n54244 , n54243 );
buf ( n54245 , n54244 );
xor ( n4925 , n54235 , n54240 );
xor ( n4926 , n4925 , n54245 );
buf ( n54248 , n4926 );
xor ( n4928 , n54235 , n54240 );
and ( n54250 , n4928 , n54245 );
and ( n54251 , n54235 , n54240 );
or ( n4931 , n54250 , n54251 );
buf ( n54253 , n4931 );
buf ( n54254 , n54123 );
buf ( n54255 , n4577 );
buf ( n54256 , n390 );
and ( n54257 , n54255 , n54256 );
buf ( n54258 , n54257 );
buf ( n54259 , n54258 );
buf ( n54260 , n4705 );
buf ( n54261 , n389 );
and ( n54262 , n54260 , n54261 );
buf ( n54263 , n54262 );
buf ( n54264 , n54263 );
xor ( n4944 , n54254 , n54259 );
xor ( n54266 , n4944 , n54264 );
buf ( n54267 , n54266 );
xor ( n54268 , n54254 , n54259 );
and ( n54269 , n54268 , n54264 );
and ( n4949 , n54254 , n54259 );
or ( n54271 , n54269 , n4949 );
buf ( n54272 , n54271 );
not ( n54273 , n54159 );
nor ( n4953 , n54273 , n53238 );
not ( n4954 , n4953 );
not ( n54276 , n4572 );
or ( n4956 , n4954 , n54276 );
or ( n4957 , n4843 , n387 );
nand ( n4958 , n4957 , n386 );
nand ( n4959 , n4956 , n4958 );
and ( n54281 , n4959 , n393 );
buf ( n4961 , n54281 );
buf ( n4962 , n54137 );
not ( n4963 , n54168 );
and ( n4964 , n4845 , n4963 );
not ( n4965 , n4845 );
not ( n4966 , n54169 );
and ( n4967 , n4965 , n4966 );
nor ( n4968 , n4964 , n4967 );
nor ( n4969 , n4968 , n53237 );
buf ( n54291 , n4969 );
xor ( n4971 , n4961 , n4962 );
xor ( n4972 , n4971 , n54291 );
buf ( n54294 , n4972 );
xor ( n4974 , n4961 , n4962 );
and ( n4975 , n4974 , n54291 );
and ( n4976 , n4961 , n4962 );
or ( n4977 , n4975 , n4976 );
buf ( n54299 , n4977 );
buf ( n54300 , n54248 );
buf ( n54301 , n54060 );
buf ( n54302 , n391 );
and ( n4982 , n54301 , n54302 );
buf ( n54304 , n4982 );
buf ( n54305 , n54304 );
buf ( n54306 , n4835 );
xor ( n54307 , n54300 , n54305 );
xor ( n54308 , n54307 , n54306 );
buf ( n54309 , n54308 );
xor ( n54310 , n54300 , n54305 );
and ( n54311 , n54310 , n54306 );
and ( n4991 , n54300 , n54305 );
or ( n4992 , n54311 , n4991 );
buf ( n54314 , n4992 );
buf ( n54315 , n54185 );
buf ( n54316 , n54267 );
buf ( n54317 , n54294 );
xor ( n4997 , n54315 , n54316 );
xor ( n54319 , n4997 , n54317 );
buf ( n54320 , n54319 );
xor ( n54321 , n54315 , n54316 );
and ( n54322 , n54321 , n54317 );
and ( n5002 , n54315 , n54316 );
or ( n5003 , n54322 , n5002 );
buf ( n54325 , n5003 );
buf ( n54326 , n54197 );
buf ( n54327 , n54309 );
buf ( n54328 , n4887 );
xor ( n5008 , n54326 , n54327 );
xor ( n54330 , n5008 , n54328 );
buf ( n54331 , n54330 );
xor ( n54332 , n54326 , n54327 );
and ( n54333 , n54332 , n54328 );
and ( n5013 , n54326 , n54327 );
or ( n5014 , n54333 , n5013 );
buf ( n54336 , n5014 );
buf ( n54337 , n54320 );
buf ( n54338 , n54219 );
buf ( n54339 , n54331 );
xor ( n5019 , n54337 , n54338 );
xor ( n54341 , n5019 , n54339 );
buf ( n54342 , n54341 );
xor ( n54343 , n54337 , n54338 );
and ( n54344 , n54343 , n54339 );
and ( n5024 , n54337 , n54338 );
or ( n5025 , n54344 , n5024 );
buf ( n54347 , n5025 );
buf ( n54348 , n53251 );
buf ( n54349 , n386 );
and ( n5029 , n54348 , n54349 );
buf ( n54351 , n5029 );
buf ( n54352 , n54351 );
buf ( n5032 , n4172 );
buf ( n5033 , n387 );
and ( n5034 , n5032 , n5033 );
buf ( n5035 , n5034 );
buf ( n54357 , n5035 );
buf ( n54358 , n4959 );
buf ( n54359 , n392 );
and ( n5039 , n54358 , n54359 );
buf ( n54361 , n5039 );
buf ( n54362 , n54361 );
xor ( n54363 , n54352 , n54357 );
xor ( n54364 , n54363 , n54362 );
buf ( n54365 , n54364 );
xor ( n5045 , n54352 , n54357 );
and ( n54367 , n5045 , n54362 );
and ( n5047 , n54352 , n54357 );
or ( n5048 , n54367 , n5047 );
buf ( n54370 , n5048 );
buf ( n5050 , n4577 );
buf ( n54372 , n5050 );
buf ( n54373 , n389 );
and ( n5053 , n54372 , n54373 );
buf ( n54375 , n5053 );
buf ( n54376 , n54375 );
buf ( n54377 , n4705 );
buf ( n54378 , n388 );
and ( n54379 , n54377 , n54378 );
buf ( n54380 , n54379 );
buf ( n54381 , n54380 );
not ( n54382 , n4968 );
and ( n54383 , n54382 , n391 );
buf ( n5063 , n54383 );
xor ( n5064 , n54376 , n54381 );
xor ( n5065 , n5064 , n5063 );
buf ( n5066 , n5065 );
xor ( n5067 , n54376 , n54381 );
and ( n5068 , n5067 , n5063 );
and ( n5069 , n54376 , n54381 );
or ( n5070 , n5068 , n5069 );
buf ( n5071 , n5070 );
and ( n54393 , n4736 , n390 );
buf ( n5073 , n54393 );
buf ( n5074 , n54253 );
buf ( n54396 , n54272 );
xor ( n54397 , n5073 , n5074 );
xor ( n54398 , n54397 , n54396 );
buf ( n54399 , n54398 );
xor ( n5079 , n5073 , n5074 );
and ( n5080 , n5079 , n54396 );
and ( n5081 , n5073 , n5074 );
or ( n54403 , n5080 , n5081 );
buf ( n54404 , n54403 );
buf ( n54405 , n54365 );
buf ( n54406 , n54299 );
buf ( n5086 , n5066 );
xor ( n5087 , n54405 , n54406 );
xor ( n5088 , n5087 , n5086 );
buf ( n5089 , n5088 );
xor ( n5090 , n54405 , n54406 );
and ( n5091 , n5090 , n5086 );
and ( n5092 , n54405 , n54406 );
or ( n5093 , n5091 , n5092 );
buf ( n5094 , n5093 );
buf ( n5095 , n54399 );
buf ( n5096 , n54314 );
buf ( n54418 , n54325 );
xor ( n54419 , n5095 , n5096 );
xor ( n54420 , n54419 , n54418 );
buf ( n54421 , n54420 );
xor ( n5101 , n5095 , n5096 );
and ( n5102 , n5101 , n54418 );
and ( n5103 , n5095 , n5096 );
or ( n5104 , n5102 , n5103 );
buf ( n54426 , n5104 );
buf ( n54427 , n5089 );
buf ( n54428 , n54421 );
buf ( n54429 , n54336 );
xor ( n5109 , n54427 , n54428 );
xor ( n5110 , n5109 , n54429 );
buf ( n54432 , n5110 );
xor ( n5112 , n54427 , n54428 );
and ( n5113 , n5112 , n54429 );
and ( n5114 , n54427 , n54428 );
or ( n5115 , n5113 , n5114 );
buf ( n54437 , n5115 );
buf ( n54438 , n53639 );
buf ( n54439 , n386 );
and ( n5119 , n54438 , n54439 );
buf ( n54441 , n5119 );
buf ( n54442 , n54441 );
buf ( n54443 , n5050 );
buf ( n5123 , n388 );
and ( n54445 , n54443 , n5123 );
buf ( n54446 , n54445 );
buf ( n54447 , n54446 );
and ( n54448 , n53691 , n387 );
buf ( n54449 , n54448 );
xor ( n5129 , n54442 , n54447 );
xor ( n5130 , n5129 , n54449 );
buf ( n54452 , n5130 );
xor ( n54453 , n54442 , n54447 );
and ( n54454 , n54453 , n54449 );
and ( n5134 , n54442 , n54447 );
or ( n54456 , n54454 , n5134 );
buf ( n54457 , n54456 );
buf ( n54458 , n4959 );
buf ( n5138 , n54458 );
buf ( n54460 , n5138 );
buf ( n54461 , n54460 );
buf ( n54462 , n391 );
and ( n5142 , n54461 , n54462 );
buf ( n54464 , n5142 );
buf ( n54465 , n54464 );
and ( n54466 , n54382 , n390 );
buf ( n5146 , n54466 );
and ( n54468 , n54060 , n389 );
buf ( n54469 , n54468 );
xor ( n5149 , n54465 , n5146 );
xor ( n54471 , n5149 , n54469 );
buf ( n54472 , n54471 );
xor ( n5152 , n54465 , n5146 );
and ( n5153 , n5152 , n54469 );
and ( n5154 , n54465 , n5146 );
or ( n54476 , n5153 , n5154 );
buf ( n54477 , n54476 );
buf ( n54478 , n54370 );
buf ( n54479 , n5071 );
buf ( n54480 , n54452 );
xor ( n5160 , n54478 , n54479 );
xor ( n54482 , n5160 , n54480 );
buf ( n54483 , n54482 );
xor ( n5163 , n54478 , n54479 );
and ( n5164 , n5163 , n54480 );
and ( n5165 , n54478 , n54479 );
or ( n54487 , n5164 , n5165 );
buf ( n54488 , n54487 );
buf ( n54489 , n54472 );
buf ( n54490 , n54404 );
buf ( n54491 , n5094 );
xor ( n5171 , n54489 , n54490 );
xor ( n54493 , n5171 , n54491 );
buf ( n54494 , n54493 );
xor ( n5174 , n54489 , n54490 );
and ( n5175 , n5174 , n54491 );
and ( n5176 , n54489 , n54490 );
or ( n54498 , n5175 , n5176 );
buf ( n54499 , n54498 );
buf ( n5179 , n54483 );
buf ( n54501 , n54494 );
buf ( n54502 , n54426 );
xor ( n5182 , n5179 , n54501 );
xor ( n54504 , n5182 , n54502 );
buf ( n54505 , n54504 );
xor ( n54506 , n5179 , n54501 );
and ( n54507 , n54506 , n54502 );
and ( n5187 , n5179 , n54501 );
or ( n54509 , n54507 , n5187 );
buf ( n54510 , n54509 );
buf ( n54511 , n54460 );
buf ( n54512 , n390 );
and ( n54513 , n54511 , n54512 );
buf ( n54514 , n54513 );
buf ( n54515 , n54514 );
buf ( n54516 , n386 );
not ( n5196 , n54516 );
buf ( n54518 , n4583 );
nor ( n54519 , n5196 , n54518 );
buf ( n54520 , n54519 );
buf ( n5200 , n54520 );
buf ( n54522 , n5050 );
buf ( n54523 , n387 );
and ( n54524 , n54522 , n54523 );
buf ( n54525 , n54524 );
buf ( n54526 , n54525 );
xor ( n54527 , n54515 , n5200 );
xor ( n54528 , n54527 , n54526 );
buf ( n54529 , n54528 );
xor ( n5209 , n54515 , n5200 );
and ( n54531 , n5209 , n54526 );
and ( n54532 , n54515 , n5200 );
or ( n5212 , n54531 , n54532 );
buf ( n54534 , n5212 );
not ( n54535 , n4968 );
and ( n5215 , n54535 , n389 );
buf ( n54537 , n5215 );
and ( n5217 , n54060 , n388 );
buf ( n54539 , n5217 );
buf ( n54540 , n54457 );
xor ( n5220 , n54537 , n54539 );
xor ( n5221 , n5220 , n54540 );
buf ( n54543 , n5221 );
xor ( n5223 , n54537 , n54539 );
and ( n5224 , n5223 , n54540 );
and ( n5225 , n54537 , n54539 );
or ( n5226 , n5224 , n5225 );
buf ( n54548 , n5226 );
buf ( n54549 , n54529 );
buf ( n54550 , n54477 );
buf ( n54551 , n54543 );
xor ( n5231 , n54549 , n54550 );
xor ( n54553 , n5231 , n54551 );
buf ( n54554 , n54553 );
xor ( n54555 , n54549 , n54550 );
and ( n5235 , n54555 , n54551 );
and ( n5236 , n54549 , n54550 );
or ( n54558 , n5235 , n5236 );
buf ( n54559 , n54558 );
buf ( n54560 , n54488 );
buf ( n54561 , n54554 );
buf ( n54562 , n54499 );
xor ( n5242 , n54560 , n54561 );
xor ( n5243 , n5242 , n54562 );
buf ( n54565 , n5243 );
xor ( n54566 , n54560 , n54561 );
and ( n54567 , n54566 , n54562 );
and ( n54568 , n54560 , n54561 );
or ( n54569 , n54567 , n54568 );
buf ( n54570 , n54569 );
buf ( n54571 , n54460 );
buf ( n5251 , n389 );
and ( n54573 , n54571 , n5251 );
buf ( n54574 , n54573 );
buf ( n54575 , n54574 );
buf ( n54576 , n5050 );
buf ( n54577 , n386 );
and ( n5257 , n54576 , n54577 );
buf ( n54579 , n5257 );
buf ( n54580 , n54579 );
buf ( n54581 , n54535 );
buf ( n54582 , n388 );
and ( n54583 , n54581 , n54582 );
buf ( n54584 , n54583 );
buf ( n54585 , n54584 );
xor ( n5265 , n54575 , n54580 );
xor ( n54587 , n5265 , n54585 );
buf ( n54588 , n54587 );
xor ( n5268 , n54575 , n54580 );
and ( n5269 , n5268 , n54585 );
and ( n5270 , n54575 , n54580 );
or ( n54592 , n5269 , n5270 );
buf ( n54593 , n54592 );
buf ( n54594 , n54060 );
buf ( n54595 , n387 );
and ( n5275 , n54594 , n54595 );
buf ( n54597 , n5275 );
buf ( n54598 , n54597 );
buf ( n54599 , n54534 );
buf ( n54600 , n54588 );
xor ( n5280 , n54598 , n54599 );
xor ( n5281 , n5280 , n54600 );
buf ( n54603 , n5281 );
xor ( n54604 , n54598 , n54599 );
and ( n54605 , n54604 , n54600 );
and ( n54606 , n54598 , n54599 );
or ( n5286 , n54605 , n54606 );
buf ( n54608 , n5286 );
buf ( n54609 , n54548 );
buf ( n54610 , n54603 );
buf ( n54611 , n54559 );
xor ( n5291 , n54609 , n54610 );
xor ( n5292 , n5291 , n54611 );
buf ( n54614 , n5292 );
xor ( n54615 , n54609 , n54610 );
and ( n54616 , n54615 , n54611 );
and ( n5296 , n54609 , n54610 );
or ( n54618 , n54616 , n5296 );
buf ( n54619 , n54618 );
buf ( n5299 , n54460 );
buf ( n5300 , n388 );
and ( n5301 , n5299 , n5300 );
buf ( n5302 , n5301 );
buf ( n54624 , n5302 );
buf ( n5304 , n54535 );
buf ( n5305 , n387 );
and ( n5306 , n5304 , n5305 );
buf ( n5307 , n5306 );
buf ( n54629 , n5307 );
buf ( n54630 , n54060 );
buf ( n54631 , n386 );
and ( n54632 , n54630 , n54631 );
buf ( n54633 , n54632 );
buf ( n54634 , n54633 );
xor ( n5314 , n54624 , n54629 );
xor ( n5315 , n5314 , n54634 );
buf ( n54637 , n5315 );
xor ( n54638 , n54624 , n54629 );
and ( n54639 , n54638 , n54634 );
and ( n5319 , n54624 , n54629 );
or ( n54641 , n54639 , n5319 );
buf ( n54642 , n54641 );
buf ( n5322 , n54593 );
buf ( n5323 , n54637 );
buf ( n54645 , n54608 );
xor ( n54646 , n5322 , n5323 );
xor ( n54647 , n54646 , n54645 );
buf ( n54648 , n54647 );
xor ( n5328 , n5322 , n5323 );
and ( n5329 , n5328 , n54645 );
and ( n5330 , n5322 , n5323 );
or ( n5331 , n5329 , n5330 );
buf ( n54653 , n5331 );
buf ( n54654 , n54460 );
not ( n54655 , n54654 );
buf ( n54656 , n53398 );
nor ( n54657 , n54655 , n54656 );
buf ( n54658 , n54657 );
buf ( n54659 , n54658 );
buf ( n54660 , n54535 );
buf ( n54661 , n386 );
and ( n5341 , n54660 , n54661 );
buf ( n54663 , n5341 );
buf ( n54664 , n54663 );
buf ( n54665 , n54642 );
xor ( n54666 , n54659 , n54664 );
xor ( n5346 , n54666 , n54665 );
buf ( n54668 , n5346 );
xor ( n54669 , n54659 , n54664 );
and ( n54670 , n54669 , n54665 );
and ( n5350 , n54659 , n54664 );
or ( n5351 , n54670 , n5350 );
buf ( n54673 , n5351 );
buf ( n54674 , n54347 );
buf ( n54675 , n54432 );
nor ( n5355 , n54674 , n54675 );
buf ( n54677 , n5355 );
buf ( n54678 , n54677 );
nand ( n54679 , n54342 , n54230 );
buf ( n5359 , n54679 );
nor ( n54681 , n54678 , n5359 );
buf ( n54682 , n54681 );
buf ( n54683 , n54437 );
buf ( n54684 , n54505 );
nor ( n5364 , n54683 , n54684 );
buf ( n54686 , n5364 );
buf ( n54687 , n54686 );
not ( n5367 , n54687 );
buf ( n54689 , n5367 );
buf ( n5369 , n54689 );
buf ( n54691 , n54437 );
buf ( n54692 , n54505 );
nand ( n5372 , n54691 , n54692 );
buf ( n54694 , n5372 );
buf ( n54695 , n54694 );
nand ( n5375 , n5369 , n54695 );
buf ( n54697 , n5375 );
buf ( n54698 , n54689 );
buf ( n54699 , n54694 );
nand ( n54700 , n54698 , n54699 );
buf ( n54701 , n54700 );
buf ( n54702 , n54679 );
buf ( n54703 , n54432 );
buf ( n54704 , n54703 );
buf ( n54705 , n54347 );
nand ( n54706 , n54704 , n54705 );
buf ( n54707 , n54706 );
buf ( n54708 , n54707 );
nand ( n5388 , n54702 , n54708 );
buf ( n54710 , n5388 );
buf ( n54711 , n54686 );
buf ( n54712 , n54677 );
nor ( n54713 , n54711 , n54712 );
buf ( n54714 , n54713 );
buf ( n54715 , n54510 );
buf ( n54716 , n54565 );
nor ( n54717 , n54715 , n54716 );
buf ( n54718 , n54717 );
buf ( n54719 , n54437 );
buf ( n54720 , n54505 );
nand ( n54721 , n54719 , n54720 );
buf ( n54722 , n54721 );
buf ( n54723 , n54432 );
buf ( n54724 , n54347 );
nand ( n5404 , n54723 , n54724 );
buf ( n5405 , n5404 );
buf ( n54727 , n54437 );
buf ( n54728 , n54505 );
nor ( n5408 , n54727 , n54728 );
buf ( n54730 , n5408 );
buf ( n54731 , n53945 );
buf ( n54732 , n53730 );
nor ( n54733 , n54731 , n54732 );
buf ( n54734 , n54733 );
buf ( n54735 , n53945 );
not ( n54736 , n54735 );
buf ( n54737 , n54736 );
buf ( n54738 , n53730 );
not ( n5418 , n54738 );
buf ( n54740 , n5418 );
buf ( n54741 , n53295 );
not ( n54742 , n54741 );
buf ( n54743 , n54742 );
not ( n54744 , n52644 );
not ( n54745 , n52457 );
and ( n54746 , n54744 , n54745 );
buf ( n54747 , n52171 );
buf ( n54748 , n52098 );
buf ( n54749 , n52093 );
xnor ( n5429 , n54748 , n54749 );
buf ( n54751 , n5429 );
buf ( n54752 , n54751 );
buf ( n54753 , n393 );
buf ( n54754 , n409 );
nand ( n54755 , n54753 , n54754 );
buf ( n54756 , n54755 );
buf ( n54757 , n54756 );
not ( n5437 , n54757 );
buf ( n54759 , n408 );
nand ( n5439 , n5437 , n54759 );
buf ( n54761 , n5439 );
buf ( n54762 , n54761 );
and ( n5442 , n54752 , n54762 );
buf ( n54764 , n408 );
not ( n54765 , n54764 );
buf ( n54766 , n54765 );
buf ( n54767 , n54766 );
not ( n5447 , n54767 );
buf ( n54769 , n54756 );
not ( n54770 , n54769 );
or ( n5450 , n5447 , n54770 );
buf ( n54772 , n417 );
nand ( n5452 , n5450 , n54772 );
buf ( n54774 , n5452 );
buf ( n54775 , n54774 );
nor ( n54776 , n5442 , n54775 );
buf ( n54777 , n54776 );
buf ( n54778 , n54777 );
not ( n5458 , n54778 );
buf ( n54780 , n52106 );
not ( n54781 , n54780 );
or ( n5461 , n5458 , n54781 );
buf ( n54783 , n52079 );
not ( n5463 , n54783 );
buf ( n54785 , n5463 );
buf ( n54786 , n54785 );
nand ( n54787 , n5461 , n54786 );
buf ( n54788 , n54787 );
buf ( n54789 , n54788 );
buf ( n54790 , n52106 );
buf ( n54791 , n54777 );
or ( n54792 , n54790 , n54791 );
buf ( n54793 , n54792 );
buf ( n54794 , n54793 );
and ( n5474 , n54747 , n54789 , n54794 );
buf ( n54796 , n5474 );
not ( n54797 , n54796 );
not ( n54798 , n52182 );
and ( n54799 , n54797 , n54798 );
buf ( n54800 , n54793 );
buf ( n54801 , n54788 );
and ( n54802 , n54800 , n54801 );
buf ( n54803 , n52171 );
nor ( n54804 , n54802 , n54803 );
buf ( n54805 , n54804 );
nor ( n54806 , n54799 , n54805 );
not ( n54807 , n54806 );
not ( n54808 , n52304 );
or ( n54809 , n54807 , n54808 );
buf ( n54810 , n52266 );
not ( n54811 , n54810 );
buf ( n54812 , n54811 );
nand ( n5492 , n54809 , n54812 );
or ( n5493 , n54806 , n52304 );
and ( n54815 , n5492 , n5493 , n52309 );
or ( n5495 , n52452 , n54815 );
not ( n5496 , n5493 );
not ( n5497 , n5492 );
or ( n5498 , n5496 , n5497 );
not ( n54820 , n52309 );
nand ( n54821 , n5498 , n54820 );
nand ( n54822 , n5495 , n54821 );
nor ( n5502 , n54746 , n54822 );
buf ( n54824 , n5502 );
buf ( n54825 , n52457 );
not ( n5505 , n54825 );
buf ( n54827 , n52644 );
not ( n54828 , n54827 );
or ( n5508 , n5505 , n54828 );
buf ( n54830 , n52649 );
not ( n54831 , n54830 );
buf ( n54832 , n54831 );
buf ( n54833 , n54832 );
nand ( n5513 , n5508 , n54833 );
buf ( n54835 , n5513 );
buf ( n54836 , n54835 );
or ( n54837 , n54824 , n54836 );
buf ( n54838 , n52821 );
nand ( n54839 , n54837 , n54838 );
buf ( n54840 , n54839 );
buf ( n54841 , n52644 );
buf ( n54842 , n52457 );
and ( n5522 , n54841 , n54842 );
buf ( n54844 , n5522 );
or ( n5524 , n5502 , n54844 );
nand ( n5525 , n5524 , n52649 );
nand ( n54847 , n54840 , n5525 );
buf ( n5527 , n54847 );
buf ( n5528 , n53059 );
nor ( n54850 , n5527 , n5528 );
buf ( n54851 , n54850 );
buf ( n54852 , n54851 );
not ( n54853 , n54852 );
buf ( n54854 , n54853 );
buf ( n54855 , n53064 );
not ( n5535 , n54855 );
buf ( n54857 , n5535 );
buf ( n54858 , n52826 );
not ( n54859 , n54858 );
buf ( n54860 , n54859 );
buf ( n54861 , n54460 );
buf ( n54862 , n386 );
nand ( n54863 , n54861 , n54862 );
buf ( n54864 , n54863 );
buf ( n54865 , n54225 );
not ( n5545 , n54865 );
buf ( n5546 , n5545 );
buf ( n54868 , n54510 );
buf ( n54869 , n54565 );
or ( n54870 , n54868 , n54869 );
buf ( n54871 , n54870 );
buf ( n54872 , n411 );
buf ( n54873 , n418 );
buf ( n54874 , n425 );
nand ( n5554 , n54873 , n54874 );
buf ( n54876 , n5554 );
buf ( n54877 , n54876 );
not ( n5557 , n54877 );
buf ( n54879 , n424 );
buf ( n54880 , n419 );
nand ( n54881 , n54879 , n54880 );
buf ( n54882 , n54881 );
buf ( n54883 , n54882 );
not ( n5563 , n54883 );
or ( n54885 , n5557 , n5563 );
buf ( n5565 , n418 );
buf ( n5566 , n421 );
xor ( n54888 , n5565 , n5566 );
buf ( n54889 , n54888 );
buf ( n54890 , n54889 );
nand ( n54891 , n54885 , n54890 );
buf ( n54892 , n54891 );
buf ( n54893 , n54892 );
buf ( n54894 , n54876 );
not ( n5574 , n54894 );
buf ( n54896 , n54882 );
not ( n54897 , n54896 );
buf ( n54898 , n54897 );
buf ( n54899 , n54898 );
nand ( n5579 , n5574 , n54899 );
buf ( n54901 , n5579 );
buf ( n54902 , n54901 );
nand ( n5582 , n54893 , n54902 );
buf ( n54904 , n5582 );
and ( n5584 , n420 , n422 );
not ( n5585 , n5584 );
and ( n54907 , n421 , n423 );
not ( n54908 , n54907 );
or ( n54909 , n5585 , n54908 );
not ( n5589 , n421 );
not ( n54911 , n422 );
or ( n54912 , n5589 , n54911 );
nand ( n54913 , n420 , n423 );
nand ( n54914 , n54912 , n54913 );
nand ( n5594 , n54909 , n54914 );
not ( n54916 , n5594 );
not ( n54917 , n370 );
nand ( n54918 , n54917 , n419 );
nand ( n54919 , n54916 , n54918 );
not ( n5599 , n54919 );
nand ( n54921 , n421 , n423 );
buf ( n54922 , n54921 );
not ( n5602 , n54922 );
nand ( n5603 , n424 , n420 );
buf ( n54925 , n5603 );
not ( n54926 , n54925 );
or ( n54927 , n5602 , n54926 );
nand ( n5605 , n419 , n425 );
not ( n5606 , n5605 );
buf ( n54930 , n5606 );
nand ( n54931 , n54927 , n54930 );
buf ( n54932 , n54931 );
buf ( n54933 , n54932 );
buf ( n54934 , n5603 );
not ( n5612 , n54934 );
buf ( n54936 , n54907 );
nand ( n5614 , n5612 , n54936 );
buf ( n54938 , n5614 );
buf ( n54939 , n54938 );
nand ( n5617 , n54933 , n54939 );
buf ( n54941 , n5617 );
not ( n54942 , n54941 );
or ( n54943 , n5599 , n54942 );
not ( n5621 , n54918 );
nand ( n54945 , n5621 , n5594 );
nand ( n54946 , n54943 , n54945 );
xor ( n54947 , n54904 , n54946 );
buf ( n54948 , n419 );
buf ( n54949 , n423 );
nand ( n54950 , n54948 , n54949 );
buf ( n54951 , n54950 );
not ( n54952 , n54951 );
not ( n5630 , n54914 );
not ( n5631 , n5630 );
or ( n54955 , n54952 , n5631 );
buf ( n54956 , n54951 );
not ( n54957 , n54956 );
buf ( n54958 , n54957 );
nand ( n5634 , n54914 , n54958 );
nand ( n54960 , n54955 , n5634 );
not ( n5636 , n424 );
nand ( n5637 , n5636 , n421 , n418 );
not ( n5638 , n421 );
nand ( n5639 , n5638 , n424 , n418 );
nand ( n5640 , n5637 , n5639 );
not ( n5641 , n5640 );
nand ( n5642 , n420 , n422 );
not ( n5643 , n5642 );
or ( n5644 , n5641 , n5643 );
not ( n5645 , n5642 );
nand ( n5646 , n5645 , n5637 , n5639 );
nand ( n5647 , n5644 , n5646 );
and ( n5648 , n54960 , n5647 );
not ( n5649 , n54960 );
not ( n5650 , n5647 );
and ( n5651 , n5649 , n5650 );
nor ( n5652 , n5648 , n5651 );
xor ( n5653 , n54947 , n5652 );
not ( n5654 , n5653 );
not ( n5655 , n54918 );
and ( n5656 , n5594 , n5655 );
not ( n5657 , n5594 );
and ( n5658 , n5657 , n54918 );
nor ( n5659 , n5656 , n5658 );
and ( n5660 , n5659 , n54941 );
not ( n5661 , n5659 );
not ( n5662 , n54941 );
and ( n5663 , n5661 , n5662 );
nor ( n5664 , n5660 , n5663 );
not ( n5665 , n5664 );
buf ( n54991 , n420 );
not ( n54992 , n54991 );
buf ( n54993 , n371 );
nor ( n54994 , n54992 , n54993 );
buf ( n54995 , n54994 );
or ( n5671 , n370 , n419 );
nand ( n5672 , n370 , n419 );
nand ( n54998 , n5671 , n5672 );
xor ( n5674 , n54995 , n54998 );
buf ( n55000 , n422 );
not ( n55001 , n55000 );
buf ( n55002 , n420 );
buf ( n55003 , n425 );
nand ( n5679 , n55002 , n55003 );
buf ( n55005 , n5679 );
buf ( n55006 , n55005 );
not ( n55007 , n55006 );
buf ( n55008 , n55007 );
buf ( n55009 , n55008 );
not ( n55010 , n55009 );
or ( n55011 , n55001 , n55010 );
buf ( n55012 , n422 );
buf ( n55013 , n423 );
nand ( n5689 , n55012 , n55013 );
buf ( n55015 , n5689 );
buf ( n55016 , n55015 );
nand ( n55017 , n55011 , n55016 );
buf ( n55018 , n55017 );
and ( n55019 , n5674 , n55018 );
and ( n5695 , n54995 , n54998 );
or ( n5696 , n55019 , n5695 );
xor ( n5697 , n54876 , n54898 );
xnor ( n55023 , n5697 , n54889 );
or ( n5699 , n5696 , n55023 );
not ( n55025 , n5699 );
or ( n55026 , n5665 , n55025 );
nand ( n5702 , n5696 , n55023 );
nand ( n55028 , n55026 , n5702 );
buf ( n55029 , n55028 );
not ( n55030 , n55029 );
buf ( n55031 , n55030 );
nand ( n55032 , n5654 , n55031 );
buf ( n55033 , n55032 );
not ( n55034 , n55033 );
buf ( n55035 , n55034 );
not ( n5711 , n55035 );
and ( n55037 , n418 , n421 );
not ( n5713 , n55037 );
nand ( n55039 , n424 , n418 );
not ( n5715 , n55039 );
not ( n55041 , n5715 );
or ( n55042 , n5713 , n55041 );
nand ( n55043 , n418 , n421 );
not ( n5719 , n55043 );
not ( n55045 , n55039 );
or ( n55046 , n5719 , n55045 );
nand ( n5722 , n55046 , n5584 );
nand ( n55048 , n55042 , n5722 );
not ( n5724 , n55048 );
not ( n55050 , n5630 );
not ( n5726 , n54958 );
or ( n5727 , n55050 , n5726 );
nand ( n55053 , n5727 , n5647 );
nand ( n5729 , n54914 , n54951 );
nand ( n55055 , n55053 , n5729 );
not ( n5731 , n55055 );
not ( n5732 , n5731 );
or ( n5733 , n5724 , n5732 );
not ( n5734 , n55048 );
nand ( n5735 , n5734 , n55055 );
nand ( n55061 , n5733 , n5735 );
xor ( n55062 , n420 , n54958 );
nand ( n5738 , n418 , n423 );
not ( n55064 , n5738 );
and ( n55065 , n419 , n422 );
xor ( n55066 , n55064 , n55065 );
nand ( n55067 , n420 , n421 );
and ( n5743 , n55066 , n55067 );
not ( n55069 , n55066 );
not ( n55070 , n55067 );
and ( n5746 , n55069 , n55070 );
nor ( n55072 , n5743 , n5746 );
xor ( n5748 , n55062 , n55072 );
and ( n55074 , n55061 , n5748 );
not ( n55075 , n55061 );
not ( n5751 , n5748 );
and ( n55077 , n55075 , n5751 );
nor ( n55078 , n55074 , n55077 );
xor ( n55079 , n54904 , n54946 );
and ( n5755 , n55079 , n5652 );
and ( n55081 , n54904 , n54946 );
or ( n5757 , n5755 , n55081 );
nor ( n55083 , n55078 , n5757 );
not ( n55084 , n5696 );
not ( n55085 , n55023 );
not ( n5761 , n55085 );
or ( n55087 , n55084 , n5761 );
not ( n55088 , n5696 );
nand ( n5764 , n55023 , n55088 );
nand ( n55090 , n55087 , n5764 );
and ( n5766 , n55090 , n5664 );
not ( n5767 , n55090 );
not ( n55093 , n5664 );
and ( n5769 , n5767 , n55093 );
nor ( n55095 , n5766 , n5769 );
buf ( n55096 , n421 );
not ( n5772 , n55096 );
buf ( n55098 , n372 );
nor ( n55099 , n5772 , n55098 );
buf ( n55100 , n55099 );
not ( n5776 , n55100 );
buf ( n55102 , n424 );
buf ( n55103 , n421 );
nand ( n5779 , n55102 , n55103 );
buf ( n55105 , n5779 );
nand ( n55106 , n5776 , n55105 );
not ( n55107 , n55106 );
xor ( n5783 , n371 , n420 );
not ( n55109 , n5783 );
not ( n5785 , n55109 );
or ( n55111 , n55107 , n5785 );
buf ( n55112 , n55100 );
not ( n5788 , n55105 );
buf ( n55114 , n5788 );
nand ( n5790 , n55112 , n55114 );
buf ( n55116 , n5790 );
nand ( n5792 , n55111 , n55116 );
buf ( n55118 , n5792 );
nand ( n5794 , n424 , n420 );
not ( n5795 , n5794 );
not ( n5796 , n5606 );
or ( n5797 , n5795 , n5796 );
not ( n55123 , n5794 );
nand ( n55124 , n55123 , n5605 );
nand ( n55125 , n5797 , n55124 );
not ( n5801 , n54921 );
and ( n55127 , n55125 , n5801 );
not ( n55128 , n55125 );
and ( n55129 , n55128 , n54921 );
nor ( n5805 , n55127 , n55129 );
buf ( n55131 , n5805 );
xor ( n55132 , n55118 , n55131 );
xor ( n55133 , n54995 , n54998 );
xor ( n55134 , n55133 , n55018 );
buf ( n55135 , n55134 );
and ( n55136 , n55132 , n55135 );
and ( n55137 , n55118 , n55131 );
or ( n5813 , n55136 , n55137 );
buf ( n55139 , n5813 );
nor ( n55140 , n55095 , n55139 );
not ( n5816 , n5748 );
not ( n55142 , n55055 );
nand ( n55143 , n55142 , n5734 );
not ( n55144 , n55143 );
or ( n5820 , n5816 , n55144 );
not ( n55146 , n55142 );
nand ( n5822 , n55146 , n55048 );
nand ( n55148 , n5820 , n5822 );
not ( n55149 , n55066 );
nand ( n5825 , n55149 , n55067 );
nand ( n5826 , n55066 , n55070 );
buf ( n55152 , n54951 );
buf ( n55153 , n420 );
nand ( n55154 , n55152 , n55153 );
buf ( n55155 , n55154 );
nand ( n55156 , n5825 , n5826 , n55155 );
buf ( n55157 , n420 );
not ( n55158 , n55157 );
buf ( n5834 , n54958 );
nand ( n5835 , n55158 , n5834 );
buf ( n5836 , n5835 );
nand ( n5837 , n55156 , n5836 );
not ( n55163 , n5837 );
nand ( n5839 , n418 , n422 );
not ( n55165 , n5839 );
nand ( n5841 , n419 , n421 );
nand ( n5842 , n55165 , n5841 , n420 );
not ( n5843 , n420 );
nand ( n55169 , n418 , n422 );
nand ( n55170 , n5843 , n5841 , n55169 );
nand ( n5846 , n5842 , n55170 );
not ( n55172 , n5846 );
not ( n5848 , n422 );
not ( n55174 , n418 );
or ( n55175 , n5848 , n55174 );
nand ( n5851 , n55175 , n420 );
not ( n55177 , n5851 );
not ( n5853 , n5841 );
nand ( n5854 , n55177 , n5853 );
not ( n5855 , n420 );
nand ( n55181 , n55165 , n5855 , n419 , n421 );
nand ( n5857 , n55172 , n5854 , n55181 );
and ( n55183 , n55064 , n55065 );
nand ( n5859 , n419 , n422 );
nand ( n5860 , n418 , n423 );
and ( n55186 , n5859 , n5860 );
nor ( n55187 , n55186 , n55067 );
nor ( n5863 , n55183 , n55187 );
and ( n5864 , n5857 , n5863 );
not ( n55190 , n5857 );
not ( n5866 , n5863 );
and ( n5867 , n55190 , n5866 );
nor ( n5868 , n5864 , n5867 );
xor ( n5869 , n55163 , n5868 );
nor ( n5870 , n55148 , n5869 );
nor ( n5871 , n55083 , n55140 , n5870 );
nand ( n5872 , n5711 , n5871 );
not ( n55198 , n5872 );
buf ( n55199 , n424 );
not ( n5875 , n55199 );
buf ( n55201 , n374 );
nor ( n55202 , n5875 , n55201 );
buf ( n55203 , n55202 );
buf ( n5879 , n55203 );
xnor ( n55205 , n422 , n373 );
buf ( n55206 , n55205 );
xor ( n55207 , n5879 , n55206 );
not ( n55208 , n424 );
nand ( n5884 , n55208 , n423 );
buf ( n55210 , n422 );
buf ( n55211 , n425 );
nand ( n55212 , n55210 , n55211 );
buf ( n55213 , n55212 );
xor ( n55214 , n5884 , n55213 );
buf ( n55215 , n55214 );
xor ( n55216 , n55207 , n55215 );
buf ( n55217 , n55216 );
buf ( n55218 , n55217 );
not ( n5894 , n55218 );
buf ( n5895 , n5894 );
buf ( n55221 , n425 );
not ( n5897 , n55221 );
buf ( n5898 , n5897 );
buf ( n55224 , n5898 );
not ( n5900 , n55224 );
not ( n55226 , n424 );
not ( n5902 , n614 );
or ( n55228 , n55226 , n5902 );
not ( n55229 , n424 );
nand ( n55230 , n55229 , n374 );
nand ( n5906 , n55228 , n55230 );
buf ( n55232 , n5906 );
not ( n55233 , n55232 );
or ( n55234 , n5900 , n55233 );
buf ( n55235 , n423 );
nand ( n5911 , n55234 , n55235 );
buf ( n55237 , n5911 );
buf ( n55238 , n55237 );
not ( n55239 , n55238 );
buf ( n55240 , n55239 );
buf ( n55241 , n55240 );
not ( n5917 , n55241 );
buf ( n5918 , n5917 );
nand ( n5919 , n5895 , n5918 );
not ( n55245 , n423 );
nor ( n5921 , n55245 , n425 );
and ( n5922 , n5906 , n5921 );
not ( n55248 , n5922 );
nor ( n5924 , n5906 , n5921 );
not ( n55250 , n5924 );
buf ( n55251 , n375 );
not ( n5927 , n55251 );
buf ( n5928 , n5927 );
and ( n55254 , n424 , n425 );
nand ( n5930 , n5928 , n55254 );
nand ( n5931 , n55248 , n55250 , n5930 );
not ( n5932 , n5931 );
buf ( n55258 , n376 );
not ( n5934 , n55258 );
and ( n5935 , n55254 , n5928 );
not ( n5936 , n55254 );
and ( n5937 , n5936 , n375 );
nor ( n5938 , n5935 , n5937 );
buf ( n55264 , n5938 );
nor ( n5940 , n5934 , n55264 );
buf ( n55266 , n5940 );
buf ( n55267 , n377 );
not ( n5943 , n55267 );
buf ( n55269 , n5943 );
or ( n5945 , n376 , n55269 );
nand ( n5946 , n5945 , n425 );
nor ( n5947 , n55266 , n5946 );
not ( n5948 , n5947 );
or ( n5949 , n5932 , n5948 );
nor ( n5950 , n5924 , n5922 );
not ( n5951 , n5950 );
not ( n5952 , n5930 );
and ( n5953 , n5951 , n5952 );
not ( n5954 , n5938 );
nor ( n5955 , n5954 , n376 );
and ( n5956 , n5931 , n5955 );
nor ( n5957 , n5953 , n5956 );
nand ( n55283 , n5949 , n5957 );
nand ( n55284 , n5919 , n55283 );
buf ( n55285 , n55217 );
buf ( n55286 , n55240 );
nand ( n5962 , n55285 , n55286 );
buf ( n55288 , n5962 );
buf ( n55289 , n421 );
not ( n5965 , n55289 );
buf ( n55291 , n372 );
not ( n5967 , n55291 );
or ( n5968 , n5965 , n5967 );
buf ( n55294 , n372 );
buf ( n55295 , n421 );
or ( n5971 , n55294 , n55295 );
nand ( n5972 , n5968 , n5971 );
buf ( n55298 , n5972 );
not ( n5974 , n55298 );
not ( n55300 , n55213 );
nand ( n5976 , n55300 , n423 );
buf ( n55302 , n424 );
buf ( n55303 , n423 );
nand ( n5979 , n55302 , n55303 );
buf ( n55305 , n5979 );
nand ( n5981 , n5976 , n55305 );
not ( n5982 , n5981 );
not ( n55308 , n5982 );
or ( n5984 , n5974 , n55308 );
not ( n5985 , n55298 );
nand ( n5986 , n5985 , n5981 );
nand ( n5987 , n5984 , n5986 );
buf ( n55313 , n421 );
buf ( n55314 , n425 );
nand ( n5990 , n55313 , n55314 );
buf ( n55316 , n5990 );
buf ( n55317 , n422 );
not ( n5993 , n55317 );
buf ( n55319 , n373 );
nor ( n55320 , n5993 , n55319 );
buf ( n55321 , n55320 );
and ( n55322 , n55316 , n55321 );
not ( n55323 , n55316 );
not ( n5999 , n373 );
nand ( n55325 , n5999 , n422 );
and ( n55326 , n55323 , n55325 );
nor ( n55327 , n55322 , n55326 );
buf ( n55328 , n424 );
buf ( n55329 , n422 );
nand ( n55330 , n55328 , n55329 );
buf ( n55331 , n55330 );
and ( n6007 , n55327 , n55331 );
not ( n55333 , n55327 );
buf ( n55334 , n55331 );
not ( n6010 , n55334 );
buf ( n6011 , n6010 );
and ( n55337 , n55333 , n6011 );
nor ( n55338 , n6007 , n55337 );
not ( n6014 , n55338 );
and ( n55340 , n5987 , n6014 );
not ( n55341 , n5987 );
and ( n6017 , n55341 , n55338 );
nor ( n55343 , n55340 , n6017 );
not ( n55344 , n55343 );
xor ( n6020 , n5879 , n55206 );
and ( n55346 , n6020 , n55215 );
and ( n55347 , n5879 , n55206 );
or ( n6023 , n55346 , n55347 );
buf ( n55349 , n6023 );
nand ( n55350 , n55344 , n55349 );
and ( n6026 , n55284 , n55288 , n55350 );
buf ( n55352 , n55349 );
not ( n55353 , n55352 );
buf ( n55354 , n55353 );
nand ( n55355 , n55343 , n55354 );
not ( n6031 , n55355 );
nor ( n6032 , n6026 , n6031 );
not ( n55358 , n6032 );
xor ( n6034 , n55118 , n55131 );
xor ( n55360 , n6034 , n55135 );
buf ( n55361 , n55360 );
buf ( n55362 , n55361 );
not ( n6038 , n55362 );
not ( n6039 , n372 );
nand ( n55365 , n6039 , n421 );
and ( n6041 , n55365 , n55105 );
not ( n55367 , n55365 );
and ( n55368 , n55367 , n5788 );
nor ( n6044 , n6041 , n55368 );
and ( n6045 , n6044 , n5783 );
not ( n6046 , n6044 );
and ( n55372 , n6046 , n55109 );
nor ( n55373 , n6045 , n55372 );
buf ( n55374 , n55316 );
not ( n6050 , n55374 );
buf ( n6051 , n6050 );
not ( n55377 , n6051 );
not ( n6053 , n6011 );
or ( n6054 , n55377 , n6053 );
buf ( n55380 , n55331 );
not ( n6056 , n55380 );
buf ( n55382 , n55316 );
not ( n55383 , n55382 );
or ( n6059 , n6056 , n55383 );
buf ( n55385 , n55321 );
nand ( n55386 , n6059 , n55385 );
buf ( n55387 , n55386 );
nand ( n55388 , n6054 , n55387 );
not ( n55389 , n55388 );
nand ( n6065 , n55373 , n55389 );
buf ( n55391 , n55015 );
buf ( n55392 , n422 );
nand ( n55393 , n55391 , n55392 );
buf ( n55394 , n55393 );
not ( n55395 , n55008 );
and ( n6071 , n55394 , n55395 );
not ( n55397 , n55394 );
not ( n6073 , n55005 );
and ( n55399 , n55397 , n6073 );
nor ( n55400 , n6071 , n55399 );
buf ( n55401 , n55400 );
and ( n6077 , n6065 , n55401 );
nor ( n55403 , n55373 , n55389 );
nor ( n55404 , n6077 , n55403 );
buf ( n55405 , n55404 );
not ( n6081 , n55405 );
buf ( n6082 , n6081 );
buf ( n55408 , n6082 );
not ( n55409 , n55408 );
and ( n6085 , n6038 , n55409 );
not ( n55411 , n55373 );
not ( n6087 , n55389 );
not ( n55413 , n55400 );
not ( n6089 , n55413 );
or ( n55415 , n6087 , n6089 );
nand ( n55416 , n55400 , n55388 );
nand ( n6092 , n55415 , n55416 );
or ( n55418 , n55411 , n6092 );
nand ( n55419 , n6092 , n55411 );
nand ( n6095 , n55418 , n55419 );
not ( n55421 , n55298 );
nand ( n6097 , n55421 , n5982 );
not ( n55423 , n6097 );
not ( n55424 , n55338 );
or ( n55425 , n55423 , n55424 );
nand ( n55426 , n55298 , n5981 );
nand ( n6102 , n55425 , n55426 );
nor ( n55428 , n6095 , n6102 );
buf ( n55429 , n55428 );
nor ( n6105 , n6085 , n55429 );
buf ( n6106 , n6105 );
not ( n55432 , n6106 );
or ( n6108 , n55358 , n55432 );
buf ( n6109 , n55361 );
buf ( n55435 , n6082 );
nand ( n55436 , n6109 , n55435 );
buf ( n55437 , n55436 );
buf ( n55438 , n55361 );
buf ( n55439 , n6082 );
or ( n6115 , n55438 , n55439 );
nand ( n6116 , n6095 , n6102 );
buf ( n55442 , n6116 );
not ( n6118 , n55442 );
buf ( n55444 , n6118 );
buf ( n55445 , n55444 );
nand ( n6121 , n6115 , n55445 );
buf ( n6122 , n6121 );
nand ( n55448 , n55437 , n6122 );
not ( n6124 , n55448 );
nand ( n55450 , n6108 , n6124 );
buf ( n6126 , n55450 );
not ( n6127 , n6126 );
buf ( n55453 , n5857 );
or ( n6129 , n55453 , n5866 );
nand ( n55455 , n6129 , n5837 );
nand ( n6131 , n55453 , n5866 );
nand ( n6132 , n55455 , n6131 );
not ( n55458 , n6132 );
nand ( n55459 , n418 , n422 );
not ( n6135 , n55459 );
not ( n55461 , n420 );
nand ( n55462 , n55461 , n418 , n422 );
not ( n55463 , n55462 );
not ( n6139 , n5853 );
or ( n55465 , n55463 , n6139 );
nand ( n6141 , n55465 , n5851 );
nand ( n55467 , n5855 , n419 );
not ( n6143 , n55467 );
nand ( n55469 , n418 , n421 );
not ( n6145 , n55469 );
and ( n55471 , n6143 , n6145 );
and ( n6147 , n55467 , n55043 );
nor ( n55473 , n55471 , n6147 );
not ( n55474 , n55473 );
and ( n6150 , n6141 , n55474 );
not ( n55476 , n6141 );
and ( n55477 , n55476 , n55473 );
or ( n6153 , n6150 , n55477 );
not ( n6154 , n6153 );
or ( n55480 , n6135 , n6154 );
or ( n55481 , n6153 , n55459 );
nand ( n6157 , n55480 , n55481 );
nand ( n55483 , n55458 , n6157 );
not ( n55484 , n55459 );
not ( n6160 , n55473 );
or ( n55486 , n55484 , n6160 );
nand ( n55487 , n55486 , n6141 );
nand ( n55488 , n55474 , n55165 );
nand ( n6164 , n55487 , n55488 );
buf ( n55490 , n418 );
buf ( n55491 , n420 );
nand ( n55492 , n55490 , n55491 );
buf ( n55493 , n55492 );
buf ( n55494 , n55493 );
not ( n55495 , n55494 );
buf ( n55496 , n55495 );
or ( n55497 , n55496 , n419 );
buf ( n55498 , n55493 );
not ( n6174 , n55498 );
buf ( n55500 , n419 );
nand ( n6176 , n6174 , n55500 );
buf ( n55502 , n6176 );
nand ( n55503 , n55497 , n55502 );
not ( n55504 , n419 );
or ( n6180 , n55504 , n420 );
nand ( n55506 , n6180 , n55037 );
xnor ( n6182 , n55503 , n55506 );
nor ( n6183 , n6164 , n6182 );
not ( n6184 , n6183 );
nand ( n6185 , n55483 , n6184 );
not ( n55511 , n6185 );
buf ( n55512 , n55511 );
buf ( n55513 , n419 );
not ( n55514 , n55513 );
buf ( n55515 , n55496 );
nand ( n6191 , n55514 , n55515 );
buf ( n55517 , n6191 );
buf ( n55518 , n55517 );
not ( n6194 , n55518 );
buf ( n6195 , n55506 );
not ( n55521 , n6195 );
buf ( n55522 , n55521 );
buf ( n55523 , n55522 );
not ( n55524 , n55523 );
or ( n55525 , n6194 , n55524 );
buf ( n55526 , n55493 );
buf ( n55527 , n419 );
nand ( n55528 , n55526 , n55527 );
buf ( n55529 , n55528 );
buf ( n55530 , n55529 );
nand ( n6206 , n55525 , n55530 );
buf ( n6207 , n6206 );
buf ( n55533 , n418 );
buf ( n55534 , n55503 );
nand ( n55535 , n55533 , n55534 );
buf ( n55536 , n55535 );
nor ( n6212 , n6207 , n55536 );
not ( n6213 , n55502 );
buf ( n55539 , n418 );
not ( n6215 , n55539 );
buf ( n55541 , n6215 );
nor ( n6217 , n6213 , n55541 );
nor ( n6218 , n6212 , n6217 );
buf ( n55544 , n6218 );
nand ( n6220 , n55512 , n55544 );
buf ( n55546 , n6220 );
buf ( n55547 , n55546 );
nor ( n6223 , n6127 , n55547 );
buf ( n55549 , n6223 );
nand ( n55550 , n55198 , n55549 );
not ( n6226 , n55028 );
buf ( n6227 , n5653 );
not ( n6228 , n6227 );
or ( n6229 , n6226 , n6228 );
nand ( n6230 , n55078 , n5757 );
nand ( n55556 , n6229 , n6230 );
not ( n6232 , n55556 );
nor ( n55558 , n6157 , n6183 );
and ( n55559 , n55558 , n6132 );
and ( n6235 , n6164 , n6182 );
nor ( n55561 , n55559 , n6235 );
buf ( n55562 , n55561 );
not ( n6238 , n55562 );
nand ( n55564 , n55148 , n5869 );
buf ( n6240 , n55564 );
buf ( n6241 , n6207 );
buf ( n6242 , n55536 );
nand ( n6243 , n6241 , n6242 );
buf ( n6244 , n6243 );
or ( n55570 , n6244 , n6217 );
buf ( n55571 , n55570 );
nand ( n6247 , n6240 , n55571 );
buf ( n55573 , n6247 );
buf ( n55574 , n55573 );
nor ( n6250 , n6238 , n55574 );
buf ( n55576 , n6250 );
buf ( n55577 , n55032 );
nand ( n6253 , n55139 , n55095 );
buf ( n55579 , n6253 );
not ( n55580 , n55579 );
buf ( n55581 , n55580 );
buf ( n55582 , n55581 );
nand ( n6258 , n55577 , n55582 );
buf ( n55584 , n6258 );
nand ( n55585 , n6232 , n55576 , n55584 );
buf ( n55586 , n55585 );
nand ( n6262 , n55561 , n5870 );
or ( n6263 , n6262 , n55573 );
nand ( n6264 , n6263 , n6218 );
not ( n6265 , n6264 );
buf ( n55591 , n6265 );
buf ( n55592 , n55561 );
buf ( n55593 , n55592 );
buf ( n55594 , n55593 );
nand ( n6270 , n6185 , n55594 , n55570 );
buf ( n55596 , n6270 );
buf ( n55597 , n55573 );
not ( n6273 , n55597 );
buf ( n55599 , n55083 );
buf ( n55600 , n55594 );
nand ( n6276 , n6273 , n55599 , n55600 );
buf ( n55602 , n6276 );
buf ( n55603 , n55602 );
nand ( n6279 , n55586 , n55591 , n55596 , n55603 );
buf ( n55605 , n6279 );
nand ( n55606 , n55550 , n55605 , n55541 );
not ( n6282 , n55606 );
not ( n55608 , n6282 );
not ( n6284 , n55608 );
buf ( n55610 , n6284 );
and ( n55611 , n54872 , n55610 );
not ( n55612 , n54872 );
not ( n6288 , n6282 );
buf ( n55614 , n6288 );
and ( n55615 , n55612 , n55614 );
nor ( n6291 , n55611 , n55615 );
buf ( n55617 , n6291 );
buf ( n55618 , n413 );
buf ( n55619 , n412 );
not ( n6295 , n55619 );
buf ( n55621 , n6295 );
buf ( n55622 , n55621 );
and ( n6298 , n55618 , n55622 );
not ( n6299 , n55618 );
buf ( n55625 , n412 );
and ( n6301 , n6299 , n55625 );
nor ( n6302 , n6298 , n6301 );
buf ( n55628 , n6302 );
buf ( n55629 , n411 );
buf ( n55630 , n412 );
and ( n6306 , n55629 , n55630 );
not ( n55632 , n55629 );
buf ( n55633 , n55621 );
and ( n55634 , n55632 , n55633 );
nor ( n6310 , n6306 , n55634 );
buf ( n6311 , n6310 );
nand ( n6312 , n55628 , n6311 );
buf ( n55638 , n6312 );
buf ( n55639 , n55628 );
nand ( n55640 , n55638 , n55639 );
buf ( n55641 , n55640 );
nand ( n55642 , n55617 , n55641 );
not ( n55643 , n55642 );
buf ( n6319 , n55643 );
not ( n6320 , n6319 );
not ( n55646 , n413 );
buf ( n6322 , n55646 );
buf ( n55648 , n6322 );
not ( n55649 , n55648 );
buf ( n55650 , n6282 );
not ( n6326 , n55650 );
or ( n6327 , n55649 , n6326 );
buf ( n55653 , n6282 );
not ( n6329 , n55653 );
buf ( n55655 , n413 );
nand ( n6331 , n6329 , n55655 );
buf ( n55657 , n6331 );
buf ( n55658 , n55657 );
nand ( n55659 , n6327 , n55658 );
buf ( n55660 , n55659 );
buf ( n55661 , n55660 );
xnor ( n6337 , n415 , n414 );
buf ( n55663 , n414 );
buf ( n55664 , n413 );
and ( n55665 , n55663 , n55664 );
not ( n6341 , n55663 );
buf ( n55667 , n55646 );
and ( n55668 , n6341 , n55667 );
nor ( n6344 , n55665 , n55668 );
buf ( n6345 , n6344 );
nand ( n55671 , n6337 , n6345 );
buf ( n55672 , n55671 );
buf ( n55673 , n6337 );
nand ( n55674 , n55672 , n55673 );
buf ( n55675 , n55674 );
buf ( n55676 , n55675 );
nand ( n6352 , n55661 , n55676 );
buf ( n55678 , n6352 );
buf ( n55679 , n55678 );
not ( n55680 , n55679 );
buf ( n55681 , n55680 );
buf ( n55682 , n55681 );
not ( n55683 , n55682 );
buf ( n55684 , n55683 );
buf ( n55685 , n55684 );
not ( n55686 , n6288 );
or ( n55687 , n410 , n411 );
nand ( n6363 , n55686 , n55687 );
buf ( n55689 , n6363 );
nand ( n6365 , n55685 , n55689 );
buf ( n55691 , n6365 );
buf ( n6367 , n55691 );
not ( n6368 , n6367 );
buf ( n6369 , n6368 );
nand ( n6370 , n6320 , n6369 );
not ( n6371 , n6370 );
not ( n6372 , n415 );
nand ( n6373 , n6372 , n55608 );
buf ( n55699 , n6282 );
buf ( n55700 , n415 );
nand ( n6376 , n55699 , n55700 );
buf ( n55702 , n6376 );
nand ( n6378 , n6373 , n55702 , n416 );
buf ( n55704 , n55608 );
not ( n6380 , n55704 );
buf ( n55706 , n416 );
not ( n55707 , n55706 );
buf ( n55708 , n55707 );
and ( n6384 , n55708 , n415 );
buf ( n55710 , n6384 );
not ( n6386 , n55710 );
buf ( n55712 , n6386 );
buf ( n55713 , n55712 );
nor ( n6389 , n6380 , n55713 );
buf ( n55715 , n6389 );
not ( n6391 , n55715 );
nand ( n6392 , n6378 , n6391 );
buf ( n55718 , n6392 );
buf ( n6394 , n55718 );
buf ( n55720 , n6394 );
not ( n6396 , n55720 );
or ( n6397 , n6371 , n6396 );
or ( n6398 , n6369 , n6320 );
nand ( n55724 , n6397 , n6398 );
buf ( n55725 , n55724 );
not ( n55726 , n55725 );
not ( n6402 , n55684 );
not ( n55728 , n6402 );
buf ( n55729 , n6363 );
not ( n55730 , n55729 );
buf ( n55731 , n55730 );
not ( n55732 , n55731 );
and ( n55733 , n55728 , n55732 );
and ( n6409 , n6402 , n55731 );
nor ( n55735 , n55733 , n6409 );
buf ( n55736 , n55735 );
not ( n6412 , n55736 );
and ( n55738 , n6363 , n55684 );
buf ( n55739 , n55720 );
not ( n55740 , n55739 );
not ( n55741 , n55643 );
buf ( n55742 , n55741 );
not ( n55743 , n55742 );
and ( n55744 , n55740 , n55743 );
buf ( n55745 , n55720 );
buf ( n55746 , n55741 );
and ( n55747 , n55745 , n55746 );
nor ( n6423 , n55744 , n55747 );
buf ( n6424 , n6423 );
or ( n55750 , n55738 , n6424 );
nand ( n6426 , n6424 , n6369 );
nand ( n55752 , n55750 , n6426 );
buf ( n55753 , n55752 );
not ( n6429 , n55753 );
buf ( n6430 , n6429 );
buf ( n55756 , n6430 );
not ( n6432 , n55756 );
or ( n55758 , n6412 , n6432 );
buf ( n6434 , n55752 );
buf ( n55760 , n55735 );
not ( n55761 , n55760 );
buf ( n55762 , n55761 );
buf ( n55763 , n55762 );
nand ( n55764 , n6434 , n55763 );
buf ( n55765 , n55764 );
buf ( n55766 , n55765 );
nand ( n6442 , n55758 , n55766 );
buf ( n6443 , n6442 );
buf ( n55769 , n6443 );
not ( n6445 , n55769 );
buf ( n55771 , n6445 );
buf ( n55772 , n55771 );
not ( n6448 , n55772 );
or ( n55774 , n55726 , n6448 );
not ( n6450 , n55724 );
buf ( n55776 , n6450 );
buf ( n55777 , n6443 );
nand ( n55778 , n55776 , n55777 );
buf ( n55779 , n55778 );
buf ( n55780 , n55779 );
nand ( n55781 , n55774 , n55780 );
buf ( n55782 , n55781 );
buf ( n55783 , n55782 );
buf ( n6459 , n6430 );
not ( n6460 , n6459 );
buf ( n55786 , n6450 );
buf ( n55787 , n55735 );
nand ( n6463 , n55786 , n55787 );
buf ( n55789 , n6463 );
buf ( n55790 , n55789 );
not ( n6466 , n55790 );
or ( n55792 , n6460 , n6466 );
buf ( n55793 , n55724 );
buf ( n55794 , n55762 );
nand ( n55795 , n55793 , n55794 );
buf ( n55796 , n55795 );
buf ( n55797 , n55796 );
nand ( n55798 , n55792 , n55797 );
buf ( n55799 , n55798 );
buf ( n6475 , n55799 );
nor ( n6476 , n55783 , n6475 );
buf ( n6477 , n6476 );
buf ( n55803 , n6477 );
not ( n6479 , n55803 );
buf ( n55805 , n55782 );
buf ( n55806 , n55799 );
nand ( n55807 , n55805 , n55806 );
buf ( n55808 , n55807 );
buf ( n55809 , n55808 );
nand ( n55810 , n6479 , n55809 );
buf ( n55811 , n55810 );
buf ( n55812 , n55811 );
not ( n55813 , n55812 );
buf ( n55814 , n55813 );
buf ( n55815 , n55814 );
not ( n6491 , n55815 );
not ( n6492 , n55140 );
not ( n6493 , n55078 );
not ( n6494 , n5757 );
nand ( n55820 , n6493 , n6494 );
and ( n6496 , n6492 , n55032 , n55820 );
buf ( n55822 , n6496 );
buf ( n55823 , n55450 );
nand ( n55824 , n55822 , n55823 );
buf ( n55825 , n55824 );
not ( n55826 , n55825 );
not ( n55827 , n6230 );
or ( n6503 , n55826 , n55827 );
buf ( n55829 , n5870 );
not ( n55830 , n55829 );
buf ( n55831 , n55830 );
buf ( n55832 , n55564 );
nand ( n55833 , n55831 , n55832 );
nand ( n6509 , n6503 , n55833 );
buf ( n55835 , n55581 );
not ( n55836 , n55835 );
buf ( n55837 , n55032 );
not ( n6513 , n55837 );
or ( n6514 , n55836 , n6513 );
nand ( n55840 , n55028 , n6227 );
buf ( n55841 , n55840 );
nand ( n6517 , n6514 , n55841 );
buf ( n6518 , n6517 );
buf ( n55844 , n6518 );
buf ( n55845 , n55820 );
nand ( n55846 , n55844 , n55845 );
buf ( n55847 , n55846 );
not ( n55848 , n55847 );
nand ( n6524 , n55848 , n55833 );
not ( n6525 , n6230 );
nor ( n6526 , n6525 , n55833 );
nand ( n55852 , n55847 , n55825 , n6526 );
and ( n6528 , n6509 , n6524 , n55852 );
not ( n55854 , n6528 );
nand ( n6530 , n410 , n411 );
not ( n55856 , n6530 );
and ( n6532 , n55854 , n55856 );
xor ( n55858 , n410 , n411 );
not ( n6534 , n55858 );
not ( n55860 , n55198 );
buf ( n6536 , n55288 );
not ( n55862 , n6536 );
buf ( n55863 , n55862 );
buf ( n55864 , n55863 );
not ( n6540 , n55864 );
buf ( n55866 , n55355 );
not ( n6542 , n55866 );
or ( n6543 , n6540 , n6542 );
buf ( n55869 , n55350 );
nand ( n6545 , n6543 , n55869 );
buf ( n55871 , n6545 );
nand ( n6547 , n6106 , n55871 );
buf ( n55873 , n55355 );
buf ( n55874 , n5919 );
buf ( n55875 , n55283 );
and ( n6551 , n55873 , n55874 , n55875 );
buf ( n55877 , n6551 );
nand ( n6553 , n6106 , n55877 );
nand ( n6554 , n6547 , n6553 , n6124 );
not ( n6555 , n6554 );
or ( n6556 , n55860 , n6555 );
nor ( n6557 , n55083 , n5870 );
not ( n55883 , n6557 );
not ( n6559 , n6518 );
or ( n55885 , n55883 , n6559 );
buf ( n6561 , n6230 );
not ( n55887 , n6561 );
buf ( n55888 , n55887 );
buf ( n55889 , n55888 );
buf ( n55890 , n55831 );
and ( n6566 , n55889 , n55890 );
not ( n6567 , n55832 );
buf ( n55893 , n6567 );
nor ( n55894 , n6566 , n55893 );
buf ( n55895 , n55894 );
nand ( n6571 , n55885 , n55895 );
buf ( n55897 , n6571 );
not ( n6573 , n55897 );
buf ( n55899 , n6573 );
nand ( n6575 , n6556 , n55899 );
or ( n6576 , n55458 , n6157 );
buf ( n55902 , n55483 );
buf ( n55903 , n55902 );
buf ( n55904 , n55903 );
nand ( n6580 , n6576 , n55904 );
not ( n55906 , n6580 );
and ( n55907 , n6575 , n55906 );
not ( n6583 , n6575 );
and ( n55909 , n6583 , n6580 );
nor ( n6585 , n55907 , n55909 );
not ( n6586 , n6585 );
buf ( n6587 , n6586 );
nor ( n6588 , n6534 , n6587 );
nor ( n6589 , n6532 , n6588 );
buf ( n6590 , n6589 );
not ( n6591 , n55671 );
not ( n55917 , n6591 );
not ( n55918 , n6322 );
buf ( n55919 , n6571 );
not ( n6594 , n6212 );
and ( n6595 , n55511 , n6594 );
and ( n6596 , n55919 , n6595 );
nor ( n6597 , n6596 , n6217 );
not ( n6598 , n6597 );
nor ( n6599 , n6185 , n6212 );
nand ( n6600 , n55198 , n6599 , n6554 );
buf ( n55927 , n6600 );
buf ( n55928 , n55594 );
not ( n6603 , n55928 );
buf ( n55930 , n6603 );
buf ( n55931 , n55930 );
buf ( n55932 , n6594 );
and ( n55933 , n55931 , n55932 );
buf ( n55934 , n6244 );
not ( n6609 , n55934 );
buf ( n6610 , n6609 );
buf ( n6611 , n6610 );
nor ( n6612 , n55933 , n6611 );
buf ( n6613 , n6612 );
buf ( n55940 , n6613 );
nand ( n55941 , n55927 , n55940 );
buf ( n55942 , n55941 );
not ( n55943 , n55942 );
buf ( n55944 , n55943 );
not ( n55945 , n55944 );
or ( n55946 , n6598 , n55945 );
not ( n55947 , n55943 );
nand ( n55948 , n55919 , n6595 );
not ( n55949 , n55948 );
or ( n6616 , n55947 , n55949 );
nand ( n55951 , n6616 , n6217 );
nand ( n6618 , n55946 , n55951 );
not ( n6619 , n6618 );
not ( n6620 , n6619 );
not ( n6621 , n6620 );
or ( n6622 , n55918 , n6621 );
not ( n6623 , n55646 );
nand ( n6624 , n6623 , n6619 );
nand ( n6625 , n6622 , n6624 );
not ( n6626 , n6625 );
or ( n6627 , n55917 , n6626 );
buf ( n55962 , n413 );
not ( n6629 , n55962 );
not ( n55964 , n418 );
not ( n55965 , n55546 );
buf ( n55966 , n55448 );
buf ( n55967 , n6106 );
buf ( n55968 , n55967 );
buf ( n55969 , n55968 );
buf ( n55970 , n55969 );
nor ( n55971 , n55966 , n55970 );
buf ( n55972 , n55971 );
not ( n55973 , n55972 );
not ( n6640 , n55448 );
not ( n55975 , n55871 );
buf ( n55976 , n55877 );
not ( n6643 , n55976 );
buf ( n55978 , n6643 );
and ( n6645 , n55975 , n55978 );
nand ( n6646 , n6640 , n6645 );
nand ( n6647 , n55965 , n55973 , n55198 , n6646 );
nand ( n6648 , n6647 , n55605 );
not ( n6649 , n6648 );
or ( n6650 , n55964 , n6649 );
nand ( n55985 , n6650 , n55608 );
buf ( n55986 , n55985 );
not ( n55987 , n55986 );
buf ( n55988 , n55987 );
not ( n55989 , n55988 );
or ( n55990 , n6629 , n55989 );
not ( n55991 , n55985 );
not ( n55992 , n55991 );
nand ( n6659 , n55992 , n6322 );
buf ( n55994 , n6659 );
nand ( n55995 , n55990 , n55994 );
buf ( n55996 , n55995 );
buf ( n55997 , n55996 );
not ( n55998 , n6337 );
buf ( n6665 , n55998 );
buf ( n56000 , n6665 );
nand ( n6667 , n55997 , n56000 );
buf ( n56002 , n6667 );
nand ( n6669 , n6627 , n56002 );
buf ( n56004 , n6669 );
xor ( n56005 , n6590 , n56004 );
not ( n56006 , n411 );
buf ( n6673 , n55511 );
not ( n56008 , n6673 );
not ( n6675 , n6571 );
or ( n56010 , n56008 , n6675 );
buf ( n56011 , n55198 );
buf ( n56012 , n6554 );
buf ( n56013 , n6673 );
and ( n6680 , n56011 , n56012 , n56013 );
buf ( n56015 , n55930 );
nor ( n6682 , n6680 , n56015 );
buf ( n56017 , n6682 );
nand ( n6684 , n56010 , n56017 );
not ( n6685 , n6244 );
nor ( n6686 , n6685 , n6212 );
not ( n6687 , n6686 );
and ( n6688 , n6684 , n6687 );
not ( n6689 , n6684 );
and ( n6690 , n6689 , n6686 );
nor ( n6691 , n6688 , n6690 );
not ( n6692 , n6691 );
not ( n6693 , n6692 );
or ( n6694 , n56006 , n6693 );
or ( n6695 , n6692 , n411 );
nand ( n56030 , n6694 , n6695 );
buf ( n56031 , n56030 );
not ( n6698 , n56031 );
buf ( n56033 , n55628 );
not ( n6700 , n56033 );
and ( n56035 , n6698 , n6700 );
not ( n56036 , n411 );
buf ( n56037 , n55904 );
not ( n56038 , n56037 );
buf ( n56039 , n6571 );
not ( n6706 , n56039 );
or ( n6707 , n56038 , n6706 );
buf ( n56042 , n55198 );
buf ( n56043 , n6554 );
buf ( n56044 , n55904 );
nand ( n6711 , n56042 , n56043 , n56044 );
buf ( n56046 , n6711 );
buf ( n56047 , n56046 );
buf ( n56048 , n6576 );
nand ( n56049 , n56047 , n56048 );
buf ( n56050 , n56049 );
buf ( n56051 , n56050 );
not ( n6718 , n56051 );
buf ( n56053 , n6718 );
buf ( n56054 , n56053 );
nand ( n6721 , n6707 , n56054 );
buf ( n56056 , n6721 );
not ( n6723 , n56056 );
not ( n6724 , n6184 );
nor ( n56059 , n6724 , n6235 );
buf ( n6726 , n56059 );
not ( n56061 , n6726 );
buf ( n56062 , n56061 );
not ( n56063 , n56062 );
and ( n56064 , n6723 , n56063 );
and ( n6731 , n56056 , n56062 );
nor ( n56066 , n56064 , n6731 );
not ( n56067 , n56066 );
or ( n6734 , n56036 , n56067 );
or ( n56069 , n56066 , n411 );
nand ( n56070 , n6734 , n56069 );
buf ( n56071 , n56070 );
not ( n56072 , n6312 );
buf ( n56073 , n56072 );
and ( n56074 , n56071 , n56073 );
nor ( n6741 , n56035 , n56074 );
buf ( n6742 , n6741 );
buf ( n56077 , n6742 );
not ( n6744 , n56077 );
buf ( n56079 , n6744 );
buf ( n56080 , n56079 );
xnor ( n6747 , n56005 , n56080 );
buf ( n56082 , n6747 );
buf ( n56083 , n56082 );
buf ( n56084 , n371 );
buf ( n56085 , n378 );
nand ( n6752 , n56084 , n56085 );
buf ( n56087 , n6752 );
buf ( n56088 , n370 );
buf ( n56089 , n379 );
nand ( n6756 , n56088 , n56089 );
buf ( n56091 , n6756 );
xor ( n6758 , n56087 , n56091 );
buf ( n56093 , n371 );
buf ( n56094 , n379 );
nand ( n6761 , n56093 , n56094 );
buf ( n56096 , n6761 );
buf ( n56097 , n56096 );
buf ( n56098 , n370 );
buf ( n56099 , n380 );
nand ( n6766 , n56098 , n56099 );
buf ( n56101 , n6766 );
buf ( n56102 , n56101 );
xor ( n6769 , n56097 , n56102 );
buf ( n56104 , n372 );
buf ( n56105 , n378 );
nand ( n6772 , n56104 , n56105 );
buf ( n56107 , n6772 );
buf ( n56108 , n56107 );
and ( n6775 , n6769 , n56108 );
and ( n6776 , n56097 , n56102 );
or ( n56111 , n6775 , n6776 );
buf ( n56112 , n56111 );
xor ( n6779 , n6758 , n56112 );
xor ( n56114 , n56097 , n56102 );
xor ( n56115 , n56114 , n56108 );
buf ( n56116 , n56115 );
not ( n56117 , n56116 );
not ( n56118 , n56117 );
buf ( n56119 , n372 );
buf ( n56120 , n379 );
nand ( n56121 , n56119 , n56120 );
buf ( n56122 , n56121 );
buf ( n56123 , n56122 );
buf ( n56124 , n370 );
buf ( n56125 , n381 );
nand ( n6792 , n56124 , n56125 );
buf ( n56127 , n6792 );
buf ( n56128 , n56127 );
xor ( n6795 , n56123 , n56128 );
buf ( n56130 , n373 );
buf ( n56131 , n378 );
nand ( n56132 , n56130 , n56131 );
buf ( n56133 , n56132 );
buf ( n56134 , n56133 );
and ( n56135 , n6795 , n56134 );
and ( n56136 , n56123 , n56128 );
or ( n6803 , n56135 , n56136 );
buf ( n56138 , n6803 );
not ( n56139 , n56138 );
not ( n6806 , n56139 );
or ( n56141 , n56118 , n6806 );
xor ( n56142 , n56123 , n56128 );
xor ( n6809 , n56142 , n56134 );
buf ( n56144 , n6809 );
not ( n6811 , n56144 );
buf ( n56146 , n371 );
buf ( n56147 , n380 );
nand ( n56148 , n56146 , n56147 );
buf ( n56149 , n56148 );
not ( n56150 , n56149 );
buf ( n6817 , n371 );
buf ( n56152 , n381 );
nand ( n56153 , n6817 , n56152 );
buf ( n56154 , n56153 );
buf ( n56155 , n56154 );
buf ( n56156 , n370 );
buf ( n56157 , n382 );
nand ( n6824 , n56156 , n56157 );
buf ( n56159 , n6824 );
buf ( n56160 , n56159 );
xor ( n6827 , n56155 , n56160 );
buf ( n56162 , n373 );
buf ( n56163 , n379 );
nand ( n6830 , n56162 , n56163 );
buf ( n56165 , n6830 );
buf ( n56166 , n56165 );
and ( n6833 , n6827 , n56166 );
and ( n6834 , n56155 , n56160 );
or ( n6835 , n6833 , n6834 );
buf ( n56170 , n6835 );
not ( n6837 , n56170 );
nand ( n56172 , n56150 , n6837 );
not ( n56173 , n56172 );
or ( n56174 , n6811 , n56173 );
nand ( n6841 , n56170 , n56149 );
nand ( n56176 , n56174 , n6841 );
nand ( n56177 , n56141 , n56176 );
nand ( n6844 , n56138 , n56116 );
nand ( n56179 , n56177 , n6844 );
not ( n6846 , n6530 );
buf ( n56181 , n6846 );
not ( n6848 , n56181 );
buf ( n56183 , n55035 );
not ( n6850 , n6492 );
buf ( n56185 , n6850 );
nor ( n6852 , n56183 , n56185 );
buf ( n56187 , n6852 );
not ( n6854 , n56187 );
not ( n56189 , n55450 );
or ( n6856 , n6854 , n56189 );
buf ( n56191 , n6518 );
not ( n56192 , n56191 );
buf ( n56193 , n56192 );
nand ( n6860 , n6856 , n56193 );
nand ( n56195 , n55820 , n6230 );
not ( n6862 , n56195 );
and ( n56197 , n6860 , n6862 );
not ( n56198 , n6860 );
and ( n6865 , n56198 , n56195 );
nor ( n56200 , n56197 , n6865 );
buf ( n56201 , n56200 );
not ( n6868 , n56201 );
or ( n56203 , n6848 , n6868 );
nand ( n56204 , n6509 , n6524 , n55852 );
buf ( n56205 , n56204 );
buf ( n56206 , n55858 );
nand ( n6873 , n56205 , n56206 );
buf ( n56208 , n6873 );
buf ( n56209 , n56208 );
nand ( n56210 , n56203 , n56209 );
buf ( n56211 , n56210 );
xor ( n6878 , n56179 , n56211 );
xor ( n6879 , n6779 , n6878 );
buf ( n56214 , n6879 );
not ( n6881 , n6846 );
nand ( n6882 , n55978 , n55975 );
not ( n6883 , n6882 );
and ( n6884 , n55969 , n6492 );
not ( n6885 , n6884 );
or ( n56220 , n6883 , n6885 );
not ( n56221 , n6122 );
not ( n6888 , n6850 );
and ( n56223 , n56221 , n6888 );
buf ( n56224 , n6850 );
buf ( n56225 , n55437 );
or ( n56226 , n56224 , n56225 );
buf ( n6893 , n6253 );
buf ( n56228 , n6893 );
nand ( n56229 , n56226 , n56228 );
buf ( n56230 , n56229 );
nor ( n56231 , n56223 , n56230 );
nand ( n6898 , n56220 , n56231 );
nand ( n56233 , n5711 , n55840 );
not ( n56234 , n56233 );
and ( n6901 , n6898 , n56234 );
not ( n56236 , n6898 );
and ( n6903 , n56236 , n56233 );
nor ( n56238 , n6901 , n6903 );
not ( n6905 , n56238 );
or ( n56240 , n6881 , n6905 );
nand ( n56241 , n55858 , n56200 );
nand ( n6908 , n56240 , n56241 );
xor ( n56243 , n56138 , n56117 );
xnor ( n6910 , n56243 , n56176 );
or ( n6911 , n6908 , n6910 );
buf ( n56246 , n372 );
buf ( n56247 , n380 );
nand ( n6914 , n56246 , n56247 );
buf ( n56249 , n6914 );
buf ( n56250 , n374 );
buf ( n56251 , n378 );
nand ( n56252 , n56250 , n56251 );
buf ( n56253 , n56252 );
xor ( n56254 , n56249 , n56253 );
nand ( n56255 , n370 , n383 );
nand ( n6922 , n372 , n381 );
or ( n56257 , n56255 , n6922 );
nand ( n56258 , n373 , n380 );
nand ( n6925 , n56257 , n56258 );
nand ( n56260 , n56255 , n6922 );
nand ( n6927 , n6925 , n56260 );
and ( n6928 , n56254 , n6927 );
and ( n6929 , n56249 , n56253 );
or ( n6930 , n6928 , n6929 );
xor ( n6931 , n56149 , n6837 );
xnor ( n6932 , n6931 , n56144 );
xor ( n56267 , n6930 , n6932 );
xor ( n56268 , n56249 , n56253 );
xor ( n6935 , n56268 , n6927 );
not ( n56270 , n6935 );
xor ( n6937 , n56155 , n56160 );
xor ( n6938 , n6937 , n56166 );
buf ( n56273 , n6938 );
not ( n6940 , n56273 );
buf ( n56275 , n374 );
buf ( n56276 , n379 );
nand ( n6943 , n56275 , n56276 );
buf ( n56278 , n6943 );
buf ( n56279 , n56278 );
buf ( n56280 , n371 );
buf ( n56281 , n382 );
nand ( n6948 , n56280 , n56281 );
buf ( n56283 , n6948 );
buf ( n6950 , n56283 );
xor ( n6951 , n56279 , n6950 );
buf ( n56286 , n375 );
buf ( n56287 , n378 );
nand ( n6954 , n56286 , n56287 );
buf ( n56289 , n6954 );
buf ( n56290 , n56289 );
and ( n56291 , n6951 , n56290 );
and ( n6958 , n56279 , n6950 );
or ( n6959 , n56291 , n6958 );
buf ( n56294 , n6959 );
not ( n6961 , n56294 );
nand ( n56296 , n6940 , n6961 );
not ( n6963 , n56296 );
or ( n6964 , n56270 , n6963 );
nand ( n6965 , n56273 , n56294 );
nand ( n6966 , n6964 , n6965 );
and ( n6967 , n56267 , n6966 );
and ( n6968 , n6930 , n6932 );
or ( n6969 , n6967 , n6968 );
nand ( n6970 , n6911 , n6969 );
buf ( n56305 , n6970 );
nand ( n6972 , n6908 , n6910 );
buf ( n56307 , n6972 );
nand ( n56308 , n56305 , n56307 );
buf ( n56309 , n56308 );
buf ( n56310 , n56309 );
xor ( n56311 , n56214 , n56310 );
buf ( n6978 , n55628 );
not ( n6979 , n6978 );
buf ( n6980 , n6979 );
not ( n56315 , n6980 );
not ( n6982 , n411 );
not ( n6983 , n6586 );
or ( n56318 , n6982 , n6983 );
or ( n6985 , n6586 , n411 );
nand ( n56320 , n56318 , n6985 );
not ( n56321 , n56320 );
or ( n6988 , n56315 , n56321 );
not ( n56323 , n411 );
not ( n6990 , n56323 );
not ( n6991 , n56204 );
or ( n6992 , n6990 , n6991 );
or ( n6993 , n56323 , n56204 );
nand ( n56328 , n6992 , n6993 );
buf ( n56329 , n56328 );
buf ( n56330 , n56072 );
nand ( n56331 , n56329 , n56330 );
buf ( n56332 , n56331 );
nand ( n56333 , n6988 , n56332 );
buf ( n56334 , n56333 );
not ( n7001 , n56334 );
not ( n7002 , n416 );
not ( n56337 , n415 );
not ( n7004 , n55991 );
or ( n56339 , n56337 , n7004 );
not ( n7006 , n415 );
nand ( n56341 , n7006 , n55985 );
nand ( n56342 , n56339 , n56341 );
not ( n7009 , n56342 );
or ( n56344 , n7002 , n7009 );
nand ( n56345 , n6618 , n415 );
nand ( n7012 , n6597 , n55944 );
nand ( n7013 , n55951 , n7012 );
not ( n56348 , n7013 );
not ( n7015 , n415 );
nand ( n7016 , n56348 , n7015 );
nand ( n7017 , n56345 , n7016 , n6384 );
nand ( n7018 , n56344 , n7017 );
buf ( n56353 , n7018 );
not ( n7020 , n56353 );
or ( n7021 , n7001 , n7020 );
or ( n56356 , n7018 , n56333 );
buf ( n56357 , n6591 );
not ( n7024 , n56357 );
and ( n56359 , n56056 , n56059 );
not ( n7026 , n56056 );
and ( n7027 , n7026 , n56062 );
nor ( n7028 , n56359 , n7027 );
xor ( n7029 , n413 , n7028 );
buf ( n56364 , n7029 );
not ( n7031 , n56364 );
or ( n56366 , n7024 , n7031 );
not ( n7033 , n55646 );
and ( n56368 , n6686 , n7033 );
not ( n7035 , n6686 );
not ( n7036 , n413 );
and ( n7037 , n7035 , n7036 );
or ( n7038 , n56368 , n7037 );
and ( n56373 , n6684 , n7038 );
not ( n7040 , n6684 );
not ( n7041 , n55646 );
and ( n56376 , n6687 , n7041 );
not ( n7043 , n6687 );
not ( n7044 , n413 );
and ( n56379 , n7043 , n7044 );
or ( n7046 , n56376 , n56379 );
and ( n7047 , n7040 , n7046 );
or ( n56382 , n56373 , n7047 );
nand ( n7049 , n56382 , n55998 );
buf ( n56384 , n7049 );
nand ( n56385 , n56366 , n56384 );
buf ( n56386 , n56385 );
nand ( n7053 , n56356 , n56386 );
buf ( n56388 , n7053 );
nand ( n56389 , n7021 , n56388 );
buf ( n56390 , n56389 );
buf ( n56391 , n56390 );
and ( n56392 , n56311 , n56391 );
and ( n56393 , n56214 , n56310 );
or ( n7060 , n56392 , n56393 );
buf ( n56395 , n7060 );
buf ( n56396 , n56395 );
xor ( n7063 , n56083 , n56396 );
xor ( n56398 , n56087 , n56091 );
xor ( n56399 , n56398 , n56112 );
and ( n7066 , n56179 , n56399 );
xor ( n7067 , n56087 , n56091 );
xor ( n7068 , n7067 , n56112 );
and ( n7069 , n56211 , n7068 );
and ( n7070 , n56179 , n56211 );
or ( n56405 , n7066 , n7069 , n7070 );
buf ( n56406 , n56405 );
xor ( n7073 , n56087 , n56091 );
and ( n7074 , n7073 , n56112 );
and ( n7075 , n56087 , n56091 );
or ( n7076 , n7074 , n7075 );
buf ( n56411 , n7076 );
buf ( n56412 , n370 );
buf ( n56413 , n378 );
nand ( n7080 , n56412 , n56413 );
buf ( n56415 , n7080 );
buf ( n7082 , n56415 );
xor ( n7083 , n56411 , n7082 );
buf ( n56418 , n7083 );
not ( n56419 , n55686 );
not ( n7086 , n55712 );
and ( n56421 , n56419 , n7086 );
and ( n56422 , n6373 , n55702 , n416 );
nor ( n7089 , n56421 , n56422 );
buf ( n56424 , n7089 );
and ( n56425 , n56418 , n56424 );
not ( n7092 , n56418 );
and ( n7093 , n7092 , n55720 );
or ( n56428 , n56425 , n7093 );
buf ( n7095 , n56428 );
xor ( n7096 , n56406 , n7095 );
not ( n56431 , n6384 );
not ( n56432 , n56342 );
or ( n7099 , n56431 , n56432 );
nand ( n7100 , n7099 , n6378 );
buf ( n7101 , n7100 );
not ( n56436 , n6591 );
not ( n7103 , n56382 );
or ( n56438 , n56436 , n7103 );
not ( n56439 , n55998 );
nor ( n56440 , n56439 , n413 );
and ( n7107 , n6620 , n56440 );
not ( n56442 , n55998 );
nor ( n7109 , n56442 , n55646 );
and ( n7110 , n6619 , n7109 );
nor ( n7111 , n7107 , n7110 );
nand ( n7112 , n56438 , n7111 );
buf ( n56447 , n7112 );
xor ( n7114 , n7101 , n56447 );
buf ( n56449 , n6980 );
not ( n7116 , n56449 );
buf ( n56451 , n56070 );
not ( n56452 , n56451 );
or ( n56453 , n7116 , n56452 );
nand ( n7120 , n56320 , n56072 );
buf ( n56455 , n7120 );
nand ( n56456 , n56453 , n56455 );
buf ( n56457 , n56456 );
buf ( n56458 , n56457 );
and ( n56459 , n7114 , n56458 );
and ( n56460 , n7101 , n56447 );
or ( n7127 , n56459 , n56460 );
buf ( n56462 , n7127 );
buf ( n7129 , n56462 );
xor ( n7130 , n7096 , n7129 );
buf ( n56465 , n7130 );
buf ( n56466 , n56465 );
xor ( n56467 , n7063 , n56466 );
buf ( n56468 , n56467 );
xor ( n56469 , n7101 , n56447 );
xor ( n56470 , n56469 , n56458 );
buf ( n56471 , n56470 );
buf ( n56472 , n56471 );
buf ( n56473 , n56472 );
buf ( n56474 , n56473 );
not ( n7141 , n56474 );
xor ( n56476 , n56214 , n56310 );
xor ( n7143 , n56476 , n56391 );
buf ( n56478 , n7143 );
buf ( n56479 , n56478 );
buf ( n7146 , n56479 );
buf ( n56481 , n7146 );
not ( n56482 , n56481 );
or ( n7149 , n7141 , n56482 );
or ( n56484 , n56481 , n56474 );
xnor ( n56485 , n6969 , n6910 );
xor ( n56486 , n56485 , n6908 );
not ( n7153 , n56486 );
buf ( n56488 , n55858 );
not ( n7155 , n56488 );
buf ( n56490 , n56238 );
not ( n56491 , n56490 );
or ( n7158 , n7155 , n56491 );
buf ( n56493 , n6846 );
not ( n56494 , n6850 );
nand ( n7161 , n56494 , n6893 );
not ( n56496 , n7161 );
not ( n7163 , n56496 );
not ( n7164 , n6554 );
not ( n56499 , n7164 );
or ( n7166 , n7163 , n56499 );
nand ( n56501 , n55973 , n6646 , n7161 );
nand ( n7168 , n7166 , n56501 );
buf ( n56503 , n7168 );
nand ( n7170 , n56493 , n56503 );
buf ( n56505 , n7170 );
buf ( n56506 , n56505 );
nand ( n7173 , n7158 , n56506 );
buf ( n56508 , n7173 );
buf ( n56509 , n56508 );
not ( n7176 , n56509 );
not ( n7177 , n6384 );
and ( n56512 , n415 , n6692 );
not ( n7179 , n415 );
not ( n56514 , n6692 );
and ( n7181 , n7179 , n56514 );
nor ( n56516 , n56512 , n7181 );
not ( n7183 , n56516 );
or ( n56518 , n7177 , n7183 );
not ( n56519 , n55708 );
not ( n7186 , n7015 );
not ( n56521 , n7013 );
or ( n7188 , n7186 , n56521 );
or ( n7189 , n7013 , n7015 );
nand ( n56524 , n7188 , n7189 );
nand ( n56525 , n56519 , n56524 );
nand ( n7192 , n56518 , n56525 );
buf ( n56527 , n7192 );
not ( n7194 , n56527 );
or ( n56529 , n7176 , n7194 );
buf ( n56530 , n7192 );
buf ( n56531 , n56508 );
or ( n56532 , n56530 , n56531 );
buf ( n56533 , n55998 );
not ( n7200 , n56533 );
buf ( n56535 , n7029 );
not ( n56536 , n56535 );
or ( n7203 , n7200 , n56536 );
not ( n7204 , n55646 );
not ( n7205 , n6585 );
or ( n7206 , n7204 , n7205 );
nand ( n56541 , n6586 , n413 );
nand ( n56542 , n7206 , n56541 );
nand ( n7209 , n56542 , n6591 );
buf ( n56544 , n7209 );
nand ( n56545 , n7203 , n56544 );
buf ( n56546 , n56545 );
buf ( n56547 , n56546 );
nand ( n7214 , n56532 , n56547 );
buf ( n7215 , n7214 );
buf ( n56550 , n7215 );
nand ( n7217 , n56529 , n56550 );
buf ( n7218 , n7217 );
buf ( n56553 , n7218 );
not ( n7220 , n56553 );
buf ( n56555 , n7220 );
not ( n56556 , n56555 );
or ( n7223 , n7153 , n56556 );
nand ( n56558 , n56328 , n6980 );
xor ( n7225 , n6930 , n6932 );
xor ( n56560 , n7225 , n6966 );
not ( n56561 , n56560 );
not ( n7228 , n56200 );
nand ( n7229 , n7228 , n411 );
not ( n7230 , n411 );
nand ( n56565 , n7230 , n56200 );
nand ( n56566 , n7229 , n56565 );
nand ( n56567 , n56566 , n56072 );
nand ( n7234 , n56558 , n56561 , n56567 );
not ( n7235 , n7234 );
nand ( n56570 , n56255 , n6922 , n56258 );
not ( n7237 , n6922 );
not ( n7238 , n56258 );
nand ( n56573 , n7237 , n7238 , n56255 );
not ( n7240 , n56255 );
nand ( n7241 , n7240 , n7237 , n56258 );
nand ( n7242 , n7240 , n7238 , n6922 );
nand ( n7243 , n56570 , n56573 , n7241 , n7242 );
buf ( n7244 , n373 );
buf ( n56579 , n381 );
nand ( n56580 , n7244 , n56579 );
buf ( n56581 , n56580 );
buf ( n56582 , n56581 );
buf ( n56583 , n375 );
buf ( n56584 , n379 );
nand ( n56585 , n56583 , n56584 );
buf ( n56586 , n56585 );
buf ( n56587 , n56586 );
or ( n56588 , n56582 , n56587 );
buf ( n56589 , n56588 );
xor ( n7256 , n7243 , n56589 );
buf ( n56591 , n371 );
buf ( n56592 , n383 );
nand ( n56593 , n56591 , n56592 );
buf ( n56594 , n56593 );
not ( n56595 , n56594 );
buf ( n56596 , n374 );
buf ( n56597 , n380 );
nand ( n56598 , n56596 , n56597 );
buf ( n56599 , n56598 );
not ( n56600 , n56599 );
or ( n56601 , n56595 , n56600 );
not ( n7268 , n56599 );
not ( n56603 , n7268 );
not ( n7270 , n56594 );
not ( n7271 , n7270 );
or ( n7272 , n56603 , n7271 );
buf ( n56607 , n376 );
buf ( n56608 , n378 );
nand ( n7275 , n56607 , n56608 );
buf ( n56610 , n7275 );
nand ( n7277 , n7272 , n56610 );
nand ( n7278 , n56601 , n7277 );
and ( n7279 , n7256 , n7278 );
and ( n7280 , n7243 , n56589 );
or ( n7281 , n7279 , n7280 );
not ( n56616 , n6961 );
not ( n56617 , n56273 );
or ( n7284 , n56616 , n56617 );
nand ( n56619 , n56294 , n6940 );
nand ( n56620 , n7284 , n56619 );
xor ( n7287 , n56620 , n6935 );
xor ( n56622 , n7281 , n7287 );
xor ( n7289 , n56279 , n6950 );
xor ( n56624 , n7289 , n56290 );
buf ( n56625 , n56624 );
buf ( n56626 , n56625 );
buf ( n56627 , n372 );
buf ( n56628 , n382 );
nand ( n7295 , n56627 , n56628 );
buf ( n56630 , n7295 );
buf ( n56631 , n56630 );
buf ( n56632 , n370 );
buf ( n56633 , n384 );
nand ( n7300 , n56632 , n56633 );
buf ( n56635 , n7300 );
buf ( n56636 , n56635 );
xor ( n7303 , n56631 , n56636 );
buf ( n56638 , n376 );
buf ( n56639 , n379 );
nand ( n7306 , n56638 , n56639 );
buf ( n56641 , n7306 );
buf ( n56642 , n56641 );
buf ( n56643 , n375 );
buf ( n56644 , n380 );
nand ( n56645 , n56643 , n56644 );
buf ( n56646 , n56645 );
buf ( n56647 , n56646 );
or ( n56648 , n56642 , n56647 );
buf ( n56649 , n377 );
buf ( n56650 , n378 );
nand ( n7317 , n56649 , n56650 );
buf ( n56652 , n7317 );
buf ( n56653 , n56652 );
nand ( n7320 , n56648 , n56653 );
buf ( n56655 , n7320 );
buf ( n56656 , n56655 );
buf ( n7323 , n56646 );
buf ( n56658 , n56641 );
nand ( n56659 , n7323 , n56658 );
buf ( n56660 , n56659 );
buf ( n56661 , n56660 );
nand ( n7328 , n56656 , n56661 );
buf ( n56663 , n7328 );
buf ( n56664 , n56663 );
and ( n7331 , n7303 , n56664 );
and ( n7332 , n56631 , n56636 );
or ( n56667 , n7331 , n7332 );
buf ( n56668 , n56667 );
buf ( n56669 , n56668 );
xor ( n56670 , n56626 , n56669 );
not ( n7337 , n7270 );
nand ( n7338 , n7337 , n56599 , n56610 );
not ( n56673 , n56610 );
nand ( n7340 , n56594 , n56673 , n7268 );
nand ( n56675 , n7270 , n56599 , n56673 );
nand ( n56676 , n7270 , n56610 , n7268 );
nand ( n7343 , n7338 , n7340 , n56675 , n56676 );
not ( n56678 , n7343 );
buf ( n7345 , n372 );
buf ( n56680 , n383 );
nand ( n7347 , n7345 , n56680 );
buf ( n7348 , n7347 );
buf ( n56683 , n7348 );
buf ( n56684 , n371 );
buf ( n56685 , n384 );
nand ( n7352 , n56684 , n56685 );
buf ( n56687 , n7352 );
buf ( n56688 , n56687 );
nor ( n56689 , n56683 , n56688 );
buf ( n56690 , n56689 );
nand ( n7357 , n56678 , n56690 );
not ( n7358 , n7357 );
buf ( n7359 , n374 );
buf ( n56694 , n381 );
nand ( n56695 , n7359 , n56694 );
buf ( n56696 , n56695 );
buf ( n56697 , n56696 );
buf ( n56698 , n373 );
buf ( n56699 , n382 );
nand ( n7366 , n56698 , n56699 );
buf ( n56701 , n7366 );
buf ( n56702 , n56701 );
xor ( n7369 , n56697 , n56702 );
buf ( n56704 , n370 );
buf ( n56705 , n385 );
nand ( n7372 , n56704 , n56705 );
buf ( n56707 , n7372 );
buf ( n56708 , n56707 );
and ( n7375 , n7369 , n56708 );
and ( n56710 , n56697 , n56702 );
or ( n7377 , n7375 , n56710 );
buf ( n56712 , n7377 );
not ( n56713 , n56712 );
or ( n7380 , n7358 , n56713 );
buf ( n56715 , n56690 );
not ( n7382 , n56715 );
buf ( n56717 , n7382 );
nand ( n7384 , n7343 , n56717 );
nand ( n7385 , n7380 , n7384 );
buf ( n56720 , n7385 );
and ( n7387 , n56670 , n56720 );
and ( n56722 , n56626 , n56669 );
or ( n56723 , n7387 , n56722 );
buf ( n56724 , n56723 );
and ( n56725 , n56622 , n56724 );
and ( n56726 , n7281 , n7287 );
or ( n7393 , n56725 , n56726 );
not ( n56728 , n7393 );
or ( n56729 , n7235 , n56728 );
not ( n7396 , n6980 );
not ( n56731 , n56328 );
or ( n7398 , n7396 , n56731 );
nand ( n7399 , n7398 , n56567 );
nand ( n56734 , n7399 , n56560 );
nand ( n7401 , n56729 , n56734 );
buf ( n56736 , n7401 );
not ( n56737 , n56736 );
buf ( n56738 , n56737 );
buf ( n56739 , n56738 );
not ( n56740 , n56739 );
buf ( n56741 , n56740 );
nand ( n7408 , n7223 , n56741 );
buf ( n56743 , n7408 );
not ( n7410 , n56486 );
nand ( n7411 , n7410 , n7218 );
buf ( n56746 , n7411 );
nand ( n7413 , n56743 , n56746 );
buf ( n56748 , n7413 );
nand ( n7415 , n56484 , n56748 );
nand ( n7416 , n7149 , n7415 );
nand ( n7417 , n56468 , n7416 );
not ( n7418 , n7417 );
buf ( n56753 , n56066 );
not ( n7420 , n56753 );
buf ( n56755 , n7420 );
and ( n7422 , n56755 , n55858 );
not ( n7423 , n6846 );
nor ( n56758 , n7423 , n6587 );
nor ( n7425 , n7422 , n56758 );
buf ( n56760 , n7425 );
buf ( n56761 , n411 );
not ( n7428 , n56761 );
buf ( n56763 , n6619 );
not ( n56764 , n56763 );
or ( n56765 , n7428 , n56764 );
buf ( n56766 , n411 );
not ( n56767 , n56766 );
buf ( n56768 , n56767 );
nand ( n56769 , n56768 , n6618 );
buf ( n56770 , n56769 );
nand ( n7437 , n56765 , n56770 );
buf ( n7438 , n7437 );
not ( n7439 , n7438 );
not ( n7440 , n6980 );
or ( n7441 , n7439 , n7440 );
not ( n7442 , n56030 );
nand ( n7443 , n7442 , n56072 );
nand ( n7444 , n7441 , n7443 );
buf ( n56779 , n7444 );
xor ( n7446 , n56760 , n56779 );
buf ( n56781 , n55720 );
xnor ( n7448 , n7446 , n56781 );
buf ( n56783 , n7448 );
buf ( n56784 , n56783 );
buf ( n56785 , n6591 );
not ( n56786 , n56785 );
buf ( n56787 , n55996 );
not ( n56788 , n56787 );
or ( n7455 , n56786 , n56788 );
buf ( n7456 , n55660 );
buf ( n56791 , n55998 );
nand ( n7458 , n7456 , n56791 );
buf ( n56793 , n7458 );
buf ( n56794 , n56793 );
nand ( n7461 , n7455 , n56794 );
buf ( n7462 , n7461 );
buf ( n56797 , n56415 );
not ( n56798 , n56797 );
buf ( n56799 , n56798 );
buf ( n56800 , n56799 );
not ( n56801 , n56800 );
buf ( n56802 , n6392 );
nand ( n56803 , n56801 , n56802 );
buf ( n56804 , n56803 );
buf ( n7471 , n56804 );
buf ( n56806 , n56799 );
not ( n56807 , n56806 );
buf ( n56808 , n7089 );
not ( n7475 , n56808 );
or ( n7476 , n56807 , n7475 );
buf ( n56811 , n7076 );
nand ( n7478 , n7476 , n56811 );
buf ( n56813 , n7478 );
buf ( n56814 , n56813 );
and ( n56815 , n7471 , n56814 );
buf ( n56816 , n56815 );
xor ( n56817 , n7462 , n56816 );
buf ( n56818 , n6589 );
not ( n7485 , n56818 );
buf ( n56820 , n6742 );
not ( n56821 , n56820 );
or ( n7488 , n7485 , n56821 );
buf ( n56823 , n6669 );
nand ( n56824 , n7488 , n56823 );
buf ( n56825 , n56824 );
buf ( n56826 , n56825 );
not ( n7493 , n6589 );
nand ( n7494 , n7493 , n56079 );
buf ( n56829 , n7494 );
nand ( n7496 , n56826 , n56829 );
buf ( n7497 , n7496 );
xnor ( n7498 , n56817 , n7497 );
buf ( n56833 , n7498 );
xor ( n7500 , n56784 , n56833 );
buf ( n56835 , n7500 );
buf ( n56836 , n56835 );
xor ( n56837 , n56406 , n7095 );
and ( n7504 , n56837 , n7129 );
and ( n56839 , n56406 , n7095 );
or ( n56840 , n7504 , n56839 );
buf ( n56841 , n56840 );
buf ( n56842 , n56841 );
and ( n56843 , n56836 , n56842 );
not ( n7510 , n56836 );
buf ( n56845 , n56841 );
not ( n56846 , n56845 );
buf ( n56847 , n56846 );
buf ( n56848 , n56847 );
and ( n56849 , n7510 , n56848 );
nor ( n7516 , n56843 , n56849 );
buf ( n56851 , n7516 );
buf ( n56852 , n56851 );
xor ( n7519 , n56083 , n56396 );
and ( n56854 , n7519 , n56466 );
and ( n7521 , n56083 , n56396 );
or ( n56856 , n56854 , n7521 );
buf ( n56857 , n56856 );
buf ( n56858 , n56857 );
nand ( n56859 , n56852 , n56858 );
buf ( n56860 , n56859 );
not ( n7527 , n56860 );
or ( n56862 , n7418 , n7527 );
buf ( n56863 , n56851 );
not ( n7530 , n56863 );
buf ( n7531 , n7530 );
buf ( n7532 , n56857 );
not ( n56867 , n7532 );
buf ( n56868 , n56867 );
nand ( n56869 , n7531 , n56868 );
nand ( n56870 , n56862 , n56869 );
not ( n7537 , n56424 );
not ( n56872 , n7425 );
and ( n56873 , n7537 , n56872 );
nand ( n7540 , n56424 , n7425 );
and ( n7541 , n7540 , n7444 );
nor ( n7542 , n56873 , n7541 );
buf ( n56877 , n7542 );
buf ( n56878 , n56825 );
not ( n7545 , n56878 );
buf ( n56880 , n7494 );
not ( n7547 , n56880 );
or ( n56882 , n7545 , n7547 );
buf ( n56883 , n7462 );
not ( n7550 , n56883 );
buf ( n56885 , n56804 );
buf ( n56886 , n56813 );
and ( n7553 , n56885 , n56886 );
buf ( n56888 , n7553 );
buf ( n56889 , n56888 );
nand ( n56890 , n7550 , n56889 );
buf ( n56891 , n56890 );
buf ( n56892 , n56891 );
nand ( n56893 , n56882 , n56892 );
buf ( n56894 , n56893 );
buf ( n56895 , n56894 );
buf ( n56896 , n56888 );
not ( n7563 , n56896 );
buf ( n56898 , n7462 );
nand ( n7565 , n7563 , n56898 );
buf ( n56900 , n7565 );
buf ( n56901 , n56900 );
and ( n7568 , n56895 , n56901 );
buf ( n56903 , n7568 );
buf ( n7570 , n56903 );
xor ( n7571 , n56877 , n7570 );
not ( n56906 , n6392 );
and ( n56907 , n55684 , n56906 );
not ( n7574 , n55684 );
not ( n56909 , n56424 );
and ( n56910 , n7574 , n56909 );
nor ( n7577 , n56907 , n56910 );
not ( n56912 , n7577 );
buf ( n56913 , n56912 );
not ( n56914 , n56913 );
buf ( n56915 , n6980 );
not ( n7582 , n56915 );
and ( n56917 , n411 , n55991 );
not ( n7584 , n411 );
and ( n56919 , n7584 , n55986 );
or ( n7586 , n56917 , n56919 );
buf ( n56921 , n7586 );
not ( n7588 , n56921 );
or ( n56923 , n7582 , n7588 );
buf ( n56924 , n7438 );
buf ( n56925 , n56072 );
nand ( n56926 , n56924 , n56925 );
buf ( n56927 , n56926 );
buf ( n56928 , n56927 );
nand ( n56929 , n56923 , n56928 );
buf ( n56930 , n56929 );
buf ( n56931 , n56930 );
buf ( n56932 , n6846 );
not ( n56933 , n56932 );
buf ( n56934 , n56755 );
not ( n7601 , n56934 );
or ( n7602 , n56933 , n7601 );
buf ( n56937 , n6691 );
not ( n56938 , n56937 );
buf ( n56939 , n55858 );
nand ( n56940 , n56938 , n56939 );
buf ( n56941 , n56940 );
buf ( n56942 , n56941 );
nand ( n7609 , n7602 , n56942 );
buf ( n56944 , n7609 );
buf ( n56945 , n56944 );
not ( n56946 , n56945 );
buf ( n56947 , n56946 );
buf ( n56948 , n56947 );
and ( n56949 , n56931 , n56948 );
not ( n7616 , n56931 );
buf ( n56951 , n56944 );
and ( n56952 , n7616 , n56951 );
nor ( n7619 , n56949 , n56952 );
buf ( n56954 , n7619 );
buf ( n56955 , n56954 );
not ( n56956 , n56955 );
and ( n56957 , n56914 , n56956 );
buf ( n56958 , n56912 );
buf ( n56959 , n56954 );
and ( n56960 , n56958 , n56959 );
nor ( n7627 , n56957 , n56960 );
buf ( n7628 , n7627 );
buf ( n56963 , n7628 );
and ( n7630 , n7571 , n56963 );
and ( n56965 , n56877 , n7570 );
or ( n56966 , n7630 , n56965 );
buf ( n56967 , n56966 );
buf ( n56968 , n56967 );
nand ( n56969 , n55684 , n56906 );
buf ( n56970 , n56969 );
not ( n7637 , n56970 );
buf ( n56972 , n7637 );
buf ( n56973 , n56972 );
buf ( n56974 , n56973 );
buf ( n56975 , n56930 );
not ( n7642 , n56975 );
buf ( n56977 , n56947 );
nand ( n7644 , n7642 , n56977 );
buf ( n56979 , n7644 );
buf ( n56980 , n56979 );
not ( n56981 , n56980 );
buf ( n56982 , n56912 );
not ( n7649 , n56982 );
or ( n56984 , n56981 , n7649 );
buf ( n7651 , n56947 );
not ( n7652 , n7651 );
buf ( n56987 , n56930 );
nand ( n56988 , n7652 , n56987 );
buf ( n56989 , n56988 );
buf ( n56990 , n56989 );
nand ( n7657 , n56984 , n56990 );
buf ( n7658 , n7657 );
buf ( n7659 , n7658 );
xor ( n7660 , n56974 , n7659 );
not ( n56995 , n6619 );
not ( n56996 , n56995 );
not ( n56997 , n55858 );
or ( n7664 , n56996 , n56997 );
buf ( n56999 , n6691 );
not ( n7666 , n56999 );
buf ( n57001 , n6846 );
nand ( n7668 , n7666 , n57001 );
buf ( n57003 , n7668 );
nand ( n57004 , n7664 , n57003 );
not ( n57005 , n6980 );
buf ( n57006 , n55617 );
buf ( n57007 , n57006 );
buf ( n57008 , n57007 );
not ( n7675 , n57008 );
or ( n57010 , n57005 , n7675 );
nand ( n57011 , n7586 , n56072 );
nand ( n7678 , n57010 , n57011 );
and ( n7679 , n57004 , n7678 );
not ( n57014 , n57004 );
buf ( n57015 , n7586 );
buf ( n57016 , n56072 );
and ( n7683 , n57015 , n57016 );
buf ( n57018 , n57008 );
buf ( n57019 , n6980 );
and ( n7686 , n57018 , n57019 );
nor ( n57021 , n7683 , n7686 );
buf ( n57022 , n57021 );
and ( n57023 , n57014 , n57022 );
or ( n7690 , n7679 , n57023 );
xor ( n57025 , n7690 , n56912 );
buf ( n57026 , n57025 );
xnor ( n7693 , n7660 , n57026 );
buf ( n7694 , n7693 );
buf ( n57029 , n7694 );
nand ( n7696 , n56968 , n57029 );
buf ( n57031 , n7696 );
buf ( n57032 , n57031 );
xor ( n7699 , n56877 , n7570 );
xor ( n7700 , n7699 , n56963 );
buf ( n57035 , n7700 );
or ( n57036 , n7498 , n56783 );
buf ( n57037 , n57036 );
buf ( n57038 , n56841 );
and ( n57039 , n57037 , n57038 );
and ( n7706 , n56784 , n56833 );
buf ( n57041 , n7706 );
buf ( n57042 , n57041 );
nor ( n57043 , n57039 , n57042 );
buf ( n57044 , n57043 );
nand ( n57045 , n57035 , n57044 );
buf ( n57046 , n57045 );
nand ( n7713 , n57032 , n57046 );
buf ( n57048 , n7713 );
or ( n57049 , n56870 , n57048 );
not ( n57050 , n57031 );
buf ( n57051 , n57035 );
buf ( n57052 , n57044 );
nor ( n57053 , n57051 , n57052 );
buf ( n57054 , n57053 );
not ( n7721 , n57054 );
or ( n7722 , n57050 , n7721 );
or ( n57057 , n7694 , n56967 );
nand ( n7724 , n7722 , n57057 );
not ( n57059 , n7724 );
nand ( n57060 , n57049 , n57059 );
buf ( n57061 , n55858 );
not ( n57062 , n57061 );
buf ( n57063 , n55986 );
not ( n7730 , n57063 );
or ( n7731 , n57062 , n7730 );
buf ( n57066 , n56995 );
buf ( n57067 , n6846 );
nand ( n57068 , n57066 , n57067 );
buf ( n57069 , n57068 );
buf ( n57070 , n57069 );
nand ( n7737 , n7731 , n57070 );
buf ( n57072 , n7737 );
buf ( n57073 , n57072 );
or ( n7740 , n57004 , n7678 );
buf ( n57075 , n7740 );
not ( n57076 , n57075 );
buf ( n57077 , n56912 );
not ( n57078 , n57077 );
or ( n7745 , n57076 , n57078 );
nand ( n57080 , n57004 , n7678 );
buf ( n57081 , n57080 );
nand ( n7748 , n7745 , n57081 );
buf ( n57083 , n7748 );
buf ( n57084 , n57083 );
xor ( n7751 , n57073 , n57084 );
and ( n7752 , n56969 , n6320 );
not ( n57087 , n56969 );
and ( n57088 , n57087 , n6319 );
nor ( n7755 , n7752 , n57088 );
and ( n57090 , n7755 , n7577 );
not ( n7757 , n7755 );
and ( n57092 , n7757 , n56912 );
nor ( n57093 , n57090 , n57092 );
buf ( n57094 , n57093 );
xor ( n57095 , n7751 , n57094 );
buf ( n57096 , n57095 );
buf ( n57097 , n57096 );
buf ( n57098 , n56973 );
not ( n57099 , n57098 );
buf ( n57100 , n57025 );
not ( n57101 , n57100 );
or ( n57102 , n57099 , n57101 );
buf ( n57103 , n7658 );
nand ( n57104 , n57102 , n57103 );
buf ( n57105 , n57104 );
buf ( n57106 , n57105 );
buf ( n57107 , n57025 );
not ( n57108 , n57107 );
buf ( n57109 , n56969 );
nand ( n7776 , n57108 , n57109 );
buf ( n57111 , n7776 );
buf ( n57112 , n57111 );
nand ( n7779 , n57106 , n57112 );
buf ( n57114 , n7779 );
buf ( n57115 , n57114 );
nor ( n7782 , n57097 , n57115 );
buf ( n57117 , n7782 );
buf ( n57118 , n57117 );
not ( n7785 , n57118 );
buf ( n57120 , n7785 );
not ( n7787 , n56424 );
buf ( n57122 , n55678 );
buf ( n57123 , n55642 );
and ( n7790 , n57122 , n57123 );
buf ( n7791 , n7790 );
buf ( n57126 , n7791 );
not ( n7793 , n57126 );
buf ( n57128 , n55643 );
buf ( n57129 , n55681 );
nand ( n7796 , n57128 , n57129 );
buf ( n57131 , n7796 );
buf ( n57132 , n57131 );
nand ( n7799 , n7793 , n57132 );
buf ( n57134 , n7799 );
not ( n7801 , n57134 );
not ( n57136 , n7801 );
or ( n7803 , n7787 , n57136 );
not ( n57138 , n56972 );
nand ( n57139 , n7803 , n57138 );
xor ( n7806 , n6363 , n57139 );
buf ( n57141 , n7791 );
not ( n57142 , n57141 );
buf ( n57143 , n57142 );
xor ( n57144 , n56424 , n57143 );
xor ( n7811 , n57144 , n7801 );
xnor ( n57146 , n7806 , n7811 );
not ( n7813 , n56912 );
not ( n57148 , n56969 );
or ( n7815 , n7813 , n57148 );
nand ( n57150 , n7815 , n6320 );
nand ( n57151 , n56424 , n56969 );
and ( n7818 , n57151 , n7801 );
not ( n57153 , n57151 );
and ( n7820 , n57153 , n57134 );
or ( n7821 , n7818 , n7820 );
buf ( n57156 , n55986 );
buf ( n57157 , n6846 );
nand ( n57158 , n57156 , n57157 );
buf ( n57159 , n57158 );
buf ( n57160 , n55686 );
buf ( n57161 , n55858 );
nand ( n7828 , n57160 , n57161 );
buf ( n7829 , n7828 );
and ( n57164 , n57159 , n7829 );
nand ( n57165 , n7821 , n57164 );
and ( n7832 , n57150 , n57165 );
nor ( n57167 , n7821 , n57164 );
nor ( n7834 , n7832 , n57167 );
nand ( n7835 , n57146 , n7834 );
buf ( n7836 , n7835 );
buf ( n57171 , n7836 );
buf ( n57172 , n57171 );
xor ( n57173 , n57073 , n57084 );
and ( n57174 , n57173 , n57094 );
and ( n7841 , n57073 , n57084 );
or ( n57176 , n57174 , n7841 );
buf ( n57177 , n57176 );
and ( n7844 , n7821 , n57164 );
not ( n7845 , n7821 );
not ( n7846 , n57164 );
and ( n57181 , n7845 , n7846 );
nor ( n57182 , n7844 , n57181 );
xor ( n7849 , n57182 , n57150 );
nor ( n57184 , n57177 , n7849 );
buf ( n57185 , n57184 );
not ( n7852 , n57185 );
buf ( n57187 , n7852 );
nand ( n7854 , n57120 , n57172 , n57187 );
buf ( n57189 , n56424 );
not ( n7856 , n57189 );
buf ( n57191 , n7791 );
not ( n57192 , n57191 );
and ( n57193 , n7856 , n57192 );
buf ( n57194 , n6320 );
not ( n57195 , n57194 );
buf ( n57196 , n57195 );
buf ( n57197 , n57196 );
nor ( n57198 , n57193 , n57197 );
buf ( n57199 , n57198 );
buf ( n57200 , n57199 );
not ( n7867 , n57200 );
buf ( n57202 , n7867 );
buf ( n57203 , n57202 );
not ( n57204 , n57203 );
buf ( n57205 , n55771 );
not ( n57206 , n57205 );
or ( n57207 , n57204 , n57206 );
buf ( n57208 , n55771 );
buf ( n57209 , n57202 );
or ( n7876 , n57208 , n57209 );
nand ( n57211 , n57207 , n7876 );
buf ( n57212 , n57211 );
not ( n7879 , n57212 );
buf ( n57214 , n55762 );
not ( n57215 , n57214 );
buf ( n57216 , n57215 );
buf ( n57217 , n57216 );
not ( n57218 , n57217 );
xnor ( n7885 , n6424 , n57143 );
buf ( n57220 , n7885 );
not ( n57221 , n57220 );
buf ( n57222 , n57221 );
buf ( n57223 , n57222 );
not ( n7890 , n57223 );
or ( n57225 , n57218 , n7890 );
buf ( n57226 , n57143 );
not ( n7893 , n57226 );
buf ( n57228 , n57134 );
not ( n57229 , n57228 );
or ( n7896 , n7893 , n57229 );
buf ( n57231 , n56424 );
nand ( n57232 , n7896 , n57231 );
buf ( n57233 , n57232 );
buf ( n57234 , n57233 );
nand ( n7901 , n57225 , n57234 );
buf ( n57236 , n7901 );
buf ( n57237 , n57236 );
buf ( n57238 , n7885 );
buf ( n57239 , n55762 );
nand ( n7906 , n57238 , n57239 );
buf ( n57241 , n7906 );
buf ( n57242 , n57241 );
nand ( n7909 , n57237 , n57242 );
buf ( n57244 , n7909 );
not ( n7911 , n57244 );
and ( n57246 , n7879 , n7911 );
buf ( n57247 , n55782 );
not ( n57248 , n55762 );
not ( n57249 , n57202 );
or ( n57250 , n57248 , n57249 );
not ( n7917 , n55735 );
not ( n57252 , n57199 );
or ( n7919 , n7917 , n57252 );
nand ( n57254 , n7919 , n6430 );
nand ( n57255 , n57250 , n57254 );
buf ( n57256 , n57255 );
nor ( n57257 , n57247 , n57256 );
buf ( n57258 , n57257 );
nor ( n7925 , n57246 , n57258 );
buf ( n57260 , n7925 );
xor ( n7927 , n55735 , n57233 );
xor ( n7928 , n7927 , n7885 );
buf ( n57263 , n7928 );
not ( n7930 , n57139 );
and ( n7931 , n7811 , n7930 );
nor ( n7932 , n7931 , n55731 );
buf ( n57267 , n7932 );
nand ( n7934 , n57263 , n57267 );
buf ( n57269 , n7934 );
buf ( n57270 , n57269 );
nand ( n57271 , n57260 , n57270 );
buf ( n57272 , n57271 );
nor ( n7939 , n7854 , n57272 );
nand ( n57274 , n57060 , n7939 );
buf ( n57275 , n57274 );
buf ( n57276 , n57048 );
not ( n57277 , n57276 );
buf ( n57278 , n56869 );
nand ( n7945 , n57277 , n57278 );
buf ( n57280 , n7945 );
buf ( n7947 , n57280 );
not ( n57282 , n56468 );
not ( n57283 , n7416 );
nand ( n7950 , n57282 , n57283 );
buf ( n57285 , n7950 );
buf ( n57286 , n57269 );
buf ( n57287 , n7835 );
nand ( n57288 , n57286 , n57287 );
buf ( n57289 , n57288 );
buf ( n57290 , n57289 );
buf ( n57291 , n57117 );
nor ( n7958 , n57290 , n57291 );
buf ( n57293 , n7958 );
buf ( n7960 , n57293 );
buf ( n57295 , n7925 );
buf ( n57296 , n57187 );
nand ( n57297 , n57285 , n7960 , n57295 , n57296 );
buf ( n57298 , n57297 );
buf ( n57299 , n57298 );
nor ( n57300 , n7947 , n57299 );
buf ( n57301 , n57300 );
buf ( n57302 , n57301 );
nand ( n57303 , n377 , n380 );
not ( n57304 , n57303 );
buf ( n57305 , n373 );
buf ( n57306 , n383 );
nand ( n57307 , n57305 , n57306 );
buf ( n57308 , n57307 );
not ( n7975 , n57308 );
buf ( n57310 , n371 );
buf ( n57311 , n385 );
nand ( n7978 , n57310 , n57311 );
buf ( n7979 , n7978 );
not ( n7980 , n7979 );
nand ( n57315 , n7975 , n7980 );
not ( n57316 , n57315 );
or ( n7983 , n57304 , n57316 );
and ( n57318 , n57308 , n7979 );
not ( n7985 , n57318 );
nand ( n57320 , n7983 , n7985 );
and ( n7987 , n7348 , n56687 );
nor ( n57322 , n7987 , n56690 );
and ( n7989 , n57320 , n57322 );
not ( n7990 , n57320 );
buf ( n57325 , n57322 );
not ( n57326 , n57325 );
buf ( n57327 , n57326 );
and ( n7994 , n7990 , n57327 );
nor ( n57329 , n7989 , n7994 );
xor ( n7996 , n56646 , n56641 );
xor ( n7997 , n7996 , n56652 );
and ( n57332 , n57329 , n7997 );
not ( n57333 , n57329 );
not ( n8000 , n7997 );
and ( n57335 , n57333 , n8000 );
nor ( n8002 , n57332 , n57335 );
not ( n57337 , n8002 );
not ( n57338 , n57337 );
buf ( n57339 , n376 );
buf ( n57340 , n382 );
nand ( n57341 , n57339 , n57340 );
buf ( n57342 , n57341 );
buf ( n57343 , n57342 );
buf ( n57344 , n56599 );
or ( n57345 , n57343 , n57344 );
buf ( n57346 , n57345 );
not ( n8013 , n57346 );
buf ( n57348 , n375 );
buf ( n57349 , n381 );
nand ( n57350 , n57348 , n57349 );
buf ( n57351 , n57350 );
buf ( n57352 , n57351 );
buf ( n57353 , n372 );
buf ( n57354 , n384 );
nand ( n8021 , n57353 , n57354 );
buf ( n57356 , n8021 );
buf ( n57357 , n57356 );
or ( n8024 , n57352 , n57357 );
buf ( n8025 , n377 );
buf ( n8026 , n379 );
nand ( n8027 , n8025 , n8026 );
buf ( n8028 , n8027 );
buf ( n57363 , n8028 );
nand ( n8030 , n8024 , n57363 );
buf ( n57365 , n8030 );
buf ( n57366 , n57365 );
buf ( n57367 , n57351 );
buf ( n57368 , n57356 );
nand ( n57369 , n57367 , n57368 );
buf ( n57370 , n57369 );
buf ( n57371 , n57370 );
nand ( n57372 , n57366 , n57371 );
buf ( n57373 , n57372 );
not ( n57374 , n57373 );
not ( n57375 , n57374 );
or ( n57376 , n8013 , n57375 );
or ( n8043 , n57374 , n57346 );
nand ( n57378 , n57376 , n8043 );
not ( n8045 , n57378 );
xor ( n57380 , n56697 , n56702 );
xor ( n8047 , n57380 , n56708 );
buf ( n57382 , n8047 );
not ( n8049 , n57382 );
not ( n8050 , n8049 );
or ( n57385 , n8045 , n8050 );
and ( n57386 , n57346 , n57373 );
not ( n8053 , n57346 );
and ( n57388 , n8053 , n57374 );
nor ( n57389 , n57386 , n57388 );
or ( n8056 , n8049 , n57389 );
nand ( n57391 , n57385 , n8056 );
not ( n57392 , n57391 );
or ( n57393 , n57338 , n57392 );
not ( n8060 , n8002 );
buf ( n57395 , n57391 );
not ( n8062 , n57395 );
buf ( n57397 , n8062 );
not ( n57398 , n57397 );
or ( n57399 , n8060 , n57398 );
xor ( n8066 , n57356 , n57351 );
xor ( n8067 , n8066 , n8028 );
not ( n57402 , n8067 );
buf ( n57403 , n376 );
buf ( n57404 , n381 );
nand ( n57405 , n57403 , n57404 );
buf ( n57406 , n57405 );
buf ( n57407 , n57406 );
buf ( n57408 , n374 );
buf ( n57409 , n383 );
nand ( n8076 , n57408 , n57409 );
buf ( n57411 , n8076 );
buf ( n57412 , n57411 );
or ( n57413 , n57407 , n57412 );
buf ( n57414 , n372 );
buf ( n57415 , n385 );
nand ( n57416 , n57414 , n57415 );
buf ( n57417 , n57416 );
buf ( n57418 , n57417 );
nand ( n57419 , n57413 , n57418 );
buf ( n57420 , n57419 );
buf ( n57421 , n57420 );
buf ( n57422 , n57406 );
buf ( n57423 , n57411 );
nand ( n57424 , n57422 , n57423 );
buf ( n57425 , n57424 );
buf ( n57426 , n57425 );
and ( n57427 , n57421 , n57426 );
buf ( n57428 , n57427 );
buf ( n57429 , n57428 );
not ( n57430 , n57429 );
buf ( n57431 , n57430 );
not ( n8098 , n57431 );
or ( n57433 , n57402 , n8098 );
not ( n57434 , n57428 );
not ( n8101 , n8067 );
not ( n57436 , n8101 );
or ( n8103 , n57434 , n57436 );
buf ( n8104 , n374 );
buf ( n57439 , n382 );
nand ( n57440 , n8104 , n57439 );
buf ( n57441 , n57440 );
buf ( n57442 , n57441 );
not ( n8109 , n57442 );
buf ( n8110 , n376 );
buf ( n57445 , n380 );
nand ( n57446 , n8110 , n57445 );
buf ( n57447 , n57446 );
buf ( n57448 , n57447 );
not ( n57449 , n57448 );
or ( n8116 , n8109 , n57449 );
buf ( n57451 , n57346 );
nand ( n57452 , n8116 , n57451 );
buf ( n57453 , n57452 );
nand ( n57454 , n8103 , n57453 );
nand ( n57455 , n57433 , n57454 );
nand ( n8122 , n57399 , n57455 );
nand ( n57457 , n57393 , n8122 );
buf ( n8124 , n57457 );
not ( n8125 , n8124 );
buf ( n57460 , n56589 );
buf ( n57461 , n56586 );
buf ( n57462 , n56581 );
nand ( n8129 , n57461 , n57462 );
buf ( n57464 , n8129 );
buf ( n57465 , n57464 );
and ( n57466 , n57460 , n57465 );
buf ( n57467 , n57466 );
xor ( n8134 , n56631 , n56636 );
xor ( n57469 , n8134 , n56664 );
buf ( n57470 , n57469 );
xor ( n57471 , n57467 , n57470 );
not ( n8138 , n57373 );
not ( n8139 , n57346 );
or ( n57474 , n8138 , n8139 );
not ( n8141 , n57374 );
nor ( n57476 , n8141 , n57346 );
or ( n8143 , n57476 , n8049 );
nand ( n57478 , n57474 , n8143 );
xor ( n8145 , n57471 , n57478 );
not ( n8146 , n8145 );
nand ( n57481 , n56712 , n7343 , n56717 );
not ( n8148 , n7357 );
nand ( n57483 , n8148 , n56712 );
not ( n8150 , n56712 );
nand ( n8151 , n8150 , n7343 , n56690 );
nor ( n8152 , n7343 , n56690 );
nand ( n8153 , n8150 , n8152 );
nand ( n8154 , n57481 , n57483 , n8151 , n8153 );
not ( n8155 , n8154 );
not ( n8156 , n57327 );
not ( n8157 , n57320 );
or ( n57492 , n8156 , n8157 );
or ( n8159 , n57327 , n57320 );
nand ( n8160 , n8159 , n7997 );
nand ( n8161 , n57492 , n8160 );
not ( n8162 , n8161 );
and ( n8163 , n8155 , n8162 );
not ( n8164 , n8155 );
and ( n8165 , n8164 , n8161 );
nor ( n8166 , n8163 , n8165 );
xor ( n8167 , n8146 , n8166 );
not ( n8168 , n8167 );
not ( n8169 , n8168 );
not ( n57504 , n8169 );
or ( n8171 , n8125 , n57504 );
not ( n57506 , n8124 );
not ( n57507 , n57506 );
not ( n8174 , n8168 );
or ( n57509 , n57507 , n8174 );
not ( n57510 , n55858 );
buf ( n57511 , n6116 );
not ( n8178 , n57511 );
buf ( n57513 , n8178 );
buf ( n57514 , n57513 );
not ( n57515 , n57514 );
or ( n57516 , n6102 , n6095 );
buf ( n57517 , n57516 );
nand ( n57518 , n57515 , n57517 );
buf ( n57519 , n57518 );
not ( n8186 , n57519 );
not ( n8187 , n8186 );
not ( n8188 , n6645 );
or ( n57523 , n8187 , n8188 );
buf ( n57524 , n6882 );
buf ( n8191 , n57519 );
nand ( n8192 , n57524 , n8191 );
buf ( n8193 , n8192 );
nand ( n8194 , n57523 , n8193 );
buf ( n8195 , n8194 );
not ( n57530 , n8195 );
or ( n8197 , n57510 , n57530 );
buf ( n57532 , n55355 );
buf ( n57533 , n55350 );
and ( n57534 , n57532 , n57533 );
buf ( n57535 , n57534 );
buf ( n57536 , n57535 );
buf ( n57537 , n55283 );
not ( n8204 , n57537 );
buf ( n57539 , n5919 );
not ( n8206 , n57539 );
or ( n57541 , n8204 , n8206 );
buf ( n57542 , n55288 );
nand ( n57543 , n57541 , n57542 );
buf ( n57544 , n57543 );
buf ( n57545 , n57544 );
and ( n57546 , n57536 , n57545 );
not ( n8213 , n57536 );
buf ( n57548 , n57544 );
not ( n8215 , n57548 );
buf ( n57550 , n8215 );
buf ( n57551 , n57550 );
and ( n57552 , n8213 , n57551 );
nor ( n57553 , n57546 , n57552 );
buf ( n57554 , n57553 );
not ( n57555 , n57554 );
or ( n8222 , n57555 , n6530 );
nand ( n8223 , n8197 , n8222 );
nand ( n8224 , n57509 , n8223 );
nand ( n8225 , n8171 , n8224 );
not ( n8226 , n8161 );
not ( n8227 , n8154 );
or ( n8228 , n8226 , n8227 );
buf ( n57563 , n8161 );
not ( n8230 , n57563 );
buf ( n57565 , n8155 );
nand ( n8232 , n8230 , n57565 );
buf ( n57567 , n8232 );
nand ( n8234 , n8146 , n57567 );
nand ( n8235 , n8228 , n8234 );
not ( n8236 , n8235 );
not ( n8237 , n8236 );
xor ( n8238 , n7243 , n56589 );
xor ( n8239 , n8238 , n7278 );
buf ( n57574 , n8239 );
buf ( n57575 , n57467 );
not ( n8242 , n57575 );
buf ( n57577 , n57470 );
not ( n8244 , n57577 );
buf ( n57579 , n8244 );
buf ( n57580 , n57579 );
not ( n8247 , n57580 );
or ( n8248 , n8242 , n8247 );
buf ( n57583 , n57478 );
nand ( n8250 , n8248 , n57583 );
buf ( n57585 , n8250 );
buf ( n57586 , n57585 );
buf ( n57587 , n57467 );
not ( n8254 , n57587 );
buf ( n57589 , n57470 );
nand ( n8256 , n8254 , n57589 );
buf ( n57591 , n8256 );
buf ( n57592 , n57591 );
nand ( n8259 , n57586 , n57592 );
buf ( n57594 , n8259 );
buf ( n57595 , n57594 );
xor ( n8262 , n57574 , n57595 );
xor ( n8263 , n56626 , n56669 );
xor ( n8264 , n8263 , n56720 );
buf ( n57599 , n8264 );
buf ( n57600 , n57599 );
xor ( n8267 , n8262 , n57600 );
buf ( n57602 , n8267 );
not ( n8269 , n57602 );
or ( n8270 , n8237 , n8269 );
not ( n8271 , n57602 );
nand ( n8272 , n8235 , n8271 );
nand ( n8273 , n8270 , n8272 );
not ( n8274 , n6846 );
not ( n8275 , n8194 );
not ( n8276 , n8275 );
not ( n8277 , n8276 );
or ( n8278 , n8274 , n8277 );
buf ( n57613 , n55361 );
buf ( n57614 , n6082 );
or ( n57615 , n57613 , n57614 );
buf ( n57616 , n57615 );
buf ( n57617 , n57616 );
buf ( n57618 , n55437 );
nand ( n57619 , n57617 , n57618 );
buf ( n57620 , n57619 );
buf ( n57621 , n57620 );
not ( n57622 , n57621 );
buf ( n57623 , n57622 );
not ( n8290 , n57623 );
buf ( n57625 , n57544 );
not ( n57626 , n57625 );
buf ( n57627 , n55428 );
buf ( n57628 , n6031 );
nor ( n57629 , n57627 , n57628 );
buf ( n57630 , n57629 );
buf ( n57631 , n57630 );
not ( n8298 , n57631 );
or ( n57633 , n57626 , n8298 );
buf ( n57634 , n57516 );
buf ( n57635 , n55350 );
not ( n57636 , n57635 );
buf ( n57637 , n57636 );
buf ( n57638 , n57637 );
and ( n8305 , n57634 , n57638 );
buf ( n57640 , n57513 );
nor ( n8307 , n8305 , n57640 );
buf ( n57642 , n8307 );
buf ( n57643 , n57642 );
nand ( n8310 , n57633 , n57643 );
buf ( n8311 , n8310 );
buf ( n57646 , n8311 );
not ( n8313 , n57646 );
buf ( n57648 , n8313 );
not ( n8315 , n57648 );
or ( n8316 , n8290 , n8315 );
buf ( n57651 , n8311 );
buf ( n57652 , n57620 );
nand ( n8319 , n57651 , n57652 );
buf ( n57654 , n8319 );
nand ( n8321 , n8316 , n57654 );
nand ( n8322 , n8321 , n55858 );
nand ( n57657 , n8278 , n8322 );
xor ( n8324 , n8273 , n57657 );
xor ( n57659 , n8225 , n8324 );
buf ( n57660 , n6980 );
not ( n8327 , n57660 );
buf ( n57662 , n411 );
buf ( n8329 , n56238 );
and ( n8330 , n57662 , n8329 );
not ( n57665 , n57662 );
buf ( n57666 , n56238 );
not ( n8333 , n57666 );
buf ( n8334 , n8333 );
buf ( n57669 , n8334 );
and ( n8336 , n57665 , n57669 );
nor ( n8337 , n8330 , n8336 );
buf ( n57672 , n8337 );
buf ( n57673 , n57672 );
not ( n8340 , n57673 );
or ( n8341 , n8327 , n8340 );
buf ( n57676 , n56072 );
buf ( n8343 , n7168 );
not ( n57678 , n8343 );
buf ( n57679 , n57678 );
and ( n57680 , n411 , n57679 );
not ( n8347 , n411 );
and ( n8348 , n8347 , n7168 );
or ( n8349 , n57680 , n8348 );
buf ( n57684 , n8349 );
nand ( n8351 , n57676 , n57684 );
buf ( n57686 , n8351 );
buf ( n57687 , n57686 );
nand ( n8354 , n8341 , n57687 );
buf ( n57689 , n8354 );
xor ( n8356 , n57659 , n57689 );
not ( n8357 , n8356 );
and ( n8358 , n57457 , n8167 );
not ( n8359 , n57457 );
and ( n57694 , n8166 , n8145 );
not ( n57695 , n8166 );
and ( n8362 , n57695 , n8146 );
nor ( n57697 , n57694 , n8362 );
and ( n8364 , n8359 , n57697 );
nor ( n8365 , n8358 , n8364 );
not ( n8366 , n8365 );
not ( n8367 , n8223 );
or ( n8368 , n8366 , n8367 );
or ( n8369 , n8223 , n8365 );
nand ( n8370 , n8368 , n8369 );
buf ( n57705 , n8370 );
buf ( n57706 , n6591 );
not ( n8373 , n57706 );
buf ( n57708 , n413 );
not ( n57709 , n57708 );
buf ( n57710 , n8334 );
not ( n57711 , n57710 );
or ( n57712 , n57709 , n57711 );
buf ( n57713 , n55646 );
buf ( n57714 , n56238 );
nand ( n57715 , n57713 , n57714 );
buf ( n57716 , n57715 );
buf ( n57717 , n57716 );
nand ( n8384 , n57712 , n57717 );
buf ( n57719 , n8384 );
buf ( n57720 , n57719 );
not ( n57721 , n57720 );
or ( n57722 , n8373 , n57721 );
not ( n8389 , n7228 );
not ( n57724 , n413 );
or ( n57725 , n8389 , n57724 );
buf ( n8392 , n56200 );
buf ( n8393 , n6322 );
nand ( n8394 , n8392 , n8393 );
buf ( n8395 , n8394 );
nand ( n57730 , n57725 , n8395 );
buf ( n57731 , n57730 );
buf ( n57732 , n6665 );
nand ( n57733 , n57731 , n57732 );
buf ( n57734 , n57733 );
buf ( n57735 , n57734 );
nand ( n8402 , n57722 , n57735 );
buf ( n57737 , n8402 );
buf ( n57738 , n57737 );
not ( n8405 , n57738 );
buf ( n57740 , n8405 );
buf ( n57741 , n57740 );
xor ( n8408 , n57705 , n57741 );
not ( n57743 , n7015 );
not ( n8410 , n6528 );
or ( n57745 , n57743 , n8410 );
or ( n8412 , n6528 , n7015 );
nand ( n57747 , n57745 , n8412 );
not ( n57748 , n57747 );
not ( n57749 , n55712 );
and ( n8416 , n57748 , n57749 );
not ( n57751 , n415 );
not ( n8418 , n6587 );
or ( n57753 , n57751 , n8418 );
or ( n57754 , n6587 , n415 );
nand ( n8421 , n57753 , n57754 );
and ( n57756 , n8421 , n416 );
nor ( n57757 , n8416 , n57756 );
buf ( n57758 , n57757 );
and ( n8425 , n8408 , n57758 );
and ( n57760 , n57705 , n57741 );
or ( n57761 , n8425 , n57760 );
buf ( n57762 , n57761 );
buf ( n57763 , n57762 );
not ( n57764 , n57763 );
buf ( n57765 , n57764 );
not ( n8432 , n57765 );
or ( n57767 , n8357 , n8432 );
buf ( n57768 , n6591 );
not ( n8435 , n57768 );
buf ( n57770 , n57730 );
not ( n57771 , n57770 );
or ( n8438 , n8435 , n57771 );
not ( n8439 , n6322 );
not ( n57774 , n6528 );
or ( n57775 , n8439 , n57774 );
and ( n8442 , n413 , n56204 );
not ( n57777 , n6665 );
nor ( n57778 , n8442 , n57777 );
nand ( n8445 , n57775 , n57778 );
buf ( n57780 , n8445 );
nand ( n57781 , n8438 , n57780 );
buf ( n57782 , n57781 );
buf ( n57783 , n8349 );
buf ( n57784 , n6980 );
and ( n57785 , n57783 , n57784 );
not ( n8452 , n411 );
not ( n57787 , n8321 );
not ( n57788 , n57787 );
or ( n8455 , n8452 , n57788 );
not ( n57790 , n8321 );
or ( n8457 , n57790 , n411 );
nand ( n8458 , n8455 , n8457 );
buf ( n57793 , n8458 );
not ( n8460 , n57793 );
buf ( n57795 , n6312 );
nor ( n8462 , n8460 , n57795 );
buf ( n57797 , n8462 );
buf ( n57798 , n57797 );
nor ( n8465 , n57785 , n57798 );
buf ( n57800 , n8465 );
buf ( n57801 , n57800 );
not ( n8468 , n57801 );
buf ( n57803 , n8468 );
not ( n8470 , n57803 );
buf ( n57805 , n374 );
buf ( n57806 , n384 );
nand ( n8473 , n57805 , n57806 );
buf ( n57808 , n8473 );
buf ( n57809 , n57808 );
not ( n57810 , n57809 );
buf ( n8477 , n375 );
buf ( n57812 , n383 );
nand ( n57813 , n8477 , n57812 );
buf ( n57814 , n57813 );
buf ( n57815 , n57814 );
not ( n57816 , n57815 );
or ( n8483 , n57810 , n57816 );
buf ( n57818 , n57814 );
buf ( n57819 , n57808 );
or ( n8486 , n57818 , n57819 );
buf ( n57821 , n377 );
buf ( n57822 , n381 );
nand ( n8489 , n57821 , n57822 );
buf ( n57824 , n8489 );
buf ( n57825 , n57824 );
nand ( n8492 , n8486 , n57825 );
buf ( n57827 , n8492 );
buf ( n57828 , n57827 );
nand ( n8495 , n8483 , n57828 );
buf ( n57830 , n8495 );
not ( n57831 , n57830 );
buf ( n8498 , n373 );
buf ( n57833 , n385 );
nand ( n57834 , n8498 , n57833 );
buf ( n57835 , n57834 );
buf ( n57836 , n57835 );
buf ( n8503 , n57342 );
or ( n8504 , n57836 , n8503 );
buf ( n57839 , n8504 );
not ( n57840 , n57839 );
nand ( n8507 , n57831 , n57840 );
not ( n57842 , n8507 );
xor ( n57843 , n57417 , n57406 );
xor ( n57844 , n57843 , n57411 );
not ( n8511 , n57844 );
or ( n57846 , n57842 , n8511 );
or ( n8513 , n57831 , n57840 );
nand ( n8514 , n57846 , n8513 );
not ( n8515 , n8514 );
not ( n8516 , n57303 );
and ( n8517 , n7980 , n57308 , n8516 );
not ( n8518 , n8517 );
and ( n57853 , n7975 , n7979 , n8516 );
not ( n8520 , n57853 );
nand ( n57855 , n57318 , n57303 );
nand ( n8522 , n7980 , n7975 , n57303 );
nand ( n8523 , n8518 , n8520 , n57855 , n8522 );
buf ( n57858 , n8523 );
not ( n8525 , n57858 );
buf ( n57860 , n373 );
buf ( n57861 , n384 );
nand ( n8528 , n57860 , n57861 );
buf ( n57863 , n8528 );
buf ( n57864 , n57863 );
not ( n8531 , n57864 );
buf ( n57866 , n375 );
buf ( n57867 , n382 );
nand ( n8534 , n57866 , n57867 );
buf ( n57869 , n8534 );
buf ( n57870 , n57869 );
not ( n8537 , n57870 );
buf ( n57872 , n8537 );
buf ( n57873 , n57872 );
nand ( n8540 , n8531 , n57873 );
buf ( n57875 , n8540 );
buf ( n57876 , n57875 );
nand ( n57877 , n377 , n380 );
buf ( n57878 , n57877 );
not ( n57879 , n57878 );
buf ( n57880 , n57879 );
buf ( n57881 , n57880 );
and ( n8548 , n57876 , n57881 );
buf ( n57883 , n57869 );
buf ( n57884 , n57863 );
and ( n8551 , n57883 , n57884 );
buf ( n57886 , n8551 );
buf ( n57887 , n57886 );
nor ( n8554 , n8548 , n57887 );
buf ( n57889 , n8554 );
buf ( n57890 , n57889 );
nand ( n8557 , n8525 , n57890 );
buf ( n57892 , n8557 );
not ( n8559 , n57892 );
or ( n8560 , n8515 , n8559 );
buf ( n57895 , n57889 );
not ( n8562 , n57895 );
buf ( n57897 , n8523 );
nand ( n8564 , n8562 , n57897 );
buf ( n57899 , n8564 );
nand ( n8566 , n8560 , n57899 );
not ( n8567 , n8566 );
and ( n57902 , n57455 , n57397 );
not ( n57903 , n57455 );
and ( n8570 , n57903 , n57391 );
or ( n57905 , n57902 , n8570 );
and ( n57906 , n57905 , n8002 );
not ( n8573 , n57905 );
and ( n57908 , n8573 , n57337 );
nor ( n8575 , n57906 , n57908 );
nand ( n8576 , n8567 , n8575 );
buf ( n57911 , n8576 );
not ( n8578 , n57911 );
and ( n8579 , n57453 , n57428 );
not ( n57914 , n57453 );
and ( n8581 , n57914 , n57431 );
or ( n8582 , n8579 , n8581 );
and ( n8583 , n8582 , n8067 );
not ( n8584 , n8582 );
and ( n8585 , n8584 , n8101 );
nor ( n8586 , n8583 , n8585 );
buf ( n57921 , n8586 );
not ( n8588 , n57921 );
not ( n8589 , n5931 );
not ( n8590 , n5947 );
or ( n8591 , n8589 , n8590 );
nand ( n8592 , n8591 , n5957 );
not ( n8593 , n8592 );
nand ( n8594 , n5919 , n55288 );
not ( n8595 , n8594 );
or ( n8596 , n8593 , n8595 );
buf ( n8597 , n55283 );
or ( n8598 , n8594 , n8597 );
nand ( n8599 , n8596 , n8598 );
buf ( n57934 , n8599 );
buf ( n8601 , n57934 );
buf ( n57936 , n8601 );
buf ( n57937 , n57936 );
buf ( n57938 , n55858 );
nand ( n8605 , n57937 , n57938 );
buf ( n57940 , n8605 );
buf ( n57941 , n57940 );
not ( n8608 , n57941 );
buf ( n57943 , n8608 );
buf ( n57944 , n57943 );
not ( n8611 , n57944 );
or ( n8612 , n8588 , n8611 );
buf ( n57947 , n8586 );
not ( n8614 , n57947 );
buf ( n57949 , n8614 );
buf ( n57950 , n57949 );
not ( n8617 , n57950 );
buf ( n57952 , n57940 );
not ( n8619 , n57952 );
or ( n8620 , n8617 , n8619 );
not ( n57955 , n8514 );
not ( n8622 , n57955 );
not ( n8623 , n8523 );
not ( n8624 , n8623 );
not ( n8625 , n57889 );
or ( n57960 , n8624 , n8625 );
or ( n8627 , n57889 , n8623 );
nand ( n57962 , n57960 , n8627 );
not ( n8629 , n57962 );
or ( n57964 , n8622 , n8629 );
or ( n57965 , n57955 , n57962 );
nand ( n57966 , n57964 , n57965 );
buf ( n57967 , n57966 );
not ( n57968 , n57967 );
buf ( n57969 , n57968 );
buf ( n57970 , n57969 );
nand ( n8637 , n8620 , n57970 );
buf ( n8638 , n8637 );
buf ( n8639 , n8638 );
nand ( n8640 , n8612 , n8639 );
buf ( n8641 , n8640 );
buf ( n57976 , n8641 );
not ( n57977 , n57976 );
or ( n8644 , n8578 , n57977 );
and ( n57979 , n57905 , n57337 );
not ( n57980 , n57905 );
not ( n8647 , n57337 );
and ( n8648 , n57980 , n8647 );
nor ( n8649 , n57979 , n8648 );
nand ( n8650 , n8649 , n8566 );
buf ( n57985 , n8650 );
nand ( n8652 , n8644 , n57985 );
buf ( n57987 , n8652 );
not ( n57988 , n57987 );
or ( n57989 , n8470 , n57988 );
not ( n8656 , n57987 );
not ( n57991 , n8656 );
not ( n8658 , n57800 );
or ( n8659 , n57991 , n8658 );
buf ( n57994 , n55858 );
not ( n57995 , n57994 );
buf ( n57996 , n57554 );
not ( n57997 , n57996 );
or ( n57998 , n57995 , n57997 );
buf ( n57999 , n8599 );
not ( n58000 , n57999 );
buf ( n58001 , n58000 );
buf ( n58002 , n58001 );
not ( n8669 , n58002 );
buf ( n58004 , n8669 );
buf ( n58005 , n58004 );
buf ( n58006 , n6846 );
nand ( n8673 , n58005 , n58006 );
buf ( n58008 , n8673 );
buf ( n58009 , n58008 );
nand ( n8676 , n57998 , n58009 );
buf ( n58011 , n8676 );
buf ( n58012 , n6980 );
not ( n8679 , n58012 );
buf ( n58014 , n8458 );
not ( n8681 , n58014 );
or ( n8682 , n8679 , n8681 );
not ( n8683 , n411 );
not ( n8684 , n8275 );
or ( n58019 , n8683 , n8684 );
not ( n8686 , n8186 );
not ( n8687 , n6645 );
or ( n8688 , n8686 , n8687 );
nand ( n58023 , n8688 , n8193 );
nand ( n8690 , n58023 , n56768 );
nand ( n58025 , n58019 , n8690 );
nand ( n58026 , n58025 , n56072 );
buf ( n58027 , n58026 );
nand ( n58028 , n8682 , n58027 );
buf ( n58029 , n58028 );
xor ( n8696 , n58011 , n58029 );
not ( n58031 , n8649 );
not ( n58032 , n8566 );
and ( n8699 , n58031 , n58032 );
and ( n8700 , n8649 , n8566 );
nor ( n8701 , n8699 , n8700 );
and ( n8702 , n8701 , n8641 );
not ( n58037 , n8701 );
not ( n8704 , n8641 );
and ( n58039 , n58037 , n8704 );
nor ( n8706 , n8702 , n58039 );
and ( n58041 , n8696 , n8706 );
and ( n8708 , n58011 , n58029 );
or ( n8709 , n58041 , n8708 );
nand ( n58044 , n8659 , n8709 );
nand ( n8711 , n57989 , n58044 );
xor ( n58046 , n57782 , n8711 );
buf ( n58047 , n416 );
not ( n58048 , n58047 );
xor ( n8715 , n415 , n7028 );
buf ( n58050 , n8715 );
not ( n58051 , n58050 );
or ( n8718 , n58048 , n58051 );
buf ( n58053 , n8421 );
buf ( n58054 , n6384 );
nand ( n8721 , n58053 , n58054 );
buf ( n58056 , n8721 );
buf ( n58057 , n58056 );
nand ( n8724 , n8718 , n58057 );
buf ( n58059 , n8724 );
xor ( n8726 , n58046 , n58059 );
buf ( n58061 , n8726 );
buf ( n58062 , n8356 );
not ( n8729 , n58062 );
buf ( n58064 , n57762 );
nand ( n8731 , n8729 , n58064 );
buf ( n58066 , n8731 );
buf ( n58067 , n58066 );
nand ( n8734 , n58061 , n58067 );
buf ( n58069 , n8734 );
nand ( n8736 , n57767 , n58069 );
buf ( n58071 , n8736 );
not ( n8738 , n58071 );
buf ( n58073 , n8738 );
not ( n8740 , n58073 );
not ( n58075 , n57657 );
nand ( n8742 , n8271 , n8236 );
not ( n8743 , n8742 );
or ( n8744 , n58075 , n8743 );
nand ( n8745 , n8235 , n57602 );
nand ( n58080 , n8744 , n8745 );
buf ( n58081 , n58080 );
buf ( n58082 , n56072 );
not ( n8749 , n58082 );
buf ( n58084 , n57672 );
not ( n58085 , n58084 );
or ( n58086 , n8749 , n58085 );
nand ( n8753 , n6980 , n56566 );
buf ( n58088 , n8753 );
nand ( n8755 , n58086 , n58088 );
buf ( n58090 , n8755 );
buf ( n58091 , n58090 );
xor ( n8758 , n58081 , n58091 );
not ( n8759 , n6665 );
not ( n8760 , n56542 );
or ( n8761 , n8759 , n8760 );
not ( n58096 , n6528 );
not ( n8763 , n413 );
or ( n8764 , n58096 , n8763 );
or ( n8765 , n413 , n6528 );
nand ( n8766 , n8764 , n8765 );
nand ( n8767 , n8766 , n6591 );
nand ( n8768 , n8761 , n8767 );
buf ( n58103 , n8768 );
xnor ( n8770 , n8758 , n58103 );
buf ( n58105 , n8770 );
buf ( n58106 , n58105 );
xor ( n58107 , n57782 , n8711 );
and ( n8774 , n58107 , n58059 );
and ( n58109 , n57782 , n8711 );
or ( n8776 , n8774 , n58109 );
buf ( n58111 , n8776 );
xor ( n58112 , n58106 , n58111 );
xor ( n8779 , n57574 , n57595 );
and ( n58114 , n8779 , n57600 );
and ( n58115 , n57574 , n57595 );
or ( n8782 , n58114 , n58115 );
buf ( n58117 , n8782 );
xor ( n58118 , n7281 , n7287 );
xor ( n8785 , n58118 , n56724 );
not ( n8786 , n8785 );
xor ( n8787 , n58117 , n8786 );
not ( n58122 , n55858 );
not ( n8789 , n7168 );
or ( n58124 , n58122 , n8789 );
nand ( n8791 , n8321 , n6846 );
nand ( n58126 , n58124 , n8791 );
xnor ( n8793 , n8787 , n58126 );
buf ( n58128 , n8793 );
buf ( n58129 , n6384 );
not ( n58130 , n58129 );
buf ( n58131 , n8715 );
not ( n58132 , n58131 );
or ( n8799 , n58130 , n58132 );
buf ( n58134 , n56516 );
buf ( n8801 , n416 );
nand ( n8802 , n58134 , n8801 );
buf ( n8803 , n8802 );
buf ( n58138 , n8803 );
nand ( n8805 , n8799 , n58138 );
buf ( n58140 , n8805 );
buf ( n58141 , n58140 );
xor ( n58142 , n58128 , n58141 );
xor ( n8809 , n8225 , n8324 );
and ( n58144 , n8809 , n57689 );
and ( n58145 , n8225 , n8324 );
or ( n8812 , n58144 , n58145 );
buf ( n58147 , n8812 );
xnor ( n8814 , n58142 , n58147 );
buf ( n58149 , n8814 );
buf ( n58150 , n58149 );
xnor ( n8817 , n58112 , n58150 );
buf ( n8818 , n8817 );
not ( n58153 , n8818 );
or ( n8820 , n8740 , n58153 );
buf ( n58155 , n57762 );
buf ( n58156 , n8356 );
nor ( n8823 , n58155 , n58156 );
buf ( n58158 , n8823 );
buf ( n58159 , n58158 );
not ( n58160 , n58159 );
buf ( n58161 , n8356 );
buf ( n58162 , n57762 );
nand ( n58163 , n58161 , n58162 );
buf ( n58164 , n58163 );
buf ( n58165 , n58164 );
nand ( n8832 , n58160 , n58165 );
buf ( n58167 , n8832 );
buf ( n58168 , n58167 );
buf ( n58169 , n8726 );
not ( n58170 , n58169 );
buf ( n58171 , n58170 );
buf ( n58172 , n58171 );
and ( n58173 , n58168 , n58172 );
not ( n8840 , n58168 );
buf ( n8841 , n8726 );
and ( n58176 , n8840 , n8841 );
nor ( n8843 , n58173 , n58176 );
buf ( n8844 , n8843 );
buf ( n8845 , n57987 );
buf ( n8846 , n57803 );
xor ( n8847 , n8845 , n8846 );
buf ( n58182 , n8709 );
xnor ( n8849 , n8847 , n58182 );
buf ( n58184 , n8849 );
buf ( n58185 , n58184 );
buf ( n58186 , n6665 );
not ( n58187 , n58186 );
buf ( n58188 , n57719 );
not ( n8855 , n58188 );
or ( n8856 , n58187 , n8855 );
buf ( n58191 , n413 );
not ( n8858 , n58191 );
buf ( n58193 , n57679 );
not ( n8860 , n58193 );
or ( n8861 , n8858 , n8860 );
buf ( n58196 , n7168 );
buf ( n58197 , n6322 );
nand ( n8864 , n58196 , n58197 );
buf ( n58199 , n8864 );
buf ( n58200 , n58199 );
nand ( n8867 , n8861 , n58200 );
buf ( n58202 , n8867 );
buf ( n58203 , n58202 );
buf ( n58204 , n6591 );
nand ( n8871 , n58203 , n58204 );
buf ( n58206 , n8871 );
buf ( n58207 , n58206 );
nand ( n8874 , n8856 , n58207 );
buf ( n58209 , n8874 );
buf ( n58210 , n58209 );
not ( n8877 , n58210 );
buf ( n58212 , n8877 );
not ( n8879 , n58212 );
buf ( n58214 , n57863 );
not ( n58215 , n58214 );
buf ( n58216 , n57872 );
not ( n8883 , n58216 );
or ( n58218 , n58215 , n8883 );
buf ( n58219 , n57863 );
buf ( n58220 , n57872 );
or ( n58221 , n58219 , n58220 );
nand ( n8888 , n58218 , n58221 );
buf ( n8889 , n8888 );
buf ( n58224 , n8889 );
buf ( n58225 , n57880 );
and ( n8892 , n58224 , n58225 );
not ( n58227 , n58224 );
buf ( n58228 , n57877 );
and ( n8895 , n58227 , n58228 );
nor ( n8896 , n8892 , n8895 );
buf ( n58231 , n8896 );
buf ( n58232 , n57824 );
buf ( n58233 , n57814 );
xor ( n8900 , n58232 , n58233 );
buf ( n58235 , n57808 );
xor ( n58236 , n8900 , n58235 );
buf ( n58237 , n58236 );
not ( n58238 , n58237 );
buf ( n58239 , n375 );
buf ( n58240 , n384 );
nand ( n58241 , n58239 , n58240 );
buf ( n58242 , n58241 );
buf ( n58243 , n58242 );
not ( n8910 , n58243 );
buf ( n58245 , n376 );
buf ( n58246 , n383 );
nand ( n58247 , n58245 , n58246 );
buf ( n58248 , n58247 );
buf ( n58249 , n58248 );
not ( n58250 , n58249 );
or ( n58251 , n8910 , n58250 );
buf ( n58252 , n58248 );
buf ( n58253 , n58242 );
or ( n58254 , n58252 , n58253 );
buf ( n58255 , n377 );
buf ( n58256 , n382 );
nand ( n8923 , n58255 , n58256 );
buf ( n58258 , n8923 );
buf ( n58259 , n58258 );
nand ( n8926 , n58254 , n58259 );
buf ( n58261 , n8926 );
buf ( n58262 , n58261 );
nand ( n8929 , n58251 , n58262 );
buf ( n58264 , n8929 );
buf ( n58265 , n58264 );
not ( n8932 , n58265 );
buf ( n58267 , n374 );
buf ( n58268 , n385 );
nand ( n58269 , n58267 , n58268 );
buf ( n58270 , n58269 );
buf ( n58271 , n58270 );
not ( n8938 , n58271 );
buf ( n58273 , n8938 );
buf ( n58274 , n58273 );
nand ( n58275 , n8932 , n58274 );
buf ( n58276 , n58275 );
not ( n58277 , n58276 );
or ( n8944 , n58238 , n58277 );
buf ( n58279 , n58264 );
buf ( n58280 , n58270 );
nand ( n58281 , n58279 , n58280 );
buf ( n58282 , n58281 );
nand ( n58283 , n8944 , n58282 );
xor ( n8950 , n58231 , n58283 );
and ( n8951 , n57840 , n57831 );
not ( n8952 , n57840 );
and ( n8953 , n8952 , n57830 );
nor ( n8954 , n8951 , n8953 );
and ( n8955 , n8954 , n57844 );
not ( n8956 , n8954 );
not ( n8957 , n57844 );
and ( n8958 , n8956 , n8957 );
nor ( n8959 , n8955 , n8958 );
and ( n58294 , n8950 , n8959 );
and ( n58295 , n58231 , n58283 );
or ( n8962 , n58294 , n58295 );
buf ( n58297 , n8962 );
not ( n58298 , n58297 );
buf ( n58299 , n58298 );
buf ( n58300 , n58299 );
not ( n8967 , n58300 );
buf ( n58302 , n8586 );
buf ( n58303 , n57966 );
xor ( n58304 , n58302 , n58303 );
buf ( n58305 , n57940 );
xnor ( n58306 , n58304 , n58305 );
buf ( n58307 , n58306 );
buf ( n58308 , n58307 );
not ( n58309 , n58308 );
or ( n8976 , n8967 , n58309 );
not ( n58311 , n57342 );
not ( n58312 , n57835 );
or ( n8979 , n58311 , n58312 );
nand ( n58314 , n8979 , n57839 );
buf ( n58315 , n58314 );
not ( n8982 , n58273 );
buf ( n58317 , n376 );
buf ( n58318 , n384 );
nand ( n8985 , n58317 , n58318 );
buf ( n8986 , n8985 );
buf ( n58321 , n8986 );
buf ( n58322 , n375 );
buf ( n58323 , n385 );
nand ( n58324 , n58322 , n58323 );
buf ( n58325 , n58324 );
buf ( n58326 , n58325 );
nor ( n8993 , n58321 , n58326 );
buf ( n58328 , n8993 );
buf ( n58329 , n58328 );
not ( n8996 , n58329 );
buf ( n58331 , n8996 );
not ( n8998 , n58331 );
or ( n58333 , n8982 , n8998 );
xor ( n9000 , n58242 , n58258 );
xor ( n58335 , n9000 , n58248 );
buf ( n58336 , n58328 );
buf ( n58337 , n58270 );
nand ( n9004 , n58336 , n58337 );
buf ( n9005 , n9004 );
nand ( n58340 , n58335 , n9005 );
nand ( n9007 , n58333 , n58340 );
buf ( n58342 , n9007 );
xor ( n58343 , n58315 , n58342 );
buf ( n58344 , n58273 );
buf ( n58345 , n58264 );
xor ( n58346 , n58344 , n58345 );
buf ( n58347 , n58237 );
xnor ( n9014 , n58346 , n58347 );
buf ( n58349 , n9014 );
buf ( n58350 , n58349 );
and ( n58351 , n58343 , n58350 );
and ( n58352 , n58315 , n58342 );
or ( n9019 , n58351 , n58352 );
buf ( n58354 , n9019 );
buf ( n58355 , n58354 );
xor ( n9022 , n58231 , n58283 );
xor ( n9023 , n9022 , n8959 );
buf ( n58358 , n9023 );
xor ( n9025 , n58355 , n58358 );
buf ( n58360 , n8599 );
buf ( n9027 , n55646 );
buf ( n58362 , n55621 );
nand ( n58363 , n9027 , n58362 );
buf ( n58364 , n58363 );
buf ( n58365 , n58364 );
and ( n58366 , n58360 , n58365 );
buf ( n58367 , n413 );
not ( n9034 , n58367 );
buf ( n58369 , n412 );
not ( n58370 , n58369 );
or ( n58371 , n9034 , n58370 );
buf ( n58372 , n411 );
nand ( n58373 , n58371 , n58372 );
buf ( n58374 , n58373 );
buf ( n58375 , n58374 );
nor ( n9042 , n58366 , n58375 );
buf ( n58377 , n9042 );
buf ( n58378 , n58377 );
and ( n9045 , n9025 , n58378 );
and ( n9046 , n58355 , n58358 );
or ( n9047 , n9045 , n9046 );
buf ( n58382 , n9047 );
buf ( n58383 , n58382 );
nand ( n9050 , n8976 , n58383 );
buf ( n58385 , n9050 );
buf ( n58386 , n58385 );
buf ( n58387 , n58307 );
not ( n9054 , n58387 );
buf ( n58389 , n8962 );
nand ( n58390 , n9054 , n58389 );
buf ( n58391 , n58390 );
buf ( n58392 , n58391 );
nand ( n58393 , n58386 , n58392 );
buf ( n58394 , n58393 );
buf ( n58395 , n58394 );
not ( n9062 , n58395 );
buf ( n58397 , n9062 );
not ( n9064 , n58397 );
and ( n9065 , n8879 , n9064 );
buf ( n58400 , n58212 );
buf ( n58401 , n58397 );
and ( n9068 , n58400 , n58401 );
xor ( n58403 , n58011 , n58029 );
xor ( n9070 , n58403 , n8706 );
buf ( n58405 , n9070 );
not ( n9072 , n58405 );
buf ( n58407 , n9072 );
buf ( n58408 , n58407 );
nor ( n9075 , n9068 , n58408 );
buf ( n58410 , n9075 );
nor ( n9077 , n9065 , n58410 );
buf ( n58412 , n9077 );
xor ( n9079 , n58185 , n58412 );
xor ( n9080 , n57705 , n57741 );
xor ( n9081 , n9080 , n57758 );
buf ( n58416 , n9081 );
buf ( n58417 , n58416 );
and ( n9084 , n9079 , n58417 );
and ( n58419 , n58185 , n58412 );
or ( n9086 , n9084 , n58419 );
buf ( n58421 , n9086 );
nand ( n9088 , n8844 , n58421 );
nand ( n58423 , n8820 , n9088 );
buf ( n58424 , n58423 );
not ( n9091 , n416 );
buf ( n58426 , n415 );
not ( n58427 , n58426 );
buf ( n58428 , n8334 );
not ( n58429 , n58428 );
or ( n58430 , n58427 , n58429 );
buf ( n58431 , n415 );
not ( n9098 , n58431 );
buf ( n58433 , n56238 );
nand ( n9100 , n9098 , n58433 );
buf ( n58435 , n9100 );
buf ( n58436 , n58435 );
nand ( n9103 , n58430 , n58436 );
buf ( n58438 , n9103 );
not ( n9105 , n58438 );
or ( n9106 , n9091 , n9105 );
buf ( n58441 , n6384 );
buf ( n58442 , n415 );
buf ( n58443 , n7168 );
and ( n9110 , n58442 , n58443 );
not ( n58445 , n58442 );
buf ( n9112 , n57679 );
and ( n58447 , n58445 , n9112 );
nor ( n9114 , n9110 , n58447 );
buf ( n9115 , n9114 );
buf ( n58450 , n9115 );
nand ( n9117 , n58441 , n58450 );
buf ( n58452 , n9117 );
nand ( n9119 , n9106 , n58452 );
not ( n58454 , n9119 );
xor ( n58455 , n58315 , n58342 );
xor ( n9122 , n58455 , n58350 );
buf ( n58457 , n9122 );
buf ( n58458 , n58457 );
not ( n9125 , n58458 );
buf ( n58460 , n58004 );
buf ( n58461 , n6980 );
nand ( n58462 , n58460 , n58461 );
buf ( n58463 , n58462 );
buf ( n58464 , n58463 );
nand ( n58465 , n9125 , n58464 );
buf ( n58466 , n58465 );
buf ( n58467 , n58466 );
not ( n58468 , n58467 );
buf ( n58469 , n58335 );
not ( n9136 , n58469 );
buf ( n58471 , n58328 );
not ( n58472 , n58471 );
buf ( n58473 , n58273 );
not ( n58474 , n58473 );
and ( n58475 , n58472 , n58474 );
buf ( n58476 , n58328 );
buf ( n58477 , n58273 );
and ( n9144 , n58476 , n58477 );
nor ( n9145 , n58475 , n9144 );
buf ( n58480 , n9145 );
buf ( n58481 , n58480 );
not ( n58482 , n58481 );
or ( n58483 , n9136 , n58482 );
buf ( n58484 , n58480 );
buf ( n58485 , n58335 );
or ( n58486 , n58484 , n58485 );
nand ( n58487 , n58483 , n58486 );
buf ( n58488 , n58487 );
buf ( n58489 , n376 );
buf ( n58490 , n385 );
nand ( n9157 , n58489 , n58490 );
buf ( n58492 , n9157 );
buf ( n58493 , n58492 );
not ( n58494 , n58493 );
buf ( n58495 , n377 );
buf ( n58496 , n383 );
nand ( n58497 , n58495 , n58496 );
buf ( n58498 , n58497 );
buf ( n58499 , n58498 );
not ( n58500 , n58499 );
or ( n9167 , n58494 , n58500 );
or ( n58502 , n58492 , n58498 );
not ( n9169 , n8986 );
not ( n9170 , n58325 );
or ( n9171 , n9169 , n9170 );
nand ( n9172 , n9171 , n58331 );
nand ( n9173 , n58502 , n9172 );
buf ( n58508 , n9173 );
nand ( n9175 , n9167 , n58508 );
buf ( n58510 , n9175 );
xor ( n9177 , n58488 , n58510 );
buf ( n58512 , n415 );
buf ( n58513 , n414 );
or ( n58514 , n58512 , n58513 );
buf ( n58515 , n58514 );
buf ( n58516 , n58515 );
not ( n58517 , n58516 );
buf ( n58518 , n8599 );
not ( n9185 , n58518 );
or ( n9186 , n58517 , n9185 );
buf ( n58521 , n414 );
buf ( n58522 , n415 );
and ( n9189 , n58521 , n58522 );
buf ( n58524 , n55646 );
nor ( n9191 , n9189 , n58524 );
buf ( n58526 , n9191 );
buf ( n58527 , n58526 );
nand ( n58528 , n9186 , n58527 );
buf ( n58529 , n58528 );
not ( n58530 , n58529 );
and ( n9197 , n9177 , n58530 );
and ( n58532 , n58488 , n58510 );
or ( n58533 , n9197 , n58532 );
buf ( n58534 , n58533 );
not ( n9201 , n58534 );
or ( n58536 , n58468 , n9201 );
buf ( n58537 , n58463 );
not ( n9204 , n58537 );
buf ( n58539 , n58457 );
nand ( n58540 , n9204 , n58539 );
buf ( n58541 , n58540 );
buf ( n58542 , n58541 );
nand ( n58543 , n58536 , n58542 );
buf ( n58544 , n58543 );
not ( n58545 , n58544 );
or ( n9212 , n58454 , n58545 );
nor ( n9213 , n9119 , n58544 );
xor ( n9214 , n58355 , n58358 );
xor ( n58549 , n9214 , n58378 );
buf ( n58550 , n58549 );
buf ( n58551 , n6980 );
not ( n9218 , n58551 );
buf ( n58553 , n411 );
buf ( n58554 , n57554 );
xor ( n9221 , n58553 , n58554 );
buf ( n58556 , n9221 );
buf ( n58557 , n58556 );
not ( n58558 , n58557 );
or ( n9225 , n9218 , n58558 );
and ( n58560 , n411 , n58001 );
not ( n58561 , n411 );
and ( n9228 , n58561 , n57936 );
or ( n58563 , n58560 , n9228 );
buf ( n9230 , n58563 );
buf ( n58565 , n56072 );
nand ( n58566 , n9230 , n58565 );
buf ( n58567 , n58566 );
buf ( n58568 , n58567 );
nand ( n9235 , n9225 , n58568 );
buf ( n58570 , n9235 );
xor ( n58571 , n58550 , n58570 );
not ( n9238 , n58571 );
not ( n9239 , n9238 );
buf ( n58574 , n55998 );
not ( n9241 , n58574 );
not ( n9242 , n413 );
not ( n9243 , n57787 );
or ( n58578 , n9242 , n9243 );
or ( n9245 , n413 , n57787 );
nand ( n58580 , n58578 , n9245 );
buf ( n58581 , n58580 );
not ( n9248 , n58581 );
or ( n58583 , n9241 , n9248 );
and ( n9250 , n8194 , n55646 );
not ( n9251 , n8194 );
and ( n58586 , n9251 , n413 );
or ( n9253 , n9250 , n58586 );
buf ( n58588 , n9253 );
buf ( n58589 , n6591 );
nand ( n9256 , n58588 , n58589 );
buf ( n9257 , n9256 );
buf ( n58592 , n9257 );
nand ( n58593 , n58583 , n58592 );
buf ( n58594 , n58593 );
not ( n58595 , n58594 );
or ( n9262 , n9239 , n58595 );
not ( n58597 , n58594 );
nand ( n58598 , n58597 , n58571 );
nand ( n9265 , n9262 , n58598 );
not ( n58600 , n9265 );
or ( n58601 , n9213 , n58600 );
nand ( n9268 , n9212 , n58601 );
not ( n58603 , n9268 );
buf ( n58604 , n6384 );
not ( n9271 , n58604 );
buf ( n58606 , n58438 );
not ( n9273 , n58606 );
or ( n9274 , n9271 , n9273 );
xor ( n58609 , n415 , n56195 );
xnor ( n9276 , n58609 , n6860 );
buf ( n58611 , n9276 );
buf ( n58612 , n416 );
nand ( n58613 , n58611 , n58612 );
buf ( n58614 , n58613 );
buf ( n58615 , n58614 );
nand ( n9282 , n9274 , n58615 );
buf ( n58617 , n9282 );
not ( n58618 , n58594 );
not ( n9285 , n58570 );
buf ( n58620 , n58550 );
not ( n9287 , n58620 );
nand ( n9288 , n9285 , n9287 );
not ( n58623 , n9288 );
or ( n9290 , n58618 , n58623 );
nand ( n58625 , n58570 , n58620 );
nand ( n9292 , n9290 , n58625 );
not ( n58627 , n9292 );
and ( n9294 , n58617 , n58627 );
not ( n9295 , n58617 );
and ( n9296 , n9295 , n9292 );
nor ( n9297 , n9294 , n9296 );
not ( n58632 , n6980 );
not ( n58633 , n58025 );
or ( n9300 , n58632 , n58633 );
buf ( n58635 , n58556 );
buf ( n58636 , n56072 );
nand ( n9303 , n58635 , n58636 );
buf ( n9304 , n9303 );
nand ( n9305 , n9300 , n9304 );
not ( n58640 , n9305 );
not ( n9307 , n58640 );
xor ( n58642 , n8962 , n58382 );
xnor ( n9309 , n58642 , n58307 );
not ( n9310 , n9309 );
not ( n9311 , n9310 );
or ( n58646 , n9307 , n9311 );
nand ( n9313 , n9305 , n9309 );
nand ( n58648 , n58646 , n9313 );
buf ( n58649 , n58202 );
buf ( n58650 , n6665 );
and ( n58651 , n58649 , n58650 );
not ( n9318 , n58580 );
nor ( n58653 , n9318 , n55671 );
buf ( n58654 , n58653 );
nor ( n9321 , n58651 , n58654 );
buf ( n58656 , n9321 );
and ( n58657 , n58648 , n58656 );
not ( n9324 , n58648 );
buf ( n58659 , n58656 );
not ( n58660 , n58659 );
buf ( n58661 , n58660 );
and ( n58662 , n9324 , n58661 );
nor ( n58663 , n58657 , n58662 );
and ( n9330 , n9297 , n58663 );
not ( n58665 , n9297 );
not ( n58666 , n58663 );
and ( n9333 , n58665 , n58666 );
nor ( n9334 , n9330 , n9333 );
nand ( n58669 , n58603 , n9334 );
not ( n58670 , n58669 );
buf ( n58671 , n416 );
not ( n9338 , n58671 );
buf ( n58673 , n9115 );
not ( n58674 , n58673 );
or ( n9341 , n9338 , n58674 );
not ( n58676 , n415 );
not ( n9343 , n57787 );
or ( n9344 , n58676 , n9343 );
or ( n58679 , n57790 , n415 );
nand ( n58680 , n9344 , n58679 );
buf ( n58681 , n58680 );
buf ( n58682 , n6384 );
nand ( n9349 , n58681 , n58682 );
buf ( n58684 , n9349 );
buf ( n58685 , n58684 );
nand ( n58686 , n9341 , n58685 );
buf ( n58687 , n58686 );
not ( n58688 , n55998 );
not ( n9355 , n9253 );
or ( n58690 , n58688 , n9355 );
buf ( n58691 , n413 );
not ( n9358 , n58691 );
buf ( n58693 , n57555 );
not ( n58694 , n58693 );
or ( n58695 , n9358 , n58694 );
buf ( n58696 , n57554 );
buf ( n58697 , n6322 );
nand ( n9364 , n58696 , n58697 );
buf ( n58699 , n9364 );
buf ( n58700 , n58699 );
nand ( n9367 , n58695 , n58700 );
buf ( n58702 , n9367 );
buf ( n58703 , n58702 );
buf ( n9370 , n6591 );
nand ( n9371 , n58703 , n9370 );
buf ( n9372 , n9371 );
nand ( n9373 , n58690 , n9372 );
nor ( n9374 , n58687 , n9373 );
buf ( n58709 , n9374 );
buf ( n58710 , n58533 );
not ( n9377 , n58710 );
and ( n58712 , n58457 , n58463 );
not ( n9379 , n58457 );
and ( n58714 , n57936 , n6980 );
and ( n9381 , n9379 , n58714 );
nor ( n9382 , n58712 , n9381 );
buf ( n58717 , n9382 );
not ( n9384 , n58717 );
and ( n9385 , n9377 , n9384 );
buf ( n58720 , n58533 );
buf ( n58721 , n9382 );
and ( n9388 , n58720 , n58721 );
nor ( n58723 , n9385 , n9388 );
buf ( n58724 , n58723 );
buf ( n58725 , n58724 );
or ( n58726 , n58709 , n58725 );
not ( n58727 , n58687 );
buf ( n58728 , n58727 );
not ( n58729 , n58728 );
buf ( n58730 , n9373 );
nand ( n9397 , n58729 , n58730 );
buf ( n58732 , n9397 );
buf ( n58733 , n58732 );
nand ( n58734 , n58726 , n58733 );
buf ( n58735 , n58734 );
not ( n9402 , n58735 );
not ( n58737 , n9402 );
xor ( n9404 , n58544 , n9265 );
xnor ( n58739 , n9404 , n9119 );
not ( n9406 , n58739 );
or ( n9407 , n58737 , n9406 );
buf ( n58742 , n416 );
not ( n9409 , n58742 );
buf ( n58744 , n58680 );
not ( n9411 , n58744 );
or ( n9412 , n9409 , n9411 );
and ( n9413 , n415 , n8195 );
not ( n9414 , n415 );
and ( n9415 , n9414 , n8275 );
nor ( n58750 , n9413 , n9415 );
buf ( n58751 , n58750 );
buf ( n58752 , n6384 );
nand ( n58753 , n58751 , n58752 );
buf ( n58754 , n58753 );
buf ( n58755 , n58754 );
nand ( n9422 , n9412 , n58755 );
buf ( n58757 , n9422 );
not ( n9424 , n58757 );
and ( n58759 , n58004 , n55646 );
not ( n58760 , n58004 );
and ( n9427 , n58760 , n413 );
nor ( n58762 , n58759 , n9427 );
not ( n9429 , n58762 );
not ( n9430 , n55671 );
and ( n58765 , n9429 , n9430 );
and ( n9432 , n58702 , n55998 );
nor ( n58767 , n58765 , n9432 );
buf ( n58768 , n58767 );
not ( n9435 , n58768 );
buf ( n58770 , n9435 );
not ( n9437 , n58770 );
or ( n58772 , n9424 , n9437 );
buf ( n58773 , n58757 );
buf ( n58774 , n58770 );
nor ( n58775 , n58773 , n58774 );
buf ( n58776 , n58775 );
xor ( n9443 , n58488 , n58510 );
not ( n58778 , n58529 );
xor ( n9445 , n9443 , n58778 );
buf ( n58780 , n9445 );
not ( n9447 , n58780 );
buf ( n58782 , n9447 );
or ( n58783 , n58776 , n58782 );
nand ( n9450 , n58772 , n58783 );
buf ( n58785 , n9450 );
not ( n9452 , n58785 );
buf ( n58787 , n9373 );
not ( n9454 , n58787 );
buf ( n58789 , n58724 );
not ( n9456 , n58789 );
or ( n9457 , n9454 , n9456 );
buf ( n58792 , n58724 );
buf ( n58793 , n9373 );
or ( n9460 , n58792 , n58793 );
nand ( n9461 , n9457 , n9460 );
buf ( n58796 , n9461 );
buf ( n58797 , n58796 );
not ( n9464 , n58797 );
buf ( n58799 , n58727 );
not ( n9466 , n58799 );
and ( n9467 , n9464 , n9466 );
buf ( n58802 , n58727 );
buf ( n58803 , n58796 );
and ( n58804 , n58802 , n58803 );
nor ( n9471 , n9467 , n58804 );
buf ( n9472 , n9471 );
buf ( n58807 , n9472 );
nand ( n9474 , n9452 , n58807 );
buf ( n58809 , n9474 );
not ( n9476 , n58809 );
buf ( n58811 , n58767 );
not ( n9478 , n58811 );
buf ( n58813 , n9445 );
not ( n9480 , n58813 );
and ( n58815 , n9478 , n9480 );
buf ( n58816 , n58767 );
buf ( n58817 , n9445 );
and ( n58818 , n58816 , n58817 );
nor ( n9485 , n58815 , n58818 );
buf ( n58820 , n9485 );
buf ( n58821 , n58820 );
not ( n58822 , n58821 );
buf ( n58823 , n58757 );
not ( n9490 , n58823 );
and ( n58825 , n58822 , n9490 );
buf ( n58826 , n58757 );
buf ( n58827 , n58820 );
and ( n9494 , n58826 , n58827 );
nor ( n9495 , n58825 , n9494 );
buf ( n58830 , n9495 );
buf ( n58831 , n58830 );
buf ( n58832 , n58498 );
buf ( n58833 , n58492 );
and ( n9500 , n58832 , n58833 );
not ( n58835 , n58832 );
buf ( n58836 , n58492 );
not ( n58837 , n58836 );
buf ( n58838 , n58837 );
buf ( n58839 , n58838 );
and ( n58840 , n58835 , n58839 );
nor ( n58841 , n9500 , n58840 );
buf ( n58842 , n58841 );
xnor ( n9509 , n9172 , n58842 );
buf ( n58844 , n9509 );
buf ( n58845 , n58004 );
buf ( n58846 , n55998 );
nand ( n58847 , n58845 , n58846 );
buf ( n58848 , n58847 );
buf ( n58849 , n58848 );
xor ( n58850 , n58844 , n58849 );
nand ( n58851 , n416 , n57936 );
buf ( n58852 , n377 );
buf ( n58853 , n384 );
nand ( n58854 , n58852 , n58853 );
buf ( n58855 , n58854 );
buf ( n58856 , n58855 );
not ( n58857 , n58856 );
buf ( n58858 , n58492 );
nand ( n58859 , n58857 , n58858 );
buf ( n58860 , n58859 );
and ( n9527 , n58851 , n58860 , n415 );
and ( n9528 , n58838 , n58855 );
nor ( n58863 , n9527 , n9528 );
buf ( n58864 , n58863 );
and ( n9531 , n58850 , n58864 );
and ( n58866 , n58844 , n58849 );
or ( n58867 , n9531 , n58866 );
buf ( n58868 , n58867 );
buf ( n58869 , n58868 );
nand ( n9536 , n58831 , n58869 );
buf ( n58871 , n9536 );
not ( n9538 , n58871 );
buf ( n58873 , n416 );
not ( n9540 , n58873 );
and ( n9541 , n415 , n57555 );
not ( n9542 , n415 );
and ( n9543 , n9542 , n57554 );
or ( n9544 , n9541 , n9543 );
buf ( n58879 , n9544 );
not ( n9546 , n58879 );
or ( n9547 , n9540 , n9546 );
buf ( n58882 , n58004 );
not ( n58883 , n58882 );
buf ( n58884 , n6384 );
nand ( n9550 , n58883 , n58884 );
buf ( n58886 , n9550 );
buf ( n58887 , n58886 );
nand ( n9553 , n9547 , n58887 );
buf ( n58889 , n9553 );
buf ( n58890 , n58889 );
xnor ( n58891 , n58855 , n58492 );
not ( n58892 , n58891 );
nand ( n58893 , n58851 , n415 );
not ( n9559 , n58893 );
or ( n58895 , n58892 , n9559 );
or ( n9561 , n58893 , n58891 );
nand ( n58897 , n58895 , n9561 );
buf ( n9563 , n58897 );
nor ( n9564 , n58890 , n9563 );
buf ( n9565 , n9564 );
buf ( n58901 , n9565 );
nand ( n58902 , n416 , n57936 );
buf ( n9566 , n58902 );
buf ( n58904 , n377 );
buf ( n58905 , n385 );
and ( n9569 , n58904 , n58905 );
buf ( n58907 , n9569 );
buf ( n9571 , n58907 );
and ( n9572 , n9566 , n9571 );
buf ( n58910 , n9572 );
buf ( n58911 , n58910 );
or ( n9575 , n58901 , n58911 );
buf ( n9576 , n58889 );
buf ( n9577 , n58897 );
nand ( n9578 , n9576 , n9577 );
buf ( n9579 , n9578 );
buf ( n58917 , n9579 );
nand ( n58918 , n9575 , n58917 );
buf ( n58919 , n58918 );
not ( n58920 , n58919 );
buf ( n58921 , n416 );
not ( n58922 , n58921 );
buf ( n58923 , n58750 );
not ( n58924 , n58923 );
or ( n58925 , n58922 , n58924 );
buf ( n58926 , n9544 );
buf ( n58927 , n6384 );
nand ( n9587 , n58926 , n58927 );
buf ( n58929 , n9587 );
buf ( n58930 , n58929 );
nand ( n9590 , n58925 , n58930 );
buf ( n58932 , n9590 );
not ( n9592 , n58932 );
or ( n58934 , n58920 , n9592 );
buf ( n58935 , n58919 );
buf ( n58936 , n58932 );
nor ( n9596 , n58935 , n58936 );
buf ( n58938 , n9596 );
xor ( n9598 , n58844 , n58849 );
xor ( n58940 , n9598 , n58864 );
buf ( n58941 , n58940 );
or ( n9601 , n58938 , n58941 );
nand ( n58943 , n58934 , n9601 );
not ( n58944 , n58943 );
or ( n58945 , n9538 , n58944 );
not ( n58946 , n58830 );
not ( n9605 , n58868 );
nand ( n58948 , n58946 , n9605 );
nand ( n9607 , n58945 , n58948 );
not ( n9608 , n9607 );
or ( n9609 , n9476 , n9608 );
buf ( n58952 , n9472 );
not ( n9611 , n58952 );
buf ( n9612 , n9450 );
buf ( n58955 , n9612 );
nand ( n58956 , n9611 , n58955 );
buf ( n58957 , n58956 );
nand ( n58958 , n9609 , n58957 );
nand ( n58959 , n9407 , n58958 );
buf ( n58960 , n58739 );
not ( n58961 , n58960 );
buf ( n58962 , n58735 );
nand ( n58963 , n58961 , n58962 );
buf ( n58964 , n58963 );
nand ( n58965 , n58959 , n58964 );
not ( n9619 , n58965 );
or ( n58967 , n58670 , n9619 );
not ( n58968 , n9334 );
nand ( n58969 , n58968 , n9268 );
nand ( n58970 , n58967 , n58969 );
not ( n58971 , n58970 );
not ( n58972 , n58663 );
or ( n58973 , n58617 , n9292 );
not ( n58974 , n58973 );
or ( n58975 , n58972 , n58974 );
buf ( n58976 , n58617 );
buf ( n58977 , n9292 );
nand ( n9624 , n58976 , n58977 );
buf ( n58979 , n9624 );
nand ( n9626 , n58975 , n58979 );
buf ( n58981 , n9626 );
not ( n58982 , n58981 );
buf ( n58983 , n58394 );
buf ( n58984 , n9070 );
xor ( n9631 , n58983 , n58984 );
buf ( n58986 , n58212 );
xnor ( n58987 , n9631 , n58986 );
buf ( n58988 , n58987 );
buf ( n58989 , n58988 );
not ( n9634 , n58989 );
buf ( n58991 , n58202 );
buf ( n58992 , n6665 );
and ( n58993 , n58991 , n58992 );
buf ( n58994 , n58653 );
nor ( n58995 , n58993 , n58994 );
buf ( n58996 , n58995 );
not ( n58997 , n58996 );
not ( n58998 , n58640 );
and ( n58999 , n58997 , n58998 );
buf ( n59000 , n9309 );
nand ( n9637 , n58996 , n58640 );
and ( n59002 , n59000 , n9637 );
nor ( n59003 , n58999 , n59002 );
buf ( n59004 , n59003 );
not ( n9641 , n59004 );
buf ( n59006 , n6384 );
not ( n59007 , n59006 );
buf ( n59008 , n9276 );
not ( n59009 , n59008 );
or ( n9646 , n59007 , n59009 );
not ( n59011 , n57747 );
nand ( n9648 , n59011 , n416 );
buf ( n59013 , n9648 );
nand ( n59014 , n9646 , n59013 );
buf ( n59015 , n59014 );
buf ( n59016 , n59015 );
not ( n9653 , n59016 );
and ( n59018 , n9641 , n9653 );
buf ( n9655 , n59003 );
buf ( n59020 , n59015 );
and ( n59021 , n9655 , n59020 );
nor ( n9658 , n59018 , n59021 );
buf ( n59023 , n9658 );
buf ( n59024 , n59023 );
not ( n59025 , n59024 );
and ( n9661 , n9634 , n59025 );
buf ( n59027 , n58988 );
buf ( n59028 , n59023 );
and ( n9664 , n59027 , n59028 );
nor ( n59030 , n9661 , n9664 );
buf ( n59031 , n59030 );
buf ( n59032 , n59031 );
nand ( n9668 , n58982 , n59032 );
buf ( n9669 , n9668 );
not ( n59035 , n9669 );
or ( n59036 , n58971 , n59035 );
buf ( n59037 , n59031 );
not ( n59038 , n59037 );
buf ( n59039 , n9626 );
nand ( n9675 , n59038 , n59039 );
buf ( n59041 , n9675 );
nand ( n9677 , n59036 , n59041 );
buf ( n59043 , n59015 );
not ( n59044 , n59043 );
buf ( n59045 , n59003 );
nand ( n9681 , n59044 , n59045 );
buf ( n9682 , n9681 );
buf ( n59048 , n9682 );
not ( n59049 , n59048 );
buf ( n59050 , n58988 );
not ( n59051 , n59050 );
or ( n59052 , n59049 , n59051 );
buf ( n59053 , n59003 );
not ( n59054 , n59053 );
buf ( n9690 , n59015 );
nand ( n9691 , n59054 , n9690 );
buf ( n9692 , n9691 );
buf ( n59058 , n9692 );
nand ( n9694 , n59052 , n59058 );
buf ( n59060 , n9694 );
buf ( n59061 , n59060 );
not ( n59062 , n59061 );
xor ( n9698 , n58185 , n58412 );
xor ( n59064 , n9698 , n58417 );
buf ( n59065 , n59064 );
buf ( n59066 , n59065 );
nand ( n59067 , n59062 , n59066 );
buf ( n59068 , n59067 );
and ( n59069 , n9677 , n59068 );
buf ( n59070 , n59060 );
not ( n9706 , n59070 );
buf ( n59072 , n59065 );
nor ( n9708 , n9706 , n59072 );
buf ( n59074 , n9708 );
nor ( n9710 , n59069 , n59074 );
buf ( n59076 , n9710 );
or ( n9712 , n58424 , n59076 );
buf ( n59078 , n8818 );
buf ( n59079 , n58073 );
nand ( n9715 , n59078 , n59079 );
buf ( n59081 , n9715 );
buf ( n59082 , n59081 );
buf ( n59083 , n8844 );
buf ( n59084 , n58421 );
nor ( n59085 , n59083 , n59084 );
buf ( n59086 , n59085 );
buf ( n59087 , n59086 );
and ( n9721 , n59082 , n59087 );
buf ( n59089 , n58073 );
buf ( n59090 , n8818 );
nor ( n59091 , n59089 , n59090 );
buf ( n59092 , n59091 );
buf ( n59093 , n59092 );
nor ( n9727 , n9721 , n59093 );
buf ( n59095 , n9727 );
buf ( n59096 , n59095 );
nand ( n9730 , n9712 , n59096 );
buf ( n9731 , n9730 );
not ( n9732 , n9731 );
buf ( n59100 , n56471 );
buf ( n59101 , n56478 );
xor ( n9735 , n59100 , n59101 );
buf ( n59103 , n56748 );
xnor ( n9737 , n9735 , n59103 );
buf ( n9738 , n9737 );
buf ( n59106 , n9738 );
not ( n9740 , n59106 );
buf ( n59108 , n56333 );
buf ( n59109 , n7018 );
buf ( n9743 , n59109 );
buf ( n59111 , n9743 );
buf ( n59112 , n59111 );
xor ( n59113 , n59108 , n59112 );
buf ( n59114 , n56386 );
xnor ( n59115 , n59113 , n59114 );
buf ( n59116 , n59115 );
buf ( n59117 , n59116 );
buf ( n59118 , n7393 );
buf ( n59119 , n56560 );
and ( n59120 , n59118 , n59119 );
not ( n9754 , n59118 );
buf ( n59122 , n56561 );
and ( n59123 , n9754 , n59122 );
nor ( n9757 , n59120 , n59123 );
buf ( n9758 , n9757 );
not ( n59126 , n9758 );
not ( n9760 , n7399 );
not ( n59128 , n9760 );
or ( n59129 , n59126 , n59128 );
not ( n9763 , n9758 );
nand ( n59131 , n9763 , n7399 );
nand ( n59132 , n59129 , n59131 );
not ( n59133 , n58126 );
not ( n9766 , n58117 );
nand ( n9767 , n9766 , n8786 );
not ( n9768 , n9767 );
or ( n59137 , n59133 , n9768 );
nand ( n9770 , n58117 , n8785 );
nand ( n9771 , n59137 , n9770 );
nor ( n9772 , n59132 , n9771 );
not ( n9773 , n9772 );
not ( n9774 , n9773 );
buf ( n59143 , n58090 );
buf ( n59144 , n8768 );
or ( n59145 , n59143 , n59144 );
buf ( n59146 , n58080 );
nand ( n9779 , n59145 , n59146 );
buf ( n9780 , n9779 );
buf ( n59149 , n8768 );
buf ( n59150 , n58090 );
nand ( n59151 , n59149 , n59150 );
buf ( n59152 , n59151 );
nand ( n9785 , n9780 , n59152 );
not ( n9786 , n9785 );
or ( n59155 , n9774 , n9786 );
nand ( n59156 , n59132 , n9771 );
nand ( n9789 , n59155 , n59156 );
buf ( n59158 , n9789 );
not ( n59159 , n59158 );
buf ( n59160 , n59159 );
buf ( n59161 , n59160 );
xor ( n59162 , n59117 , n59161 );
buf ( n59163 , n56555 );
not ( n9796 , n59163 );
not ( n59165 , n7410 );
not ( n59166 , n56738 );
or ( n59167 , n59165 , n59166 );
or ( n9800 , n56738 , n7410 );
nand ( n59169 , n59167 , n9800 );
buf ( n59170 , n59169 );
not ( n9803 , n59170 );
and ( n59172 , n9796 , n9803 );
buf ( n59173 , n56555 );
buf ( n59174 , n59169 );
and ( n59175 , n59173 , n59174 );
nor ( n9808 , n59172 , n59175 );
buf ( n9809 , n9808 );
buf ( n59178 , n9809 );
and ( n9811 , n59162 , n59178 );
and ( n59180 , n59117 , n59161 );
or ( n59181 , n9811 , n59180 );
buf ( n59182 , n59181 );
buf ( n59183 , n59182 );
not ( n59184 , n59183 );
or ( n59185 , n9740 , n59184 );
xor ( n9816 , n59117 , n59161 );
xor ( n9817 , n9816 , n59178 );
buf ( n59188 , n9817 );
buf ( n59189 , n56508 );
not ( n59190 , n59189 );
buf ( n59191 , n59190 );
xor ( n9822 , n56546 , n59191 );
buf ( n59193 , n7192 );
buf ( n59194 , n59193 );
buf ( n59195 , n59194 );
not ( n59196 , n59195 );
and ( n9827 , n9822 , n59196 );
not ( n59198 , n9822 );
and ( n59199 , n59198 , n59195 );
nor ( n9830 , n9827 , n59199 );
not ( n9831 , n9830 );
not ( n59202 , n9772 );
nand ( n9833 , n59202 , n59156 );
not ( n9834 , n9833 );
not ( n59205 , n9785 );
not ( n9836 , n59205 );
or ( n59207 , n9834 , n9836 );
or ( n9838 , n59205 , n9833 );
nand ( n59209 , n59207 , n9838 );
nand ( n59210 , n9831 , n59209 );
not ( n9841 , n8793 );
buf ( n59212 , n58140 );
not ( n59213 , n59212 );
buf ( n59214 , n59213 );
nand ( n59215 , n9841 , n59214 );
not ( n59216 , n59215 );
not ( n9847 , n8812 );
or ( n59218 , n59216 , n9847 );
buf ( n59219 , n59214 );
not ( n9850 , n59219 );
buf ( n59221 , n8793 );
nand ( n59222 , n9850 , n59221 );
buf ( n59223 , n59222 );
nand ( n9854 , n59218 , n59223 );
and ( n59225 , n59210 , n9854 );
not ( n9856 , n9830 );
nor ( n9857 , n9856 , n59209 );
nor ( n59228 , n59225 , n9857 );
nand ( n9859 , n59188 , n59228 );
buf ( n59230 , n9859 );
nand ( n59231 , n59185 , n59230 );
buf ( n59232 , n59231 );
buf ( n59233 , n58105 );
not ( n9864 , n59233 );
buf ( n59235 , n58149 );
not ( n9866 , n59235 );
or ( n9867 , n9864 , n9866 );
buf ( n59238 , n8776 );
nand ( n59239 , n9867 , n59238 );
buf ( n59240 , n59239 );
buf ( n59241 , n59240 );
buf ( n59242 , n58149 );
buf ( n59243 , n58105 );
or ( n59244 , n59242 , n59243 );
buf ( n59245 , n59244 );
buf ( n59246 , n59245 );
nand ( n9877 , n59241 , n59246 );
buf ( n59248 , n9877 );
buf ( n59249 , n59248 );
xor ( n59250 , n9830 , n9854 );
not ( n59251 , n59209 );
xor ( n9882 , n59250 , n59251 );
buf ( n59253 , n9882 );
nor ( n59254 , n59249 , n59253 );
buf ( n59255 , n59254 );
nor ( n59256 , n59232 , n59255 );
not ( n59257 , n59256 );
or ( n9888 , n9732 , n59257 );
buf ( n59259 , n59232 );
not ( n9890 , n59259 );
buf ( n59261 , n9890 );
buf ( n59262 , n9882 );
buf ( n59263 , n59248 );
and ( n59264 , n59262 , n59263 );
buf ( n59265 , n59264 );
and ( n59266 , n59261 , n59265 );
buf ( n9897 , n9738 );
buf ( n59268 , n59182 );
nand ( n59269 , n9897 , n59268 );
buf ( n59270 , n59269 );
buf ( n59271 , n59270 );
not ( n59272 , n59271 );
buf ( n59273 , n59272 );
buf ( n59274 , n59273 );
buf ( n59275 , n59188 );
not ( n9906 , n59275 );
buf ( n59277 , n9906 );
not ( n9908 , n59228 );
nand ( n9909 , n59277 , n9908 );
buf ( n59280 , n9909 );
or ( n59281 , n59274 , n59280 );
buf ( n59282 , n9738 );
buf ( n59283 , n59182 );
or ( n59284 , n59282 , n59283 );
buf ( n59285 , n59284 );
buf ( n59286 , n59285 );
nand ( n59287 , n59281 , n59286 );
buf ( n59288 , n59287 );
nor ( n9919 , n59266 , n59288 );
nand ( n59290 , n9888 , n9919 );
buf ( n9921 , n59290 );
nand ( n9922 , n57302 , n9921 );
buf ( n9923 , n9922 );
buf ( n59294 , n9923 );
buf ( n59295 , n57272 );
not ( n9926 , n59295 );
buf ( n59297 , n57172 );
not ( n9928 , n59297 );
buf ( n59299 , n57184 );
buf ( n59300 , n57114 );
buf ( n59301 , n57096 );
nand ( n9932 , n59300 , n59301 );
buf ( n59303 , n9932 );
buf ( n59304 , n59303 );
or ( n9935 , n59299 , n59304 );
nand ( n59306 , n57177 , n7849 );
buf ( n59307 , n59306 );
nand ( n59308 , n9935 , n59307 );
buf ( n59309 , n59308 );
buf ( n59310 , n59309 );
not ( n59311 , n59310 );
or ( n9942 , n9928 , n59311 );
or ( n59313 , n7834 , n57146 );
buf ( n59314 , n59313 );
nand ( n9945 , n9942 , n59314 );
buf ( n59316 , n9945 );
buf ( n59317 , n59316 );
nand ( n9948 , n9926 , n59317 );
buf ( n59319 , n9948 );
buf ( n59320 , n59319 );
buf ( n59321 , n7925 );
not ( n9952 , n59321 );
buf ( n59323 , n9952 );
buf ( n59324 , n59323 );
not ( n9955 , n59324 );
buf ( n59326 , n7928 );
buf ( n9957 , n7932 );
or ( n9958 , n59326 , n9957 );
buf ( n59329 , n9958 );
buf ( n59330 , n59329 );
not ( n9961 , n59330 );
and ( n9962 , n9955 , n9961 );
buf ( n59333 , n57212 );
buf ( n59334 , n57244 );
and ( n9965 , n59333 , n59334 );
buf ( n59336 , n55782 );
buf ( n59337 , n57255 );
and ( n9968 , n59336 , n59337 );
nor ( n59339 , n9965 , n9968 );
buf ( n59340 , n59339 );
buf ( n59341 , n59340 );
buf ( n59342 , n57258 );
or ( n9973 , n59341 , n59342 );
buf ( n59344 , n55808 );
nand ( n9975 , n9973 , n59344 );
buf ( n59346 , n9975 );
buf ( n59347 , n59346 );
nor ( n59348 , n9962 , n59347 );
buf ( n59349 , n59348 );
buf ( n59350 , n59349 );
nand ( n9981 , n57275 , n59294 , n59320 , n59350 );
buf ( n59352 , n9981 );
buf ( n59353 , n59352 );
not ( n59354 , n59353 );
buf ( n59355 , n59354 );
buf ( n59356 , n59355 );
not ( n9987 , n59356 );
or ( n9988 , n6491 , n9987 );
buf ( n59359 , n59352 );
buf ( n59360 , n55811 );
nand ( n59361 , n59359 , n59360 );
buf ( n59362 , n59361 );
buf ( n59363 , n59362 );
nand ( n9994 , n9988 , n59363 );
buf ( n59365 , n9994 );
buf ( n59366 , n59365 );
not ( n59367 , n59366 );
not ( n59368 , n382 );
buf ( n59369 , n381 );
not ( n59370 , n59369 );
buf ( n59371 , n59370 );
not ( n10002 , n59371 );
or ( n10003 , n59368 , n10002 );
not ( n59374 , n382 );
nand ( n59375 , n59374 , n381 );
nand ( n10005 , n10003 , n59375 );
not ( n59377 , n10005 );
buf ( n59378 , n59377 );
not ( n59379 , n59378 );
not ( n59380 , n380 );
and ( n10010 , n59380 , n59371 );
and ( n59382 , n380 , n381 );
nor ( n59383 , n10010 , n59382 , n10005 );
not ( n59384 , n59383 );
buf ( n59385 , n59384 );
not ( n10015 , n59385 );
or ( n10016 , n59379 , n10015 );
buf ( n59388 , n380 );
nand ( n10018 , n10016 , n59388 );
buf ( n59390 , n10018 );
buf ( n59391 , n59390 );
buf ( n59392 , n59391 );
not ( n59393 , n59392 );
buf ( n59394 , n59393 );
buf ( n59395 , n59394 );
nor ( n10025 , n59367 , n59395 );
buf ( n59397 , n10025 );
not ( n59398 , n59397 );
buf ( n59399 , n379 );
not ( n10029 , n59399 );
buf ( n59401 , n10029 );
not ( n59402 , n59401 );
not ( n10032 , n378 );
and ( n59404 , n59402 , n10032 );
and ( n59405 , n59401 , n378 );
nor ( n59406 , n59404 , n59405 );
not ( n10036 , n380 );
not ( n59408 , n59401 );
or ( n59409 , n10036 , n59408 );
not ( n59410 , n380 );
nand ( n10040 , n59410 , n379 );
nand ( n59412 , n59409 , n10040 );
or ( n59413 , n59406 , n59412 );
not ( n10043 , n59413 );
not ( n59415 , n59412 );
not ( n59416 , n59415 );
or ( n10046 , n10043 , n59416 );
nand ( n10047 , n10046 , n378 );
not ( n59419 , n10047 );
not ( n59420 , n59365 );
buf ( n59421 , n59420 );
buf ( n59422 , n59394 );
nand ( n59423 , n59421 , n59422 );
buf ( n59424 , n59423 );
nand ( n10054 , n59419 , n59424 );
nand ( n10055 , n59398 , n10054 );
buf ( n59427 , n10055 );
not ( n59428 , n59427 );
buf ( n59429 , n10047 );
not ( n59430 , n59429 );
buf ( n59431 , n59430 );
xor ( n59432 , n59431 , n59394 );
not ( n10062 , n59432 );
nor ( n59434 , n10062 , n59394 );
and ( n10064 , n59431 , n59394 );
or ( n59436 , n59434 , n10064 );
buf ( n10066 , n59436 );
nand ( n10067 , n59428 , n10066 );
buf ( n59439 , n10067 );
buf ( n59440 , n59439 );
not ( n59441 , n59440 );
buf ( n59442 , n59394 );
buf ( n59443 , n59431 );
nor ( n10073 , n59442 , n59443 );
buf ( n59445 , n10073 );
buf ( n59446 , n59445 );
not ( n59447 , n59446 );
buf ( n59448 , n59447 );
not ( n59449 , n59448 );
buf ( n59450 , n10047 );
not ( n10080 , n59374 );
not ( n59452 , n383 );
or ( n59453 , n10080 , n59452 );
not ( n59454 , n383 );
nand ( n10084 , n59454 , n382 );
nand ( n59456 , n59453 , n10084 );
not ( n10086 , n383 );
buf ( n59458 , n384 );
not ( n59459 , n59458 );
buf ( n59460 , n59459 );
not ( n59461 , n59460 );
or ( n10091 , n10086 , n59461 );
nand ( n10092 , n59454 , n384 );
nand ( n10093 , n10091 , n10092 );
not ( n10094 , n10093 );
nand ( n10095 , n59456 , n10094 );
not ( n10096 , n10095 );
not ( n10097 , n10094 );
or ( n10098 , n10096 , n10097 );
nand ( n10099 , n10098 , n382 );
buf ( n59471 , n10099 );
nand ( n10101 , n59450 , n59471 );
buf ( n59473 , n10101 );
not ( n10103 , n59473 );
not ( n10104 , n59365 );
not ( n10105 , n10104 );
or ( n10106 , n10103 , n10105 );
buf ( n59478 , n10099 );
not ( n10108 , n59478 );
buf ( n59480 , n10108 );
buf ( n59481 , n59480 );
buf ( n59482 , n59431 );
nand ( n10112 , n59481 , n59482 );
buf ( n59484 , n10112 );
nand ( n10114 , n10106 , n59484 );
not ( n10115 , n10114 );
or ( n10116 , n59449 , n10115 );
buf ( n59488 , n59431 );
buf ( n59489 , n59394 );
nand ( n10119 , n59488 , n59489 );
buf ( n59491 , n10119 );
nand ( n10121 , n10116 , n59491 );
buf ( n59493 , n10121 );
not ( n10123 , n59493 );
buf ( n59495 , n59432 );
buf ( n10125 , n10104 );
buf ( n59497 , n10125 );
and ( n10127 , n59495 , n59497 );
not ( n10128 , n59495 );
not ( n10129 , n10125 );
buf ( n59501 , n10129 );
and ( n10131 , n10128 , n59501 );
or ( n10132 , n10127 , n10131 );
buf ( n59504 , n10132 );
buf ( n59505 , n59504 );
nand ( n10135 , n10123 , n59505 );
buf ( n59507 , n10135 );
buf ( n59508 , n59507 );
not ( n10138 , n59508 );
not ( n10139 , n59480 );
and ( n10140 , n10114 , n59432 );
not ( n10141 , n10114 );
not ( n10142 , n59432 );
and ( n10143 , n10141 , n10142 );
nor ( n10144 , n10140 , n10143 );
not ( n10145 , n10144 );
not ( n10146 , n10145 );
or ( n10147 , n10139 , n10146 );
buf ( n59519 , n59420 );
buf ( n59520 , n10099 );
and ( n59521 , n59519 , n59520 );
buf ( n59522 , n59521 );
buf ( n59523 , n59522 );
not ( n59524 , n59523 );
buf ( n59525 , n59524 );
not ( n10155 , n59525 );
not ( n10156 , n59394 );
or ( n10157 , n10155 , n10156 );
not ( n10158 , n59391 );
not ( n10159 , n59522 );
or ( n10160 , n10158 , n10159 );
buf ( n59532 , n59445 );
buf ( n59533 , n384 );
or ( n10163 , n59532 , n59533 );
buf ( n59535 , n59491 );
nand ( n10165 , n10163 , n59535 );
buf ( n59537 , n10165 );
nand ( n10167 , n10160 , n59537 );
nand ( n10168 , n10157 , n10167 );
nand ( n10169 , n10147 , n10168 );
buf ( n59541 , n10169 );
nand ( n10171 , n10144 , n10099 );
buf ( n59543 , n10171 );
nand ( n10173 , n59541 , n59543 );
buf ( n59545 , n10173 );
buf ( n59546 , n59545 );
not ( n10176 , n59546 );
or ( n59548 , n10138 , n10176 );
buf ( n59549 , n59504 );
not ( n10179 , n59549 );
buf ( n59551 , n10121 );
nand ( n10181 , n10179 , n59551 );
buf ( n59553 , n10181 );
buf ( n59554 , n59553 );
nand ( n10184 , n59548 , n59554 );
buf ( n59556 , n10184 );
buf ( n59557 , n59556 );
not ( n10187 , n59557 );
or ( n59559 , n59441 , n10187 );
buf ( n59560 , n59436 );
not ( n10190 , n59560 );
buf ( n59562 , n10055 );
nand ( n10192 , n10190 , n59562 );
buf ( n59564 , n10192 );
buf ( n59565 , n59564 );
nand ( n10195 , n59559 , n59565 );
buf ( n59567 , n10195 );
buf ( n59568 , n59567 );
buf ( n10198 , n59568 );
buf ( n59570 , n10198 );
buf ( n59571 , n59570 );
not ( n10201 , n59571 );
buf ( n10202 , n10201 );
buf ( n59574 , n10202 );
buf ( n59575 , n57008 );
not ( n59576 , n59575 );
buf ( n59577 , n59576 );
buf ( n59578 , n59577 );
buf ( n59579 , n6312 );
or ( n59580 , n59578 , n59579 );
buf ( n59581 , n55628 );
buf ( n59582 , n56768 );
or ( n59583 , n59581 , n59582 );
nand ( n59584 , n59580 , n59583 );
buf ( n59585 , n59584 );
xor ( n59586 , n59585 , n6363 );
buf ( n59587 , n55731 );
buf ( n59588 , n55675 );
buf ( n59589 , n413 );
nand ( n10219 , n59588 , n59589 );
buf ( n59591 , n10219 );
buf ( n59592 , n59591 );
xor ( n10222 , n59587 , n59592 );
buf ( n59594 , n57196 );
and ( n10224 , n10222 , n59594 );
and ( n59596 , n59587 , n59592 );
or ( n10226 , n10224 , n59596 );
buf ( n59598 , n10226 );
and ( n10228 , n59586 , n59598 );
and ( n10229 , n59585 , n6363 );
or ( n10230 , n10228 , n10229 );
buf ( n59602 , n10230 );
buf ( n59603 , n55641 );
buf ( n59604 , n411 );
nand ( n10234 , n59603 , n59604 );
buf ( n59606 , n10234 );
buf ( n59607 , n59606 );
and ( n10237 , n59602 , n59607 );
buf ( n59609 , n10237 );
buf ( n59610 , n59609 );
not ( n10240 , n59610 );
buf ( n59612 , n10230 );
buf ( n59613 , n59606 );
or ( n10243 , n59612 , n59613 );
buf ( n59615 , n10243 );
buf ( n59616 , n59615 );
nand ( n10246 , n10240 , n59616 );
buf ( n59618 , n10246 );
xor ( n10248 , n59587 , n59592 );
xor ( n10249 , n10248 , n59594 );
buf ( n59621 , n10249 );
xor ( n10251 , n59621 , n55731 );
buf ( n59623 , n6363 );
buf ( n59624 , n415 );
nor ( n59625 , n59623 , n59624 );
buf ( n59626 , n59625 );
buf ( n59627 , n59626 );
buf ( n59628 , n55660 );
not ( n59629 , n59628 );
buf ( n59630 , n59629 );
buf ( n59631 , n59630 );
buf ( n59632 , n55671 );
or ( n10262 , n59631 , n59632 );
buf ( n59634 , n6337 );
buf ( n59635 , n6322 );
or ( n10264 , n59634 , n59635 );
nand ( n10265 , n10262 , n10264 );
buf ( n59638 , n10265 );
buf ( n59639 , n59638 );
xor ( n59640 , n59627 , n59639 );
buf ( n59641 , n57196 );
and ( n10270 , n59640 , n59641 );
and ( n59643 , n59627 , n59639 );
or ( n59644 , n10270 , n59643 );
buf ( n59645 , n59644 );
and ( n59646 , n10251 , n59645 );
and ( n59647 , n59621 , n55731 );
or ( n59648 , n59646 , n59647 );
xor ( n59649 , n59585 , n6363 );
xor ( n10278 , n59649 , n59598 );
and ( n59651 , n59648 , n10278 );
buf ( n59652 , n7791 );
buf ( n59653 , n415 );
buf ( n59654 , n55731 );
and ( n59655 , n59653 , n59654 );
not ( n10284 , n59653 );
buf ( n59657 , n6363 );
and ( n59658 , n10284 , n59657 );
nor ( n10287 , n59655 , n59658 );
buf ( n59660 , n10287 );
buf ( n59661 , n59660 );
or ( n59662 , n59652 , n59661 );
buf ( n59663 , n57131 );
nand ( n10292 , n59662 , n59663 );
buf ( n10293 , n10292 );
buf ( n59666 , n10293 );
buf ( n59667 , n6363 );
xor ( n10296 , n59666 , n59667 );
xor ( n10297 , n59627 , n59639 );
xor ( n10298 , n10297 , n59641 );
buf ( n59671 , n10298 );
buf ( n59672 , n59671 );
and ( n59673 , n10296 , n59672 );
and ( n59674 , n59666 , n59667 );
or ( n10301 , n59673 , n59674 );
buf ( n59676 , n10301 );
xor ( n10303 , n59621 , n55731 );
xor ( n10304 , n10303 , n59645 );
and ( n10305 , n59676 , n10304 );
buf ( n59680 , n6370 );
not ( n10307 , n59680 );
buf ( n59682 , n10307 );
buf ( n59683 , n59682 );
buf ( n59684 , n415 );
buf ( n59685 , n416 );
and ( n10312 , n59684 , n59685 );
buf ( n59687 , n55715 );
nor ( n10314 , n10312 , n59687 );
buf ( n10315 , n10314 );
buf ( n59690 , n10315 );
or ( n10317 , n59683 , n59690 );
buf ( n59692 , n6398 );
nand ( n10319 , n10317 , n59692 );
buf ( n59694 , n10319 );
buf ( n59695 , n59694 );
buf ( n59696 , n55691 );
xor ( n59697 , n59695 , n59696 );
xnor ( n59698 , n59660 , n7801 );
buf ( n59699 , n59698 );
xor ( n59700 , n59697 , n59699 );
buf ( n59701 , n59700 );
buf ( n59702 , n55789 );
not ( n10329 , n59702 );
buf ( n59704 , n10329 );
buf ( n59705 , n59704 );
buf ( n59706 , n10315 );
buf ( n59707 , n57196 );
and ( n10334 , n59706 , n59707 );
not ( n10335 , n59706 );
buf ( n59710 , n6320 );
and ( n10337 , n10335 , n59710 );
nor ( n10338 , n10334 , n10337 );
buf ( n59713 , n10338 );
buf ( n59714 , n59713 );
not ( n10341 , n59714 );
buf ( n59716 , n55691 );
not ( n10343 , n59716 );
and ( n59718 , n10341 , n10343 );
buf ( n59719 , n59713 );
buf ( n59720 , n55691 );
and ( n10347 , n59719 , n59720 );
nor ( n59722 , n59718 , n10347 );
buf ( n59723 , n59722 );
buf ( n59724 , n59723 );
or ( n59725 , n59705 , n59724 );
buf ( n59726 , n55796 );
nand ( n59727 , n59725 , n59726 );
buf ( n59728 , n59727 );
nor ( n59729 , n59701 , n59728 );
xor ( n59730 , n59695 , n59696 );
and ( n10357 , n59730 , n59699 );
and ( n59732 , n59695 , n59696 );
or ( n59733 , n10357 , n59732 );
buf ( n59734 , n59733 );
xor ( n59735 , n59666 , n59667 );
xor ( n59736 , n59735 , n59672 );
buf ( n59737 , n59736 );
nor ( n59738 , n59734 , n59737 );
not ( n59739 , n6477 );
buf ( n59740 , n59352 );
buf ( n59741 , n59740 );
buf ( n59742 , n59741 );
buf ( n59743 , n59723 );
buf ( n59744 , n57216 );
xor ( n10371 , n59743 , n59744 );
buf ( n59746 , n10371 );
buf ( n59747 , n59746 );
not ( n59748 , n59747 );
buf ( n59749 , n6450 );
not ( n59750 , n59749 );
and ( n59751 , n59748 , n59750 );
buf ( n59752 , n59746 );
buf ( n59753 , n6450 );
and ( n59754 , n59752 , n59753 );
nor ( n10381 , n59751 , n59754 );
buf ( n59756 , n10381 );
buf ( n10383 , n59756 );
buf ( n59758 , n55799 );
not ( n10385 , n59758 );
buf ( n10386 , n10385 );
buf ( n59761 , n10386 );
nand ( n10388 , n10383 , n59761 );
buf ( n59763 , n10388 );
nand ( n10390 , n59739 , n59742 , n59763 );
or ( n59765 , n59729 , n59738 , n10390 );
buf ( n59766 , n59756 );
buf ( n59767 , n10386 );
nor ( n10394 , n59766 , n59767 );
buf ( n59769 , n10394 );
nor ( n10396 , n59729 , n59738 );
and ( n10397 , n59769 , n10396 );
nand ( n10398 , n59701 , n59728 );
or ( n10399 , n10398 , n59738 );
nand ( n10400 , n59734 , n59737 );
nand ( n10401 , n10399 , n10400 );
nor ( n10402 , n10397 , n10401 );
nand ( n10403 , n59765 , n10402 );
xor ( n10404 , n59621 , n55731 );
xor ( n10405 , n10404 , n59645 );
and ( n10406 , n10403 , n10405 );
and ( n10407 , n59676 , n10403 );
or ( n10408 , n10305 , n10406 , n10407 );
xor ( n10409 , n59585 , n6363 );
xor ( n10410 , n10409 , n59598 );
and ( n10411 , n10408 , n10410 );
and ( n10412 , n59648 , n10408 );
or ( n10413 , n59651 , n10411 , n10412 );
xnor ( n10414 , n59618 , n10413 );
buf ( n59789 , n10414 );
nand ( n59790 , n59574 , n59789 );
buf ( n59791 , n59790 );
buf ( n59792 , n59791 );
buf ( n59793 , n10414 );
not ( n10420 , n59793 );
buf ( n59795 , n59570 );
nand ( n10422 , n10420 , n59795 );
buf ( n59797 , n10422 );
buf ( n59798 , n59797 );
nand ( n10425 , n59792 , n59798 );
buf ( n59800 , n10425 );
buf ( n59801 , n59800 );
buf ( n59802 , n59800 );
not ( n10429 , n59802 );
buf ( n59804 , n10429 );
buf ( n59805 , n59804 );
xor ( n10432 , n59585 , n6363 );
xor ( n10433 , n10432 , n59598 );
xor ( n59808 , n59648 , n10408 );
xor ( n10435 , n10433 , n59808 );
buf ( n59810 , n10435 );
not ( n10437 , n59810 );
buf ( n59812 , n59567 );
nand ( n59813 , n10437 , n59812 );
buf ( n59814 , n59813 );
not ( n10441 , n59814 );
buf ( n59816 , n59397 );
not ( n10443 , n59816 );
buf ( n59818 , n59424 );
nand ( n10445 , n10443 , n59818 );
buf ( n59820 , n10445 );
not ( n10447 , n59820 );
buf ( n59822 , n10447 );
not ( n10449 , n59822 );
buf ( n59824 , n55814 );
not ( n10451 , n59824 );
buf ( n59826 , n59355 );
not ( n10453 , n59826 );
or ( n10454 , n10451 , n10453 );
buf ( n59829 , n59362 );
nand ( n10456 , n10454 , n59829 );
buf ( n59831 , n10456 );
buf ( n59832 , n59831 );
buf ( n59833 , n59394 );
nand ( n10460 , n59832 , n59833 );
buf ( n59835 , n10460 );
buf ( n59836 , n59835 );
not ( n10463 , n59836 );
or ( n10464 , n10449 , n10463 );
buf ( n59839 , n59480 );
buf ( n59840 , n384 );
nand ( n10467 , n59839 , n59840 );
buf ( n10468 , n10467 );
buf ( n59843 , n10468 );
buf ( n59844 , n59431 );
buf ( n59845 , n384 );
nand ( n59846 , n59844 , n59845 );
buf ( n59847 , n59846 );
buf ( n59848 , n59847 );
nand ( n59849 , n59843 , n59848 );
buf ( n59850 , n59849 );
buf ( n59851 , n59850 );
buf ( n59852 , n59484 );
not ( n59853 , n59852 );
buf ( n59854 , n59853 );
buf ( n59855 , n59854 );
or ( n59856 , n59851 , n59855 );
buf ( n59857 , n59856 );
buf ( n59858 , n59857 );
nand ( n10485 , n10464 , n59858 );
buf ( n59860 , n10485 );
buf ( n59861 , n59860 );
not ( n59862 , n59861 );
buf ( n59863 , n59862 );
buf ( n59864 , n384 );
buf ( n59865 , n10047 );
and ( n59866 , n59864 , n59865 );
not ( n59867 , n59864 );
buf ( n59868 , n59431 );
and ( n59869 , n59867 , n59868 );
nor ( n59870 , n59866 , n59869 );
buf ( n59871 , n59870 );
buf ( n59872 , n59871 );
buf ( n59873 , n59391 );
and ( n10500 , n59872 , n59873 );
buf ( n59875 , n59871 );
not ( n10502 , n59875 );
buf ( n59877 , n10502 );
buf ( n59878 , n59877 );
buf ( n59879 , n59394 );
and ( n10506 , n59878 , n59879 );
nor ( n59881 , n10500 , n10506 );
buf ( n59882 , n59881 );
xor ( n10509 , n59863 , n59882 );
buf ( n59884 , n59473 );
buf ( n59885 , n384 );
and ( n10512 , n59884 , n59885 );
buf ( n59887 , n59854 );
nor ( n10514 , n10512 , n59887 );
buf ( n59889 , n10514 );
buf ( n59890 , n59889 );
buf ( n59891 , n59835 );
xor ( n10518 , n59890 , n59891 );
not ( n10519 , n10099 );
nand ( n10520 , n10519 , n10129 );
and ( n10521 , n10520 , n59525 );
buf ( n59896 , n10521 );
xor ( n10523 , n10518 , n59896 );
buf ( n59898 , n10523 );
xor ( n10525 , n10509 , n59898 );
buf ( n59900 , n10525 );
not ( n10527 , n59900 );
buf ( n59902 , n59857 );
not ( n10529 , n59902 );
buf ( n59904 , n59835 );
not ( n10531 , n59904 );
or ( n10532 , n10529 , n10531 );
buf ( n59907 , n59857 );
buf ( n59908 , n59835 );
or ( n10535 , n59907 , n59908 );
nand ( n10536 , n10532 , n10535 );
buf ( n59911 , n10536 );
buf ( n59912 , n59911 );
not ( n59913 , n59912 );
buf ( n59914 , n10447 );
not ( n59915 , n59914 );
or ( n10542 , n59913 , n59915 );
buf ( n59917 , n10447 );
buf ( n59918 , n59911 );
or ( n10545 , n59917 , n59918 );
nand ( n10546 , n10542 , n10545 );
buf ( n59921 , n10546 );
buf ( n59922 , n59921 );
not ( n59923 , n59922 );
buf ( n59924 , n59871 );
buf ( n59925 , n59480 );
and ( n10552 , n59924 , n59925 );
buf ( n59927 , n59877 );
buf ( n59928 , n10099 );
and ( n10555 , n59927 , n59928 );
nor ( n10556 , n10552 , n10555 );
buf ( n59931 , n10556 );
buf ( n59932 , n59931 );
nand ( n10559 , n59923 , n59932 );
buf ( n59934 , n10559 );
not ( n10561 , n59934 );
not ( n59936 , n59863 );
or ( n10563 , n10561 , n59936 );
buf ( n59938 , n59921 );
buf ( n59939 , n59931 );
not ( n10566 , n59939 );
buf ( n59941 , n10566 );
buf ( n59942 , n59941 );
nand ( n10569 , n59938 , n59942 );
buf ( n59944 , n10569 );
nand ( n59945 , n10563 , n59944 );
buf ( n59946 , n59945 );
not ( n10573 , n59946 );
buf ( n59948 , n10573 );
buf ( n59949 , n59948 );
nand ( n10576 , n10527 , n59949 );
buf ( n10577 , n10576 );
buf ( n59952 , n10577 );
buf ( n59953 , n59525 );
buf ( n59954 , n59537 );
not ( n59955 , n59954 );
buf ( n59956 , n59391 );
not ( n10583 , n59956 );
and ( n10584 , n59955 , n10583 );
buf ( n59959 , n59537 );
buf ( n59960 , n59391 );
and ( n10587 , n59959 , n59960 );
nor ( n10588 , n10584 , n10587 );
buf ( n59963 , n10588 );
buf ( n59964 , n59963 );
xor ( n10591 , n59953 , n59964 );
buf ( n59966 , n10591 );
xor ( n10593 , n59890 , n59891 );
and ( n10594 , n10593 , n59896 );
and ( n10595 , n59890 , n59891 );
or ( n10596 , n10594 , n10595 );
buf ( n59971 , n10596 );
xor ( n59972 , n59966 , n59971 );
xnor ( n10599 , n10521 , n10047 );
xnor ( n10600 , n59972 , n10599 );
not ( n59975 , n10600 );
not ( n59976 , n59898 );
not ( n10603 , n59882 );
and ( n59978 , n59976 , n10603 );
buf ( n59979 , n59898 );
buf ( n59980 , n59882 );
nand ( n59981 , n59979 , n59980 );
buf ( n59982 , n59981 );
and ( n10609 , n59982 , n59863 );
nor ( n59984 , n59978 , n10609 );
nand ( n10611 , n59975 , n59984 );
buf ( n59986 , n10611 );
and ( n10613 , n59952 , n59986 );
buf ( n59988 , n10613 );
buf ( n10615 , n10055 );
not ( n10616 , n10615 );
buf ( n10617 , n59436 );
not ( n10618 , n10617 );
and ( n10619 , n10616 , n10618 );
buf ( n59994 , n10055 );
buf ( n59995 , n59436 );
and ( n59996 , n59994 , n59995 );
nor ( n10623 , n10619 , n59996 );
buf ( n10624 , n10623 );
or ( n59999 , n59556 , n10624 );
nand ( n60000 , n59556 , n10624 );
not ( n10627 , n59729 );
and ( n60002 , n10627 , n10398 );
not ( n60003 , n60002 );
not ( n10630 , n59769 );
nand ( n60005 , n10630 , n10390 );
not ( n60006 , n60005 );
or ( n10633 , n60003 , n60006 );
or ( n10634 , n60005 , n60002 );
nand ( n10635 , n10633 , n10634 );
nand ( n60010 , n59999 , n60000 , n10635 );
xor ( n60011 , n59504 , n10121 );
buf ( n10638 , n59545 );
and ( n10639 , n60011 , n10638 );
not ( n10640 , n60011 );
not ( n60015 , n10638 );
and ( n60016 , n10640 , n60015 );
nor ( n10643 , n10639 , n60016 );
buf ( n60018 , n59769 );
not ( n60019 , n60018 );
buf ( n60020 , n59763 );
nand ( n60021 , n60019 , n60020 );
buf ( n60022 , n60021 );
buf ( n60023 , n60022 );
not ( n60024 , n60023 );
buf ( n60025 , n59742 );
not ( n60026 , n60025 );
or ( n60027 , n60024 , n60026 );
buf ( n60028 , n59742 );
buf ( n60029 , n60022 );
or ( n60030 , n60028 , n60029 );
nand ( n10657 , n60027 , n60030 );
buf ( n10658 , n10657 );
buf ( n10659 , n10658 );
not ( n10660 , n10659 );
buf ( n10661 , n10660 );
nand ( n60036 , n10643 , n10661 );
and ( n10663 , n60010 , n60036 );
xor ( n60038 , n59621 , n55731 );
xor ( n60039 , n60038 , n59645 );
xor ( n10666 , n59676 , n10403 );
xor ( n10667 , n60039 , n10666 );
buf ( n60042 , n10667 );
not ( n10669 , n60042 );
buf ( n60044 , n59567 );
nand ( n60045 , n10669 , n60044 );
buf ( n60046 , n60045 );
not ( n60047 , n10627 );
not ( n10674 , n60005 );
or ( n60049 , n60047 , n10674 );
nand ( n10676 , n60049 , n10398 );
not ( n60051 , n10400 );
nor ( n60052 , n60051 , n59738 );
and ( n10679 , n10676 , n60052 );
not ( n60054 , n10676 );
xnor ( n60055 , n59737 , n59734 );
and ( n10682 , n60054 , n60055 );
nor ( n60057 , n10679 , n10682 );
buf ( n60058 , n60057 );
not ( n10685 , n60058 );
buf ( n60060 , n59567 );
nand ( n60061 , n10685 , n60060 );
buf ( n60062 , n60061 );
and ( n10689 , n60046 , n60062 );
xor ( n60064 , n59432 , n10099 );
xor ( n60065 , n60064 , n10114 );
xnor ( n10692 , n60065 , n10168 );
not ( n10693 , n59966 );
not ( n60068 , n10599 );
or ( n10695 , n10693 , n60068 );
or ( n60070 , n10599 , n59966 );
nand ( n10697 , n60070 , n59971 );
nand ( n10698 , n10695 , n10697 );
nand ( n10699 , n10692 , n10698 );
and ( n10700 , n59988 , n10663 , n10689 , n10699 );
not ( n10701 , n10700 );
buf ( n60076 , n10099 );
buf ( n60077 , n59391 );
nor ( n10704 , n60076 , n60077 );
buf ( n60079 , n10704 );
buf ( n60080 , n60079 );
buf ( n60081 , n59941 );
xor ( n10708 , n60080 , n60081 );
buf ( n60083 , n59820 );
and ( n10710 , n10708 , n60083 );
and ( n10711 , n60080 , n60081 );
or ( n60086 , n10710 , n10711 );
buf ( n60087 , n60086 );
xor ( n60088 , n59931 , n60087 );
not ( n60089 , n59921 );
xnor ( n10716 , n60088 , n60089 );
buf ( n60091 , n59480 );
buf ( n60092 , n59391 );
and ( n60093 , n60091 , n60092 );
buf ( n60094 , n59394 );
buf ( n60095 , n10099 );
and ( n60096 , n60094 , n60095 );
nor ( n60097 , n60093 , n60096 );
buf ( n60098 , n60097 );
buf ( n60099 , n60098 );
buf ( n60100 , n59431 );
buf ( n60101 , n384 );
nor ( n10728 , n60100 , n60101 );
buf ( n60103 , n10728 );
buf ( n60104 , n60103 );
or ( n60105 , n60099 , n60104 );
buf ( n60106 , n59847 );
nand ( n10733 , n60105 , n60106 );
buf ( n10734 , n10733 );
not ( n60109 , n10734 );
buf ( n60110 , n60098 );
not ( n10737 , n60110 );
buf ( n60112 , n10737 );
buf ( n60113 , n60112 );
buf ( n60114 , n59871 );
or ( n60115 , n60113 , n60114 );
buf ( n60116 , n60098 );
buf ( n60117 , n59877 );
or ( n60118 , n60116 , n60117 );
nand ( n60119 , n60115 , n60118 );
buf ( n60120 , n60119 );
buf ( n60121 , n60120 );
buf ( n60122 , n60079 );
not ( n10749 , n60122 );
buf ( n60124 , n59491 );
buf ( n60125 , n59484 );
nand ( n10752 , n10749 , n60124 , n60125 );
buf ( n60127 , n10752 );
buf ( n60128 , n60127 );
xor ( n10755 , n60121 , n60128 );
buf ( n60130 , n60079 );
buf ( n60131 , n384 );
xor ( n10758 , n60130 , n60131 );
buf ( n60133 , n60112 );
buf ( n60134 , n10047 );
or ( n10761 , n60133 , n60134 );
buf ( n60136 , n60098 );
buf ( n60137 , n59431 );
or ( n10764 , n60136 , n60137 );
nand ( n60139 , n10761 , n10764 );
buf ( n60140 , n60139 );
buf ( n60141 , n60140 );
and ( n60142 , n10758 , n60141 );
and ( n60143 , n60130 , n60131 );
or ( n10770 , n60142 , n60143 );
buf ( n60145 , n10770 );
buf ( n60146 , n60145 );
and ( n10773 , n10755 , n60146 );
and ( n60148 , n60121 , n60128 );
or ( n10775 , n10773 , n60148 );
buf ( n60150 , n10775 );
not ( n10777 , n60150 );
or ( n60152 , n60109 , n10777 );
not ( n60153 , n10734 );
not ( n10780 , n60150 );
and ( n10781 , n60153 , n10780 );
not ( n60156 , n10781 );
xor ( n60157 , n60080 , n60081 );
xor ( n10784 , n60157 , n60083 );
buf ( n60159 , n10784 );
nand ( n60160 , n60156 , n60159 );
nand ( n10787 , n60152 , n60160 );
not ( n10788 , n10787 );
and ( n10789 , n10716 , n10788 );
not ( n10790 , n60159 );
xor ( n60165 , n60153 , n10780 );
and ( n10792 , n10790 , n60165 );
not ( n10793 , n10790 );
not ( n60168 , n60165 );
and ( n10795 , n10793 , n60168 );
or ( n60170 , n10792 , n10795 );
xor ( n60171 , n60121 , n60128 );
xor ( n10798 , n60171 , n60146 );
buf ( n60173 , n10798 );
not ( n60174 , n60173 );
xor ( n60175 , n60130 , n60131 );
xor ( n10802 , n60175 , n60141 );
buf ( n60177 , n10802 );
buf ( n60178 , n60177 );
buf ( n60179 , n59850 );
xor ( n10806 , n60178 , n60179 );
buf ( n60181 , n10468 );
not ( n10808 , n60181 );
buf ( n60183 , n10808 );
buf ( n60184 , n60183 );
buf ( n60185 , n59871 );
and ( n60186 , n60184 , n60185 );
buf ( n60187 , n10468 );
buf ( n60188 , n59877 );
and ( n10815 , n60187 , n60188 );
nor ( n60190 , n60186 , n10815 );
buf ( n60191 , n60190 );
buf ( n60192 , n60191 );
buf ( n60193 , n60098 );
or ( n10820 , n60192 , n60193 );
buf ( n60195 , n60191 );
buf ( n60196 , n60098 );
and ( n10823 , n60195 , n60196 );
buf ( n60198 , n384 );
buf ( n60199 , n10099 );
and ( n60200 , n60198 , n60199 );
not ( n10827 , n60198 );
buf ( n60202 , n59480 );
and ( n60203 , n10827 , n60202 );
nor ( n10830 , n60200 , n60203 );
buf ( n10831 , n10830 );
buf ( n60206 , n10831 );
not ( n10833 , n60206 );
buf ( n60208 , n60183 );
nor ( n10835 , n10833 , n60208 );
buf ( n60210 , n10835 );
buf ( n60211 , n60210 );
buf ( n60212 , n59391 );
or ( n10839 , n60211 , n60212 );
buf ( n60214 , n10839 );
buf ( n60215 , n60214 );
nor ( n10842 , n10823 , n60215 );
buf ( n60217 , n10842 );
buf ( n60218 , n60217 );
not ( n10845 , n60218 );
buf ( n60220 , n10845 );
buf ( n60221 , n60220 );
nand ( n10848 , n10820 , n60221 );
buf ( n60223 , n10848 );
buf ( n60224 , n60223 );
and ( n10851 , n10806 , n60224 );
and ( n60226 , n60178 , n60179 );
or ( n10853 , n10851 , n60226 );
buf ( n60228 , n10853 );
not ( n10855 , n60228 );
or ( n10856 , n60174 , n10855 );
or ( n10857 , n60228 , n60173 );
nand ( n10858 , n10857 , n10129 );
nand ( n10859 , n10856 , n10858 );
nor ( n10860 , n60170 , n10859 );
nor ( n10861 , n10789 , n10860 );
buf ( n60236 , n10861 );
not ( n10863 , n60236 );
buf ( n60238 , n57120 );
not ( n60239 , n60238 );
not ( n60240 , n56468 );
nand ( n60241 , n60240 , n57283 );
buf ( n60242 , n60241 );
not ( n60243 , n60242 );
buf ( n60244 , n57280 );
nor ( n60245 , n60243 , n60244 );
buf ( n60246 , n60245 );
not ( n10873 , n60246 );
not ( n60248 , n59290 );
or ( n60249 , n10873 , n60248 );
buf ( n60250 , n57060 );
not ( n60251 , n60250 );
buf ( n60252 , n60251 );
nand ( n10879 , n60249 , n60252 );
buf ( n60254 , n10879 );
not ( n60255 , n60254 );
or ( n10882 , n60239 , n60255 );
buf ( n60257 , n59303 );
nand ( n60258 , n10882 , n60257 );
buf ( n60259 , n60258 );
buf ( n60260 , n60259 );
buf ( n60261 , n59306 );
buf ( n60262 , n57187 );
nand ( n10889 , n60261 , n60262 );
buf ( n60264 , n10889 );
buf ( n60265 , n60264 );
xnor ( n60266 , n60260 , n60265 );
buf ( n60267 , n60266 );
buf ( n60268 , n60267 );
buf ( n60269 , n10831 );
not ( n10896 , n60269 );
buf ( n60271 , n59394 );
not ( n10898 , n60271 );
buf ( n60273 , n10468 );
not ( n10900 , n60273 );
or ( n60275 , n10898 , n10900 );
buf ( n60276 , n10468 );
buf ( n60277 , n59394 );
or ( n60278 , n60276 , n60277 );
nand ( n60279 , n60275 , n60278 );
buf ( n60280 , n60279 );
buf ( n60281 , n60280 );
not ( n10908 , n60281 );
or ( n60283 , n10896 , n10908 );
buf ( n60284 , n60280 );
buf ( n60285 , n10831 );
or ( n60286 , n60284 , n60285 );
nand ( n10913 , n60283 , n60286 );
buf ( n10914 , n10913 );
buf ( n60289 , n10914 );
not ( n10916 , n60289 );
buf ( n60291 , n60214 );
nand ( n10918 , n10916 , n60291 );
buf ( n60293 , n10918 );
buf ( n60294 , n60293 );
nand ( n10921 , n60268 , n60294 );
buf ( n60296 , n10921 );
buf ( n60297 , n60191 );
buf ( n60298 , n60098 );
and ( n60299 , n60297 , n60298 );
not ( n10926 , n60297 );
buf ( n60301 , n60112 );
and ( n60302 , n10926 , n60301 );
nor ( n10929 , n60299 , n60302 );
buf ( n10930 , n10929 );
buf ( n60305 , n10930 );
buf ( n60306 , n60214 );
and ( n10933 , n60305 , n60306 );
buf ( n60308 , n10930 );
buf ( n60309 , n60214 );
nor ( n10936 , n60308 , n60309 );
buf ( n60311 , n10936 );
buf ( n60312 , n60311 );
nor ( n10939 , n10933 , n60312 );
buf ( n60314 , n10939 );
or ( n10941 , n54653 , n54668 );
not ( n10942 , n54673 );
nand ( n10943 , n10942 , n54864 );
and ( n60318 , n10941 , n10943 );
not ( n10945 , n60318 );
not ( n60320 , n54570 );
not ( n60321 , n54614 );
and ( n10948 , n60320 , n60321 );
nor ( n60323 , n10948 , n54718 );
or ( n60324 , n54648 , n54619 );
and ( n10951 , n54714 , n60323 , n60324 );
not ( n10952 , n10951 );
not ( n10953 , n4188 );
not ( n10954 , n10953 );
nand ( n10955 , n10954 , n53300 );
not ( n10956 , n10955 );
not ( n10957 , n53300 );
nand ( n10958 , n10957 , n10953 );
not ( n10959 , n53059 );
not ( n60334 , n54847 );
or ( n60335 , n10959 , n60334 );
nand ( n60336 , n60335 , n54860 );
not ( n10963 , n60336 );
not ( n60338 , n54854 );
or ( n60339 , n10963 , n60338 );
nand ( n10966 , n60339 , n54857 );
nor ( n60341 , n54851 , n54857 );
not ( n60342 , n60341 );
not ( n10969 , n60336 );
or ( n10970 , n60342 , n10969 );
nand ( n60345 , n10970 , n54743 );
nand ( n10972 , n10958 , n10966 , n60345 );
not ( n10973 , n10972 );
or ( n60348 , n10956 , n10973 );
not ( n60349 , n53725 );
not ( n10976 , n53513 );
nand ( n60351 , n60349 , n10976 );
nand ( n60352 , n60348 , n60351 );
not ( n10979 , n53730 );
not ( n60354 , n53945 );
or ( n60355 , n10979 , n60354 );
buf ( n60356 , n53513 );
nand ( n10983 , n60356 , n53725 );
nand ( n60358 , n60355 , n10983 );
not ( n10985 , n60358 );
nand ( n10986 , n60352 , n10985 );
nor ( n10987 , n4777 , n53950 );
nor ( n10988 , n10987 , n54734 );
not ( n60363 , n54225 );
not ( n10990 , n4782 );
nand ( n60365 , n60363 , n10990 );
nand ( n10992 , n10986 , n10988 , n60365 );
not ( n10993 , n10992 );
not ( n10994 , n54342 );
not ( n10995 , n10994 );
not ( n10996 , n54230 );
not ( n10997 , n10996 );
and ( n10998 , n10995 , n10997 );
not ( n10999 , n4782 );
not ( n11000 , n54225 );
or ( n11001 , n10999 , n11000 );
nand ( n11002 , n4777 , n53950 );
nand ( n11003 , n11001 , n11002 );
nand ( n11004 , n5546 , n10990 );
and ( n60379 , n11003 , n11004 );
nor ( n11006 , n10998 , n60379 );
not ( n60381 , n11006 );
or ( n11008 , n10993 , n60381 );
not ( n11009 , n54342 );
nand ( n11010 , n11009 , n10996 );
nand ( n11011 , n11008 , n11010 );
not ( n11012 , n11011 );
not ( n60387 , n11012 );
or ( n11014 , n10952 , n60387 );
not ( n60389 , n60323 );
or ( n60390 , n54730 , n5405 );
nand ( n11017 , n60390 , n54722 );
not ( n11018 , n11017 );
or ( n11019 , n60389 , n11018 );
not ( n11020 , n54570 );
not ( n11021 , n54614 );
and ( n11022 , n11020 , n11021 );
nand ( n11023 , n54565 , n54510 );
nor ( n60398 , n11022 , n11023 );
and ( n11025 , n54570 , n54614 );
nor ( n60400 , n60398 , n11025 );
nand ( n60401 , n11019 , n60400 );
buf ( n11028 , n60324 );
and ( n60403 , n60401 , n11028 );
and ( n60404 , n54619 , n54648 );
nor ( n11031 , n60403 , n60404 );
nand ( n11032 , n11014 , n11031 );
not ( n11033 , n11032 );
or ( n11034 , n10945 , n11033 );
not ( n60409 , n54864 );
nand ( n60410 , n60409 , n54673 );
not ( n11037 , n60410 );
not ( n60412 , n10943 );
nand ( n60413 , n54653 , n54668 );
nor ( n11040 , n60412 , n60413 );
nor ( n60415 , n11037 , n11040 );
nand ( n60416 , n11034 , n60415 );
and ( n60417 , n60416 , n378 );
xor ( n11044 , n60314 , n60417 );
buf ( n60419 , n59313 );
buf ( n60420 , n57172 );
nand ( n60421 , n60419 , n60420 );
buf ( n60422 , n60421 );
buf ( n60423 , n60422 );
not ( n60424 , n60423 );
and ( n60425 , n57120 , n57187 );
buf ( n60426 , n60425 );
not ( n11053 , n60426 );
buf ( n60428 , n10879 );
not ( n11055 , n60428 );
or ( n60430 , n11053 , n11055 );
buf ( n60431 , n59306 );
not ( n60432 , n60431 );
buf ( n60433 , n59303 );
not ( n60434 , n60433 );
or ( n11061 , n60432 , n60434 );
buf ( n60436 , n57187 );
nand ( n11063 , n11061 , n60436 );
buf ( n60438 , n11063 );
buf ( n60439 , n60438 );
nand ( n11066 , n60430 , n60439 );
buf ( n60441 , n11066 );
buf ( n60442 , n60441 );
not ( n11069 , n60442 );
or ( n11070 , n60424 , n11069 );
buf ( n60445 , n60441 );
buf ( n60446 , n60422 );
or ( n60447 , n60445 , n60446 );
nand ( n60448 , n11070 , n60447 );
buf ( n60449 , n60448 );
xnor ( n60450 , n11044 , n60449 );
not ( n60451 , n60450 );
nand ( n11078 , n60296 , n60451 );
buf ( n11079 , n11078 );
not ( n11080 , n11079 );
buf ( n11081 , n378 );
and ( n11082 , n10943 , n60410 );
not ( n60457 , n10941 );
not ( n60458 , n11032 );
or ( n11085 , n60457 , n60458 );
nand ( n11086 , n11085 , n60413 );
xor ( n60461 , n11082 , n11086 );
buf ( n60462 , n60461 );
not ( n60463 , n60462 );
buf ( n60464 , n60463 );
buf ( n60465 , n60464 );
not ( n60466 , n60465 );
buf ( n60467 , n60466 );
buf ( n11094 , n60467 );
and ( n11095 , n11081 , n11094 );
buf ( n60470 , n11095 );
buf ( n60471 , n60293 );
buf ( n60472 , n60267 );
xor ( n11099 , n60471 , n60472 );
buf ( n60474 , n11099 );
xor ( n11101 , n60470 , n60474 );
not ( n60476 , n59413 );
buf ( n60477 , n60476 );
not ( n60478 , n60477 );
not ( n11105 , n378 );
buf ( n60480 , n11105 );
not ( n11107 , n60480 );
buf ( n60482 , n60416 );
not ( n11109 , n60482 );
or ( n11110 , n11107 , n11109 );
buf ( n60485 , n60416 );
not ( n11112 , n60485 );
buf ( n60487 , n11112 );
buf ( n60488 , n60487 );
buf ( n11115 , n378 );
nand ( n11116 , n60488 , n11115 );
buf ( n60491 , n11116 );
buf ( n60492 , n60491 );
nand ( n11119 , n11110 , n60492 );
buf ( n60494 , n11119 );
buf ( n60495 , n60494 );
not ( n11122 , n60495 );
or ( n11123 , n60478 , n11122 );
not ( n60498 , n59415 );
buf ( n60499 , n60498 );
buf ( n60500 , n378 );
nand ( n60501 , n60499 , n60500 );
buf ( n60502 , n60501 );
buf ( n60503 , n60502 );
nand ( n11130 , n11123 , n60503 );
buf ( n60505 , n11130 );
and ( n60506 , n11101 , n60505 );
and ( n11133 , n60470 , n60474 );
or ( n11134 , n60506 , n11133 );
buf ( n60509 , n11134 );
not ( n11136 , n60509 );
or ( n60511 , n11080 , n11136 );
not ( n60512 , n60296 );
nand ( n11139 , n60512 , n60450 );
buf ( n60514 , n11139 );
nand ( n60515 , n60511 , n60514 );
buf ( n60516 , n60515 );
not ( n11143 , n60516 );
not ( n11144 , n60417 );
not ( n60519 , n60449 );
or ( n11146 , n11144 , n60519 );
not ( n60521 , n60417 );
not ( n11148 , n60521 );
buf ( n60523 , n60449 );
not ( n60524 , n60523 );
buf ( n60525 , n60524 );
not ( n11152 , n60525 );
or ( n60527 , n11148 , n11152 );
buf ( n60528 , n60314 );
not ( n11155 , n60528 );
buf ( n11156 , n11155 );
nand ( n60531 , n60527 , n11156 );
nand ( n60532 , n11146 , n60531 );
xor ( n11159 , n60178 , n60179 );
xor ( n60534 , n11159 , n60224 );
buf ( n60535 , n60534 );
buf ( n60536 , n60535 );
buf ( n60537 , n60441 );
buf ( n60538 , n57172 );
and ( n60539 , n60537 , n60538 );
buf ( n60540 , n59313 );
not ( n60541 , n60540 );
buf ( n60542 , n60541 );
buf ( n60543 , n60542 );
nor ( n60544 , n60539 , n60543 );
buf ( n60545 , n60544 );
buf ( n60546 , n60545 );
buf ( n11173 , n59329 );
buf ( n11174 , n57269 );
nand ( n11175 , n11173 , n11174 );
buf ( n11176 , n11175 );
buf ( n60551 , n11176 );
xor ( n11178 , n60546 , n60551 );
buf ( n11179 , n11178 );
buf ( n60554 , n11179 );
not ( n11181 , n60554 );
buf ( n60556 , n11181 );
buf ( n60557 , n60556 );
and ( n11184 , n60536 , n60557 );
not ( n11185 , n60536 );
buf ( n60560 , n11179 );
and ( n11187 , n11185 , n60560 );
nor ( n11188 , n11184 , n11187 );
buf ( n60563 , n11188 );
xor ( n11190 , n60532 , n60563 );
nand ( n11191 , n11143 , n11190 );
buf ( n60566 , n11191 );
not ( n11193 , n60532 );
buf ( n60568 , n60535 );
not ( n11195 , n60568 );
buf ( n60570 , n60556 );
nand ( n11197 , n11195 , n60570 );
buf ( n60572 , n11197 );
not ( n60573 , n60572 );
or ( n60574 , n11193 , n60573 );
buf ( n60575 , n11179 );
buf ( n60576 , n60535 );
nand ( n60577 , n60575 , n60576 );
buf ( n60578 , n60577 );
nand ( n60579 , n60574 , n60578 );
buf ( n60580 , n60579 );
not ( n11207 , n10129 );
not ( n11208 , n60228 );
not ( n11209 , n60173 );
not ( n11210 , n11209 );
and ( n11211 , n11208 , n11210 );
and ( n11212 , n60228 , n11209 );
nor ( n11213 , n11211 , n11212 );
not ( n11214 , n11213 );
or ( n11215 , n11207 , n11214 );
or ( n11216 , n10129 , n11213 );
nand ( n11217 , n11215 , n11216 );
buf ( n60592 , n11217 );
nor ( n11219 , n60580 , n60592 );
buf ( n60594 , n11219 );
buf ( n60595 , n60594 );
not ( n60596 , n60595 );
buf ( n60597 , n60596 );
buf ( n60598 , n60597 );
nand ( n11225 , n60566 , n60598 );
buf ( n60600 , n11225 );
buf ( n60601 , n60600 );
nor ( n11228 , n10863 , n60601 );
buf ( n60603 , n11228 );
not ( n11230 , n59941 );
not ( n11231 , n59921 );
or ( n11232 , n11230 , n11231 );
nand ( n11233 , n60089 , n59931 );
nand ( n60608 , n11232 , n11233 );
xnor ( n60609 , n59863 , n60608 );
not ( n11236 , n60609 );
buf ( n60611 , n59934 );
buf ( n60612 , n60087 );
nand ( n11239 , n60611 , n60612 );
buf ( n60614 , n11239 );
and ( n11241 , n59944 , n60614 );
nand ( n11242 , n11236 , n11241 );
and ( n11243 , n60603 , n11242 );
not ( n11244 , n11243 );
buf ( n60619 , n60476 );
not ( n11246 , n60619 );
buf ( n60621 , n378 );
not ( n11248 , n54570 );
not ( n11249 , n54614 );
and ( n11250 , n11248 , n11249 );
nor ( n11251 , n11250 , n11025 );
buf ( n60626 , n11251 );
not ( n11253 , n54871 );
not ( n11254 , n11017 );
or ( n11255 , n11253 , n11254 );
buf ( n11256 , n11023 );
nand ( n11257 , n11255 , n11256 );
not ( n11258 , n11257 );
not ( n11259 , n10992 );
not ( n11260 , n11259 );
buf ( n11261 , n11006 );
nand ( n11262 , n11260 , n11261 );
not ( n11263 , n54677 );
not ( n11264 , n54730 );
and ( n11265 , n11263 , n11264 , n11010 );
nand ( n11266 , n11262 , n11265 , n54871 );
nand ( n11267 , n11258 , n11266 );
buf ( n60642 , n11267 );
xor ( n11269 , n60626 , n60642 );
buf ( n60644 , n11269 );
buf ( n60645 , n60644 );
xor ( n11272 , n60621 , n60645 );
buf ( n60647 , n11272 );
buf ( n60648 , n60647 );
not ( n11275 , n60648 );
or ( n11276 , n11246 , n11275 );
buf ( n60651 , n378 );
and ( n11278 , n54714 , n60323 );
not ( n11279 , n11278 );
not ( n11280 , n11012 );
or ( n11281 , n11279 , n11280 );
not ( n60656 , n60401 );
nand ( n11283 , n11281 , n60656 );
not ( n60658 , n54619 );
not ( n60659 , n54648 );
or ( n11286 , n60658 , n60659 );
nand ( n60661 , n11286 , n60324 );
not ( n11288 , n60661 );
and ( n60663 , n11283 , n11288 );
not ( n60664 , n11283 );
and ( n11291 , n60664 , n60661 );
nor ( n60666 , n60663 , n11291 );
buf ( n60667 , n60666 );
xor ( n11294 , n60651 , n60667 );
buf ( n60669 , n11294 );
buf ( n60670 , n60669 );
buf ( n60671 , n60498 );
nand ( n60672 , n60670 , n60671 );
buf ( n60673 , n60672 );
buf ( n60674 , n60673 );
nand ( n60675 , n11276 , n60674 );
buf ( n60676 , n60675 );
buf ( n60677 , n60676 );
not ( n60678 , n10095 );
not ( n11305 , n60678 );
not ( n60680 , n59374 );
not ( n60681 , n60416 );
or ( n11308 , n60680 , n60681 );
or ( n60683 , n60416 , n59374 );
nand ( n60684 , n11308 , n60683 );
not ( n11311 , n60684 );
or ( n60686 , n11305 , n11311 );
nand ( n60687 , n10093 , n382 );
nand ( n60688 , n60686 , n60687 );
buf ( n60689 , n60688 );
xor ( n60690 , n60677 , n60689 );
buf ( n60691 , n10005 );
not ( n11318 , n60691 );
not ( n11319 , n380 );
not ( n11320 , n60464 );
or ( n11321 , n11319 , n11320 );
nand ( n11322 , n60461 , n59380 );
nand ( n11323 , n11321 , n11322 );
buf ( n60698 , n11323 );
not ( n11325 , n60698 );
or ( n11326 , n11318 , n11325 );
and ( n11327 , n10941 , n60413 );
xor ( n11328 , n11327 , n11032 );
and ( n11329 , n11328 , n59380 );
not ( n11330 , n11328 );
and ( n11331 , n11330 , n380 );
or ( n11332 , n11329 , n11331 );
not ( n11333 , n59384 );
nand ( n11334 , n11332 , n11333 );
buf ( n60709 , n11334 );
nand ( n11336 , n11326 , n60709 );
buf ( n60711 , n11336 );
buf ( n60712 , n60711 );
xor ( n11339 , n60690 , n60712 );
buf ( n60714 , n11339 );
buf ( n60715 , n60714 );
nor ( n11342 , n54710 , n54701 );
not ( n11343 , n54342 );
nand ( n11344 , n11343 , n10996 );
not ( n11345 , n11003 );
not ( n11346 , n11004 );
or ( n11347 , n11345 , n11346 );
nand ( n11348 , n11347 , n10992 );
nand ( n11349 , n11344 , n11348 );
nand ( n11350 , n11342 , n11349 );
not ( n11351 , n11349 );
not ( n11352 , n54703 );
not ( n11353 , n54347 );
nand ( n11354 , n11352 , n11353 );
and ( n11355 , n54701 , n11354 );
nand ( n11356 , n11351 , n11355 );
not ( n11357 , n54701 );
not ( n11358 , n11354 );
and ( n11359 , n11357 , n11358 );
not ( n11360 , n54682 );
nand ( n11361 , n11360 , n54707 );
and ( n11362 , n11361 , n54697 );
nor ( n11363 , n11359 , n11362 );
nand ( n11364 , n11350 , n11356 , n11363 );
and ( n60739 , n11364 , n378 );
not ( n11366 , n384 );
buf ( n60741 , n7417 );
buf ( n60742 , n60241 );
nand ( n11369 , n60741 , n60742 );
buf ( n60744 , n11369 );
not ( n60745 , n60744 );
not ( n11372 , n59290 );
or ( n60747 , n60745 , n11372 );
or ( n60748 , n60744 , n59290 );
nand ( n60749 , n60747 , n60748 );
buf ( n60750 , n60749 );
not ( n60751 , n60750 );
buf ( n60752 , n60751 );
not ( n11379 , n60752 );
or ( n11380 , n11366 , n11379 );
buf ( n60755 , n384 );
not ( n11382 , n60755 );
buf ( n60757 , n60749 );
nand ( n60758 , n11382 , n60757 );
buf ( n60759 , n60758 );
nand ( n60760 , n11380 , n60759 );
or ( n60761 , n60739 , n60760 );
nand ( n11388 , n11354 , n54707 );
xor ( n60763 , n11388 , n11011 );
buf ( n60764 , n60763 );
buf ( n60765 , n378 );
nand ( n60766 , n60764 , n60765 );
buf ( n60767 , n60766 );
buf ( n60768 , n60767 );
not ( n60769 , n60768 );
buf ( n60770 , n60769 );
buf ( n60771 , n9859 );
buf ( n11398 , n60771 );
buf ( n11399 , n11398 );
not ( n11400 , n11399 );
buf ( n60775 , n59255 );
not ( n11402 , n60775 );
buf ( n60777 , n11402 );
not ( n11404 , n60777 );
not ( n11405 , n9731 );
or ( n11406 , n11404 , n11405 );
buf ( n60781 , n59265 );
not ( n11408 , n60781 );
buf ( n60783 , n11408 );
nand ( n60784 , n11406 , n60783 );
not ( n11411 , n60784 );
or ( n60786 , n11400 , n11411 );
buf ( n60787 , n9909 );
buf ( n11414 , n60787 );
buf ( n60789 , n11414 );
nand ( n60790 , n60786 , n60789 );
not ( n11417 , n59273 );
nand ( n60792 , n11417 , n59285 );
not ( n60793 , n60792 );
and ( n11420 , n60790 , n60793 );
not ( n60795 , n60790 );
and ( n11422 , n60795 , n60792 );
nor ( n11423 , n11420 , n11422 );
or ( n60798 , n60770 , n11423 );
not ( n11425 , n60784 );
not ( n60800 , n11425 );
nand ( n11427 , n60789 , n11399 );
not ( n11428 , n11427 );
not ( n11429 , n11428 );
or ( n11430 , n60800 , n11429 );
nand ( n11431 , n60784 , n11427 );
nand ( n11432 , n11430 , n11431 );
not ( n60807 , n51459 );
not ( n60808 , n2467 );
not ( n11435 , n2449 );
nand ( n60810 , n11435 , n51268 );
nor ( n11437 , n60810 , n2477 );
nand ( n11438 , n60808 , n11437 );
buf ( n11439 , n11438 );
not ( n11440 , n11439 );
not ( n11441 , n52006 );
and ( n11442 , n52045 , n11441 , n1907 );
nand ( n11443 , n11440 , n11442 );
nor ( n11444 , n11443 , n2442 );
not ( n60819 , n11444 );
or ( n11446 , n60807 , n60819 );
not ( n60821 , n11443 );
not ( n11448 , n51748 );
not ( n11449 , n2563 );
or ( n11450 , n11448 , n11449 );
and ( n11451 , n2673 , n51981 );
nor ( n11452 , n11451 , n51832 );
nand ( n11453 , n11450 , n11452 );
and ( n11454 , n60821 , n11453 );
not ( n11455 , n11442 );
not ( n11456 , n52029 );
or ( n60831 , n11455 , n11456 );
nand ( n11458 , n60831 , n52036 );
nor ( n11459 , n11454 , n11458 );
nand ( n11460 , n11446 , n11459 );
nand ( n11461 , n11432 , n11460 );
buf ( n60836 , n11461 );
not ( n60837 , n60836 );
buf ( n60838 , n60837 );
nand ( n11465 , n60798 , n60838 );
nand ( n60840 , n60770 , n11423 );
nand ( n60841 , n11465 , n60840 );
nand ( n11468 , n60761 , n60841 );
buf ( n60843 , n11468 );
nand ( n60844 , n60760 , n60739 );
buf ( n60845 , n60844 );
nand ( n11472 , n60843 , n60845 );
buf ( n11473 , n11472 );
buf ( n11474 , n60749 );
buf ( n60849 , n11474 );
buf ( n60850 , n60849 );
nand ( n60851 , n60850 , n384 );
nand ( n60852 , n54871 , n11256 );
not ( n11479 , n60852 );
not ( n60854 , n11348 );
not ( n11481 , n11265 );
or ( n11482 , n60854 , n11481 );
buf ( n11483 , n11017 );
not ( n11484 , n54714 );
buf ( n11485 , n54679 );
nor ( n11486 , n11484 , n11485 );
nor ( n11487 , n11483 , n11486 );
nand ( n11488 , n11482 , n11487 );
not ( n11489 , n11488 );
not ( n11490 , n11489 );
or ( n60865 , n11479 , n11490 );
not ( n11492 , n60852 );
nand ( n60867 , n11492 , n11488 );
nand ( n11494 , n60865 , n60867 );
not ( n11495 , n11494 );
nand ( n60870 , n11495 , n378 );
and ( n60871 , n60851 , n60870 );
not ( n11498 , n60851 );
buf ( n60873 , n60870 );
not ( n11500 , n60873 );
buf ( n60875 , n11500 );
and ( n60876 , n11498 , n60875 );
nor ( n11503 , n60871 , n60876 );
buf ( n60878 , n56869 );
buf ( n11505 , n60878 );
buf ( n11506 , n11505 );
buf ( n60881 , n11506 );
buf ( n60882 , n56860 );
nand ( n11509 , n60881 , n60882 );
buf ( n60884 , n11509 );
and ( n11511 , n60884 , n384 );
not ( n11512 , n60884 );
and ( n11513 , n11512 , n59460 );
or ( n11514 , n11511 , n11513 );
buf ( n60889 , n59290 );
buf ( n60890 , n60241 );
and ( n11517 , n60889 , n60890 );
buf ( n60892 , n11517 );
buf ( n60893 , n60892 );
not ( n60894 , n60893 );
buf ( n60895 , n7417 );
nand ( n60896 , n60894 , n60895 );
buf ( n60897 , n60896 );
xor ( n11524 , n11514 , n60897 );
buf ( n11525 , n11524 );
and ( n11526 , n11503 , n11525 );
not ( n11527 , n11503 );
not ( n11528 , n11524 );
and ( n11529 , n11527 , n11528 );
nor ( n11530 , n11526 , n11529 );
xor ( n11531 , n11473 , n11530 );
buf ( n60906 , n60498 );
not ( n11533 , n60906 );
buf ( n11534 , n60647 );
not ( n11535 , n11534 );
or ( n11536 , n11533 , n11535 );
not ( n11537 , n378 );
not ( n11538 , n11494 );
or ( n11539 , n11537 , n11538 );
not ( n11540 , n11488 );
nand ( n11541 , n11540 , n60852 );
nand ( n60916 , n11541 , n60867 , n11105 );
nand ( n60917 , n11539 , n60916 );
buf ( n60918 , n60917 );
buf ( n60919 , n60476 );
nand ( n60920 , n60918 , n60919 );
buf ( n60921 , n60920 );
buf ( n60922 , n60921 );
nand ( n60923 , n11536 , n60922 );
buf ( n60924 , n60923 );
buf ( n60925 , n60924 );
not ( n60926 , n10005 );
not ( n11553 , n11332 );
or ( n60928 , n60926 , n11553 );
not ( n11555 , n59380 );
and ( n60930 , n11288 , n11555 );
not ( n60931 , n11288 );
not ( n11558 , n380 );
and ( n60933 , n60931 , n11558 );
or ( n11560 , n60930 , n60933 );
and ( n11561 , n11283 , n11560 );
not ( n11562 , n11283 );
not ( n11563 , n59380 );
and ( n11564 , n60661 , n11563 );
not ( n11565 , n60661 );
not ( n60940 , n380 );
and ( n60941 , n11565 , n60940 );
or ( n11568 , n11564 , n60941 );
and ( n60943 , n11562 , n11568 );
or ( n11570 , n11561 , n60943 );
buf ( n60945 , n11570 );
buf ( n60946 , n11333 );
nand ( n60947 , n60945 , n60946 );
buf ( n60948 , n60947 );
nand ( n60949 , n60928 , n60948 );
buf ( n60950 , n60949 );
xor ( n11577 , n60925 , n60950 );
not ( n11578 , n60678 );
buf ( n60953 , n382 );
not ( n60954 , n60953 );
buf ( n60955 , n60464 );
not ( n11582 , n60955 );
or ( n60957 , n60954 , n11582 );
nand ( n60958 , n60461 , n59374 );
buf ( n60959 , n60958 );
nand ( n60960 , n60957 , n60959 );
buf ( n60961 , n60960 );
not ( n60962 , n60961 );
or ( n60963 , n11578 , n60962 );
not ( n11590 , n10094 );
nand ( n60965 , n11590 , n60684 );
nand ( n60966 , n60963 , n60965 );
buf ( n60967 , n60966 );
and ( n11594 , n11577 , n60967 );
and ( n60969 , n60925 , n60950 );
or ( n11596 , n11594 , n60969 );
buf ( n60971 , n11596 );
xor ( n60972 , n11531 , n60971 );
buf ( n60973 , n60972 );
xor ( n11600 , n60715 , n60973 );
not ( n11601 , n10005 );
not ( n11602 , n11570 );
or ( n11603 , n11601 , n11602 );
not ( n11604 , n380 );
not ( n60979 , n60644 );
not ( n11606 , n60979 );
or ( n60981 , n11604 , n11606 );
nand ( n11608 , n60644 , n59380 );
nand ( n11609 , n60981 , n11608 );
nand ( n11610 , n11609 , n11333 );
nand ( n11611 , n11603 , n11610 );
not ( n11612 , n10093 );
buf ( n60987 , n382 );
not ( n11614 , n60987 );
buf ( n60989 , n60464 );
not ( n11616 , n60989 );
or ( n11617 , n11614 , n11616 );
buf ( n60992 , n60958 );
nand ( n11619 , n11617 , n60992 );
buf ( n60994 , n11619 );
not ( n11621 , n60994 );
or ( n11622 , n11612 , n11621 );
not ( n11623 , n59374 );
not ( n11624 , n11328 );
or ( n11625 , n11623 , n11624 );
or ( n11626 , n11328 , n59374 );
nand ( n61001 , n11625 , n11626 );
nand ( n11628 , n61001 , n60678 );
nand ( n61003 , n11622 , n11628 );
xor ( n61004 , n11611 , n61003 );
buf ( n61005 , n385 );
not ( n61006 , n61005 );
buf ( n61007 , n61006 );
and ( n11634 , n61007 , n384 );
not ( n61009 , n11634 );
and ( n11636 , n384 , n60487 );
not ( n61011 , n384 );
and ( n11638 , n61011 , n60416 );
or ( n11639 , n11636 , n11638 );
not ( n61014 , n11639 );
or ( n11641 , n61009 , n61014 );
buf ( n61016 , n384 );
buf ( n61017 , n385 );
nand ( n11644 , n61016 , n61017 );
buf ( n61019 , n11644 );
nand ( n61020 , n11641 , n61019 );
and ( n61021 , n61004 , n61020 );
and ( n11648 , n11611 , n61003 );
or ( n61023 , n61021 , n11648 );
not ( n61024 , n61023 );
nand ( n11651 , n11344 , n54679 );
not ( n61026 , n11651 );
not ( n61027 , n61026 );
not ( n11654 , n11348 );
not ( n61029 , n11654 );
or ( n61030 , n61027 , n61029 );
or ( n11657 , n11654 , n61026 );
nand ( n61032 , n61030 , n11657 );
and ( n11659 , n61032 , n378 );
not ( n11660 , n11659 );
nand ( n61035 , n52045 , n11441 );
nor ( n11662 , n11439 , n61035 );
not ( n61037 , n11662 );
not ( n11664 , n11453 );
or ( n61039 , n61037 , n11664 );
not ( n61040 , n51747 );
and ( n11667 , n51933 , n51935 );
not ( n61042 , n2709 );
not ( n11669 , n51268 );
or ( n11670 , n61042 , n11669 );
and ( n11671 , n52014 , n1971 );
nand ( n11672 , n11670 , n11671 );
nor ( n11673 , n11667 , n11672 );
not ( n11674 , n11673 );
or ( n11675 , n61040 , n11674 );
not ( n11676 , n52030 );
nand ( n11677 , n11676 , n61035 );
nand ( n11678 , n11675 , n11677 );
not ( n11679 , n11678 );
not ( n11680 , n51321 );
not ( n11681 , n11680 );
nand ( n11682 , n51409 , n2153 );
not ( n11683 , n11682 );
and ( n11684 , n11681 , n11683 );
buf ( n11685 , n2497 );
buf ( n11686 , n51935 );
and ( n11687 , n11685 , n11686 );
nor ( n61062 , n11684 , n11687 );
nor ( n11689 , n51333 , n11672 );
nand ( n61064 , n61062 , n11689 , n51410 );
not ( n11691 , n52018 );
nand ( n11692 , n11691 , n11438 , n2629 );
nand ( n11693 , n11679 , n61064 , n11692 , n2717 );
nand ( n11694 , n61039 , n11693 );
not ( n11695 , n1907 );
nor ( n11696 , n11695 , n51211 );
buf ( n11697 , n11696 );
and ( n11698 , n11694 , n11697 );
not ( n11699 , n11694 );
not ( n11700 , n11696 );
and ( n11701 , n11699 , n11700 );
nor ( n11702 , n11698 , n11701 );
buf ( n61077 , n9731 );
buf ( n11704 , n61077 );
buf ( n61079 , n11704 );
buf ( n61080 , n59255 );
not ( n11707 , n61080 );
buf ( n61082 , n60783 );
nand ( n11709 , n11707 , n61082 );
buf ( n61084 , n11709 );
not ( n11711 , n61084 );
and ( n61086 , n61079 , n11711 );
not ( n11713 , n61079 );
and ( n61088 , n11713 , n61084 );
nor ( n11715 , n61086 , n61088 );
nand ( n11716 , n11702 , n11715 );
not ( n61091 , n11716 );
not ( n61092 , n61091 );
or ( n11719 , n11660 , n61092 );
not ( n61094 , n11659 );
not ( n11721 , n61094 );
not ( n61096 , n11716 );
or ( n11723 , n11721 , n61096 );
not ( n61098 , n11460 );
not ( n11725 , n61098 );
not ( n11726 , n11432 );
or ( n11727 , n11725 , n11726 );
not ( n11728 , n11432 );
nand ( n61103 , n11728 , n11460 );
nand ( n11730 , n11727 , n61103 );
nand ( n11731 , n11723 , n11730 );
nand ( n61106 , n11719 , n11731 );
not ( n61107 , n61106 );
not ( n11734 , n61107 );
not ( n61109 , n60767 );
not ( n61110 , n11461 );
or ( n11737 , n61109 , n61110 );
nand ( n61112 , n60838 , n60770 );
nand ( n11739 , n11737 , n61112 );
and ( n61114 , n11739 , n11423 );
not ( n11741 , n11739 );
not ( n61116 , n11423 );
and ( n11743 , n11741 , n61116 );
nor ( n11744 , n61114 , n11743 );
not ( n11745 , n11744 );
or ( n11746 , n11734 , n11745 );
nand ( n11747 , n60917 , n60498 );
nand ( n11748 , n11356 , n11350 , n11363 );
not ( n11749 , n11748 );
and ( n11750 , n11749 , n11105 );
not ( n61125 , n11749 );
and ( n61126 , n61125 , n378 );
nor ( n11753 , n11750 , n61126 );
nand ( n61128 , n11753 , n60476 );
nand ( n61129 , n11747 , n61128 );
nand ( n11756 , n11746 , n61129 );
not ( n61131 , n61107 );
not ( n61132 , n11744 );
nand ( n11759 , n61131 , n61132 );
nand ( n61134 , n11756 , n11759 );
buf ( n61135 , n61134 );
not ( n11762 , n61135 );
xor ( n11763 , n60739 , n60760 );
xnor ( n11764 , n11763 , n60841 );
buf ( n61139 , n11764 );
nand ( n11766 , n11762 , n61139 );
buf ( n61141 , n11766 );
not ( n11768 , n61141 );
or ( n11769 , n61024 , n11768 );
not ( n11770 , n11764 );
nand ( n11771 , n11770 , n61134 );
nand ( n61146 , n11769 , n11771 );
buf ( n61147 , n61146 );
xor ( n11774 , n11600 , n61147 );
buf ( n61149 , n11774 );
buf ( n61150 , n61149 );
xor ( n11777 , n60925 , n60950 );
xor ( n61152 , n11777 , n60967 );
buf ( n61153 , n61152 );
buf ( n11780 , n61153 );
nand ( n61155 , n11753 , n60498 );
buf ( n61156 , n60763 );
not ( n61157 , n61156 );
buf ( n61158 , n61157 );
and ( n61159 , n11105 , n61158 );
not ( n11786 , n11105 );
buf ( n61161 , n60763 );
buf ( n11788 , n61161 );
buf ( n61163 , n11788 );
and ( n11790 , n11786 , n61163 );
nor ( n11791 , n61159 , n11790 );
nand ( n11792 , n11791 , n60476 );
nand ( n11793 , n61155 , n11792 );
buf ( n61168 , n11793 );
not ( n11795 , n61168 );
not ( n11796 , n10005 );
not ( n11797 , n11609 );
or ( n11798 , n11796 , n11797 );
xor ( n61173 , n380 , n60852 );
buf ( n11800 , n11488 );
xnor ( n61175 , n61173 , n11800 );
nand ( n11802 , n11333 , n61175 );
nand ( n61177 , n11798 , n11802 );
buf ( n61178 , n61177 );
not ( n11805 , n61178 );
or ( n61180 , n11795 , n11805 );
or ( n11807 , n61177 , n11793 );
buf ( n61182 , n9710 );
not ( n11809 , n61182 );
buf ( n61184 , n11809 );
buf ( n61185 , n61184 );
not ( n61186 , n61185 );
buf ( n61187 , n8844 );
buf ( n61188 , n58421 );
nor ( n11815 , n61187 , n61188 );
buf ( n61190 , n11815 );
not ( n11817 , n61190 );
nand ( n11818 , n11817 , n9088 );
buf ( n11819 , n11818 );
not ( n11820 , n11819 );
or ( n11821 , n61186 , n11820 );
buf ( n61196 , n61184 );
buf ( n61197 , n11818 );
or ( n11824 , n61196 , n61197 );
nand ( n61199 , n11821 , n11824 );
buf ( n61200 , n61199 );
buf ( n61201 , n61200 );
not ( n61202 , n61201 );
not ( n11829 , n58970 );
not ( n11830 , n9669 );
or ( n61205 , n11829 , n11830 );
nand ( n61206 , n61205 , n59041 );
not ( n61207 , n61206 );
buf ( n61208 , n59065 );
not ( n11835 , n61208 );
buf ( n61210 , n59060 );
nand ( n11837 , n11835 , n61210 );
buf ( n61212 , n11837 );
nand ( n61213 , n61207 , n59068 , n61212 );
not ( n61214 , n61213 );
not ( n11841 , n59068 );
not ( n61216 , n61212 );
or ( n11843 , n11841 , n61216 );
nand ( n11844 , n11843 , n61206 );
not ( n11845 , n11844 );
or ( n11846 , n61214 , n11845 );
nand ( n11847 , n10972 , n10955 );
not ( n11848 , n11847 );
not ( n61223 , n10976 );
not ( n11850 , n53725 );
not ( n61225 , n11850 );
or ( n61226 , n61223 , n61225 );
nand ( n61227 , n61226 , n10983 );
not ( n11854 , n61227 );
not ( n61229 , n11854 );
or ( n11856 , n11848 , n61229 );
not ( n11857 , n11847 );
nand ( n61232 , n11857 , n61227 );
nand ( n61233 , n11856 , n61232 );
not ( n11860 , n61233 );
not ( n11861 , n11860 );
nor ( n61236 , n11861 , n11105 );
nand ( n61237 , n11846 , n61236 );
buf ( n61238 , n61237 );
nor ( n61239 , n61202 , n61238 );
buf ( n61240 , n61239 );
buf ( n61241 , n61240 );
buf ( n11868 , n9088 );
and ( n11869 , n61184 , n11868 );
buf ( n61244 , n61190 );
nor ( n11871 , n11869 , n61244 );
not ( n61246 , n11871 );
buf ( n61247 , n59081 );
not ( n61248 , n61247 );
buf ( n61249 , n59092 );
nor ( n11876 , n61248 , n61249 );
buf ( n61251 , n11876 );
not ( n61252 , n61251 );
or ( n61253 , n61246 , n61252 );
or ( n11880 , n61251 , n11871 );
nand ( n61255 , n61253 , n11880 );
buf ( n61256 , n61255 );
and ( n11883 , n61241 , n61256 );
buf ( n61258 , n11883 );
not ( n61259 , n61258 );
buf ( n61260 , n378 );
not ( n11887 , n10986 );
and ( n61262 , n54740 , n54737 );
nor ( n61263 , n61262 , n10987 );
not ( n11890 , n61263 );
or ( n61265 , n11887 , n11890 );
buf ( n61266 , n11002 );
nand ( n11893 , n61265 , n61266 );
not ( n11894 , n4782 );
not ( n11895 , n54225 );
or ( n61270 , n11894 , n11895 );
nand ( n61271 , n61270 , n11004 );
not ( n11898 , n61271 );
and ( n61273 , n11893 , n11898 );
not ( n11900 , n11893 );
and ( n11901 , n11900 , n61271 );
nor ( n11902 , n61273 , n11901 );
buf ( n61277 , n11902 );
and ( n11904 , n61260 , n61277 );
buf ( n61279 , n11904 );
not ( n11906 , n61279 );
nand ( n11907 , n61259 , n11906 );
not ( n11908 , n11907 );
not ( n11909 , n60476 );
nand ( n11910 , n11651 , n11348 );
nand ( n11911 , n61026 , n11654 );
nand ( n11912 , n11910 , n11911 );
and ( n61287 , n11105 , n11912 );
not ( n11914 , n11105 );
not ( n61289 , n61032 );
and ( n11916 , n11914 , n61289 );
or ( n11917 , n61287 , n11916 );
not ( n61292 , n11917 );
or ( n11919 , n11909 , n61292 );
and ( n61294 , n60763 , n60498 , n11105 );
or ( n11921 , n59415 , n11105 );
nor ( n11922 , n61163 , n11921 );
nor ( n61297 , n61294 , n11922 );
nand ( n61298 , n11919 , n61297 );
not ( n11925 , n61298 );
or ( n61300 , n11908 , n11925 );
not ( n11927 , n61259 );
nand ( n61302 , n11927 , n61279 );
nand ( n61303 , n61300 , n61302 );
nand ( n11930 , n11807 , n61303 );
buf ( n61305 , n11930 );
nand ( n61306 , n61180 , n61305 );
buf ( n61307 , n61306 );
buf ( n61308 , n61307 );
not ( n61309 , n60498 );
not ( n11936 , n60917 );
or ( n61311 , n61309 , n11936 );
nand ( n61312 , n61311 , n61128 );
xor ( n11939 , n61106 , n61312 );
and ( n11940 , n11939 , n61132 );
not ( n11941 , n11939 );
and ( n11942 , n11941 , n11744 );
nor ( n11943 , n11940 , n11942 );
buf ( n61318 , n11943 );
xor ( n11945 , n61308 , n61318 );
xor ( n11946 , n11659 , n11716 );
xnor ( n61321 , n11946 , n11730 );
buf ( n61322 , n61321 );
not ( n11949 , n10093 );
not ( n61324 , n61001 );
or ( n61325 , n11949 , n61324 );
not ( n11952 , n382 );
buf ( n61327 , n60666 );
not ( n61328 , n61327 );
buf ( n61329 , n61328 );
not ( n61330 , n61329 );
or ( n61331 , n11952 , n61330 );
not ( n11958 , n382 );
nand ( n11959 , n11958 , n60666 );
nand ( n61334 , n61331 , n11959 );
nand ( n61335 , n61334 , n60678 );
nand ( n11962 , n61325 , n61335 );
buf ( n61337 , n11962 );
xor ( n11964 , n61322 , n61337 );
not ( n11965 , n11333 );
and ( n61340 , n11356 , n11350 , n11363 );
not ( n11967 , n61340 );
and ( n61342 , n380 , n11967 );
not ( n61343 , n380 );
and ( n11970 , n61343 , n61340 );
nor ( n61345 , n61342 , n11970 );
not ( n11972 , n61345 );
or ( n61347 , n11965 , n11972 );
nand ( n11974 , n61175 , n10005 );
nand ( n61349 , n61347 , n11974 );
not ( n61350 , n61349 );
not ( n11977 , n10985 );
not ( n61352 , n60352 );
or ( n11979 , n11977 , n61352 );
nand ( n11980 , n54740 , n54737 );
nand ( n61355 , n11979 , n11980 );
not ( n11982 , n53950 );
not ( n61357 , n11982 );
not ( n11984 , n4777 );
not ( n61359 , n11984 );
or ( n61360 , n61357 , n61359 );
nand ( n11987 , n61360 , n11002 );
and ( n61362 , n61355 , n11987 );
not ( n61363 , n61355 );
not ( n11990 , n11987 );
and ( n61365 , n61363 , n11990 );
nor ( n61366 , n61362 , n61365 );
buf ( n61367 , n61366 );
buf ( n61368 , n61367 );
buf ( n61369 , n61368 );
buf ( n61370 , n61369 );
buf ( n61371 , n378 );
nand ( n61372 , n61370 , n61371 );
buf ( n61373 , n61372 );
not ( n61374 , n61373 );
not ( n61375 , n52006 );
nand ( n12002 , n61375 , n52012 );
nor ( n12003 , n11439 , n52048 );
not ( n12004 , n12003 );
not ( n12005 , n51748 );
not ( n12006 , n2563 );
or ( n12007 , n12005 , n12006 );
nand ( n61382 , n12007 , n11452 );
not ( n12009 , n61382 );
or ( n61384 , n12004 , n12009 );
not ( n12011 , n51748 );
not ( n61386 , n11438 );
not ( n12013 , n61386 );
or ( n61388 , n12011 , n12013 );
not ( n12015 , n52052 );
not ( n61390 , n52061 );
or ( n12017 , n12015 , n61390 );
and ( n61392 , n52052 , n51800 , n51811 );
nand ( n12019 , n51803 , n61392 );
nand ( n12020 , n12017 , n12019 );
nand ( n12021 , n61388 , n12020 );
and ( n12022 , n12020 , n2613 );
nor ( n12023 , n12022 , n52048 );
nand ( n12024 , n12021 , n51970 , n12023 );
nand ( n12025 , n61384 , n12024 );
xor ( n12026 , n12002 , n12025 );
not ( n12027 , n12026 );
or ( n12028 , n61374 , n12027 );
xor ( n12029 , n61241 , n61256 );
buf ( n61404 , n12029 );
nand ( n61405 , n12028 , n61404 );
not ( n12032 , n12026 );
not ( n61407 , n61373 );
nand ( n12034 , n12032 , n61407 );
nand ( n61409 , n61405 , n12034 );
not ( n12036 , n61409 );
not ( n12037 , n11715 );
not ( n61412 , n11702 );
or ( n61413 , n12037 , n61412 );
not ( n12040 , n11715 );
nand ( n61415 , n12040 , n61412 );
nand ( n61416 , n61413 , n61415 );
nand ( n12043 , n12036 , n61416 );
not ( n61418 , n12043 );
or ( n61419 , n61350 , n61418 );
not ( n12046 , n61416 );
nand ( n12047 , n61409 , n12046 );
nand ( n61422 , n61419 , n12047 );
buf ( n61423 , n61422 );
and ( n12050 , n11964 , n61423 );
and ( n61425 , n61322 , n61337 );
or ( n61426 , n12050 , n61425 );
buf ( n61427 , n61426 );
buf ( n61428 , n61427 );
and ( n61429 , n11945 , n61428 );
and ( n12056 , n61308 , n61318 );
or ( n61431 , n61429 , n12056 );
buf ( n61432 , n61431 );
buf ( n61433 , n61432 );
xor ( n12060 , n11780 , n61433 );
buf ( n12061 , n11764 );
and ( n12062 , n61134 , n12061 );
not ( n61437 , n61134 );
not ( n12064 , n11764 );
and ( n12065 , n61437 , n12064 );
nor ( n12066 , n12062 , n12065 );
not ( n61441 , n61023 );
and ( n61442 , n12066 , n61441 );
not ( n12069 , n12066 );
and ( n61444 , n12069 , n61023 );
nor ( n61445 , n61442 , n61444 );
buf ( n61446 , n61445 );
and ( n61447 , n12060 , n61446 );
and ( n61448 , n11780 , n61433 );
or ( n12075 , n61447 , n61448 );
buf ( n61450 , n12075 );
buf ( n61451 , n61450 );
nor ( n12078 , n61150 , n61451 );
buf ( n61453 , n12078 );
buf ( n61454 , n61453 );
not ( n61455 , n61454 );
buf ( n61456 , n61455 );
xor ( n12083 , n60715 , n60973 );
and ( n12084 , n12083 , n61147 );
and ( n12085 , n60715 , n60973 );
or ( n12086 , n12084 , n12085 );
buf ( n61461 , n12086 );
not ( n12088 , n61461 );
and ( n12089 , n60621 , n60645 );
buf ( n61464 , n12089 );
buf ( n61465 , n61464 );
buf ( n61466 , n60498 );
not ( n61467 , n61466 );
and ( n12094 , n11328 , n11105 );
not ( n12095 , n11328 );
and ( n12096 , n12095 , n378 );
or ( n12097 , n12094 , n12096 );
buf ( n61472 , n12097 );
not ( n12099 , n61472 );
or ( n12100 , n61467 , n12099 );
buf ( n61475 , n60669 );
buf ( n61476 , n60476 );
nand ( n12103 , n61475 , n61476 );
buf ( n61478 , n12103 );
buf ( n61479 , n61478 );
nand ( n61480 , n12100 , n61479 );
buf ( n61481 , n61480 );
buf ( n61482 , n61481 );
xor ( n61483 , n61465 , n61482 );
not ( n12110 , n11333 );
not ( n61485 , n11323 );
or ( n12112 , n12110 , n61485 );
not ( n12113 , n380 );
not ( n12114 , n60487 );
or ( n12115 , n12113 , n12114 );
nand ( n12116 , n60416 , n59380 );
nand ( n12117 , n12115 , n12116 );
nand ( n12118 , n12117 , n10005 );
nand ( n12119 , n12112 , n12118 );
buf ( n61494 , n12119 );
xor ( n12121 , n61483 , n61494 );
buf ( n61496 , n12121 );
buf ( n61497 , n61496 );
xor ( n12124 , n11473 , n11530 );
and ( n12125 , n12124 , n60971 );
and ( n61500 , n11473 , n11530 );
or ( n12127 , n12125 , n61500 );
buf ( n61502 , n12127 );
xor ( n12129 , n61497 , n61502 );
buf ( n61504 , n60851 );
buf ( n61505 , n60870 );
nand ( n12132 , n61504 , n61505 );
buf ( n61507 , n12132 );
buf ( n61508 , n61507 );
not ( n61509 , n61508 );
buf ( n61510 , n11524 );
not ( n12137 , n61510 );
or ( n61512 , n61509 , n12137 );
not ( n61513 , n60851 );
nand ( n12140 , n61513 , n60875 );
buf ( n61515 , n12140 );
nand ( n61516 , n61512 , n61515 );
buf ( n61517 , n61516 );
buf ( n61518 , n57054 );
not ( n12145 , n61518 );
buf ( n61520 , n12145 );
buf ( n12147 , n57045 );
nand ( n12148 , n61520 , n12147 );
not ( n12149 , n12148 );
not ( n12150 , n11506 );
not ( n12151 , n60892 );
or ( n12152 , n12150 , n12151 );
nand ( n12153 , n12152 , n56870 );
not ( n12154 , n12153 );
not ( n12155 , n12154 );
or ( n12156 , n12149 , n12155 );
not ( n12157 , n12148 );
nand ( n12158 , n12157 , n12153 );
nand ( n12159 , n12156 , n12158 );
xor ( n12160 , n10831 , n12159 );
not ( n12161 , n60884 );
not ( n12162 , n60897 );
or ( n12163 , n12161 , n12162 );
or ( n61538 , n60897 , n60884 );
nand ( n12165 , n12163 , n61538 );
buf ( n61540 , n12165 );
buf ( n61541 , n384 );
nand ( n61542 , n61540 , n61541 );
buf ( n61543 , n61542 );
xor ( n61544 , n12160 , n61543 );
xor ( n12171 , n61517 , n61544 );
xor ( n61546 , n60677 , n60689 );
and ( n12173 , n61546 , n60712 );
and ( n12174 , n60677 , n60689 );
or ( n61549 , n12173 , n12174 );
buf ( n61550 , n61549 );
xnor ( n61551 , n12171 , n61550 );
buf ( n61552 , n61551 );
xor ( n61553 , n12129 , n61552 );
buf ( n61554 , n61553 );
not ( n12181 , n61554 );
nand ( n12182 , n12088 , n12181 );
xor ( n61557 , n11611 , n61003 );
xor ( n12184 , n61557 , n61020 );
xor ( n61559 , n61308 , n61318 );
xor ( n61560 , n61559 , n61428 );
buf ( n61561 , n61560 );
xor ( n12188 , n12184 , n61561 );
buf ( n61563 , n385 );
not ( n61564 , n61563 );
buf ( n61565 , n11639 );
not ( n61566 , n61565 );
or ( n61567 , n61564 , n61566 );
not ( n61568 , n384 );
not ( n12195 , n60464 );
or ( n61570 , n61568 , n12195 );
buf ( n61571 , n384 );
not ( n12198 , n61571 );
buf ( n61573 , n60461 );
nand ( n61574 , n12198 , n61573 );
buf ( n61575 , n61574 );
nand ( n12202 , n61570 , n61575 );
nand ( n61577 , n12202 , n11634 );
buf ( n61578 , n61577 );
nand ( n61579 , n61567 , n61578 );
buf ( n61580 , n61579 );
nand ( n12207 , n61155 , n11792 );
buf ( n61582 , n12207 );
buf ( n61583 , n61303 );
xor ( n61584 , n61582 , n61583 );
buf ( n61585 , n61177 );
xor ( n12212 , n61584 , n61585 );
buf ( n61587 , n12212 );
xor ( n61588 , n61580 , n61587 );
xor ( n12215 , n61322 , n61337 );
xor ( n61590 , n12215 , n61423 );
buf ( n61591 , n61590 );
and ( n61592 , n61588 , n61591 );
and ( n12219 , n61580 , n61587 );
or ( n61594 , n61592 , n12219 );
and ( n61595 , n12188 , n61594 );
and ( n12222 , n12184 , n61561 );
or ( n61597 , n61595 , n12222 );
not ( n12224 , n61597 );
buf ( n61599 , n12224 );
buf ( n61600 , n61153 );
buf ( n61601 , n61432 );
xor ( n12228 , n61600 , n61601 );
buf ( n61603 , n61445 );
xnor ( n12230 , n12228 , n61603 );
buf ( n61605 , n12230 );
buf ( n61606 , n61605 );
nand ( n12233 , n61599 , n61606 );
buf ( n61608 , n12233 );
xor ( n12235 , n12184 , n61561 );
xor ( n12236 , n12235 , n61594 );
buf ( n61611 , n12236 );
not ( n12238 , n61611 );
buf ( n61613 , n12238 );
buf ( n61614 , n61613 );
buf ( n61615 , n385 );
not ( n12242 , n61615 );
buf ( n61617 , n12202 );
not ( n12244 , n61617 );
or ( n61619 , n12242 , n12244 );
not ( n12246 , n59460 );
not ( n61621 , n11328 );
or ( n12248 , n12246 , n61621 );
or ( n12249 , n11328 , n59460 );
nand ( n12250 , n12248 , n12249 );
buf ( n61625 , n12250 );
buf ( n61626 , n11634 );
nand ( n12253 , n61625 , n61626 );
buf ( n61628 , n12253 );
buf ( n61629 , n61628 );
nand ( n61630 , n61619 , n61629 );
buf ( n61631 , n61630 );
not ( n12258 , n61631 );
not ( n61633 , n12036 );
not ( n12260 , n12046 );
or ( n12261 , n61633 , n12260 );
nand ( n12262 , n61409 , n61416 );
nand ( n61637 , n12261 , n12262 );
and ( n61638 , n61637 , n61349 );
not ( n12265 , n61637 );
not ( n61640 , n61349 );
and ( n12267 , n12265 , n61640 );
nor ( n61642 , n61638 , n12267 );
not ( n12269 , n61642 );
or ( n12270 , n12258 , n12269 );
buf ( n61645 , n61631 );
not ( n12272 , n61645 );
buf ( n61647 , n12272 );
not ( n12274 , n61647 );
and ( n12275 , n61637 , n61640 );
not ( n12276 , n61637 );
and ( n12277 , n12276 , n61349 );
nor ( n61652 , n12275 , n12277 );
not ( n12279 , n61652 );
or ( n61654 , n12274 , n12279 );
not ( n61655 , n10005 );
not ( n12282 , n61345 );
or ( n61657 , n61655 , n12282 );
and ( n61658 , n380 , n60763 );
not ( n12285 , n380 );
and ( n61660 , n12285 , n61158 );
nor ( n12287 , n61658 , n61660 );
nand ( n12288 , n12287 , n11333 );
nand ( n61663 , n61657 , n12288 );
buf ( n61664 , n61663 );
not ( n12291 , n61664 );
buf ( n61666 , n12291 );
buf ( n61667 , n61666 );
not ( n61668 , n61667 );
not ( n61669 , n10093 );
buf ( n61670 , n382 );
buf ( n61671 , n60644 );
xor ( n12298 , n61670 , n61671 );
buf ( n61673 , n12298 );
not ( n12300 , n61673 );
or ( n12301 , n61669 , n12300 );
not ( n12302 , n382 );
nand ( n12303 , n12302 , n11494 );
not ( n12304 , n11494 );
nand ( n12305 , n12304 , n382 );
nand ( n12306 , n12303 , n12305 , n60678 );
nand ( n12307 , n12301 , n12306 );
not ( n12308 , n12307 );
buf ( n61683 , n12308 );
not ( n12310 , n61683 );
or ( n12311 , n61668 , n12310 );
buf ( n61686 , n60498 );
not ( n12313 , n61686 );
xor ( n61688 , n61260 , n61277 );
buf ( n61689 , n61688 );
buf ( n61690 , n61689 );
not ( n12317 , n61690 );
or ( n12318 , n12313 , n12317 );
and ( n12319 , n61366 , n11105 );
not ( n61694 , n61366 );
and ( n61695 , n61694 , n378 );
or ( n12322 , n12319 , n61695 );
buf ( n61697 , n12322 );
buf ( n61698 , n60476 );
nand ( n12325 , n61697 , n61698 );
buf ( n61700 , n12325 );
buf ( n61701 , n61700 );
nand ( n12328 , n12318 , n61701 );
buf ( n61703 , n12328 );
buf ( n61704 , n61227 );
not ( n12331 , n61704 );
buf ( n61706 , n59380 );
buf ( n61707 , n59401 );
nand ( n12334 , n61706 , n61707 );
buf ( n12335 , n12334 );
not ( n12336 , n12335 );
buf ( n12337 , n11847 );
nor ( n12338 , n12336 , n12337 );
nand ( n12339 , n12331 , n12338 );
nand ( n12340 , n61704 , n12337 , n12335 );
buf ( n61715 , n379 );
buf ( n61716 , n380 );
and ( n12343 , n61715 , n61716 );
buf ( n61718 , n11105 );
nor ( n12345 , n12343 , n61718 );
buf ( n61720 , n12345 );
nand ( n12347 , n12339 , n12340 , n61720 );
not ( n61722 , n12347 );
not ( n12349 , n61722 );
not ( n12350 , n395 );
not ( n12351 , n9268 );
not ( n61726 , n58968 );
or ( n61727 , n12351 , n61726 );
nand ( n12354 , n61727 , n58669 );
buf ( n12355 , n58965 );
xnor ( n12356 , n12354 , n12355 );
not ( n61731 , n12356 );
or ( n61732 , n12350 , n61731 );
buf ( n61733 , n12356 );
buf ( n61734 , n395 );
nor ( n61735 , n61733 , n61734 );
buf ( n61736 , n61735 );
not ( n12363 , n61736 );
nand ( n12364 , n12363 , n11860 , n60498 );
nand ( n61739 , n61732 , n12364 );
not ( n61740 , n61739 );
or ( n12367 , n12349 , n61740 );
not ( n12368 , n12347 );
not ( n12369 , n61739 );
not ( n12370 , n12369 );
or ( n12371 , n12368 , n12370 );
not ( n12372 , n394 );
buf ( n61747 , n58970 );
buf ( n61748 , n61747 );
buf ( n61749 , n61748 );
buf ( n61750 , n59041 );
buf ( n12377 , n9669 );
nand ( n12378 , n61750 , n12377 );
buf ( n61753 , n12378 );
not ( n12380 , n61753 );
and ( n61755 , n61749 , n12380 );
not ( n61756 , n61749 );
and ( n61757 , n61756 , n61753 );
nor ( n12384 , n61755 , n61757 );
buf ( n61759 , n12384 );
not ( n12386 , n61759 );
buf ( n61761 , n12386 );
not ( n61762 , n61761 );
or ( n61763 , n12372 , n61762 );
not ( n12390 , n394 );
nand ( n61765 , n12390 , n12384 );
nand ( n61766 , n61763 , n61765 );
nand ( n12393 , n12371 , n61766 );
nand ( n61768 , n12367 , n12393 );
not ( n61769 , n61768 );
nand ( n12396 , n11860 , n378 );
not ( n12397 , n12396 );
nand ( n12398 , n11844 , n61213 );
not ( n12399 , n12398 );
or ( n61774 , n12397 , n12399 );
nand ( n12401 , n11844 , n61213 , n11860 , n378 );
nand ( n12402 , n61774 , n12401 );
not ( n61777 , n12402 );
buf ( n61778 , n61777 );
buf ( n61779 , n61761 );
not ( n61780 , n61779 );
buf ( n12407 , n394 );
nand ( n12408 , n61780 , n12407 );
buf ( n12409 , n12408 );
buf ( n61784 , n12409 );
nand ( n12411 , n61778 , n61784 );
buf ( n12412 , n12411 );
not ( n61787 , n12412 );
or ( n61788 , n61769 , n61787 );
not ( n12415 , n61777 );
buf ( n61790 , n12409 );
not ( n12417 , n61790 );
buf ( n61792 , n12417 );
nand ( n12419 , n12415 , n61792 );
nand ( n12420 , n61788 , n12419 );
xor ( n12421 , n61703 , n12420 );
not ( n12422 , n10005 );
not ( n12423 , n12287 );
or ( n12424 , n12422 , n12423 );
not ( n12425 , n380 );
not ( n12426 , n61289 );
or ( n12427 , n12425 , n12426 );
not ( n12428 , n11911 );
not ( n12429 , n11910 );
or ( n12430 , n12428 , n12429 );
nand ( n12431 , n12430 , n59380 );
nand ( n12432 , n12427 , n12431 );
nand ( n61807 , n12432 , n59383 );
nand ( n61808 , n12424 , n61807 );
and ( n61809 , n12421 , n61808 );
and ( n12433 , n61703 , n12420 );
or ( n12434 , n61809 , n12433 );
buf ( n12435 , n12434 );
buf ( n61813 , n12435 );
nand ( n12437 , n12311 , n61813 );
buf ( n61815 , n12437 );
nand ( n12439 , n12307 , n61663 );
nand ( n12440 , n61815 , n12439 );
nand ( n12441 , n61654 , n12440 );
nand ( n12442 , n12270 , n12441 );
not ( n12443 , n12442 );
buf ( n61821 , n12443 );
not ( n12445 , n60678 );
not ( n12446 , n61673 );
or ( n12447 , n12445 , n12446 );
nand ( n12448 , n61334 , n10093 );
nand ( n12449 , n12447 , n12448 );
xor ( n12450 , n61279 , n61259 );
xnor ( n12451 , n12450 , n61298 );
or ( n12452 , n12449 , n12451 );
buf ( n61830 , n60498 );
not ( n12454 , n61830 );
buf ( n61832 , n11917 );
not ( n12456 , n61832 );
or ( n12457 , n12454 , n12456 );
buf ( n61835 , n61689 );
buf ( n61836 , n60476 );
nand ( n12460 , n61835 , n61836 );
buf ( n61838 , n12460 );
buf ( n61839 , n61838 );
nand ( n12463 , n12457 , n61839 );
buf ( n61841 , n12463 );
or ( n61842 , n61184 , n11818 );
nand ( n61843 , n61184 , n11818 );
nand ( n12467 , n61842 , n61843 );
xor ( n61845 , n61237 , n12467 );
not ( n61846 , n11105 );
not ( n12470 , n54740 );
not ( n12471 , n54737 );
or ( n61849 , n12470 , n12471 );
nand ( n12473 , n53730 , n53945 );
nand ( n61851 , n61849 , n12473 );
nand ( n61852 , n60352 , n10983 );
xor ( n12476 , n61851 , n61852 );
not ( n12477 , n12476 );
nand ( n61855 , n61846 , n12477 );
nand ( n61856 , n61845 , n61855 );
not ( n12480 , n61856 );
nand ( n12481 , n52045 , n51960 );
not ( n61859 , n12481 );
not ( n61860 , n11439 );
nand ( n12484 , n61860 , n2677 );
not ( n61862 , n11439 );
nand ( n61863 , n61862 , n2665 , n51914 );
not ( n12487 , n52029 );
nand ( n12488 , n12484 , n61863 , n12487 );
not ( n12489 , n12488 );
or ( n12490 , n61859 , n12489 );
not ( n12491 , n12481 );
nand ( n12492 , n12491 , n12484 , n61863 , n12487 );
nand ( n12493 , n12490 , n12492 );
not ( n61871 , n12493 );
or ( n12495 , n12480 , n61871 );
or ( n61873 , n61845 , n61855 );
nand ( n12497 , n12495 , n61873 );
xor ( n12498 , n61841 , n12497 );
xor ( n12499 , n61407 , n12026 );
buf ( n61877 , n61404 );
not ( n12501 , n61877 );
buf ( n61879 , n12501 );
and ( n12503 , n12499 , n61879 );
not ( n61881 , n12499 );
and ( n12505 , n61881 , n61404 );
nor ( n12506 , n12503 , n12505 );
and ( n61884 , n12498 , n12506 );
and ( n61885 , n61841 , n12497 );
or ( n12509 , n61884 , n61885 );
nand ( n12510 , n12452 , n12509 );
nand ( n61888 , n12449 , n12451 );
nand ( n12512 , n12510 , n61888 );
buf ( n61890 , n12512 );
not ( n61891 , n61890 );
buf ( n61892 , n61891 );
buf ( n12516 , n61892 );
nand ( n12517 , n61821 , n12516 );
buf ( n12518 , n12517 );
not ( n61896 , n12518 );
xor ( n12520 , n61580 , n61587 );
xor ( n61898 , n12520 , n61591 );
not ( n61899 , n61898 );
or ( n12523 , n61896 , n61899 );
buf ( n61901 , n12443 );
buf ( n61902 , n61892 );
or ( n12526 , n61901 , n61902 );
buf ( n61904 , n12526 );
nand ( n61905 , n12523 , n61904 );
buf ( n61906 , n61905 );
not ( n61907 , n61906 );
buf ( n61908 , n61907 );
buf ( n61909 , n61908 );
nand ( n12533 , n61614 , n61909 );
buf ( n61911 , n12533 );
and ( n12535 , n61456 , n12182 , n61608 , n61911 );
not ( n12536 , n61200 );
xor ( n12537 , n61855 , n12536 );
xnor ( n12538 , n12537 , n61237 );
and ( n61916 , n12538 , n12493 );
not ( n61917 , n12538 );
not ( n12541 , n12493 );
and ( n61919 , n61917 , n12541 );
nor ( n12543 , n61916 , n61919 );
not ( n61921 , n60498 );
not ( n61922 , n12322 );
or ( n12546 , n61921 , n61922 );
not ( n61924 , n378 );
not ( n61925 , n12476 );
or ( n12549 , n61924 , n61925 );
or ( n61927 , n12476 , n378 );
nand ( n61928 , n12549 , n61927 );
buf ( n61929 , n61928 );
buf ( n61930 , n60476 );
nand ( n12554 , n61929 , n61930 );
buf ( n61932 , n12554 );
nand ( n12556 , n12546 , n61932 );
xor ( n12557 , n12556 , n2591 );
not ( n61935 , n61768 );
not ( n61936 , n12409 );
not ( n12560 , n61777 );
or ( n12561 , n61936 , n12560 );
nand ( n12562 , n12402 , n61792 );
nand ( n61940 , n12561 , n12562 );
not ( n12564 , n61940 );
or ( n61942 , n61935 , n12564 );
or ( n12566 , n61768 , n61940 );
nand ( n12567 , n61942 , n12566 );
and ( n61945 , n12557 , n12567 );
and ( n12569 , n12556 , n2591 );
or ( n12570 , n61945 , n12569 );
xor ( n12571 , n12543 , n12570 );
buf ( n61949 , n60678 );
not ( n61950 , n61949 );
not ( n61951 , n382 );
not ( n12575 , n11749 );
or ( n61953 , n61951 , n12575 );
not ( n61954 , n382 );
nand ( n61955 , n61954 , n11364 );
nand ( n61956 , n61953 , n61955 );
buf ( n61957 , n61956 );
not ( n61958 , n61957 );
or ( n61959 , n61950 , n61958 );
nand ( n12583 , n12303 , n12305 , n10093 );
buf ( n61961 , n12583 );
nand ( n61962 , n61959 , n61961 );
buf ( n61963 , n61962 );
xor ( n61964 , n12571 , n61963 );
xor ( n12588 , n12556 , n2591 );
xor ( n61966 , n12588 , n12567 );
buf ( n61967 , n61966 );
not ( n12591 , n61967 );
buf ( n61969 , n396 );
not ( n61970 , n58739 );
not ( n61971 , n9402 );
or ( n12595 , n61970 , n61971 );
nand ( n61973 , n12595 , n58964 );
xnor ( n12597 , n61973 , n58958 );
buf ( n61975 , n12597 );
and ( n61976 , n61969 , n61975 );
buf ( n61977 , n61976 );
buf ( n61978 , n61233 );
not ( n61979 , n61978 );
nand ( n61980 , n61979 , n60498 );
xor ( n12604 , n395 , n12356 );
or ( n61982 , n61980 , n12604 );
not ( n12606 , n60498 );
not ( n12607 , n61979 );
or ( n12608 , n12606 , n12607 );
nand ( n12609 , n12608 , n12604 );
nand ( n12610 , n61982 , n12609 );
xor ( n12611 , n61977 , n12610 );
buf ( n61989 , n397 );
buf ( n61990 , n58957 );
buf ( n61991 , n58809 );
nand ( n12615 , n61990 , n61991 );
buf ( n61993 , n12615 );
buf ( n12617 , n61993 );
buf ( n12618 , n9607 );
xnor ( n12619 , n12617 , n12618 );
buf ( n12620 , n12619 );
buf ( n61998 , n12620 );
and ( n12622 , n61989 , n61998 );
buf ( n62000 , n12622 );
buf ( n62001 , n62000 );
xor ( n12625 , n61969 , n61975 );
buf ( n62003 , n12625 );
buf ( n62004 , n62003 );
xor ( n62005 , n62001 , n62004 );
buf ( n62006 , n382 );
not ( n12630 , n62006 );
buf ( n62008 , n59371 );
nand ( n62009 , n12630 , n62008 );
buf ( n62010 , n62009 );
buf ( n62011 , n62010 );
not ( n62012 , n62011 );
buf ( n62013 , n11860 );
not ( n12637 , n62013 );
or ( n62015 , n62012 , n12637 );
buf ( n62016 , n381 );
buf ( n62017 , n382 );
and ( n12641 , n62016 , n62017 );
buf ( n62019 , n59380 );
nor ( n12643 , n12641 , n62019 );
buf ( n62021 , n12643 );
buf ( n62022 , n62021 );
nand ( n62023 , n62015 , n62022 );
buf ( n62024 , n62023 );
buf ( n62025 , n62024 );
not ( n12645 , n62025 );
buf ( n62027 , n12645 );
buf ( n62028 , n62027 );
and ( n12648 , n62005 , n62028 );
and ( n12649 , n62001 , n62004 );
or ( n12650 , n12648 , n12649 );
buf ( n62032 , n12650 );
and ( n12652 , n12611 , n62032 );
and ( n12653 , n61977 , n12610 );
or ( n12654 , n12652 , n12653 );
not ( n12655 , n12654 );
not ( n12656 , n12655 );
nand ( n62038 , n2677 , n51788 );
nand ( n62039 , n51807 , n62038 , n51976 );
xor ( n62040 , n52041 , n62039 );
not ( n12657 , n62040 );
or ( n12658 , n12656 , n12657 );
not ( n12659 , n10093 );
buf ( n62044 , n61163 );
not ( n12661 , n62044 );
buf ( n62046 , n12661 );
nand ( n12663 , n62046 , n382 );
nand ( n62048 , n61163 , n59374 );
nand ( n12665 , n12663 , n62048 );
not ( n12666 , n12665 );
or ( n62051 , n12659 , n12666 );
not ( n62052 , n382 );
buf ( n62053 , n11912 );
not ( n62054 , n62053 );
buf ( n62055 , n62054 );
not ( n12672 , n62055 );
or ( n62057 , n62052 , n12672 );
buf ( n62058 , n382 );
not ( n12675 , n62058 );
buf ( n62060 , n11912 );
nand ( n12677 , n12675 , n62060 );
buf ( n62062 , n12677 );
nand ( n12679 , n62057 , n62062 );
nand ( n12680 , n12679 , n60678 );
nand ( n12681 , n62051 , n12680 );
nand ( n12682 , n12658 , n12681 );
not ( n12683 , n62040 );
nand ( n62068 , n12683 , n12654 );
nand ( n12685 , n12682 , n62068 );
not ( n12686 , n12685 );
or ( n12687 , n12591 , n12686 );
buf ( n12688 , n12685 );
or ( n12689 , n61967 , n12688 );
not ( n12690 , n11634 );
buf ( n62075 , n384 );
not ( n12692 , n62075 );
buf ( n62077 , n11494 );
not ( n12694 , n62077 );
or ( n12695 , n12692 , n12694 );
not ( n12696 , n60852 );
and ( n12697 , n11800 , n12696 );
not ( n12698 , n11800 );
and ( n62083 , n12698 , n60852 );
nor ( n12700 , n12697 , n62083 );
nand ( n62085 , n12700 , n59460 );
buf ( n62086 , n62085 );
nand ( n62087 , n12695 , n62086 );
buf ( n62088 , n62087 );
not ( n62089 , n62088 );
or ( n12706 , n12690 , n62089 );
and ( n12707 , n384 , n60979 );
not ( n62092 , n384 );
and ( n62093 , n62092 , n60644 );
or ( n12710 , n12707 , n62093 );
nand ( n62095 , n12710 , n385 );
nand ( n62096 , n12706 , n62095 );
nand ( n12713 , n12689 , n62096 );
nand ( n62098 , n12687 , n12713 );
xor ( n62099 , n61964 , n62098 );
xor ( n12716 , n61703 , n12420 );
xor ( n12717 , n12716 , n61808 );
not ( n62102 , n12717 );
not ( n62103 , n11634 );
not ( n12720 , n12710 );
or ( n62105 , n62103 , n12720 );
not ( n62106 , n384 );
not ( n12723 , n61329 );
or ( n12724 , n62106 , n12723 );
not ( n62109 , n384 );
nand ( n62110 , n62109 , n60666 );
nand ( n12727 , n12724 , n62110 );
nand ( n62112 , n12727 , n385 );
nand ( n62113 , n62105 , n62112 );
not ( n12730 , n62113 );
not ( n12731 , n12730 );
or ( n62116 , n62102 , n12731 );
not ( n12733 , n12717 );
nand ( n62118 , n12733 , n62113 );
nand ( n62119 , n62116 , n62118 );
not ( n12736 , n10093 );
not ( n62121 , n61956 );
or ( n62122 , n12736 , n62121 );
not ( n12739 , n62048 );
not ( n12740 , n12663 );
or ( n12741 , n12739 , n12740 );
nand ( n12742 , n12741 , n60678 );
nand ( n12743 , n62122 , n12742 );
not ( n12744 , n12743 );
not ( n12745 , n10005 );
not ( n62130 , n12432 );
or ( n12747 , n12745 , n62130 );
buf ( n62132 , n380 );
buf ( n12749 , n11902 );
xor ( n12750 , n62132 , n12749 );
buf ( n62135 , n12750 );
buf ( n62136 , n62135 );
buf ( n62137 , n11333 );
nand ( n12754 , n62136 , n62137 );
buf ( n62139 , n12754 );
nand ( n12756 , n12747 , n62139 );
not ( n12757 , n12756 );
nand ( n12758 , n12744 , n12757 );
not ( n12759 , n12758 );
buf ( n62144 , n60498 );
not ( n12761 , n62144 );
buf ( n62146 , n61928 );
not ( n12763 , n62146 );
or ( n12764 , n12761 , n12763 );
not ( n12765 , n11105 );
not ( n12766 , n61979 );
or ( n12767 , n12765 , n12766 );
buf ( n62152 , n11860 );
not ( n62153 , n62152 );
buf ( n62154 , n62153 );
nand ( n12771 , n62154 , n378 );
nand ( n62156 , n12767 , n12771 );
buf ( n62157 , n62156 );
buf ( n62158 , n60476 );
nand ( n12775 , n62157 , n62158 );
buf ( n12776 , n12775 );
buf ( n62161 , n12776 );
nand ( n12778 , n12764 , n62161 );
buf ( n62163 , n12778 );
xor ( n62164 , n12347 , n61739 );
not ( n12781 , n61766 );
xor ( n62166 , n62164 , n12781 );
xor ( n12783 , n62163 , n62166 );
buf ( n62168 , n11333 );
not ( n62169 , n62168 );
and ( n62170 , n61366 , n59380 );
not ( n12787 , n61366 );
and ( n62172 , n12787 , n380 );
or ( n62173 , n62170 , n62172 );
buf ( n62174 , n62173 );
not ( n62175 , n62174 );
or ( n12792 , n62169 , n62175 );
buf ( n62177 , n62135 );
buf ( n62178 , n10005 );
nand ( n12795 , n62177 , n62178 );
buf ( n62180 , n12795 );
buf ( n12797 , n62180 );
nand ( n12798 , n12792 , n12797 );
buf ( n12799 , n12798 );
and ( n62184 , n12783 , n12799 );
and ( n62185 , n62163 , n62166 );
or ( n12802 , n62184 , n62185 );
not ( n62187 , n12802 );
or ( n12804 , n12759 , n62187 );
nand ( n62189 , n12743 , n12756 );
nand ( n62190 , n12804 , n62189 );
and ( n12807 , n62119 , n62190 );
not ( n62192 , n62119 );
not ( n62193 , n62190 );
and ( n12810 , n62192 , n62193 );
nor ( n12811 , n12807 , n12810 );
xor ( n62196 , n62099 , n12811 );
not ( n62197 , n62196 );
not ( n62198 , n12685 );
xor ( n12815 , n61966 , n62198 );
xor ( n62200 , n12815 , n62096 );
not ( n62201 , n62200 );
not ( n12818 , n62201 );
xor ( n62203 , n12756 , n12802 );
xnor ( n12820 , n62203 , n12743 );
not ( n12821 , n12820 );
not ( n62206 , n12821 );
or ( n62207 , n12818 , n62206 );
not ( n12824 , n12820 );
not ( n62209 , n62200 );
or ( n12826 , n12824 , n62209 );
not ( n62211 , n385 );
not ( n62212 , n62088 );
or ( n12829 , n62211 , n62212 );
not ( n62214 , n384 );
not ( n62215 , n61340 );
or ( n12832 , n62214 , n62215 );
nand ( n12833 , n59460 , n11364 );
nand ( n12834 , n12832 , n12833 );
nand ( n62219 , n11634 , n12834 );
nand ( n62220 , n12829 , n62219 );
not ( n12837 , n62220 );
xor ( n12838 , n62163 , n62166 );
xor ( n12839 , n12838 , n12799 );
not ( n12840 , n12839 );
not ( n12841 , n12840 );
not ( n12842 , n12841 );
or ( n62227 , n12837 , n12842 );
nand ( n12844 , n62088 , n385 );
nand ( n62229 , n12840 , n62219 , n12844 );
not ( n12846 , n10005 );
not ( n62231 , n62173 );
or ( n12848 , n12846 , n62231 );
buf ( n62233 , n380 );
not ( n62234 , n62233 );
buf ( n62235 , n12476 );
not ( n12852 , n62235 );
or ( n62237 , n62234 , n12852 );
nand ( n62238 , n12477 , n59380 );
buf ( n62239 , n62238 );
nand ( n62240 , n62237 , n62239 );
buf ( n62241 , n62240 );
buf ( n62242 , n62241 );
buf ( n62243 , n59383 );
nand ( n62244 , n62242 , n62243 );
buf ( n62245 , n62244 );
nand ( n62246 , n12848 , n62245 );
not ( n62247 , n62246 );
or ( n12864 , n2466 , n2461 );
not ( n12865 , n12864 );
not ( n62250 , n2677 );
or ( n12867 , n12865 , n62250 );
and ( n62252 , n2665 , n51914 , n12864 );
not ( n12869 , n51802 );
not ( n12870 , n12869 );
nor ( n12871 , n62252 , n12870 );
nand ( n12872 , n12867 , n12871 );
not ( n12873 , n2477 );
nand ( n12874 , n12873 , n51800 );
and ( n12875 , n12872 , n12874 );
not ( n12876 , n12872 );
not ( n12877 , n12874 );
and ( n12878 , n12876 , n12877 );
nor ( n62263 , n12875 , n12878 );
not ( n12880 , n62263 );
not ( n12881 , n12880 );
or ( n12882 , n62247 , n12881 );
not ( n12883 , n62246 );
not ( n12884 , n12883 );
not ( n12885 , n62263 );
or ( n12886 , n12884 , n12885 );
xor ( n12887 , n61977 , n12610 );
xor ( n12888 , n12887 , n62032 );
nand ( n12889 , n12886 , n12888 );
nand ( n62274 , n12882 , n12889 );
nand ( n12891 , n62229 , n62274 );
nand ( n12892 , n62227 , n12891 );
nand ( n62277 , n12826 , n12892 );
nand ( n12894 , n62207 , n62277 );
not ( n62279 , n12894 );
nand ( n12896 , n62197 , n62279 );
nand ( n62281 , n12733 , n12730 );
and ( n12898 , n62190 , n62281 );
buf ( n12899 , n12717 );
and ( n12900 , n12899 , n62113 );
nor ( n62285 , n12898 , n12900 );
not ( n62286 , n62285 );
not ( n12903 , n61663 );
not ( n12904 , n12434 );
not ( n62289 , n12904 );
or ( n12906 , n12903 , n62289 );
buf ( n62291 , n12434 );
buf ( n62292 , n61666 );
nand ( n62293 , n62291 , n62292 );
buf ( n62294 , n62293 );
nand ( n12911 , n12906 , n62294 );
and ( n62296 , n12911 , n12307 );
not ( n12913 , n12911 );
and ( n12914 , n12913 , n12308 );
nor ( n12915 , n62296 , n12914 );
not ( n12916 , n12915 );
or ( n62301 , n62286 , n12916 );
not ( n62302 , n12915 );
not ( n62303 , n62285 );
nand ( n12920 , n62302 , n62303 );
nand ( n62305 , n62301 , n12920 );
not ( n12922 , n385 );
not ( n62307 , n12250 );
or ( n62308 , n12922 , n62307 );
nand ( n12925 , n12727 , n11634 );
nand ( n62310 , n62308 , n12925 );
xor ( n12927 , n61841 , n12497 );
xor ( n12928 , n12927 , n12506 );
xor ( n62313 , n62310 , n12928 );
xor ( n62314 , n12543 , n12570 );
and ( n12931 , n62314 , n61963 );
and ( n62316 , n12543 , n12570 );
or ( n12933 , n12931 , n62316 );
xor ( n62318 , n62313 , n12933 );
not ( n62319 , n62318 );
and ( n12936 , n62305 , n62319 );
not ( n62321 , n62305 );
and ( n62322 , n62321 , n62318 );
nor ( n12939 , n12936 , n62322 );
xor ( n62324 , n61964 , n62098 );
and ( n62325 , n62324 , n12811 );
and ( n12942 , n61964 , n62098 );
or ( n62327 , n62325 , n12942 );
buf ( n62328 , n62327 );
not ( n62329 , n62328 );
buf ( n62330 , n62329 );
nand ( n12947 , n12939 , n62330 );
nand ( n12948 , n12896 , n12947 );
not ( n12949 , n12948 );
not ( n12950 , n12949 );
not ( n62335 , n385 );
buf ( n62336 , n384 );
not ( n12953 , n62336 );
buf ( n62338 , n62046 );
not ( n12955 , n62338 );
or ( n12956 , n12953 , n12955 );
buf ( n62341 , n61163 );
buf ( n62342 , n59460 );
nand ( n12959 , n62341 , n62342 );
buf ( n12960 , n12959 );
buf ( n62345 , n12960 );
nand ( n12962 , n12956 , n62345 );
buf ( n62347 , n12962 );
not ( n12964 , n62347 );
or ( n62349 , n62335 , n12964 );
and ( n12966 , n384 , n62055 );
not ( n12967 , n384 );
and ( n62352 , n12967 , n11912 );
or ( n62353 , n12966 , n62352 );
nand ( n12970 , n62353 , n11634 );
nand ( n12971 , n62349 , n12970 );
not ( n12972 , n12971 );
not ( n62357 , n12972 );
buf ( n62358 , n58941 );
buf ( n62359 , n58932 );
xor ( n12976 , n62358 , n62359 );
buf ( n62361 , n12976 );
buf ( n62362 , n62361 );
buf ( n62363 , n58919 );
xnor ( n62364 , n62362 , n62363 );
buf ( n62365 , n62364 );
nand ( n12982 , n62365 , n399 );
not ( n12983 , n12982 );
not ( n62368 , n12983 );
buf ( n62369 , n58943 );
not ( n62370 , n62369 );
buf ( n62371 , n58948 );
buf ( n62372 , n58871 );
nand ( n62373 , n62371 , n62372 );
buf ( n62374 , n62373 );
buf ( n62375 , n62374 );
not ( n12992 , n62375 );
or ( n62377 , n62370 , n12992 );
buf ( n62378 , n62374 );
buf ( n62379 , n58943 );
or ( n62380 , n62378 , n62379 );
nand ( n62381 , n62377 , n62380 );
buf ( n62382 , n62381 );
not ( n12999 , n62382 );
not ( n13000 , n398 );
nand ( n13001 , n12999 , n13000 );
not ( n13002 , n13001 );
or ( n13003 , n62368 , n13002 );
nand ( n13004 , n398 , n62382 );
nand ( n13005 , n13003 , n13004 );
xor ( n13006 , n61989 , n61998 );
buf ( n62391 , n13006 );
xor ( n13008 , n13005 , n62391 );
nor ( n13009 , n61978 , n59377 );
xor ( n13010 , n13008 , n13009 );
not ( n13011 , n51459 );
not ( n13012 , n52057 );
or ( n13013 , n13011 , n13012 );
nand ( n62398 , n13013 , n52002 );
nand ( n62399 , n2521 , n51829 );
nand ( n13016 , n62399 , n2394 );
xnor ( n62401 , n62398 , n13016 );
xor ( n13018 , n13010 , n62401 );
not ( n13019 , n10093 );
not ( n13020 , n382 );
buf ( n62405 , n61369 );
not ( n13022 , n62405 );
buf ( n62407 , n13022 );
not ( n13024 , n62407 );
or ( n62409 , n13020 , n13024 );
buf ( n62410 , n382 );
not ( n62411 , n62410 );
buf ( n62412 , n61369 );
nand ( n62413 , n62411 , n62412 );
buf ( n62414 , n62413 );
nand ( n13031 , n62409 , n62414 );
not ( n62416 , n13031 );
or ( n13033 , n13019 , n62416 );
buf ( n62418 , n382 );
not ( n13035 , n62418 );
buf ( n62420 , n12476 );
not ( n62421 , n62420 );
or ( n13038 , n13035 , n62421 );
not ( n62423 , n382 );
nand ( n62424 , n62423 , n12477 );
buf ( n62425 , n62424 );
nand ( n13042 , n13038 , n62425 );
buf ( n62427 , n13042 );
nand ( n62428 , n62427 , n60678 );
nand ( n13045 , n13033 , n62428 );
and ( n13046 , n13018 , n13045 );
and ( n62431 , n13010 , n62401 );
or ( n13048 , n13046 , n62431 );
not ( n13049 , n13048 );
or ( n62434 , n62357 , n13049 );
or ( n62435 , n13048 , n12972 );
nand ( n62436 , n62434 , n62435 );
buf ( n62437 , n62436 );
not ( n13054 , n62437 );
not ( n62439 , n2665 );
not ( n62440 , n51459 );
or ( n13057 , n62439 , n62440 );
nand ( n13058 , n13057 , n51987 );
nand ( n13059 , n12864 , n12869 );
xnor ( n13060 , n13058 , n13059 );
buf ( n62445 , n13060 );
not ( n62446 , n10093 );
buf ( n62447 , n382 );
buf ( n62448 , n11902 );
buf ( n62449 , n62448 );
buf ( n62450 , n62449 );
buf ( n62451 , n62450 );
and ( n62452 , n62447 , n62451 );
not ( n13069 , n62447 );
buf ( n62454 , n62450 );
not ( n62455 , n62454 );
buf ( n62456 , n62455 );
buf ( n13073 , n62456 );
and ( n62458 , n13069 , n13073 );
nor ( n13075 , n62452 , n62458 );
buf ( n62460 , n13075 );
not ( n13077 , n62460 );
or ( n62462 , n62446 , n13077 );
nand ( n62463 , n13031 , n60678 );
nand ( n62464 , n62462 , n62463 );
buf ( n62465 , n62464 );
xor ( n62466 , n62445 , n62465 );
xor ( n62467 , n13005 , n62391 );
and ( n13084 , n62467 , n13009 );
and ( n62469 , n13005 , n62391 );
or ( n62470 , n13084 , n62469 );
buf ( n62471 , n62470 );
xor ( n62472 , n62001 , n62004 );
xor ( n62473 , n62472 , n62028 );
buf ( n62474 , n62473 );
buf ( n62475 , n62474 );
xor ( n62476 , n62471 , n62475 );
buf ( n62477 , n10005 );
not ( n13094 , n62477 );
buf ( n62479 , n62241 );
not ( n13096 , n62479 );
or ( n62481 , n13094 , n13096 );
buf ( n62482 , n380 );
not ( n13099 , n62482 );
buf ( n62484 , n62154 );
not ( n62485 , n62484 );
or ( n13102 , n13099 , n62485 );
buf ( n62487 , n62154 );
not ( n13104 , n62487 );
buf ( n62489 , n13104 );
buf ( n62490 , n62489 );
buf ( n62491 , n59380 );
nand ( n13108 , n62490 , n62491 );
buf ( n62493 , n13108 );
buf ( n13110 , n62493 );
nand ( n62495 , n13102 , n13110 );
buf ( n62496 , n62495 );
buf ( n62497 , n62496 );
buf ( n62498 , n59383 );
nand ( n62499 , n62497 , n62498 );
buf ( n62500 , n62499 );
buf ( n62501 , n62500 );
nand ( n62502 , n62481 , n62501 );
buf ( n62503 , n62502 );
buf ( n62504 , n62503 );
xor ( n13121 , n62476 , n62504 );
buf ( n13122 , n13121 );
buf ( n62507 , n13122 );
xnor ( n13124 , n62466 , n62507 );
buf ( n62509 , n13124 );
buf ( n62510 , n62509 );
not ( n13127 , n62510 );
and ( n13128 , n13054 , n13127 );
buf ( n62513 , n62509 );
buf ( n62514 , n62436 );
and ( n13131 , n62513 , n62514 );
nor ( n13132 , n13128 , n13131 );
buf ( n62517 , n13132 );
buf ( n62518 , n62517 );
nand ( n62519 , n12982 , n62382 , n13000 );
nand ( n13136 , n12999 , n12982 , n398 );
nand ( n13137 , n12999 , n12983 , n13000 );
not ( n13138 , n12999 );
nand ( n62523 , n13138 , n12983 , n398 );
nand ( n13140 , n62519 , n13136 , n13137 , n62523 );
buf ( n62525 , n13140 );
not ( n62526 , n62525 );
buf ( n62527 , n384 );
not ( n13144 , n62527 );
buf ( n62529 , n59454 );
nand ( n13146 , n13144 , n62529 );
buf ( n62531 , n13146 );
buf ( n62532 , n62531 );
not ( n13149 , n62532 );
buf ( n62534 , n62489 );
not ( n13151 , n62534 );
or ( n13152 , n13149 , n13151 );
buf ( n62537 , n383 );
buf ( n62538 , n384 );
and ( n62539 , n62537 , n62538 );
buf ( n62540 , n59374 );
nor ( n62541 , n62539 , n62540 );
buf ( n62542 , n62541 );
buf ( n62543 , n62542 );
nand ( n13160 , n13152 , n62543 );
buf ( n62545 , n13160 );
buf ( n62546 , n62545 );
nand ( n13163 , n62526 , n62546 );
buf ( n62548 , n13163 );
not ( n13165 , n62548 );
not ( n62550 , n10093 );
not ( n62551 , n62427 );
or ( n13168 , n62550 , n62551 );
and ( n62553 , n59374 , n62154 );
not ( n13170 , n59374 );
and ( n13171 , n13170 , n62489 );
nor ( n13172 , n62553 , n13171 );
nand ( n13173 , n13172 , n60678 );
nand ( n13174 , n13168 , n13173 );
not ( n13175 , n13174 );
or ( n13176 , n13165 , n13175 );
buf ( n62561 , n62545 );
not ( n13178 , n62561 );
buf ( n62563 , n13140 );
nand ( n13180 , n13178 , n62563 );
buf ( n62565 , n13180 );
nand ( n62566 , n13176 , n62565 );
not ( n13183 , n62566 );
not ( n62568 , n385 );
not ( n13185 , n62353 );
or ( n62570 , n62568 , n13185 );
buf ( n62571 , n11634 );
and ( n13188 , n384 , n62450 );
not ( n13189 , n384 );
and ( n13190 , n13189 , n62456 );
nor ( n13191 , n13188 , n13190 );
buf ( n62576 , n13191 );
nand ( n13193 , n62571 , n62576 );
buf ( n62578 , n13193 );
nand ( n62579 , n62570 , n62578 );
not ( n13196 , n62579 );
nand ( n62581 , n13183 , n13196 );
not ( n13198 , n62581 );
not ( n13199 , n11634 );
not ( n13200 , n384 );
not ( n13201 , n62407 );
or ( n13202 , n13200 , n13201 );
buf ( n62587 , n384 );
not ( n62588 , n62587 );
buf ( n62589 , n61369 );
nand ( n13206 , n62588 , n62589 );
buf ( n62591 , n13206 );
nand ( n13208 , n13202 , n62591 );
not ( n62593 , n13208 );
or ( n13210 , n13199 , n62593 );
nand ( n62595 , n13191 , n385 );
nand ( n62596 , n13210 , n62595 );
not ( n13213 , n62596 );
not ( n62598 , n2625 );
buf ( n62599 , n62598 );
nand ( n13216 , n13213 , n62599 );
not ( n13217 , n13216 );
not ( n13218 , n399 );
not ( n62603 , n13218 );
not ( n62604 , n62365 );
or ( n13221 , n62603 , n62604 );
or ( n62606 , n62365 , n13218 );
nand ( n62607 , n13221 , n62606 );
buf ( n62608 , n62607 );
buf ( n62609 , n11860 );
buf ( n62610 , n10093 );
and ( n13227 , n62609 , n62610 );
buf ( n62612 , n13227 );
buf ( n62613 , n62612 );
xor ( n62614 , n62608 , n62613 );
buf ( n62615 , n58910 );
not ( n62616 , n62615 );
buf ( n62617 , n62616 );
buf ( n62618 , n62617 );
not ( n13235 , n62618 );
buf ( n62620 , n9565 );
not ( n13237 , n62620 );
buf ( n62622 , n9579 );
nand ( n62623 , n13237 , n62622 );
buf ( n62624 , n62623 );
buf ( n62625 , n62624 );
not ( n13242 , n62625 );
or ( n13243 , n13235 , n13242 );
buf ( n62628 , n62624 );
buf ( n62629 , n62617 );
or ( n62630 , n62628 , n62629 );
nand ( n13247 , n13243 , n62630 );
buf ( n62632 , n13247 );
buf ( n62633 , n62632 );
not ( n62634 , n62633 );
buf ( n62635 , n62634 );
buf ( n62636 , n400 );
not ( n13253 , n62636 );
buf ( n62638 , n13253 );
and ( n62639 , n62635 , n62638 );
nor ( n62640 , n62639 , n59460 );
not ( n13257 , n62640 );
buf ( n62642 , n11860 );
buf ( n62643 , n385 );
nand ( n13260 , n62642 , n62643 );
buf ( n13261 , n13260 );
not ( n62646 , n13261 );
or ( n62647 , n13257 , n62646 );
nand ( n13264 , n62632 , n400 );
nand ( n13265 , n62647 , n13264 );
buf ( n62650 , n13265 );
and ( n13267 , n62614 , n62650 );
and ( n62652 , n62608 , n62613 );
or ( n62653 , n13267 , n62652 );
buf ( n62654 , n62653 );
not ( n13271 , n62654 );
or ( n62656 , n13217 , n13271 );
not ( n13273 , n62599 );
buf ( n62658 , n13273 );
buf ( n62659 , n62596 );
nand ( n13276 , n62658 , n62659 );
buf ( n62661 , n13276 );
nand ( n62662 , n62656 , n62661 );
not ( n13279 , n62662 );
or ( n13280 , n13198 , n13279 );
not ( n13281 , n13196 );
nand ( n13282 , n13281 , n62566 );
nand ( n62667 , n13280 , n13282 );
buf ( n62668 , n62667 );
not ( n13285 , n62668 );
buf ( n62670 , n13285 );
buf ( n62671 , n62670 );
nand ( n13288 , n62518 , n62671 );
buf ( n62673 , n13288 );
buf ( n62674 , n62673 );
not ( n62675 , n62674 );
xor ( n62676 , n62608 , n62613 );
xor ( n13293 , n62676 , n62650 );
buf ( n62678 , n13293 );
buf ( n13295 , n62678 );
not ( n62680 , n385 );
not ( n13297 , n13208 );
or ( n62682 , n62680 , n13297 );
not ( n62683 , n384 );
not ( n13300 , n12477 );
or ( n62685 , n62683 , n13300 );
or ( n13302 , n384 , n12477 );
nand ( n62687 , n62685 , n13302 );
buf ( n62688 , n62687 );
not ( n13305 , n62688 );
buf ( n62690 , n11634 );
nand ( n13307 , n13305 , n62690 );
buf ( n62692 , n13307 );
nand ( n13309 , n62682 , n62692 );
buf ( n62694 , n13309 );
xor ( n62695 , n13295 , n62694 );
buf ( n62696 , n401 );
not ( n62697 , n62696 );
buf ( n62698 , n58902 );
buf ( n62699 , n58907 );
or ( n62700 , n62698 , n62699 );
buf ( n62701 , n62617 );
nand ( n13318 , n62700 , n62701 );
buf ( n13319 , n13318 );
buf ( n62704 , n13319 );
not ( n13321 , n62704 );
or ( n62706 , n62697 , n13321 );
buf ( n62707 , n13261 );
buf ( n62708 , n13319 );
buf ( n62709 , n401 );
nor ( n13326 , n62708 , n62709 );
buf ( n13327 , n13326 );
buf ( n62712 , n13327 );
or ( n13329 , n62707 , n62712 );
nand ( n62714 , n62706 , n13329 );
buf ( n62715 , n62714 );
buf ( n62716 , n62715 );
nand ( n13333 , n13261 , n384 );
buf ( n13334 , n13333 );
xor ( n13335 , n62635 , n62638 );
buf ( n62720 , n13335 );
xnor ( n13337 , n13334 , n62720 );
buf ( n62722 , n13337 );
buf ( n13339 , n62722 );
xor ( n13340 , n62716 , n13339 );
buf ( n62725 , n11634 );
not ( n13342 , n62725 );
buf ( n62727 , n62154 );
not ( n62728 , n62727 );
or ( n62729 , n13342 , n62728 );
buf ( n62730 , n62687 );
buf ( n62731 , n61007 );
or ( n13348 , n62730 , n62731 );
nand ( n13349 , n62729 , n13348 );
buf ( n62734 , n13349 );
buf ( n62735 , n62734 );
and ( n13352 , n13340 , n62735 );
and ( n13353 , n62716 , n13339 );
or ( n13354 , n13352 , n13353 );
buf ( n62739 , n13354 );
buf ( n62740 , n62739 );
and ( n13357 , n62695 , n62740 );
and ( n62742 , n13295 , n62694 );
or ( n13359 , n13357 , n62742 );
buf ( n62744 , n13359 );
not ( n13361 , n62744 );
buf ( n62746 , n62654 );
buf ( n62747 , n62598 );
and ( n13364 , n62746 , n62747 );
not ( n13365 , n62746 );
buf ( n62750 , n2625 );
and ( n13367 , n13365 , n62750 );
nor ( n13368 , n13364 , n13367 );
buf ( n62753 , n13368 );
buf ( n62754 , n62753 );
not ( n13371 , n62754 );
buf ( n62756 , n62596 );
not ( n62757 , n62756 );
and ( n13374 , n13371 , n62757 );
buf ( n13375 , n62596 );
buf ( n62760 , n62753 );
and ( n62761 , n13375 , n62760 );
nor ( n13378 , n13374 , n62761 );
buf ( n62763 , n13378 );
buf ( n62764 , n62763 );
xor ( n62765 , n62545 , n13140 );
xor ( n62766 , n62765 , n13174 );
buf ( n62767 , n62766 );
nand ( n13384 , n62764 , n62767 );
buf ( n62769 , n13384 );
not ( n13386 , n62769 );
or ( n62771 , n13361 , n13386 );
buf ( n62772 , n62763 );
not ( n13389 , n62772 );
buf ( n13390 , n13389 );
buf ( n62775 , n62766 );
not ( n13392 , n62775 );
buf ( n62777 , n13392 );
nand ( n62778 , n13390 , n62777 );
nand ( n13395 , n62771 , n62778 );
xor ( n13396 , n13010 , n62401 );
xor ( n13397 , n13396 , n13045 );
nor ( n13398 , n13395 , n13397 );
xor ( n13399 , n62579 , n62566 );
not ( n13400 , n13399 );
not ( n13401 , n62662 );
or ( n13402 , n13400 , n13401 );
or ( n13403 , n62662 , n13399 );
nand ( n62788 , n13402 , n13403 );
or ( n13405 , n13398 , n62788 );
nand ( n62790 , n13395 , n13397 );
nand ( n13407 , n13405 , n62790 );
buf ( n62792 , n13407 );
not ( n13409 , n62792 );
or ( n13410 , n62675 , n13409 );
buf ( n62795 , n62517 );
not ( n13412 , n62795 );
buf ( n62797 , n13412 );
buf ( n62798 , n62797 );
buf ( n62799 , n62667 );
nand ( n13416 , n62798 , n62799 );
buf ( n62801 , n13416 );
buf ( n62802 , n62801 );
nand ( n13419 , n13410 , n62802 );
buf ( n62804 , n13419 );
not ( n13421 , n62804 );
buf ( n62806 , n62464 );
buf ( n62807 , n13060 );
or ( n13424 , n62806 , n62807 );
buf ( n62809 , n13122 );
nand ( n13426 , n13424 , n62809 );
buf ( n62811 , n13426 );
buf ( n62812 , n62811 );
buf ( n62813 , n13060 );
buf ( n62814 , n62464 );
nand ( n13431 , n62813 , n62814 );
buf ( n62816 , n13431 );
buf ( n62817 , n62816 );
nand ( n13434 , n62812 , n62817 );
buf ( n62819 , n13434 );
not ( n13436 , n12883 );
and ( n13437 , n12888 , n62263 );
not ( n13438 , n12888 );
and ( n13439 , n13438 , n12880 );
nor ( n13440 , n13437 , n13439 );
not ( n13441 , n13440 );
not ( n13442 , n13441 );
or ( n13443 , n13436 , n13442 );
nand ( n13444 , n13440 , n62246 );
nand ( n13445 , n13443 , n13444 );
xor ( n13446 , n62819 , n13445 );
xor ( n13447 , n62471 , n62475 );
and ( n13448 , n13447 , n62504 );
and ( n13449 , n62471 , n62475 );
or ( n13450 , n13448 , n13449 );
buf ( n62835 , n13450 );
buf ( n13452 , n62835 );
not ( n13453 , n10093 );
not ( n62838 , n12679 );
or ( n62839 , n13453 , n62838 );
buf ( n62840 , n60678 );
buf ( n62841 , n62460 );
nand ( n13458 , n62840 , n62841 );
buf ( n62843 , n13458 );
nand ( n13460 , n62839 , n62843 );
buf ( n62845 , n13460 );
xor ( n13462 , n13452 , n62845 );
not ( n13463 , n385 );
not ( n13464 , n12834 );
or ( n13465 , n13463 , n13464 );
nand ( n13466 , n62347 , n11634 );
nand ( n13467 , n13465 , n13466 );
buf ( n62852 , n13467 );
xor ( n13469 , n13462 , n62852 );
buf ( n62854 , n13469 );
xor ( n13471 , n13446 , n62854 );
not ( n13472 , n13471 );
buf ( n62857 , n13048 );
not ( n13474 , n62857 );
buf ( n13475 , n12972 );
nand ( n13476 , n13474 , n13475 );
buf ( n13477 , n13476 );
buf ( n62862 , n13477 );
not ( n13479 , n62862 );
buf ( n62864 , n62509 );
not ( n13481 , n62864 );
buf ( n62866 , n13481 );
buf ( n62867 , n62866 );
not ( n13484 , n62867 );
or ( n13485 , n13479 , n13484 );
buf ( n62870 , n12971 );
buf ( n62871 , n13048 );
nand ( n13488 , n62870 , n62871 );
buf ( n62873 , n13488 );
buf ( n62874 , n62873 );
nand ( n13491 , n13485 , n62874 );
buf ( n62876 , n13491 );
not ( n62877 , n62876 );
nand ( n13494 , n13472 , n62877 );
not ( n13495 , n13494 );
or ( n62880 , n13421 , n13495 );
nand ( n13497 , n62876 , n13471 );
nand ( n62882 , n62880 , n13497 );
not ( n13499 , n62882 );
not ( n13500 , n12892 );
not ( n13501 , n12820 );
or ( n62886 , n13500 , n13501 );
or ( n13503 , n12892 , n12820 );
nand ( n62888 , n62886 , n13503 );
xor ( n62889 , n62888 , n62200 );
xor ( n13506 , n12654 , n62040 );
xnor ( n62891 , n13506 , n12681 );
xor ( n13508 , n13452 , n62845 );
and ( n13509 , n13508 , n62852 );
and ( n13510 , n13452 , n62845 );
or ( n13511 , n13509 , n13510 );
buf ( n62896 , n13511 );
xor ( n13513 , n62891 , n62896 );
not ( n13514 , n62274 );
not ( n13515 , n12840 );
or ( n13516 , n13514 , n13515 );
buf ( n62901 , n62274 );
not ( n13518 , n62901 );
buf ( n62903 , n13518 );
buf ( n62904 , n62903 );
buf ( n62905 , n12839 );
nand ( n13522 , n62904 , n62905 );
buf ( n62907 , n13522 );
nand ( n62908 , n13516 , n62907 );
not ( n13525 , n385 );
not ( n62910 , n62088 );
or ( n62911 , n13525 , n62910 );
nand ( n13528 , n62911 , n62219 );
and ( n62913 , n62908 , n13528 );
not ( n13530 , n62908 );
not ( n62915 , n13528 );
and ( n13532 , n13530 , n62915 );
nor ( n62917 , n62913 , n13532 );
and ( n13534 , n13513 , n62917 );
and ( n62919 , n62891 , n62896 );
or ( n13536 , n13534 , n62919 );
buf ( n62921 , n13536 );
not ( n62922 , n62921 );
buf ( n62923 , n62922 );
nand ( n13540 , n62889 , n62923 );
xor ( n62925 , n62891 , n62896 );
xor ( n13542 , n62925 , n62917 );
not ( n13543 , n13542 );
buf ( n62928 , n13543 );
xor ( n13545 , n62819 , n13445 );
and ( n13546 , n13545 , n62854 );
and ( n13547 , n62819 , n13445 );
or ( n13548 , n13546 , n13547 );
buf ( n62933 , n13548 );
not ( n13550 , n62933 );
buf ( n62935 , n13550 );
buf ( n62936 , n62935 );
nand ( n13553 , n62928 , n62936 );
buf ( n13554 , n13553 );
and ( n62939 , n13540 , n13554 );
not ( n62940 , n62939 );
or ( n13557 , n13499 , n62940 );
buf ( n62942 , n13542 );
buf ( n62943 , n13548 );
and ( n13560 , n62942 , n62943 );
buf ( n62945 , n13560 );
not ( n13562 , n62945 );
not ( n13563 , n13540 );
or ( n13564 , n13562 , n13563 );
not ( n13565 , n62889 );
buf ( n62950 , n62923 );
not ( n13567 , n62950 );
buf ( n62952 , n13567 );
nand ( n13569 , n13565 , n62952 );
nand ( n13570 , n13564 , n13569 );
not ( n13571 , n13570 );
nand ( n13572 , n13557 , n13571 );
not ( n13573 , n13572 );
or ( n13574 , n12950 , n13573 );
and ( n13575 , n62196 , n12894 );
not ( n62960 , n13575 );
not ( n13576 , n12947 );
or ( n62962 , n62960 , n13576 );
not ( n13578 , n12939 );
nand ( n62964 , n13578 , n62327 );
nand ( n13580 , n62962 , n62964 );
not ( n62966 , n13580 );
nand ( n13582 , n13574 , n62966 );
not ( n13583 , n13582 );
not ( n13584 , n61892 );
not ( n13585 , n12443 );
or ( n62971 , n13584 , n13585 );
nand ( n62972 , n12512 , n12442 );
nand ( n13588 , n62971 , n62972 );
and ( n62974 , n13588 , n61898 );
not ( n13590 , n13588 );
not ( n62976 , n61898 );
and ( n62977 , n13590 , n62976 );
nor ( n62978 , n62974 , n62977 );
xor ( n13594 , n62310 , n12928 );
and ( n62980 , n13594 , n12933 );
and ( n62981 , n62310 , n12928 );
or ( n13597 , n62980 , n62981 );
xor ( n13598 , n12451 , n12449 );
xor ( n62984 , n13598 , n12509 );
or ( n13600 , n13597 , n62984 );
not ( n62986 , n61647 );
not ( n13602 , n61642 );
or ( n62988 , n62986 , n13602 );
nand ( n13604 , n61652 , n61631 );
nand ( n62990 , n62988 , n13604 );
not ( n62991 , n12440 );
and ( n13607 , n62990 , n62991 );
not ( n62993 , n62990 );
and ( n62994 , n62993 , n12440 );
nor ( n13610 , n13607 , n62994 );
not ( n13611 , n13610 );
and ( n13612 , n13600 , n13611 );
and ( n13613 , n62984 , n13597 );
nor ( n13614 , n13612 , n13613 );
nand ( n13615 , n62978 , n13614 );
not ( n63001 , n62303 );
buf ( n13617 , n12915 );
not ( n13618 , n13617 );
nand ( n63004 , n62319 , n13618 );
not ( n13620 , n63004 );
or ( n63006 , n63001 , n13620 );
nand ( n13622 , n13617 , n62318 );
nand ( n63008 , n63006 , n13622 );
not ( n13624 , n63008 );
xor ( n63010 , n62984 , n13597 );
and ( n13626 , n63010 , n13611 );
not ( n13627 , n63010 );
and ( n13628 , n13627 , n13610 );
nor ( n13629 , n13626 , n13628 );
not ( n63015 , n13629 );
nand ( n13631 , n13624 , n63015 );
and ( n13632 , n13615 , n13631 );
not ( n13633 , n13632 );
or ( n13634 , n13583 , n13633 );
buf ( n63020 , n13629 );
buf ( n63021 , n63008 );
and ( n63022 , n63020 , n63021 );
buf ( n63023 , n63022 );
not ( n63024 , n63023 );
not ( n63025 , n13615 );
or ( n63026 , n63024 , n63025 );
buf ( n63027 , n13614 );
not ( n63028 , n63027 );
buf ( n63029 , n63028 );
not ( n63030 , n62978 );
nand ( n13646 , n63029 , n63030 );
nand ( n13647 , n63026 , n13646 );
not ( n13648 , n13647 );
nand ( n13649 , n13634 , n13648 );
and ( n63035 , n60651 , n60667 );
buf ( n63036 , n63035 );
buf ( n63037 , n63036 );
not ( n13653 , n60210 );
nand ( n63039 , n57057 , n57031 );
not ( n63040 , n63039 );
nand ( n13656 , n63040 , n12154 , n61520 );
and ( n13657 , n12147 , n63039 );
nand ( n63043 , n12153 , n13657 );
and ( n63044 , n63039 , n61520 );
not ( n63045 , n63039 );
not ( n13661 , n12147 );
nand ( n13662 , n13661 , n61520 );
and ( n63048 , n63045 , n13662 );
or ( n13664 , n63044 , n63048 );
nand ( n13665 , n13656 , n63043 , n13664 );
xor ( n63051 , n13653 , n13665 );
buf ( n63052 , n63051 );
xor ( n63053 , n63037 , n63052 );
buf ( n63054 , n60498 );
not ( n13670 , n63054 );
xor ( n63056 , n11081 , n11094 );
buf ( n63057 , n63056 );
buf ( n63058 , n63057 );
not ( n63059 , n63058 );
or ( n63060 , n13670 , n63059 );
buf ( n63061 , n12097 );
buf ( n63062 , n60476 );
nand ( n63063 , n63061 , n63062 );
buf ( n63064 , n63063 );
buf ( n63065 , n63064 );
nand ( n63066 , n63060 , n63065 );
buf ( n63067 , n63066 );
buf ( n63068 , n63067 );
xor ( n13684 , n63053 , n63068 );
buf ( n63070 , n13684 );
not ( n63071 , n63070 );
not ( n13687 , n11333 );
not ( n63073 , n12117 );
or ( n63074 , n13687 , n63073 );
buf ( n63075 , n10005 );
buf ( n63076 , n380 );
nand ( n63077 , n63075 , n63076 );
buf ( n63078 , n63077 );
nand ( n13694 , n63074 , n63078 );
xor ( n13695 , n10831 , n12159 );
and ( n63081 , n13695 , n61543 );
and ( n63082 , n10831 , n12159 );
or ( n63083 , n63081 , n63082 );
xor ( n63084 , n13694 , n63083 );
xor ( n13699 , n61465 , n61482 );
and ( n63086 , n13699 , n61494 );
and ( n63087 , n61465 , n61482 );
or ( n13702 , n63086 , n63087 );
buf ( n63089 , n13702 );
xnor ( n13704 , n63084 , n63089 );
not ( n13705 , n13704 );
not ( n13706 , n13705 );
or ( n63093 , n63071 , n13706 );
not ( n63094 , n63070 );
nand ( n13709 , n63094 , n13704 );
nand ( n63096 , n63093 , n13709 );
buf ( n63097 , n61517 );
not ( n13712 , n63097 );
buf ( n63099 , n13712 );
buf ( n63100 , n63099 );
not ( n13715 , n63100 );
buf ( n63102 , n61550 );
not ( n63103 , n63102 );
buf ( n63104 , n63103 );
buf ( n63105 , n63104 );
not ( n63106 , n63105 );
or ( n13721 , n13715 , n63106 );
buf ( n63108 , n61544 );
not ( n13723 , n63108 );
buf ( n63110 , n13723 );
buf ( n63111 , n63110 );
nand ( n63112 , n13721 , n63111 );
buf ( n63113 , n63112 );
nand ( n63114 , n61517 , n61550 );
nand ( n63115 , n63113 , n63114 );
not ( n63116 , n63115 );
and ( n13726 , n63096 , n63116 );
not ( n63118 , n63096 );
nand ( n13728 , n63113 , n63114 );
and ( n63120 , n63118 , n13728 );
nor ( n13730 , n13726 , n63120 );
xor ( n13731 , n61497 , n61502 );
and ( n13732 , n13731 , n61552 );
and ( n13733 , n61497 , n61502 );
or ( n13734 , n13732 , n13733 );
buf ( n63126 , n13734 );
buf ( n63127 , n63126 );
not ( n63128 , n63127 );
buf ( n63129 , n63128 );
nand ( n13739 , n13730 , n63129 );
buf ( n63131 , n57120 );
buf ( n63132 , n59303 );
nand ( n63133 , n63131 , n63132 );
buf ( n63134 , n63133 );
not ( n63135 , n63134 );
and ( n13745 , n10879 , n63135 );
not ( n63137 , n10879 );
and ( n13747 , n63137 , n63134 );
nor ( n63139 , n13745 , n13747 );
xor ( n63140 , n10914 , n63139 );
and ( n13750 , n11328 , n378 );
and ( n63142 , n63140 , n13750 );
and ( n63143 , n10914 , n63139 );
or ( n13753 , n63142 , n63143 );
not ( n63145 , n13753 );
xor ( n63146 , n60470 , n60474 );
xor ( n13756 , n63146 , n60505 );
not ( n13757 , n13756 );
nand ( n63149 , n63145 , n13757 );
not ( n13759 , n63149 );
and ( n13760 , n13653 , n13665 );
buf ( n63152 , n13760 );
not ( n63153 , n63152 );
buf ( n63154 , n60498 );
not ( n63155 , n63154 );
buf ( n63156 , n60494 );
not ( n63157 , n63156 );
or ( n63158 , n63155 , n63157 );
buf ( n63159 , n63057 );
buf ( n63160 , n60476 );
nand ( n63161 , n63159 , n63160 );
buf ( n63162 , n63161 );
buf ( n63163 , n63162 );
nand ( n63164 , n63158 , n63163 );
buf ( n63165 , n63164 );
not ( n63166 , n63165 );
or ( n63167 , n63153 , n63166 );
or ( n13777 , n63165 , n63152 );
xor ( n63169 , n10914 , n63139 );
xor ( n13779 , n63169 , n13750 );
buf ( n13780 , n13779 );
nand ( n63172 , n13777 , n13780 );
nand ( n63173 , n63167 , n63172 );
not ( n13783 , n63173 );
or ( n13784 , n13759 , n13783 );
nand ( n63176 , n13753 , n13756 );
nand ( n63177 , n13784 , n63176 );
not ( n13787 , n63177 );
not ( n13788 , n60450 );
not ( n13789 , n60512 );
or ( n63181 , n13788 , n13789 );
nand ( n63182 , n60296 , n60451 );
nand ( n13792 , n63181 , n63182 );
or ( n13793 , n11134 , n13792 );
nand ( n63185 , n13792 , n11134 );
nand ( n63186 , n13793 , n63185 );
not ( n13796 , n63186 );
nand ( n63188 , n13787 , n13796 );
not ( n63189 , n13753 );
xor ( n13799 , n63189 , n63173 );
xnor ( n63191 , n13799 , n13757 );
xor ( n63192 , n63037 , n63052 );
and ( n13802 , n63192 , n63068 );
and ( n13803 , n63037 , n63052 );
or ( n63195 , n13802 , n13803 );
buf ( n63196 , n63195 );
buf ( n63197 , n63196 );
not ( n63198 , n63197 );
buf ( n63199 , n63198 );
not ( n13809 , n63199 );
buf ( n63201 , n13694 );
not ( n63202 , n63201 );
buf ( n63203 , n63202 );
buf ( n63204 , n63203 );
buf ( n63205 , n63083 );
nand ( n13815 , n63204 , n63205 );
buf ( n13816 , n13815 );
buf ( n63208 , n13816 );
not ( n63209 , n63208 );
buf ( n63210 , n63089 );
not ( n13820 , n63210 );
or ( n63212 , n63209 , n13820 );
buf ( n63213 , n63203 );
buf ( n63214 , n63083 );
or ( n63215 , n63213 , n63214 );
buf ( n63216 , n63215 );
buf ( n63217 , n63216 );
nand ( n63218 , n63212 , n63217 );
buf ( n63219 , n63218 );
not ( n63220 , n63219 );
not ( n13830 , n63220 );
or ( n63222 , n13809 , n13830 );
xor ( n63223 , n13779 , n63152 );
xor ( n63224 , n63223 , n63165 );
nand ( n13834 , n63222 , n63224 );
buf ( n63226 , n63219 );
buf ( n13836 , n63196 );
nand ( n13837 , n63226 , n13836 );
buf ( n63229 , n13837 );
nand ( n63230 , n63191 , n13834 , n63229 );
xor ( n13840 , n63196 , n63224 );
xor ( n13841 , n13840 , n63220 );
not ( n63233 , n63114 );
not ( n63234 , n63113 );
or ( n13844 , n63233 , n63234 );
buf ( n63236 , n13704 );
nand ( n13846 , n13844 , n63236 );
buf ( n63238 , n63115 );
buf ( n63239 , n63236 );
or ( n63240 , n63238 , n63239 );
buf ( n63241 , n63070 );
nand ( n13851 , n63240 , n63241 );
buf ( n13852 , n13851 );
nand ( n63244 , n13841 , n13846 , n13852 );
and ( n13854 , n13739 , n63188 , n63230 , n63244 );
nand ( n13855 , n12535 , n13649 , n13854 );
not ( n13856 , n13855 );
not ( n63248 , n13856 );
or ( n63249 , n11244 , n63248 );
buf ( n63250 , n61149 );
buf ( n63251 , n61450 );
nand ( n13861 , n63250 , n63251 );
buf ( n63253 , n13861 );
xor ( n63254 , n11780 , n61433 );
xor ( n13864 , n63254 , n61446 );
buf ( n63256 , n13864 );
buf ( n63257 , n63256 );
buf ( n63258 , n61597 );
nand ( n63259 , n63257 , n63258 );
buf ( n63260 , n63259 );
buf ( n13870 , n61461 );
buf ( n63262 , n61554 );
nand ( n63263 , n13870 , n63262 );
buf ( n63264 , n63263 );
and ( n13874 , n63253 , n63260 , n63264 );
not ( n63266 , n61605 );
not ( n63267 , n12224 );
or ( n13877 , n63266 , n63267 );
buf ( n63269 , n12236 );
buf ( n63270 , n61905 );
and ( n63271 , n63269 , n63270 );
buf ( n63272 , n63271 );
nand ( n63273 , n13877 , n63272 );
nand ( n63274 , n13874 , n63273 );
not ( n13884 , n61461 );
nand ( n63276 , n13884 , n12181 );
nand ( n63277 , n63276 , n63244 , n63188 );
nand ( n13887 , n63229 , n13834 , n63191 );
nand ( n63279 , n13739 , n13887 );
nor ( n63280 , n63277 , n63279 );
nand ( n13890 , n63264 , n61453 );
nand ( n63282 , n63274 , n63280 , n13890 );
not ( n63283 , n63282 );
buf ( n63284 , n13852 );
buf ( n63285 , n13846 );
nand ( n13895 , n63284 , n63285 );
buf ( n63287 , n13895 );
buf ( n63288 , n63287 );
buf ( n63289 , n13841 );
not ( n63290 , n63289 );
buf ( n63291 , n63290 );
buf ( n63292 , n63291 );
nor ( n13902 , n63288 , n63292 );
buf ( n63294 , n13902 );
not ( n13904 , n63229 );
not ( n13905 , n13834 );
or ( n63297 , n13904 , n13905 );
not ( n13907 , n63191 );
nand ( n63299 , n63297 , n13907 );
and ( n63300 , n63294 , n63299 );
nand ( n13910 , n63188 , n13887 );
nor ( n63302 , n63300 , n13910 );
not ( n13912 , n63302 );
not ( n13913 , n13730 );
nand ( n13914 , n13913 , n63126 );
buf ( n63306 , n63287 );
buf ( n13916 , n63291 );
nand ( n13917 , n63306 , n13916 );
buf ( n13918 , n13917 );
nand ( n63310 , n13914 , n13918 , n63299 );
not ( n13920 , n63310 );
or ( n13921 , n13912 , n13920 );
not ( n13922 , n11242 );
buf ( n63314 , n60594 );
buf ( n63315 , n11190 );
nor ( n63316 , n63314 , n63315 );
buf ( n63317 , n63316 );
nand ( n63318 , n63317 , n60516 );
buf ( n63319 , n60579 );
buf ( n63320 , n11217 );
nand ( n13930 , n63319 , n63320 );
buf ( n13931 , n13930 );
nor ( n13932 , n10790 , n60165 );
nor ( n13933 , n60159 , n60168 );
or ( n63325 , n13932 , n13933 );
nand ( n13935 , n63325 , n10859 );
nand ( n63327 , n63318 , n13931 , n13935 );
not ( n13937 , n63327 );
not ( n63329 , n10861 );
or ( n13939 , n13937 , n63329 );
not ( n63331 , n10716 );
nand ( n13941 , n63331 , n10787 );
nand ( n13942 , n13939 , n13941 );
not ( n63334 , n13942 );
or ( n13944 , n13922 , n63334 );
not ( n63336 , n11241 );
nand ( n13946 , n63336 , n60609 );
nand ( n63338 , n13944 , n13946 );
nand ( n63339 , n63177 , n63186 );
not ( n13949 , n63339 );
nor ( n63341 , n63338 , n13949 );
nand ( n63342 , n13921 , n63341 );
or ( n13952 , n63283 , n63342 );
or ( n63344 , n11243 , n63338 );
nand ( n13954 , n13952 , n63344 );
nand ( n63346 , n63249 , n13954 );
not ( n63347 , n63346 );
or ( n63348 , n10701 , n63347 );
nand ( n63349 , n10689 , n10663 );
not ( n63350 , n63349 );
not ( n63351 , n63350 );
not ( n63352 , n10699 );
not ( n13959 , n10611 );
and ( n63354 , n10525 , n59945 );
not ( n63355 , n63354 );
or ( n13962 , n13959 , n63355 );
not ( n63357 , n59984 );
nand ( n63358 , n63357 , n10600 );
nand ( n63359 , n13962 , n63358 );
not ( n13966 , n63359 );
or ( n63361 , n63352 , n13966 );
or ( n63362 , n10692 , n10698 );
nand ( n63363 , n63361 , n63362 );
not ( n63364 , n63363 );
or ( n13971 , n63351 , n63364 );
not ( n63366 , n60046 );
buf ( n63367 , n60062 );
not ( n63368 , n63367 );
not ( n13975 , n60015 );
or ( n13976 , n59504 , n10121 , n10661 );
nand ( n13977 , n59504 , n10121 , n10658 );
nand ( n63372 , n13976 , n13977 );
not ( n13979 , n63372 );
or ( n63374 , n13975 , n13979 );
not ( n63375 , n10661 );
nand ( n13982 , n63375 , n10638 , n60011 );
nand ( n13983 , n63374 , n13982 );
not ( n63378 , n13983 );
not ( n13985 , n60010 );
or ( n63380 , n63378 , n13985 );
not ( n13987 , n10635 );
not ( n63382 , n10624 );
or ( n63383 , n63382 , n59556 );
nand ( n63384 , n63382 , n59556 );
nand ( n63385 , n13987 , n63383 , n63384 );
nand ( n13992 , n63380 , n63385 );
buf ( n63387 , n13992 );
not ( n63388 , n63387 );
or ( n13995 , n63368 , n63388 );
buf ( n63390 , n59567 );
not ( n63391 , n63390 );
buf ( n63392 , n63391 );
buf ( n63393 , n63392 );
buf ( n14000 , n60057 );
nand ( n14001 , n63393 , n14000 );
buf ( n63396 , n14001 );
buf ( n63397 , n63396 );
nand ( n14004 , n13995 , n63397 );
buf ( n63399 , n14004 );
not ( n14006 , n63399 );
or ( n14007 , n63366 , n14006 );
nand ( n63402 , n63392 , n10667 );
nand ( n14009 , n14007 , n63402 );
not ( n63404 , n14009 );
nand ( n14011 , n13971 , n63404 );
not ( n14012 , n14011 );
nand ( n63407 , n63348 , n14012 );
not ( n63408 , n63407 );
or ( n14015 , n10441 , n63408 );
buf ( n63410 , n63392 );
buf ( n63411 , n10435 );
nand ( n14018 , n63410 , n63411 );
buf ( n63413 , n14018 );
buf ( n63414 , n63413 );
buf ( n14021 , n63414 );
buf ( n63416 , n14021 );
nand ( n14023 , n14015 , n63416 );
buf ( n63418 , n14023 );
and ( n14025 , n63418 , n59805 );
not ( n14026 , n63418 );
and ( n14027 , n14026 , n59801 );
nor ( n14028 , n14025 , n14027 );
buf ( n63423 , n14028 );
buf ( n63424 , n60046 );
buf ( n63425 , n63402 );
nand ( n14032 , n63424 , n63425 );
buf ( n63427 , n14032 );
buf ( n63428 , n63427 );
buf ( n63429 , n63427 );
not ( n63430 , n63429 );
buf ( n63431 , n63430 );
buf ( n63432 , n63431 );
buf ( n63433 , n60062 );
not ( n14040 , n63433 );
buf ( n63435 , n10663 );
not ( n14042 , n63435 );
nand ( n14043 , n10699 , n59988 );
buf ( n63438 , n14043 );
nor ( n14045 , n14042 , n63438 );
buf ( n63440 , n14045 );
not ( n14047 , n63440 );
not ( n14048 , n63346 );
or ( n14049 , n14047 , n14048 );
buf ( n63444 , n10663 );
not ( n14051 , n63444 );
buf ( n63446 , n63363 );
not ( n14053 , n63446 );
or ( n63448 , n14051 , n14053 );
buf ( n63449 , n13992 );
not ( n63450 , n63449 );
buf ( n63451 , n63450 );
buf ( n63452 , n63451 );
nand ( n63453 , n63448 , n63452 );
buf ( n63454 , n63453 );
buf ( n63455 , n63454 );
not ( n63456 , n63455 );
buf ( n63457 , n63456 );
nand ( n14060 , n14049 , n63457 );
buf ( n63459 , n14060 );
not ( n14062 , n63459 );
or ( n14063 , n14040 , n14062 );
buf ( n63462 , n63396 );
nand ( n14065 , n14063 , n63462 );
buf ( n63464 , n14065 );
buf ( n63465 , n63464 );
and ( n14068 , n63465 , n63432 );
not ( n14069 , n63465 );
and ( n63468 , n14069 , n63428 );
nor ( n63469 , n14068 , n63468 );
buf ( n63470 , n63469 );
buf ( n63471 , n59570 );
buf ( n63472 , n10202 );
buf ( n63473 , n59797 );
buf ( n63474 , n59814 );
and ( n63475 , n63473 , n63474 );
buf ( n63476 , n63475 );
buf ( n63477 , n63476 );
buf ( n63478 , n59570 );
buf ( n63479 , n10413 );
buf ( n63480 , n59615 );
and ( n63481 , n63479 , n63480 );
buf ( n63482 , n59609 );
nor ( n63483 , n63481 , n63482 );
buf ( n63484 , n63483 );
buf ( n63485 , n55731 );
buf ( n63486 , n6530 );
nand ( n63487 , n63485 , n63486 );
buf ( n63488 , n63487 );
xor ( n63489 , n63484 , n63488 );
buf ( n63490 , n63489 );
nand ( n63491 , n63478 , n63490 );
buf ( n63492 , n63491 );
buf ( n63493 , n63492 );
nand ( n63494 , n63477 , n63493 );
buf ( n63495 , n63494 );
buf ( n63496 , n63495 );
buf ( n63497 , n63349 );
nor ( n14072 , n63496 , n63497 );
buf ( n63499 , n14072 );
not ( n14074 , n63499 );
not ( n14075 , n11243 );
not ( n14076 , n13856 );
or ( n14077 , n14075 , n14076 );
nand ( n63504 , n14077 , n13954 );
buf ( n63505 , n14043 );
not ( n14080 , n63505 );
buf ( n63507 , n14080 );
and ( n14082 , n63504 , n63507 );
not ( n63509 , n14082 );
or ( n63510 , n14074 , n63509 );
not ( n63511 , n63476 );
not ( n14086 , n14011 );
or ( n63513 , n63511 , n14086 );
buf ( n63514 , n59791 );
buf ( n63515 , n63413 );
and ( n14090 , n63514 , n63515 );
buf ( n63517 , n14090 );
nand ( n14092 , n63513 , n63517 );
buf ( n63519 , n14092 );
buf ( n63520 , n63492 );
and ( n14095 , n63519 , n63520 );
buf ( n63522 , n63489 );
buf ( n63523 , n59570 );
nor ( n14098 , n63522 , n63523 );
buf ( n14099 , n14098 );
buf ( n63526 , n14099 );
nor ( n14101 , n14095 , n63526 );
buf ( n63528 , n14101 );
nand ( n14103 , n63510 , n63528 );
buf ( n63530 , n14103 );
and ( n63531 , n63530 , n63472 );
not ( n14106 , n63530 );
and ( n63533 , n14106 , n63471 );
nor ( n63534 , n63531 , n63533 );
buf ( n63535 , n63534 );
buf ( n63536 , n10699 );
buf ( n63537 , n63362 );
nand ( n14112 , n63536 , n63537 );
buf ( n63539 , n14112 );
buf ( n63540 , n63539 );
buf ( n63541 , n63539 );
not ( n63542 , n63541 );
buf ( n63543 , n63542 );
buf ( n63544 , n63543 );
not ( n14119 , n59988 );
not ( n14120 , n63346 );
or ( n63547 , n14119 , n14120 );
buf ( n14122 , n63359 );
not ( n63549 , n14122 );
buf ( n63550 , n63549 );
nand ( n63551 , n63547 , n63550 );
buf ( n63552 , n63551 );
and ( n63553 , n63552 , n63544 );
not ( n14128 , n63552 );
and ( n63555 , n14128 , n63540 );
nor ( n63556 , n63553 , n63555 );
buf ( n63557 , n63556 );
buf ( n63558 , n63358 );
buf ( n63559 , n10611 );
nand ( n14134 , n63558 , n63559 );
buf ( n63561 , n14134 );
buf ( n63562 , n63561 );
buf ( n14137 , n63561 );
not ( n63564 , n14137 );
buf ( n63565 , n63564 );
buf ( n63566 , n63565 );
buf ( n63567 , n10577 );
not ( n63568 , n63567 );
buf ( n63569 , n63504 );
not ( n63570 , n63569 );
or ( n63571 , n63568 , n63570 );
not ( n63572 , n63354 );
buf ( n63573 , n63572 );
nand ( n63574 , n63571 , n63573 );
buf ( n63575 , n63574 );
buf ( n63576 , n63575 );
and ( n63577 , n63576 , n63566 );
not ( n14152 , n63576 );
and ( n63579 , n14152 , n63562 );
nor ( n14154 , n63577 , n63579 );
buf ( n63581 , n14154 );
buf ( n63582 , n13946 );
buf ( n63583 , n11242 );
nand ( n14158 , n63582 , n63583 );
buf ( n63585 , n14158 );
buf ( n63586 , n63585 );
buf ( n14161 , n63585 );
not ( n14162 , n14161 );
buf ( n14163 , n14162 );
buf ( n63590 , n14163 );
buf ( n63591 , n60603 );
not ( n14166 , n63591 );
not ( n14167 , n63283 );
buf ( n14168 , n13856 );
not ( n14169 , n14168 );
buf ( n14170 , n14169 );
not ( n63597 , n63310 );
not ( n14172 , n63302 );
or ( n63599 , n63597 , n14172 );
nand ( n63600 , n63599 , n63339 );
buf ( n63601 , n63600 );
not ( n14176 , n63601 );
buf ( n63603 , n14176 );
nand ( n14178 , n14167 , n14170 , n63603 );
buf ( n63605 , n14178 );
not ( n14180 , n63605 );
or ( n63607 , n14166 , n14180 );
buf ( n14182 , n13942 );
not ( n14183 , n14182 );
buf ( n14184 , n14183 );
buf ( n63611 , n14184 );
nand ( n14186 , n63607 , n63611 );
buf ( n63613 , n14186 );
buf ( n63614 , n63613 );
and ( n14189 , n63614 , n63590 );
not ( n14190 , n63614 );
and ( n14191 , n14190 , n63586 );
nor ( n14192 , n14189 , n14191 );
buf ( n63619 , n14192 );
buf ( n63620 , n60597 );
buf ( n63621 , n13931 );
nand ( n14196 , n63620 , n63621 );
buf ( n63623 , n14196 );
buf ( n63624 , n63623 );
buf ( n63625 , n63623 );
not ( n63626 , n63625 );
buf ( n63627 , n63626 );
buf ( n14202 , n63627 );
not ( n14203 , n11191 );
not ( n63630 , n14178 );
or ( n63631 , n14203 , n63630 );
not ( n14206 , n11190 );
nand ( n63633 , n14206 , n60516 );
nand ( n63634 , n63631 , n63633 );
buf ( n63635 , n63634 );
and ( n63636 , n63635 , n14202 );
not ( n14211 , n63635 );
and ( n63638 , n14211 , n63624 );
nor ( n14213 , n63636 , n63638 );
buf ( n63640 , n14213 );
buf ( n63641 , n63294 );
buf ( n14216 , n63641 );
buf ( n14217 , n14216 );
buf ( n63644 , n14217 );
not ( n14219 , n63644 );
buf ( n63646 , n13918 );
nand ( n63647 , n14219 , n63646 );
buf ( n63648 , n63647 );
buf ( n63649 , n63648 );
buf ( n63650 , n63648 );
not ( n14225 , n63650 );
buf ( n14226 , n14225 );
buf ( n63653 , n14226 );
buf ( n63654 , n13739 );
buf ( n63655 , n63654 );
not ( n63656 , n63655 );
buf ( n63657 , n63260 );
buf ( n63658 , n63657 );
buf ( n63659 , n63658 );
and ( n63660 , n63273 , n63659 );
buf ( n63661 , n63253 );
buf ( n63662 , n63661 );
buf ( n14237 , n63662 );
buf ( n63664 , n14237 );
buf ( n63665 , n63264 );
nand ( n14240 , n63660 , n63664 , n63665 );
buf ( n63667 , n63276 );
nand ( n63668 , n63667 , n13890 );
not ( n63669 , n63668 );
nand ( n63670 , n14240 , n63669 );
not ( n14245 , n61461 );
not ( n14246 , n61554 );
and ( n14247 , n14245 , n14246 );
nor ( n14248 , n14247 , n61453 );
and ( n14249 , n61911 , n61608 );
nand ( n63676 , n14248 , n14249 , n13649 );
nand ( n14251 , n63670 , n63676 );
buf ( n63678 , n14251 );
not ( n63679 , n63678 );
or ( n63680 , n63656 , n63679 );
buf ( n63681 , n13914 );
buf ( n14256 , n63681 );
buf ( n63683 , n14256 );
buf ( n63684 , n63683 );
nand ( n14259 , n63680 , n63684 );
buf ( n63686 , n14259 );
buf ( n63687 , n63686 );
and ( n14262 , n63687 , n63653 );
not ( n14263 , n63687 );
and ( n14264 , n14263 , n63649 );
nor ( n14265 , n14262 , n14264 );
buf ( n63692 , n14265 );
nand ( n14267 , n63299 , n63230 );
buf ( n63694 , n14267 );
buf ( n63695 , n14267 );
not ( n14270 , n63695 );
buf ( n63697 , n14270 );
buf ( n63698 , n63697 );
not ( n14273 , n63654 );
nor ( n14274 , n14273 , n14217 );
not ( n14275 , n14274 );
not ( n14276 , n14251 );
or ( n14277 , n14275 , n14276 );
not ( n14278 , n14217 );
buf ( n63705 , n13918 );
buf ( n63706 , n63683 );
nand ( n14281 , n63705 , n63706 );
buf ( n63708 , n14281 );
nand ( n14283 , n14278 , n63708 );
nand ( n14284 , n14277 , n14283 );
buf ( n63711 , n14284 );
and ( n14286 , n63711 , n63698 );
not ( n14287 , n63711 );
and ( n14288 , n14287 , n63694 );
nor ( n14289 , n14286 , n14288 );
buf ( n63716 , n14289 );
buf ( n63717 , n10577 );
buf ( n63718 , n63572 );
nand ( n14293 , n63717 , n63718 );
buf ( n63720 , n14293 );
buf ( n63721 , n63720 );
buf ( n63722 , n63504 );
buf ( n63723 , n63722 );
buf ( n63724 , n63723 );
buf ( n63725 , n63724 );
buf ( n63726 , n63720 );
buf ( n63727 , n63724 );
not ( n14302 , n63721 );
not ( n63729 , n63725 );
or ( n14304 , n14302 , n63729 );
or ( n14305 , n63726 , n63727 );
nand ( n14306 , n14304 , n14305 );
buf ( n63733 , n14306 );
buf ( n63734 , n63667 );
buf ( n63735 , n63665 );
nand ( n14310 , n63734 , n63735 );
buf ( n63737 , n14310 );
buf ( n63738 , n63737 );
buf ( n63739 , n63737 );
not ( n14314 , n63739 );
buf ( n63741 , n14314 );
buf ( n63742 , n63741 );
buf ( n63743 , n61456 );
not ( n14318 , n63743 );
not ( n63745 , n14249 );
not ( n14319 , n13632 );
not ( n14320 , n13582 );
or ( n63748 , n14319 , n14320 );
nand ( n63749 , n63748 , n13648 );
not ( n63750 , n63749 );
or ( n63751 , n63745 , n63750 );
nand ( n63752 , n63751 , n63660 );
buf ( n63753 , n63752 );
not ( n63754 , n63753 );
or ( n63755 , n14318 , n63754 );
buf ( n63756 , n63664 );
nand ( n63757 , n63755 , n63756 );
buf ( n63758 , n63757 );
buf ( n63759 , n63758 );
and ( n63760 , n63759 , n63742 );
not ( n63761 , n63759 );
and ( n63762 , n63761 , n63738 );
nor ( n63763 , n63760 , n63762 );
buf ( n63764 , n63763 );
buf ( n63765 , n61456 );
buf ( n63766 , n63664 );
nand ( n14321 , n63765 , n63766 );
buf ( n63768 , n14321 );
buf ( n63769 , n63768 );
buf ( n14324 , n63768 );
not ( n14325 , n14324 );
buf ( n63772 , n14325 );
buf ( n63773 , n63772 );
buf ( n63774 , n63752 );
and ( n14329 , n63774 , n63773 );
not ( n14330 , n63774 );
and ( n14331 , n14330 , n63769 );
nor ( n14332 , n14329 , n14331 );
buf ( n63779 , n14332 );
buf ( n63780 , n61605 );
buf ( n63781 , n12224 );
nand ( n14336 , n63780 , n63781 );
buf ( n63783 , n14336 );
buf ( n63784 , n63783 );
buf ( n63785 , n63659 );
nand ( n14340 , n63784 , n63785 );
buf ( n63787 , n14340 );
buf ( n63788 , n63787 );
buf ( n63789 , n63787 );
not ( n14344 , n63789 );
buf ( n14345 , n14344 );
buf ( n63792 , n14345 );
buf ( n63793 , n61911 );
not ( n14347 , n63793 );
buf ( n63795 , n63749 );
not ( n14349 , n63795 );
or ( n14350 , n14347 , n14349 );
buf ( n14351 , n63272 );
not ( n14352 , n14351 );
buf ( n63800 , n14352 );
nand ( n14354 , n14350 , n63800 );
buf ( n63802 , n14354 );
buf ( n63803 , n63802 );
and ( n63804 , n63803 , n63792 );
not ( n63805 , n63803 );
and ( n63806 , n63805 , n63788 );
nor ( n14360 , n63804 , n63806 );
buf ( n14361 , n14360 );
nand ( n63809 , n62964 , n12947 );
buf ( n63810 , n63809 );
buf ( n63811 , n63809 );
not ( n63812 , n63811 );
buf ( n63813 , n63812 );
buf ( n63814 , n63813 );
buf ( n63815 , n12896 );
buf ( n63816 , n63815 );
buf ( n63817 , n63816 );
buf ( n63818 , n63817 );
not ( n63819 , n63818 );
not ( n63820 , n62882 );
not ( n63821 , n62939 );
or ( n63822 , n63820 , n63821 );
nand ( n63823 , n63822 , n13571 );
buf ( n63824 , n63823 );
not ( n63825 , n63824 );
or ( n63826 , n63819 , n63825 );
not ( n63827 , n13575 );
buf ( n63828 , n63827 );
nand ( n63829 , n63826 , n63828 );
buf ( n63830 , n63829 );
buf ( n63831 , n63830 );
and ( n63832 , n63831 , n63814 );
not ( n63833 , n63831 );
and ( n63834 , n63833 , n63810 );
nor ( n63835 , n63832 , n63834 );
buf ( n63836 , n63835 );
not ( n63837 , n63023 );
buf ( n63838 , n13631 );
nand ( n63839 , n63837 , n63838 );
buf ( n63840 , n63839 );
not ( n14369 , n63840 );
buf ( n63842 , n14369 );
nand ( n14371 , n13569 , n13540 );
buf ( n63844 , n14371 );
buf ( n63845 , n13554 );
buf ( n14374 , n63845 );
buf ( n63847 , n14374 );
buf ( n63848 , n63847 );
not ( n63849 , n63848 );
buf ( n63850 , n62882 );
buf ( n63851 , n63850 );
buf ( n63852 , n63851 );
buf ( n63853 , n63852 );
not ( n63854 , n63853 );
or ( n63855 , n63849 , n63854 );
buf ( n63856 , n62945 );
not ( n63857 , n63856 );
buf ( n63858 , n63857 );
buf ( n63859 , n63858 );
nand ( n63860 , n63855 , n63859 );
buf ( n63861 , n63860 );
buf ( n63862 , n63861 );
buf ( n63863 , n14371 );
buf ( n63864 , n63861 );
not ( n63865 , n63844 );
not ( n63866 , n63862 );
or ( n63867 , n63865 , n63866 );
or ( n63868 , n63863 , n63864 );
nand ( n63869 , n63867 , n63868 );
buf ( n63870 , n63869 );
buf ( n63871 , n63858 );
buf ( n63872 , n63847 );
nand ( n63873 , n63871 , n63872 );
buf ( n63874 , n63873 );
buf ( n63875 , n63874 );
buf ( n63876 , n63852 );
buf ( n63877 , n63874 );
buf ( n63878 , n63852 );
not ( n63879 , n63875 );
not ( n63880 , n63876 );
or ( n14394 , n63879 , n63880 );
or ( n63882 , n63877 , n63878 );
nand ( n63883 , n14394 , n63882 );
buf ( n63884 , n63883 );
buf ( n63885 , n14099 );
not ( n63886 , n63885 );
buf ( n63887 , n63492 );
nand ( n63888 , n63886 , n63887 );
buf ( n63889 , n63888 );
buf ( n63890 , n63889 );
not ( n14399 , n63890 );
buf ( n14400 , n14399 );
buf ( n14401 , n13407 );
buf ( n14402 , n14401 );
buf ( n14403 , n14402 );
buf ( n63896 , n14403 );
buf ( n14405 , n62801 );
buf ( n14406 , n62673 );
nand ( n14407 , n14405 , n14406 );
buf ( n14408 , n14407 );
buf ( n63901 , n14408 );
buf ( n63902 , n14403 );
buf ( n63903 , n14408 );
not ( n63904 , n63896 );
not ( n63905 , n63901 );
or ( n14414 , n63904 , n63905 );
or ( n63907 , n63902 , n63903 );
nand ( n63908 , n14414 , n63907 );
buf ( n63909 , n63908 );
not ( n63910 , n13983 );
nand ( n63911 , n63910 , n60036 );
buf ( n63912 , n63911 );
not ( n63913 , n63912 );
buf ( n63914 , n63913 );
xor ( n63915 , n13295 , n62694 );
xor ( n14421 , n63915 , n62740 );
buf ( n63917 , n14421 );
xor ( n63918 , n62716 , n13339 );
xor ( n63919 , n63918 , n62735 );
buf ( n63920 , n63919 );
buf ( n63921 , n59814 );
buf ( n63922 , n63416 );
nand ( n63923 , n63921 , n63922 );
buf ( n63924 , n63923 );
buf ( n63925 , n62778 );
buf ( n63926 , n62769 );
and ( n14432 , n63925 , n63926 );
buf ( n63928 , n14432 );
buf ( n63929 , n63928 );
buf ( n63930 , n62744 );
xor ( n63931 , n63929 , n63930 );
buf ( n63932 , n63931 );
not ( n14438 , n63363 );
and ( n63934 , n60609 , n59945 );
not ( n63935 , n60609 );
and ( n14441 , n63935 , n59948 );
nor ( n63937 , n63934 , n14441 );
and ( n63938 , n63504 , n63937 );
not ( n63939 , n63504 );
not ( n14445 , n63937 );
and ( n63941 , n63939 , n14445 );
nor ( n63942 , n63938 , n63941 );
buf ( n14448 , n63942 );
and ( n63944 , n13931 , n63318 );
nand ( n63945 , n63339 , n63188 );
not ( n63946 , n63945 );
not ( n63947 , n63676 );
buf ( n63948 , n13854 );
not ( n63949 , n63948 );
buf ( n63950 , n60600 );
nor ( n63951 , n63949 , n63950 );
buf ( n63952 , n63951 );
buf ( n63953 , n10860 );
not ( n63954 , n63953 );
nand ( n63955 , n63947 , n63952 , n63954 );
not ( n63956 , n63274 );
nor ( n14457 , n63956 , n63668 );
nand ( n63958 , n63954 , n63952 , n14457 );
not ( n63959 , n60600 );
nand ( n63960 , n63954 , n63600 , n63959 );
not ( n63961 , n13935 );
nor ( n63962 , n63944 , n63953 );
nor ( n63963 , n63961 , n63962 );
nand ( n14462 , n63955 , n63958 , n63960 , n63963 );
not ( n63965 , n10788 );
not ( n14464 , n10716 );
or ( n14465 , n63965 , n14464 );
nand ( n63968 , n14465 , n13941 );
not ( n14467 , n63968 );
and ( n14468 , n14462 , n14467 );
not ( n63971 , n14462 );
and ( n63972 , n63971 , n63968 );
nor ( n63973 , n14468 , n63972 );
not ( n14472 , n14457 );
not ( n63975 , n63947 );
and ( n63976 , n14472 , n63975 );
not ( n63977 , n63952 );
nor ( n14476 , n63976 , n63977 );
not ( n63979 , n63476 );
not ( n63980 , n63407 );
or ( n63981 , n63979 , n63980 );
nand ( n14480 , n63981 , n63517 );
and ( n63983 , n14480 , n14400 );
not ( n63984 , n14480 );
and ( n63985 , n63984 , n63889 );
nor ( n14484 , n63983 , n63985 );
not ( n14485 , n63945 );
nand ( n63988 , n14485 , n63299 );
or ( n14487 , n14284 , n63988 );
not ( n14488 , n13887 );
nor ( n63991 , n14488 , n63946 );
nand ( n14490 , n14284 , n63991 );
not ( n14491 , n63946 );
not ( n14492 , n63299 );
and ( n14493 , n14491 , n14492 );
nor ( n14494 , n63945 , n13887 );
and ( n14495 , n14494 , n63299 );
nor ( n63998 , n14493 , n14495 );
nand ( n63999 , n14487 , n14490 , n63998 );
buf ( n64000 , n63407 );
not ( n14496 , n63924 );
and ( n14497 , n64000 , n14496 );
not ( n14498 , n64000 );
and ( n64004 , n14498 , n63924 );
nor ( n64005 , n14497 , n64004 );
buf ( n14501 , n13471 );
not ( n64007 , n62804 );
not ( n14503 , n13494 );
not ( n14504 , n13497 );
nand ( n14505 , n63954 , n13935 );
buf ( n64011 , n63600 );
buf ( n64012 , n63959 );
nand ( n64013 , n64011 , n64012 );
buf ( n64014 , n64013 );
nand ( n14507 , n63944 , n64014 );
or ( n14508 , n14476 , n14507 );
nand ( n14509 , n14508 , n14505 );
not ( n14510 , n14476 );
nor ( n14511 , n14507 , n14505 );
nand ( n14512 , n14510 , n14511 );
nand ( n64021 , n14509 , n14512 );
not ( n14513 , n60036 );
not ( n14514 , n63507 );
not ( n14515 , n63504 );
or ( n14516 , n14514 , n14515 );
nand ( n14517 , n14516 , n14438 );
not ( n14518 , n14517 );
or ( n14519 , n14513 , n14518 );
buf ( n14520 , n63910 );
nand ( n14521 , n14519 , n14520 );
nand ( n14522 , n63385 , n60010 );
not ( n14523 , n14522 );
and ( n64033 , n14521 , n14523 );
not ( n14524 , n14521 );
and ( n14525 , n14524 , n14522 );
nor ( n14526 , n64033 , n14525 );
and ( n14527 , n14517 , n63914 );
not ( n14528 , n14517 );
and ( n64039 , n14528 , n63911 );
nor ( n64040 , n14527 , n64039 );
not ( n64041 , n64007 );
and ( n64042 , n14501 , n62877 );
not ( n14529 , n14501 );
and ( n14530 , n14529 , n62876 );
or ( n14531 , n64042 , n14530 );
not ( n14532 , n14531 );
or ( n14533 , n64041 , n14532 );
not ( n14534 , n64007 );
and ( n14535 , n14534 , n14503 );
and ( n14536 , n14504 , n62804 );
nor ( n14537 , n14535 , n14536 );
nand ( n14538 , n14533 , n14537 );
nand ( n14539 , n63817 , n63827 );
not ( n14540 , n14539 );
nand ( n14541 , n63396 , n60062 );
not ( n14542 , n14541 );
and ( n14543 , n14060 , n14542 );
not ( n14544 , n14060 );
and ( n14545 , n14544 , n14541 );
nor ( n14546 , n14543 , n14545 );
not ( n14547 , n12949 );
not ( n14548 , n63823 );
or ( n14549 , n14547 , n14548 );
nand ( n14550 , n14549 , n62966 );
and ( n14551 , n14550 , n63838 );
nor ( n14552 , n14551 , n63023 );
nand ( n14553 , n13646 , n13615 );
and ( n14554 , n14552 , n14553 );
not ( n64069 , n14552 );
not ( n64070 , n14553 );
and ( n14555 , n64069 , n64070 );
nor ( n14556 , n14554 , n14555 );
nand ( n14557 , n14352 , n61911 );
nand ( n14558 , n63633 , n11191 );
not ( n14559 , n14558 );
and ( n14560 , n14178 , n14559 );
not ( n64077 , n14178 );
and ( n64078 , n64077 , n14558 );
nor ( n14561 , n14560 , n64078 );
xor ( n14562 , n13319 , n401 );
not ( n14563 , n14562 );
not ( n14564 , n13261 );
or ( n14565 , n14563 , n14564 );
or ( n14566 , n13261 , n14562 );
nand ( n14567 , n14565 , n14566 );
or ( n14568 , n62790 , n62788 );
xor ( n14569 , n13395 , n13397 );
and ( n14570 , n62788 , n14569 );
not ( n14571 , n62788 );
and ( n14572 , n14571 , n13398 );
nor ( n14573 , n14570 , n14572 );
nand ( n14574 , n14568 , n14573 );
and ( n14575 , n63823 , n14540 );
not ( n14576 , n63823 );
and ( n14577 , n14576 , n14539 );
nor ( n14578 , n14575 , n14577 );
nand ( n14579 , n63654 , n63683 );
not ( n14580 , n14579 );
and ( n14581 , n14251 , n14580 );
not ( n14582 , n14251 );
and ( n14583 , n14582 , n14579 );
nor ( n14584 , n14581 , n14583 );
buf ( n64103 , n63839 );
buf ( n64104 , n63842 );
buf ( n64105 , n14550 );
and ( n14588 , n64105 , n64104 );
not ( n14589 , n64105 );
and ( n14590 , n14589 , n64103 );
nor ( n14591 , n14588 , n14590 );
buf ( n64110 , n14591 );
xnor ( n14593 , n63749 , n14557 );
endmodule

