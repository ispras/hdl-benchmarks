//NOTE: no-implementation module stub

module GtCLK_OA21 (
    output Z,
    input A,
    input B,
    input C
);

endmodule
